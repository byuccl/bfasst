module top (O, I);
    input I;
    output O;

    BUFG bufg1 (O, I);

endmodule 