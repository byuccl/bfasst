// Reading file 'mem_b_extracted.asc'..

module chip (output \data_out[1] , output \data_out[0] , output \data_out[11] , output \data_out[15] , output \data_out[10] , output \data_out[17] , output \data_out[12] , output \data_out[13] , output \data_out[14] , output \data_out[16] , output \data_out[18] , output \data_out[19] , output \data_out[22] , output \data_out[2] , output \data_out[20] , output \data_out[21] , output \data_out[23] , output \data_out[24] , output \data_out[27] , output \data_out[25] , output \data_out[26] , output \data_out[29] , output \data_out[28] , output \data_out[3] , input read_clk, output \data_out[30] , input write_clk, output \data_out[31] , output \data_out[4] , output \data_out[5] , output \data_out[9] , output \data_out[6] , output \data_out[7] , output \data_out[8] , input rd_en, input \read_address[0] , input \read_address[1] , input \read_address[2] , input \read_address[3] , input \read_address[4] , input \read_address[5] , input wr_en, input \write_address[0] , input \write_address[1] , input \write_address[2] , input \write_address[3] , input \write_address[4] , input \write_address[5] , input \data_in[20] , input \data_in[0] , input \data_in[9] , input \data_in[8] , input \data_in[21] , input \data_in[7] , input \data_in[6] , input \data_in[4] , input \data_in[5] , input \data_in[22] , input \data_in[23] , input \data_in[3] , input \data_in[2] , input \data_in[25] , input \data_in[24] , input \data_in[15] , input \data_in[13] , input \data_in[26] , input \data_in[14] , input \data_in[27] , input \data_in[17] , input \data_in[19] , input \data_in[28] , input \data_in[18] , input \data_in[12] , input \data_in[11] , input \data_in[29] , input \data_in[31] , input \data_in[30] , input \data_in[16] , input \data_in[10] , input \data_in[1] , input \write_address[6] , input \read_address[6] , input \write_address[7] , input \read_address[7] );

wire \data_out[1] ;
// (0, 2, 'span4_vert_t_13')
// (0, 3, 'io_1/D_OUT_0')
// (0, 3, 'io_1/PAD')
// (0, 3, 'local_g0_5')
// (0, 3, 'span4_vert_b_13')
// (0, 4, 'span4_vert_b_9')
// (0, 5, 'span4_vert_b_5')
// (0, 6, 'span4_horz_7')
// (0, 6, 'span4_vert_b_1')
// (1, 6, 'sp4_h_r_18')
// (2, 6, 'sp4_h_r_31')
// (3, 6, 'sp4_h_r_42')
// (4, 6, 'sp4_h_l_42')
// (4, 6, 'sp4_h_r_4')
// (5, 6, 'sp4_h_r_17')
// (6, 6, 'sp4_h_r_28')
// (7, 6, 'sp4_h_r_41')
// (7, 7, 'sp4_r_v_b_47')
// (7, 8, 'sp4_r_v_b_34')
// (7, 9, 'sp4_r_v_b_23')
// (7, 10, 'sp4_r_v_b_10')
// (7, 25, 'neigh_op_tnr_6')
// (7, 26, 'neigh_op_rgt_6')
// (7, 27, 'neigh_op_bnr_6')
// (8, 6, 'sp4_h_l_41')
// (8, 6, 'sp4_v_t_47')
// (8, 7, 'sp4_v_b_47')
// (8, 8, 'sp12_v_t_23')
// (8, 8, 'sp4_v_b_34')
// (8, 9, 'sp12_v_b_23')
// (8, 9, 'sp4_v_b_23')
// (8, 10, 'sp12_v_b_20')
// (8, 10, 'sp4_v_b_10')
// (8, 11, 'sp12_v_b_19')
// (8, 12, 'sp12_v_b_16')
// (8, 13, 'sp12_v_b_15')
// (8, 14, 'sp12_v_b_12')
// (8, 15, 'sp12_v_b_11')
// (8, 16, 'sp12_v_b_8')
// (8, 17, 'sp12_v_b_7')
// (8, 18, 'sp12_v_b_4')
// (8, 19, 'sp12_v_b_3')
// (8, 20, 'sp12_v_b_0')
// (8, 20, 'sp12_v_t_23')
// (8, 21, 'sp12_v_b_23')
// (8, 22, 'sp12_v_b_20')
// (8, 23, 'sp12_v_b_19')
// (8, 24, 'sp12_v_b_16')
// (8, 25, 'neigh_op_top_6')
// (8, 25, 'sp12_v_b_15')
// (8, 26, 'ram/RDATA_1')
// (8, 26, 'sp12_v_b_12')
// (8, 27, 'neigh_op_bot_6')
// (8, 27, 'sp12_v_b_11')
// (8, 28, 'sp12_v_b_8')
// (8, 29, 'sp12_v_b_7')
// (8, 30, 'sp12_v_b_4')
// (8, 31, 'sp12_v_b_3')
// (8, 32, 'sp12_v_b_0')
// (9, 25, 'neigh_op_tnl_6')
// (9, 26, 'neigh_op_lft_6')
// (9, 27, 'neigh_op_bnl_6')

wire \data_out[0] ;
// (0, 3, 'io_0/D_OUT_0')
// (0, 3, 'io_0/PAD')
// (0, 3, 'local_g0_0')
// (0, 3, 'span4_horz_40')
// (1, 3, 'sp4_h_l_40')
// (1, 3, 'sp4_h_r_9')
// (2, 3, 'sp4_h_r_20')
// (3, 3, 'sp4_h_r_33')
// (4, 3, 'sp4_h_r_44')
// (4, 4, 'sp4_r_v_b_44')
// (4, 5, 'sp4_r_v_b_33')
// (4, 6, 'sp4_r_v_b_20')
// (4, 7, 'sp4_r_v_b_9')
// (5, 2, 'sp12_v_t_22')
// (5, 3, 'sp12_v_b_22')
// (5, 3, 'sp4_h_l_44')
// (5, 3, 'sp4_v_t_44')
// (5, 4, 'sp12_v_b_21')
// (5, 4, 'sp4_v_b_44')
// (5, 5, 'sp12_v_b_18')
// (5, 5, 'sp4_v_b_33')
// (5, 6, 'sp12_v_b_17')
// (5, 6, 'sp4_v_b_20')
// (5, 7, 'sp12_v_b_14')
// (5, 7, 'sp4_v_b_9')
// (5, 8, 'sp12_v_b_13')
// (5, 9, 'sp12_v_b_10')
// (5, 10, 'sp12_v_b_9')
// (5, 11, 'sp12_v_b_6')
// (5, 12, 'sp12_v_b_5')
// (5, 13, 'sp12_v_b_2')
// (5, 14, 'sp12_v_b_1')
// (5, 14, 'sp12_v_t_22')
// (5, 15, 'sp12_v_b_22')
// (5, 16, 'sp12_v_b_21')
// (5, 17, 'sp12_v_b_18')
// (5, 18, 'sp12_v_b_17')
// (5, 19, 'sp12_v_b_14')
// (5, 20, 'sp12_v_b_13')
// (5, 21, 'sp12_v_b_10')
// (5, 22, 'sp12_v_b_9')
// (5, 23, 'sp12_v_b_6')
// (5, 24, 'sp12_v_b_5')
// (5, 25, 'sp12_v_b_2')
// (5, 26, 'sp12_h_r_1')
// (5, 26, 'sp12_v_b_1')
// (6, 26, 'sp12_h_r_2')
// (7, 25, 'neigh_op_tnr_7')
// (7, 26, 'neigh_op_rgt_7')
// (7, 26, 'sp12_h_r_5')
// (7, 27, 'neigh_op_bnr_7')
// (8, 25, 'neigh_op_top_7')
// (8, 26, 'ram/RDATA_0')
// (8, 26, 'sp12_h_r_6')
// (8, 27, 'neigh_op_bot_7')
// (9, 25, 'neigh_op_tnl_7')
// (9, 26, 'neigh_op_lft_7')
// (9, 26, 'sp12_h_r_9')
// (9, 27, 'neigh_op_bnl_7')
// (10, 26, 'sp12_h_r_10')
// (11, 26, 'sp12_h_r_13')
// (12, 26, 'sp12_h_r_14')
// (13, 26, 'sp12_h_r_17')
// (14, 26, 'sp12_h_r_18')
// (15, 26, 'sp12_h_r_21')
// (16, 26, 'sp12_h_r_22')
// (17, 26, 'sp12_h_l_22')

wire \data_out[11] ;
// (0, 3, 'span4_horz_7')
// (0, 3, 'span4_vert_t_13')
// (0, 4, 'io_1/D_OUT_0')
// (0, 4, 'io_1/PAD')
// (0, 4, 'local_g0_5')
// (0, 4, 'span4_vert_b_13')
// (0, 5, 'span4_vert_b_9')
// (0, 6, 'span4_vert_b_5')
// (0, 7, 'span4_vert_b_1')
// (1, 3, 'sp4_h_r_18')
// (2, 3, 'sp4_h_r_31')
// (3, 3, 'sp4_h_r_42')
// (4, 3, 'sp4_h_l_42')
// (4, 3, 'sp4_h_r_4')
// (5, 3, 'sp4_h_r_17')
// (6, 3, 'sp4_h_r_28')
// (7, 3, 'sp4_h_r_41')
// (7, 4, 'sp4_r_v_b_47')
// (7, 5, 'sp4_r_v_b_34')
// (7, 6, 'sp4_r_v_b_23')
// (7, 7, 'sp4_r_v_b_10')
// (7, 24, 'neigh_op_tnr_4')
// (7, 25, 'neigh_op_rgt_4')
// (7, 26, 'neigh_op_bnr_4')
// (8, 3, 'sp4_h_l_41')
// (8, 3, 'sp4_v_t_47')
// (8, 4, 'sp4_v_b_47')
// (8, 5, 'sp12_v_t_23')
// (8, 5, 'sp4_v_b_34')
// (8, 6, 'sp12_v_b_23')
// (8, 6, 'sp4_v_b_23')
// (8, 7, 'sp12_v_b_20')
// (8, 7, 'sp4_v_b_10')
// (8, 8, 'sp12_v_b_19')
// (8, 9, 'sp12_v_b_16')
// (8, 10, 'sp12_v_b_15')
// (8, 11, 'sp12_v_b_12')
// (8, 12, 'sp12_v_b_11')
// (8, 13, 'sp12_v_b_8')
// (8, 14, 'sp12_v_b_7')
// (8, 15, 'sp12_v_b_4')
// (8, 16, 'sp12_v_b_3')
// (8, 17, 'sp12_v_b_0')
// (8, 17, 'sp12_v_t_23')
// (8, 18, 'sp12_v_b_23')
// (8, 19, 'sp12_v_b_20')
// (8, 20, 'sp12_v_b_19')
// (8, 21, 'sp12_v_b_16')
// (8, 22, 'sp12_v_b_15')
// (8, 23, 'sp12_v_b_12')
// (8, 24, 'neigh_op_top_4')
// (8, 24, 'sp12_v_b_11')
// (8, 25, 'ram/RDATA_11')
// (8, 25, 'sp12_v_b_8')
// (8, 26, 'neigh_op_bot_4')
// (8, 26, 'sp12_v_b_7')
// (8, 27, 'sp12_v_b_4')
// (8, 28, 'sp12_v_b_3')
// (8, 29, 'sp12_v_b_0')
// (9, 24, 'neigh_op_tnl_4')
// (9, 25, 'neigh_op_lft_4')
// (9, 26, 'neigh_op_bnl_4')

wire \data_out[15] ;
// (0, 3, 'span4_vert_t_12')
// (0, 4, 'span4_vert_b_12')
// (0, 5, 'span4_vert_b_8')
// (0, 6, 'io_1/D_OUT_0')
// (0, 6, 'io_1/PAD')
// (0, 6, 'local_g1_4')
// (0, 6, 'span4_vert_b_4')
// (0, 7, 'span4_horz_1')
// (0, 7, 'span4_vert_b_0')
// (1, 7, 'sp4_h_r_12')
// (2, 7, 'sp4_h_r_25')
// (3, 7, 'sp4_h_r_36')
// (3, 8, 'sp4_r_v_b_36')
// (3, 9, 'sp4_r_v_b_25')
// (3, 10, 'sp4_r_v_b_12')
// (3, 11, 'sp4_r_v_b_1')
// (3, 12, 'sp4_r_v_b_47')
// (3, 13, 'sp4_r_v_b_34')
// (3, 14, 'sp4_r_v_b_23')
// (3, 15, 'sp4_r_v_b_10')
// (4, 7, 'sp4_h_l_36')
// (4, 7, 'sp4_v_t_36')
// (4, 8, 'sp4_v_b_36')
// (4, 9, 'sp4_v_b_25')
// (4, 10, 'sp4_v_b_12')
// (4, 11, 'sp4_v_b_1')
// (4, 11, 'sp4_v_t_47')
// (4, 12, 'sp4_v_b_47')
// (4, 13, 'sp12_v_t_23')
// (4, 13, 'sp4_v_b_34')
// (4, 14, 'sp12_v_b_23')
// (4, 14, 'sp4_v_b_23')
// (4, 15, 'sp12_v_b_20')
// (4, 15, 'sp4_v_b_10')
// (4, 16, 'sp12_v_b_19')
// (4, 17, 'sp12_v_b_16')
// (4, 18, 'sp12_v_b_15')
// (4, 19, 'sp12_v_b_12')
// (4, 20, 'sp12_v_b_11')
// (4, 21, 'sp12_v_b_8')
// (4, 22, 'sp12_v_b_7')
// (4, 23, 'sp12_v_b_4')
// (4, 24, 'sp12_v_b_3')
// (4, 25, 'sp12_h_r_0')
// (4, 25, 'sp12_v_b_0')
// (5, 25, 'sp12_h_r_3')
// (6, 25, 'sp12_h_r_4')
// (7, 24, 'neigh_op_tnr_0')
// (7, 25, 'neigh_op_rgt_0')
// (7, 25, 'sp12_h_r_7')
// (7, 26, 'neigh_op_bnr_0')
// (8, 24, 'neigh_op_top_0')
// (8, 25, 'ram/RDATA_15')
// (8, 25, 'sp12_h_r_8')
// (8, 26, 'neigh_op_bot_0')
// (9, 24, 'neigh_op_tnl_0')
// (9, 25, 'neigh_op_lft_0')
// (9, 25, 'sp12_h_r_11')
// (9, 26, 'neigh_op_bnl_0')
// (10, 25, 'sp12_h_r_12')
// (11, 25, 'sp12_h_r_15')
// (12, 25, 'sp12_h_r_16')
// (13, 25, 'sp12_h_r_19')
// (14, 25, 'sp12_h_r_20')
// (15, 25, 'sp12_h_r_23')
// (16, 25, 'sp12_h_l_23')

wire \data_out[10] ;
// (0, 4, 'io_0/D_OUT_0')
// (0, 4, 'io_0/PAD')
// (0, 4, 'local_g0_2')
// (0, 4, 'span4_horz_18')
// (1, 4, 'sp4_h_r_31')
// (2, 4, 'sp4_h_r_42')
// (3, 4, 'sp4_h_l_42')
// (3, 4, 'sp4_h_r_11')
// (4, 4, 'sp4_h_r_22')
// (5, 4, 'sp4_h_r_35')
// (6, 1, 'sp4_r_v_b_46')
// (6, 2, 'sp4_r_v_b_35')
// (6, 3, 'sp4_r_v_b_22')
// (6, 4, 'sp4_h_r_46')
// (6, 4, 'sp4_r_v_b_11')
// (7, 0, 'span4_vert_46')
// (7, 1, 'sp12_v_t_22')
// (7, 1, 'sp4_v_b_46')
// (7, 2, 'sp12_v_b_22')
// (7, 2, 'sp4_v_b_35')
// (7, 3, 'sp12_v_b_21')
// (7, 3, 'sp4_v_b_22')
// (7, 4, 'sp12_v_b_18')
// (7, 4, 'sp4_h_l_46')
// (7, 4, 'sp4_v_b_11')
// (7, 5, 'sp12_v_b_17')
// (7, 6, 'sp12_v_b_14')
// (7, 7, 'sp12_v_b_13')
// (7, 8, 'sp12_v_b_10')
// (7, 9, 'sp12_v_b_9')
// (7, 10, 'sp12_v_b_6')
// (7, 11, 'sp12_v_b_5')
// (7, 12, 'sp12_v_b_2')
// (7, 13, 'sp12_v_b_1')
// (7, 13, 'sp12_v_t_22')
// (7, 14, 'sp12_v_b_22')
// (7, 15, 'sp12_v_b_21')
// (7, 16, 'sp12_v_b_18')
// (7, 17, 'sp12_v_b_17')
// (7, 18, 'sp12_v_b_14')
// (7, 19, 'sp12_v_b_13')
// (7, 20, 'sp12_v_b_10')
// (7, 21, 'sp12_v_b_9')
// (7, 22, 'sp12_v_b_6')
// (7, 23, 'sp12_v_b_5')
// (7, 24, 'neigh_op_tnr_5')
// (7, 24, 'sp12_v_b_2')
// (7, 25, 'neigh_op_rgt_5')
// (7, 25, 'sp12_h_r_1')
// (7, 25, 'sp12_v_b_1')
// (7, 26, 'neigh_op_bnr_5')
// (8, 24, 'neigh_op_top_5')
// (8, 25, 'ram/RDATA_10')
// (8, 25, 'sp12_h_r_2')
// (8, 26, 'neigh_op_bot_5')
// (9, 24, 'neigh_op_tnl_5')
// (9, 25, 'neigh_op_lft_5')
// (9, 25, 'sp12_h_r_5')
// (9, 26, 'neigh_op_bnl_5')
// (10, 25, 'sp12_h_r_6')
// (11, 25, 'sp12_h_r_9')
// (12, 25, 'sp12_h_r_10')
// (13, 25, 'sp12_h_r_13')
// (14, 25, 'sp12_h_r_14')
// (15, 25, 'sp12_h_r_17')
// (16, 25, 'sp12_h_r_18')
// (17, 25, 'sp12_h_r_21')
// (18, 25, 'sp12_h_r_22')
// (19, 25, 'sp12_h_l_22')

wire \data_out[17] ;
// (0, 4, 'span4_horz_7')
// (0, 4, 'span4_vert_t_13')
// (0, 5, 'span4_vert_b_13')
// (0, 6, 'span4_vert_b_9')
// (0, 7, 'io_1/D_OUT_0')
// (0, 7, 'io_1/PAD')
// (0, 7, 'local_g0_5')
// (0, 7, 'span4_vert_b_5')
// (0, 8, 'span4_vert_b_1')
// (1, 4, 'sp4_h_r_18')
// (2, 4, 'sp4_h_r_31')
// (3, 4, 'sp4_h_r_42')
// (4, 4, 'sp4_h_l_42')
// (4, 4, 'sp4_h_r_4')
// (5, 4, 'sp4_h_r_17')
// (6, 4, 'sp4_h_r_28')
// (7, 4, 'sp4_h_r_41')
// (7, 5, 'sp4_r_v_b_47')
// (7, 6, 'sp4_r_v_b_34')
// (7, 7, 'sp4_r_v_b_23')
// (7, 8, 'sp4_r_v_b_10')
// (7, 23, 'neigh_op_tnr_6')
// (7, 24, 'neigh_op_rgt_6')
// (7, 25, 'neigh_op_bnr_6')
// (8, 4, 'sp4_h_l_41')
// (8, 4, 'sp4_v_t_47')
// (8, 5, 'sp4_v_b_47')
// (8, 6, 'sp12_v_t_23')
// (8, 6, 'sp4_v_b_34')
// (8, 7, 'sp12_v_b_23')
// (8, 7, 'sp4_v_b_23')
// (8, 8, 'sp12_v_b_20')
// (8, 8, 'sp4_v_b_10')
// (8, 9, 'sp12_v_b_19')
// (8, 10, 'sp12_v_b_16')
// (8, 11, 'sp12_v_b_15')
// (8, 12, 'sp12_v_b_12')
// (8, 13, 'sp12_v_b_11')
// (8, 14, 'sp12_v_b_8')
// (8, 15, 'sp12_v_b_7')
// (8, 16, 'sp12_v_b_4')
// (8, 17, 'sp12_v_b_3')
// (8, 18, 'sp12_v_b_0')
// (8, 18, 'sp12_v_t_23')
// (8, 19, 'sp12_v_b_23')
// (8, 20, 'sp12_v_b_20')
// (8, 21, 'sp12_v_b_19')
// (8, 22, 'sp12_v_b_16')
// (8, 23, 'neigh_op_top_6')
// (8, 23, 'sp12_v_b_15')
// (8, 24, 'ram/RDATA_1')
// (8, 24, 'sp12_v_b_12')
// (8, 25, 'neigh_op_bot_6')
// (8, 25, 'sp12_v_b_11')
// (8, 26, 'sp12_v_b_8')
// (8, 27, 'sp12_v_b_7')
// (8, 28, 'sp12_v_b_4')
// (8, 29, 'sp12_v_b_3')
// (8, 30, 'sp12_v_b_0')
// (9, 23, 'neigh_op_tnl_6')
// (9, 24, 'neigh_op_lft_6')
// (9, 25, 'neigh_op_bnl_6')

wire \data_out[12] ;
// (0, 5, 'io_0/D_OUT_0')
// (0, 5, 'io_0/PAD')
// (0, 5, 'local_g0_0')
// (0, 5, 'span4_horz_0')
// (1, 5, 'sp4_h_r_13')
// (2, 5, 'sp4_h_r_24')
// (3, 5, 'sp4_h_r_37')
// (4, 5, 'sp4_h_l_37')
// (4, 5, 'sp4_h_r_9')
// (5, 5, 'sp4_h_r_20')
// (6, 5, 'sp4_h_r_33')
// (7, 5, 'sp4_h_r_44')
// (7, 6, 'sp4_r_v_b_44')
// (7, 7, 'sp4_r_v_b_33')
// (7, 8, 'sp4_r_v_b_20')
// (7, 9, 'sp4_r_v_b_9')
// (7, 24, 'neigh_op_tnr_3')
// (7, 25, 'neigh_op_rgt_3')
// (7, 26, 'neigh_op_bnr_3')
// (8, 4, 'sp12_v_t_22')
// (8, 5, 'sp12_v_b_22')
// (8, 5, 'sp4_h_l_44')
// (8, 5, 'sp4_v_t_44')
// (8, 6, 'sp12_v_b_21')
// (8, 6, 'sp4_v_b_44')
// (8, 7, 'sp12_v_b_18')
// (8, 7, 'sp4_v_b_33')
// (8, 8, 'sp12_v_b_17')
// (8, 8, 'sp4_v_b_20')
// (8, 9, 'sp12_v_b_14')
// (8, 9, 'sp4_v_b_9')
// (8, 10, 'sp12_v_b_13')
// (8, 11, 'sp12_v_b_10')
// (8, 12, 'sp12_v_b_9')
// (8, 13, 'sp12_v_b_6')
// (8, 14, 'sp12_v_b_5')
// (8, 15, 'sp12_v_b_2')
// (8, 16, 'sp12_v_b_1')
// (8, 16, 'sp12_v_t_22')
// (8, 17, 'sp12_v_b_22')
// (8, 18, 'sp12_v_b_21')
// (8, 19, 'sp12_v_b_18')
// (8, 20, 'sp12_v_b_17')
// (8, 21, 'sp12_v_b_14')
// (8, 22, 'sp12_v_b_13')
// (8, 23, 'sp12_v_b_10')
// (8, 24, 'neigh_op_top_3')
// (8, 24, 'sp12_v_b_9')
// (8, 25, 'ram/RDATA_12')
// (8, 25, 'sp12_v_b_6')
// (8, 26, 'neigh_op_bot_3')
// (8, 26, 'sp12_v_b_5')
// (8, 27, 'sp12_v_b_2')
// (8, 28, 'sp12_v_b_1')
// (9, 24, 'neigh_op_tnl_3')
// (9, 25, 'neigh_op_lft_3')
// (9, 26, 'neigh_op_bnl_3')

wire \data_out[13] ;
// (0, 5, 'io_1/D_OUT_0')
// (0, 5, 'io_1/PAD')
// (0, 5, 'local_g0_1')
// (0, 5, 'span4_horz_1')
// (1, 5, 'sp4_h_r_12')
// (2, 5, 'sp4_h_r_25')
// (3, 5, 'sp4_h_r_36')
// (4, 5, 'sp4_h_l_36')
// (4, 5, 'sp4_h_r_10')
// (5, 5, 'sp4_h_r_23')
// (6, 5, 'sp4_h_r_34')
// (7, 2, 'sp4_r_v_b_47')
// (7, 3, 'sp4_r_v_b_34')
// (7, 4, 'sp4_r_v_b_23')
// (7, 5, 'sp4_h_r_47')
// (7, 5, 'sp4_r_v_b_10')
// (7, 24, 'neigh_op_tnr_2')
// (7, 25, 'neigh_op_rgt_2')
// (7, 26, 'neigh_op_bnr_2')
// (8, 1, 'sp4_v_t_47')
// (8, 2, 'sp4_v_b_47')
// (8, 3, 'sp12_v_t_23')
// (8, 3, 'sp4_v_b_34')
// (8, 4, 'sp12_v_b_23')
// (8, 4, 'sp4_v_b_23')
// (8, 5, 'sp12_v_b_20')
// (8, 5, 'sp4_h_l_47')
// (8, 5, 'sp4_v_b_10')
// (8, 6, 'sp12_v_b_19')
// (8, 7, 'sp12_v_b_16')
// (8, 8, 'sp12_v_b_15')
// (8, 9, 'sp12_v_b_12')
// (8, 10, 'sp12_v_b_11')
// (8, 11, 'sp12_v_b_8')
// (8, 12, 'sp12_v_b_7')
// (8, 13, 'sp12_v_b_4')
// (8, 14, 'sp12_v_b_3')
// (8, 15, 'sp12_v_b_0')
// (8, 15, 'sp12_v_t_23')
// (8, 16, 'sp12_v_b_23')
// (8, 17, 'sp12_v_b_20')
// (8, 18, 'sp12_v_b_19')
// (8, 19, 'sp12_v_b_16')
// (8, 20, 'sp12_v_b_15')
// (8, 21, 'sp12_v_b_12')
// (8, 22, 'sp12_v_b_11')
// (8, 23, 'sp12_v_b_8')
// (8, 24, 'neigh_op_top_2')
// (8, 24, 'sp12_v_b_7')
// (8, 25, 'ram/RDATA_13')
// (8, 25, 'sp12_v_b_4')
// (8, 26, 'neigh_op_bot_2')
// (8, 26, 'sp12_v_b_3')
// (8, 27, 'sp12_v_b_0')
// (9, 24, 'neigh_op_tnl_2')
// (9, 25, 'neigh_op_lft_2')
// (9, 26, 'neigh_op_bnl_2')

wire \data_out[14] ;
// (0, 6, 'io_0/D_OUT_0')
// (0, 6, 'io_0/PAD')
// (0, 6, 'local_g0_0')
// (0, 6, 'span4_horz_16')
// (1, 6, 'sp4_h_r_29')
// (2, 6, 'sp4_h_r_40')
// (2, 7, 'sp4_r_v_b_40')
// (2, 8, 'sp4_r_v_b_29')
// (2, 9, 'sp4_r_v_b_16')
// (2, 10, 'sp4_r_v_b_5')
// (3, 1, 'sp12_v_t_22')
// (3, 2, 'sp12_v_b_22')
// (3, 3, 'sp12_v_b_21')
// (3, 4, 'sp12_v_b_18')
// (3, 5, 'sp12_v_b_17')
// (3, 6, 'sp12_v_b_14')
// (3, 6, 'sp4_h_l_40')
// (3, 6, 'sp4_v_t_40')
// (3, 7, 'sp12_v_b_13')
// (3, 7, 'sp4_v_b_40')
// (3, 8, 'sp12_v_b_10')
// (3, 8, 'sp4_v_b_29')
// (3, 9, 'sp12_v_b_9')
// (3, 9, 'sp4_v_b_16')
// (3, 10, 'sp12_v_b_6')
// (3, 10, 'sp4_v_b_5')
// (3, 11, 'sp12_v_b_5')
// (3, 12, 'sp12_v_b_2')
// (3, 13, 'sp12_v_b_1')
// (3, 13, 'sp12_v_t_22')
// (3, 14, 'sp12_v_b_22')
// (3, 15, 'sp12_v_b_21')
// (3, 16, 'sp12_v_b_18')
// (3, 17, 'sp12_v_b_17')
// (3, 18, 'sp12_v_b_14')
// (3, 19, 'sp12_v_b_13')
// (3, 20, 'sp12_v_b_10')
// (3, 21, 'sp12_v_b_9')
// (3, 22, 'sp12_v_b_6')
// (3, 23, 'sp12_v_b_5')
// (3, 24, 'sp12_v_b_2')
// (3, 25, 'sp12_h_r_1')
// (3, 25, 'sp12_v_b_1')
// (4, 25, 'sp12_h_r_2')
// (5, 25, 'sp12_h_r_5')
// (6, 25, 'sp12_h_r_6')
// (7, 24, 'neigh_op_tnr_1')
// (7, 25, 'neigh_op_rgt_1')
// (7, 25, 'sp12_h_r_9')
// (7, 26, 'neigh_op_bnr_1')
// (8, 24, 'neigh_op_top_1')
// (8, 25, 'ram/RDATA_14')
// (8, 25, 'sp12_h_r_10')
// (8, 26, 'neigh_op_bot_1')
// (9, 24, 'neigh_op_tnl_1')
// (9, 25, 'neigh_op_lft_1')
// (9, 25, 'sp12_h_r_13')
// (9, 26, 'neigh_op_bnl_1')
// (10, 25, 'sp12_h_r_14')
// (11, 25, 'sp12_h_r_17')
// (12, 25, 'sp12_h_r_18')
// (13, 25, 'sp12_h_r_21')
// (14, 25, 'sp12_h_r_22')
// (15, 25, 'sp12_h_l_22')

wire \data_out[16] ;
// (0, 7, 'io_0/D_OUT_0')
// (0, 7, 'io_0/PAD')
// (0, 7, 'local_g1_1')
// (0, 7, 'span12_horz_9')
// (1, 7, 'sp12_h_r_10')
// (2, 7, 'sp12_h_r_13')
// (3, 7, 'sp12_h_r_14')
// (4, 7, 'sp12_h_r_17')
// (5, 7, 'sp12_h_r_18')
// (6, 7, 'sp12_h_r_21')
// (7, 7, 'sp12_h_r_22')
// (7, 23, 'neigh_op_tnr_7')
// (7, 24, 'neigh_op_rgt_7')
// (7, 25, 'neigh_op_bnr_7')
// (8, 7, 'sp12_h_l_22')
// (8, 7, 'sp12_v_t_22')
// (8, 8, 'sp12_v_b_22')
// (8, 9, 'sp12_v_b_21')
// (8, 10, 'sp12_v_b_18')
// (8, 11, 'sp12_v_b_17')
// (8, 12, 'sp12_v_b_14')
// (8, 13, 'sp12_v_b_13')
// (8, 14, 'sp12_v_b_10')
// (8, 15, 'sp12_v_b_9')
// (8, 16, 'sp12_v_b_6')
// (8, 17, 'sp12_v_b_5')
// (8, 18, 'sp12_v_b_2')
// (8, 19, 'sp12_v_b_1')
// (8, 19, 'sp12_v_t_22')
// (8, 20, 'sp12_v_b_22')
// (8, 21, 'sp12_v_b_21')
// (8, 22, 'sp12_v_b_18')
// (8, 23, 'neigh_op_top_7')
// (8, 23, 'sp12_v_b_17')
// (8, 24, 'ram/RDATA_0')
// (8, 24, 'sp12_v_b_14')
// (8, 25, 'neigh_op_bot_7')
// (8, 25, 'sp12_v_b_13')
// (8, 26, 'sp12_v_b_10')
// (8, 27, 'sp12_v_b_9')
// (8, 28, 'sp12_v_b_6')
// (8, 29, 'sp12_v_b_5')
// (8, 30, 'sp12_v_b_2')
// (8, 31, 'sp12_v_b_1')
// (9, 23, 'neigh_op_tnl_7')
// (9, 24, 'neigh_op_lft_7')
// (9, 25, 'neigh_op_bnl_7')

wire \data_out[18] ;
// (0, 8, 'io_0/D_OUT_0')
// (0, 8, 'io_0/PAD')
// (0, 8, 'local_g0_0')
// (0, 8, 'span4_horz_0')
// (1, 8, 'sp4_h_r_13')
// (2, 8, 'sp4_h_r_24')
// (3, 8, 'sp4_h_r_37')
// (4, 8, 'sp4_h_l_37')
// (4, 8, 'sp4_h_r_4')
// (5, 8, 'sp4_h_r_17')
// (6, 8, 'sp4_h_r_28')
// (7, 5, 'sp4_r_v_b_46')
// (7, 6, 'sp4_r_v_b_35')
// (7, 7, 'sp4_r_v_b_22')
// (7, 8, 'sp4_h_r_41')
// (7, 8, 'sp4_r_v_b_11')
// (7, 23, 'neigh_op_tnr_5')
// (7, 24, 'neigh_op_rgt_5')
// (7, 25, 'neigh_op_bnr_5')
// (8, 4, 'sp4_v_t_46')
// (8, 5, 'sp12_v_t_22')
// (8, 5, 'sp4_v_b_46')
// (8, 6, 'sp12_v_b_22')
// (8, 6, 'sp4_v_b_35')
// (8, 7, 'sp12_v_b_21')
// (8, 7, 'sp4_v_b_22')
// (8, 8, 'sp12_v_b_18')
// (8, 8, 'sp4_h_l_41')
// (8, 8, 'sp4_v_b_11')
// (8, 9, 'sp12_v_b_17')
// (8, 10, 'sp12_v_b_14')
// (8, 11, 'sp12_v_b_13')
// (8, 12, 'sp12_v_b_10')
// (8, 13, 'sp12_v_b_9')
// (8, 14, 'sp12_v_b_6')
// (8, 15, 'sp12_v_b_5')
// (8, 16, 'sp12_v_b_2')
// (8, 17, 'sp12_v_b_1')
// (8, 17, 'sp12_v_t_22')
// (8, 18, 'sp12_v_b_22')
// (8, 19, 'sp12_v_b_21')
// (8, 20, 'sp12_v_b_18')
// (8, 21, 'sp12_v_b_17')
// (8, 22, 'sp12_v_b_14')
// (8, 23, 'neigh_op_top_5')
// (8, 23, 'sp12_v_b_13')
// (8, 24, 'ram/RDATA_2')
// (8, 24, 'sp12_v_b_10')
// (8, 25, 'neigh_op_bot_5')
// (8, 25, 'sp12_v_b_9')
// (8, 26, 'sp12_v_b_6')
// (8, 27, 'sp12_v_b_5')
// (8, 28, 'sp12_v_b_2')
// (8, 29, 'sp12_v_b_1')
// (9, 23, 'neigh_op_tnl_5')
// (9, 24, 'neigh_op_lft_5')
// (9, 25, 'neigh_op_bnl_5')

wire \data_out[19] ;
// (0, 8, 'io_1/D_OUT_0')
// (0, 8, 'io_1/PAD')
// (0, 8, 'local_g0_1')
// (0, 8, 'span4_horz_1')
// (1, 8, 'sp4_h_r_12')
// (2, 8, 'sp4_h_r_25')
// (3, 8, 'sp4_h_r_36')
// (4, 8, 'sp4_h_l_36')
// (4, 8, 'sp4_h_r_1')
// (5, 8, 'sp4_h_r_12')
// (6, 8, 'sp4_h_r_25')
// (7, 5, 'sp4_r_v_b_45')
// (7, 6, 'sp4_r_v_b_32')
// (7, 7, 'sp4_r_v_b_21')
// (7, 8, 'sp4_h_r_36')
// (7, 8, 'sp4_r_v_b_8')
// (7, 23, 'neigh_op_tnr_4')
// (7, 24, 'neigh_op_rgt_4')
// (7, 25, 'neigh_op_bnr_4')
// (8, 4, 'sp12_v_t_23')
// (8, 4, 'sp4_v_t_45')
// (8, 5, 'sp12_v_b_23')
// (8, 5, 'sp4_v_b_45')
// (8, 6, 'sp12_v_b_20')
// (8, 6, 'sp4_v_b_32')
// (8, 7, 'sp12_v_b_19')
// (8, 7, 'sp4_v_b_21')
// (8, 8, 'sp12_v_b_16')
// (8, 8, 'sp4_h_l_36')
// (8, 8, 'sp4_v_b_8')
// (8, 9, 'sp12_v_b_15')
// (8, 10, 'sp12_v_b_12')
// (8, 11, 'sp12_v_b_11')
// (8, 12, 'sp12_v_b_8')
// (8, 13, 'sp12_v_b_7')
// (8, 14, 'sp12_v_b_4')
// (8, 15, 'sp12_v_b_3')
// (8, 16, 'sp12_v_b_0')
// (8, 16, 'sp12_v_t_23')
// (8, 17, 'sp12_v_b_23')
// (8, 18, 'sp12_v_b_20')
// (8, 19, 'sp12_v_b_19')
// (8, 20, 'sp12_v_b_16')
// (8, 21, 'sp12_v_b_15')
// (8, 22, 'sp12_v_b_12')
// (8, 23, 'neigh_op_top_4')
// (8, 23, 'sp12_v_b_11')
// (8, 24, 'ram/RDATA_3')
// (8, 24, 'sp12_v_b_8')
// (8, 25, 'neigh_op_bot_4')
// (8, 25, 'sp12_v_b_7')
// (8, 26, 'sp12_v_b_4')
// (8, 27, 'sp12_v_b_3')
// (8, 28, 'sp12_v_b_0')
// (9, 23, 'neigh_op_tnl_4')
// (9, 24, 'neigh_op_lft_4')
// (9, 25, 'neigh_op_bnl_4')

wire \data_out[22] ;
// (0, 8, 'span4_vert_t_13')
// (0, 9, 'span4_vert_b_13')
// (0, 10, 'io_1/D_OUT_0')
// (0, 10, 'io_1/PAD')
// (0, 10, 'local_g0_1')
// (0, 10, 'span4_vert_b_9')
// (0, 11, 'span4_vert_b_5')
// (0, 12, 'span4_horz_7')
// (0, 12, 'span4_vert_b_1')
// (1, 12, 'sp4_h_r_18')
// (2, 12, 'sp4_h_r_31')
// (3, 12, 'sp4_h_r_42')
// (4, 12, 'sp4_h_l_42')
// (4, 12, 'sp4_h_r_11')
// (5, 12, 'sp4_h_r_22')
// (6, 12, 'sp4_h_r_35')
// (7, 12, 'sp4_h_r_46')
// (7, 13, 'sp4_r_v_b_46')
// (7, 14, 'sp4_r_v_b_35')
// (7, 15, 'sp4_r_v_b_22')
// (7, 16, 'sp4_r_v_b_11')
// (7, 23, 'neigh_op_tnr_1')
// (7, 24, 'neigh_op_rgt_1')
// (7, 25, 'neigh_op_bnr_1')
// (8, 12, 'sp4_h_l_46')
// (8, 12, 'sp4_v_t_46')
// (8, 13, 'sp12_v_t_22')
// (8, 13, 'sp4_v_b_46')
// (8, 14, 'sp12_v_b_22')
// (8, 14, 'sp4_v_b_35')
// (8, 15, 'sp12_v_b_21')
// (8, 15, 'sp4_v_b_22')
// (8, 16, 'sp12_v_b_18')
// (8, 16, 'sp4_v_b_11')
// (8, 17, 'sp12_v_b_17')
// (8, 18, 'sp12_v_b_14')
// (8, 19, 'sp12_v_b_13')
// (8, 20, 'sp12_v_b_10')
// (8, 21, 'sp12_v_b_9')
// (8, 22, 'sp12_v_b_6')
// (8, 23, 'neigh_op_top_1')
// (8, 23, 'sp12_v_b_5')
// (8, 24, 'ram/RDATA_6')
// (8, 24, 'sp12_v_b_2')
// (8, 25, 'neigh_op_bot_1')
// (8, 25, 'sp12_v_b_1')
// (9, 23, 'neigh_op_tnl_1')
// (9, 24, 'neigh_op_lft_1')
// (9, 25, 'neigh_op_bnl_1')

wire \data_out[2] ;
// (0, 9, 'io_0/D_OUT_0')
// (0, 9, 'io_0/PAD')
// (0, 9, 'local_g0_0')
// (0, 9, 'span4_horz_16')
// (1, 9, 'sp4_h_r_29')
// (2, 9, 'sp4_h_r_40')
// (2, 10, 'sp4_r_v_b_40')
// (2, 11, 'sp4_r_v_b_29')
// (2, 12, 'sp4_r_v_b_16')
// (2, 13, 'sp4_r_v_b_5')
// (3, 9, 'sp4_h_l_40')
// (3, 9, 'sp4_v_t_40')
// (3, 10, 'sp4_v_b_40')
// (3, 11, 'sp4_v_b_29')
// (3, 12, 'sp4_v_b_16')
// (3, 13, 'sp4_h_r_5')
// (3, 13, 'sp4_v_b_5')
// (4, 13, 'sp4_h_r_16')
// (5, 13, 'sp4_h_r_29')
// (6, 13, 'sp4_h_r_40')
// (6, 14, 'sp4_r_v_b_46')
// (6, 15, 'sp4_r_v_b_35')
// (6, 16, 'sp4_r_v_b_22')
// (6, 17, 'sp4_r_v_b_11')
// (7, 13, 'sp4_h_l_40')
// (7, 13, 'sp4_v_t_46')
// (7, 14, 'sp12_v_t_22')
// (7, 14, 'sp4_v_b_46')
// (7, 15, 'sp12_v_b_22')
// (7, 15, 'sp4_v_b_35')
// (7, 16, 'sp12_v_b_21')
// (7, 16, 'sp4_v_b_22')
// (7, 17, 'sp12_v_b_18')
// (7, 17, 'sp4_v_b_11')
// (7, 18, 'sp12_v_b_17')
// (7, 19, 'sp12_v_b_14')
// (7, 20, 'sp12_v_b_13')
// (7, 21, 'sp12_v_b_10')
// (7, 22, 'sp12_v_b_9')
// (7, 23, 'sp12_v_b_6')
// (7, 24, 'sp12_v_b_5')
// (7, 25, 'neigh_op_tnr_5')
// (7, 25, 'sp12_v_b_2')
// (7, 26, 'neigh_op_rgt_5')
// (7, 26, 'sp12_h_r_1')
// (7, 26, 'sp12_v_b_1')
// (7, 27, 'neigh_op_bnr_5')
// (8, 25, 'neigh_op_top_5')
// (8, 26, 'ram/RDATA_2')
// (8, 26, 'sp12_h_r_2')
// (8, 27, 'neigh_op_bot_5')
// (9, 25, 'neigh_op_tnl_5')
// (9, 26, 'neigh_op_lft_5')
// (9, 26, 'sp12_h_r_5')
// (9, 27, 'neigh_op_bnl_5')
// (10, 26, 'sp12_h_r_6')
// (11, 26, 'sp12_h_r_9')
// (12, 26, 'sp12_h_r_10')
// (13, 26, 'sp12_h_r_13')
// (14, 26, 'sp12_h_r_14')
// (15, 26, 'sp12_h_r_17')
// (16, 26, 'sp12_h_r_18')
// (17, 26, 'sp12_h_r_21')
// (18, 26, 'sp12_h_r_22')
// (19, 26, 'sp12_h_l_22')

wire \data_out[20] ;
// (0, 9, 'io_1/D_OUT_0')
// (0, 9, 'io_1/PAD')
// (0, 9, 'local_g0_3')
// (0, 9, 'span4_horz_43')
// (1, 9, 'sp4_h_l_43')
// (1, 9, 'sp4_v_t_37')
// (1, 10, 'sp4_v_b_37')
// (1, 11, 'sp4_v_b_24')
// (1, 12, 'sp12_v_t_22')
// (1, 12, 'sp4_v_b_13')
// (1, 13, 'sp12_v_b_22')
// (1, 13, 'sp4_v_b_0')
// (1, 13, 'sp4_v_t_44')
// (1, 14, 'sp12_v_b_21')
// (1, 14, 'sp4_v_b_44')
// (1, 15, 'sp12_v_b_18')
// (1, 15, 'sp4_v_b_33')
// (1, 16, 'sp12_v_b_17')
// (1, 16, 'sp4_v_b_20')
// (1, 17, 'sp12_v_b_14')
// (1, 17, 'sp4_v_b_9')
// (1, 18, 'sp12_v_b_13')
// (1, 19, 'sp12_v_b_10')
// (1, 20, 'sp12_v_b_9')
// (1, 21, 'sp12_v_b_6')
// (1, 22, 'sp12_v_b_5')
// (1, 23, 'sp12_v_b_2')
// (1, 24, 'sp12_h_r_1')
// (1, 24, 'sp12_v_b_1')
// (2, 24, 'sp12_h_r_2')
// (3, 24, 'sp12_h_r_5')
// (4, 24, 'sp12_h_r_6')
// (5, 24, 'sp12_h_r_9')
// (6, 24, 'sp12_h_r_10')
// (7, 23, 'neigh_op_tnr_3')
// (7, 24, 'neigh_op_rgt_3')
// (7, 24, 'sp12_h_r_13')
// (7, 25, 'neigh_op_bnr_3')
// (8, 23, 'neigh_op_top_3')
// (8, 24, 'ram/RDATA_4')
// (8, 24, 'sp12_h_r_14')
// (8, 25, 'neigh_op_bot_3')
// (9, 23, 'neigh_op_tnl_3')
// (9, 24, 'neigh_op_lft_3')
// (9, 24, 'sp12_h_r_17')
// (9, 25, 'neigh_op_bnl_3')
// (10, 24, 'sp12_h_r_18')
// (11, 24, 'sp12_h_r_21')
// (12, 24, 'sp12_h_r_22')
// (13, 24, 'sp12_h_l_22')

wire \data_out[21] ;
// (0, 10, 'io_0/D_OUT_0')
// (0, 10, 'io_0/PAD')
// (0, 10, 'local_g0_0')
// (0, 10, 'span12_horz_8')
// (1, 10, 'sp12_h_r_11')
// (2, 10, 'sp12_h_r_12')
// (3, 10, 'sp12_h_r_15')
// (4, 10, 'sp12_h_r_16')
// (5, 10, 'sp12_h_r_19')
// (6, 10, 'sp12_h_r_20')
// (7, 10, 'sp12_h_r_23')
// (7, 23, 'neigh_op_tnr_2')
// (7, 24, 'neigh_op_rgt_2')
// (7, 25, 'neigh_op_bnr_2')
// (8, 10, 'sp12_h_l_23')
// (8, 10, 'sp12_v_t_23')
// (8, 11, 'sp12_v_b_23')
// (8, 12, 'sp12_v_b_20')
// (8, 13, 'sp12_v_b_19')
// (8, 14, 'sp12_v_b_16')
// (8, 15, 'sp12_v_b_15')
// (8, 16, 'sp12_v_b_12')
// (8, 17, 'sp12_v_b_11')
// (8, 18, 'sp12_v_b_8')
// (8, 19, 'sp12_v_b_7')
// (8, 20, 'sp12_v_b_4')
// (8, 21, 'sp12_v_b_3')
// (8, 22, 'sp12_v_b_0')
// (8, 22, 'sp12_v_t_23')
// (8, 23, 'neigh_op_top_2')
// (8, 23, 'sp12_v_b_23')
// (8, 24, 'ram/RDATA_5')
// (8, 24, 'sp12_v_b_20')
// (8, 25, 'neigh_op_bot_2')
// (8, 25, 'sp12_v_b_19')
// (8, 26, 'sp12_v_b_16')
// (8, 27, 'sp12_v_b_15')
// (8, 28, 'sp12_v_b_12')
// (8, 29, 'sp12_v_b_11')
// (8, 30, 'sp12_v_b_8')
// (8, 31, 'sp12_v_b_7')
// (8, 32, 'sp12_v_b_4')
// (8, 33, 'span12_vert_3')
// (9, 23, 'neigh_op_tnl_2')
// (9, 24, 'neigh_op_lft_2')
// (9, 25, 'neigh_op_bnl_2')

wire \data_out[23] ;
// (0, 10, 'span4_horz_1')
// (0, 10, 'span4_vert_t_12')
// (0, 11, 'io_0/D_OUT_0')
// (0, 11, 'io_0/PAD')
// (0, 11, 'local_g0_4')
// (0, 11, 'span4_vert_b_12')
// (0, 12, 'span4_vert_b_8')
// (0, 13, 'span4_vert_b_4')
// (0, 14, 'span4_vert_b_0')
// (1, 10, 'sp4_h_r_12')
// (2, 10, 'sp4_h_r_25')
// (3, 10, 'sp4_h_r_36')
// (4, 10, 'sp4_h_l_36')
// (4, 10, 'sp4_h_r_10')
// (5, 10, 'sp4_h_r_23')
// (6, 10, 'sp4_h_r_34')
// (7, 10, 'sp4_h_r_47')
// (7, 11, 'sp4_r_v_b_47')
// (7, 12, 'sp4_r_v_b_34')
// (7, 13, 'sp4_r_v_b_23')
// (7, 14, 'sp4_r_v_b_10')
// (7, 23, 'neigh_op_tnr_0')
// (7, 24, 'neigh_op_rgt_0')
// (7, 25, 'neigh_op_bnr_0')
// (8, 10, 'sp4_h_l_47')
// (8, 10, 'sp4_v_t_47')
// (8, 11, 'sp4_v_b_47')
// (8, 12, 'sp12_v_t_23')
// (8, 12, 'sp4_v_b_34')
// (8, 13, 'sp12_v_b_23')
// (8, 13, 'sp4_v_b_23')
// (8, 14, 'sp12_v_b_20')
// (8, 14, 'sp4_v_b_10')
// (8, 15, 'sp12_v_b_19')
// (8, 16, 'sp12_v_b_16')
// (8, 17, 'sp12_v_b_15')
// (8, 18, 'sp12_v_b_12')
// (8, 19, 'sp12_v_b_11')
// (8, 20, 'sp12_v_b_8')
// (8, 21, 'sp12_v_b_7')
// (8, 22, 'sp12_v_b_4')
// (8, 23, 'neigh_op_top_0')
// (8, 23, 'sp12_v_b_3')
// (8, 24, 'ram/RDATA_7')
// (8, 24, 'sp12_v_b_0')
// (8, 25, 'neigh_op_bot_0')
// (9, 23, 'neigh_op_tnl_0')
// (9, 24, 'neigh_op_lft_0')
// (9, 25, 'neigh_op_bnl_0')

wire \data_out[24] ;
// (0, 11, 'io_1/D_OUT_0')
// (0, 11, 'io_1/PAD')
// (0, 11, 'local_g1_6')
// (0, 11, 'span12_horz_14')
// (1, 11, 'sp12_h_r_17')
// (2, 11, 'sp12_h_r_18')
// (3, 11, 'sp12_h_r_21')
// (4, 11, 'sp12_h_r_22')
// (5, 11, 'sp12_h_l_22')
// (5, 11, 'sp12_v_t_22')
// (5, 12, 'sp12_v_b_22')
// (5, 13, 'sp12_v_b_21')
// (5, 14, 'sp12_v_b_18')
// (5, 15, 'sp12_v_b_17')
// (5, 16, 'sp12_v_b_14')
// (5, 17, 'sp12_v_b_13')
// (5, 18, 'sp12_v_b_10')
// (5, 19, 'sp12_v_b_9')
// (5, 20, 'sp12_v_b_6')
// (5, 21, 'sp12_v_b_5')
// (5, 22, 'sp12_v_b_2')
// (5, 23, 'sp12_h_r_1')
// (5, 23, 'sp12_v_b_1')
// (6, 23, 'sp12_h_r_2')
// (7, 22, 'neigh_op_tnr_7')
// (7, 23, 'neigh_op_rgt_7')
// (7, 23, 'sp12_h_r_5')
// (7, 24, 'neigh_op_bnr_7')
// (8, 22, 'neigh_op_top_7')
// (8, 23, 'ram/RDATA_8')
// (8, 23, 'sp12_h_r_6')
// (8, 24, 'neigh_op_bot_7')
// (9, 22, 'neigh_op_tnl_7')
// (9, 23, 'neigh_op_lft_7')
// (9, 23, 'sp12_h_r_9')
// (9, 24, 'neigh_op_bnl_7')
// (10, 23, 'sp12_h_r_10')
// (11, 23, 'sp12_h_r_13')
// (12, 23, 'sp12_h_r_14')
// (13, 23, 'sp12_h_r_17')
// (14, 23, 'sp12_h_r_18')
// (15, 23, 'sp12_h_r_21')
// (16, 23, 'sp12_h_r_22')
// (17, 23, 'sp12_h_l_22')

wire \data_out[27] ;
// (0, 11, 'span4_vert_t_12')
// (0, 12, 'span4_vert_b_12')
// (0, 13, 'io_0/D_OUT_0')
// (0, 13, 'io_0/PAD')
// (0, 13, 'local_g0_0')
// (0, 13, 'span4_vert_b_8')
// (0, 14, 'span4_vert_b_4')
// (0, 15, 'span4_horz_1')
// (0, 15, 'span4_vert_b_0')
// (1, 15, 'sp4_h_r_12')
// (2, 15, 'sp4_h_r_25')
// (3, 15, 'sp4_h_r_36')
// (3, 16, 'sp4_r_v_b_36')
// (3, 17, 'sp4_r_v_b_25')
// (3, 18, 'sp4_r_v_b_12')
// (3, 19, 'sp4_r_v_b_1')
// (4, 15, 'sp4_h_l_36')
// (4, 15, 'sp4_v_t_36')
// (4, 16, 'sp4_v_b_36')
// (4, 17, 'sp4_v_b_25')
// (4, 18, 'sp4_v_b_12')
// (4, 19, 'sp4_h_r_8')
// (4, 19, 'sp4_v_b_1')
// (5, 19, 'sp4_h_r_21')
// (6, 19, 'sp4_h_r_32')
// (7, 19, 'sp4_h_r_45')
// (7, 20, 'sp4_r_v_b_45')
// (7, 21, 'sp4_r_v_b_32')
// (7, 22, 'neigh_op_tnr_4')
// (7, 22, 'sp4_r_v_b_21')
// (7, 23, 'neigh_op_rgt_4')
// (7, 23, 'sp4_r_v_b_8')
// (7, 24, 'neigh_op_bnr_4')
// (8, 19, 'sp4_h_l_45')
// (8, 19, 'sp4_v_t_45')
// (8, 20, 'sp4_v_b_45')
// (8, 21, 'sp4_v_b_32')
// (8, 22, 'neigh_op_top_4')
// (8, 22, 'sp4_v_b_21')
// (8, 23, 'ram/RDATA_11')
// (8, 23, 'sp4_v_b_8')
// (8, 24, 'neigh_op_bot_4')
// (9, 22, 'neigh_op_tnl_4')
// (9, 23, 'neigh_op_lft_4')
// (9, 24, 'neigh_op_bnl_4')

wire \data_out[25] ;
// (0, 12, 'io_0/D_OUT_0')
// (0, 12, 'io_0/PAD')
// (0, 12, 'local_g0_0')
// (0, 12, 'span4_horz_0')
// (1, 12, 'sp4_h_r_13')
// (2, 12, 'sp4_h_r_24')
// (3, 12, 'sp4_h_r_37')
// (3, 13, 'sp4_r_v_b_37')
// (3, 14, 'sp4_r_v_b_24')
// (3, 15, 'sp4_r_v_b_13')
// (3, 16, 'sp4_r_v_b_0')
// (3, 17, 'sp4_r_v_b_37')
// (3, 18, 'sp4_r_v_b_24')
// (3, 19, 'sp4_r_v_b_13')
// (3, 20, 'sp4_r_v_b_0')
// (4, 12, 'sp4_h_l_37')
// (4, 12, 'sp4_v_t_37')
// (4, 13, 'sp4_v_b_37')
// (4, 14, 'sp4_v_b_24')
// (4, 15, 'sp4_v_b_13')
// (4, 16, 'sp4_v_b_0')
// (4, 16, 'sp4_v_t_37')
// (4, 17, 'sp4_v_b_37')
// (4, 18, 'sp4_v_b_24')
// (4, 19, 'sp4_v_b_13')
// (4, 20, 'sp4_h_r_7')
// (4, 20, 'sp4_v_b_0')
// (5, 20, 'sp4_h_r_18')
// (6, 20, 'sp4_h_r_31')
// (7, 20, 'sp4_h_r_42')
// (7, 21, 'sp4_r_v_b_36')
// (7, 22, 'neigh_op_tnr_6')
// (7, 22, 'sp4_r_v_b_25')
// (7, 23, 'neigh_op_rgt_6')
// (7, 23, 'sp4_r_v_b_12')
// (7, 24, 'neigh_op_bnr_6')
// (7, 24, 'sp4_r_v_b_1')
// (8, 20, 'sp4_h_l_42')
// (8, 20, 'sp4_v_t_36')
// (8, 21, 'sp4_v_b_36')
// (8, 22, 'neigh_op_top_6')
// (8, 22, 'sp4_v_b_25')
// (8, 23, 'ram/RDATA_9')
// (8, 23, 'sp4_v_b_12')
// (8, 24, 'neigh_op_bot_6')
// (8, 24, 'sp4_v_b_1')
// (9, 22, 'neigh_op_tnl_6')
// (9, 23, 'neigh_op_lft_6')
// (9, 24, 'neigh_op_bnl_6')

wire \data_out[26] ;
// (0, 12, 'io_1/D_OUT_0')
// (0, 12, 'io_1/PAD')
// (0, 12, 'local_g0_3')
// (0, 12, 'span4_horz_19')
// (1, 12, 'sp4_h_r_30')
// (2, 12, 'sp4_h_r_43')
// (3, 12, 'sp4_h_l_43')
// (3, 12, 'sp4_h_r_3')
// (4, 12, 'sp4_h_r_14')
// (5, 12, 'sp4_h_r_27')
// (6, 12, 'sp4_h_r_38')
// (6, 13, 'sp4_r_v_b_44')
// (6, 14, 'sp4_r_v_b_33')
// (6, 15, 'sp4_r_v_b_20')
// (6, 16, 'sp4_r_v_b_9')
// (7, 11, 'sp12_v_t_22')
// (7, 12, 'sp12_v_b_22')
// (7, 12, 'sp4_h_l_38')
// (7, 12, 'sp4_v_t_44')
// (7, 13, 'sp12_v_b_21')
// (7, 13, 'sp4_v_b_44')
// (7, 14, 'sp12_v_b_18')
// (7, 14, 'sp4_v_b_33')
// (7, 15, 'sp12_v_b_17')
// (7, 15, 'sp4_v_b_20')
// (7, 16, 'sp12_v_b_14')
// (7, 16, 'sp4_v_b_9')
// (7, 17, 'sp12_v_b_13')
// (7, 18, 'sp12_v_b_10')
// (7, 19, 'sp12_v_b_9')
// (7, 20, 'sp12_v_b_6')
// (7, 21, 'sp12_v_b_5')
// (7, 22, 'neigh_op_tnr_5')
// (7, 22, 'sp12_v_b_2')
// (7, 23, 'neigh_op_rgt_5')
// (7, 23, 'sp12_h_r_1')
// (7, 23, 'sp12_v_b_1')
// (7, 24, 'neigh_op_bnr_5')
// (8, 22, 'neigh_op_top_5')
// (8, 23, 'ram/RDATA_10')
// (8, 23, 'sp12_h_r_2')
// (8, 24, 'neigh_op_bot_5')
// (9, 22, 'neigh_op_tnl_5')
// (9, 23, 'neigh_op_lft_5')
// (9, 23, 'sp12_h_r_5')
// (9, 24, 'neigh_op_bnl_5')
// (10, 23, 'sp12_h_r_6')
// (11, 23, 'sp12_h_r_9')
// (12, 23, 'sp12_h_r_10')
// (13, 23, 'sp12_h_r_13')
// (14, 23, 'sp12_h_r_14')
// (15, 23, 'sp12_h_r_17')
// (16, 23, 'sp12_h_r_18')
// (17, 23, 'sp12_h_r_21')
// (18, 23, 'sp12_h_r_22')
// (19, 23, 'sp12_h_l_22')

wire \data_out[29] ;
// (0, 12, 'span4_vert_t_12')
// (0, 13, 'span4_vert_b_12')
// (0, 14, 'io_0/D_OUT_0')
// (0, 14, 'io_0/PAD')
// (0, 14, 'local_g0_0')
// (0, 14, 'span4_vert_b_8')
// (0, 15, 'span4_vert_b_4')
// (0, 16, 'span4_horz_1')
// (0, 16, 'span4_vert_b_0')
// (1, 16, 'sp4_h_r_12')
// (2, 16, 'sp4_h_r_25')
// (3, 16, 'sp4_h_r_36')
// (4, 16, 'sp4_h_l_36')
// (4, 16, 'sp4_h_r_5')
// (5, 16, 'sp4_h_r_16')
// (6, 16, 'sp4_h_r_29')
// (7, 16, 'sp4_h_r_40')
// (7, 17, 'sp4_r_v_b_40')
// (7, 18, 'sp4_r_v_b_29')
// (7, 19, 'sp4_r_v_b_16')
// (7, 20, 'sp4_r_v_b_5')
// (7, 21, 'sp4_r_v_b_44')
// (7, 22, 'neigh_op_tnr_2')
// (7, 22, 'sp4_r_v_b_33')
// (7, 23, 'neigh_op_rgt_2')
// (7, 23, 'sp4_r_v_b_20')
// (7, 24, 'neigh_op_bnr_2')
// (7, 24, 'sp4_r_v_b_9')
// (8, 16, 'sp4_h_l_40')
// (8, 16, 'sp4_v_t_40')
// (8, 17, 'sp4_v_b_40')
// (8, 18, 'sp4_v_b_29')
// (8, 19, 'sp4_v_b_16')
// (8, 20, 'sp4_v_b_5')
// (8, 20, 'sp4_v_t_44')
// (8, 21, 'sp4_v_b_44')
// (8, 22, 'neigh_op_top_2')
// (8, 22, 'sp4_v_b_33')
// (8, 23, 'ram/RDATA_13')
// (8, 23, 'sp4_v_b_20')
// (8, 24, 'neigh_op_bot_2')
// (8, 24, 'sp4_v_b_9')
// (9, 22, 'neigh_op_tnl_2')
// (9, 23, 'neigh_op_lft_2')
// (9, 24, 'neigh_op_bnl_2')

wire \data_out[28] ;
// (0, 13, 'io_1/D_OUT_0')
// (0, 13, 'io_1/PAD')
// (0, 13, 'local_g0_1')
// (0, 13, 'span4_horz_1')
// (1, 13, 'sp4_h_r_12')
// (2, 13, 'sp4_h_r_25')
// (3, 13, 'sp4_h_r_36')
// (4, 13, 'sp4_h_l_36')
// (4, 13, 'sp4_h_r_5')
// (5, 13, 'sp4_h_r_16')
// (6, 13, 'sp4_h_r_29')
// (7, 13, 'sp4_h_r_40')
// (7, 14, 'sp4_r_v_b_46')
// (7, 15, 'sp4_r_v_b_35')
// (7, 16, 'sp4_r_v_b_22')
// (7, 17, 'sp4_r_v_b_11')
// (7, 22, 'neigh_op_tnr_3')
// (7, 23, 'neigh_op_rgt_3')
// (7, 24, 'neigh_op_bnr_3')
// (8, 13, 'sp4_h_l_40')
// (8, 13, 'sp4_v_t_46')
// (8, 14, 'sp12_v_t_22')
// (8, 14, 'sp4_v_b_46')
// (8, 15, 'sp12_v_b_22')
// (8, 15, 'sp4_v_b_35')
// (8, 16, 'sp12_v_b_21')
// (8, 16, 'sp4_v_b_22')
// (8, 17, 'sp12_v_b_18')
// (8, 17, 'sp4_v_b_11')
// (8, 18, 'sp12_v_b_17')
// (8, 19, 'sp12_v_b_14')
// (8, 20, 'sp12_v_b_13')
// (8, 21, 'sp12_v_b_10')
// (8, 22, 'neigh_op_top_3')
// (8, 22, 'sp12_v_b_9')
// (8, 23, 'ram/RDATA_12')
// (8, 23, 'sp12_v_b_6')
// (8, 24, 'neigh_op_bot_3')
// (8, 24, 'sp12_v_b_5')
// (8, 25, 'sp12_v_b_2')
// (8, 26, 'sp12_v_b_1')
// (9, 22, 'neigh_op_tnl_3')
// (9, 23, 'neigh_op_lft_3')
// (9, 24, 'neigh_op_bnl_3')

wire \data_out[3] ;
// (0, 14, 'io_1/D_OUT_0')
// (0, 14, 'io_1/PAD')
// (0, 14, 'local_g1_0')
// (0, 14, 'span12_horz_0')
// (0, 26, 'span12_horz_0')
// (1, 14, 'sp12_h_r_3')
// (1, 26, 'sp12_h_r_3')
// (2, 14, 'sp12_h_r_4')
// (2, 26, 'sp12_h_r_4')
// (3, 14, 'sp12_h_r_7')
// (3, 26, 'sp12_h_r_7')
// (4, 14, 'sp12_h_r_8')
// (4, 26, 'sp12_h_r_8')
// (5, 14, 'sp12_h_r_11')
// (5, 26, 'sp12_h_r_11')
// (6, 14, 'sp12_h_r_12')
// (6, 26, 'sp12_h_r_12')
// (7, 14, 'sp12_h_r_15')
// (7, 25, 'neigh_op_tnr_4')
// (7, 26, 'neigh_op_rgt_4')
// (7, 26, 'sp12_h_r_15')
// (7, 27, 'neigh_op_bnr_4')
// (8, 14, 'sp12_h_r_16')
// (8, 25, 'neigh_op_top_4')
// (8, 26, 'ram/RDATA_3')
// (8, 26, 'sp12_h_r_16')
// (8, 27, 'neigh_op_bot_4')
// (9, 14, 'sp12_h_r_19')
// (9, 25, 'neigh_op_tnl_4')
// (9, 26, 'neigh_op_lft_4')
// (9, 26, 'sp12_h_r_19')
// (9, 27, 'neigh_op_bnl_4')
// (10, 14, 'sp12_h_r_20')
// (10, 26, 'sp12_h_r_20')
// (11, 14, 'sp12_h_r_23')
// (11, 26, 'sp12_h_r_23')
// (12, 14, 'sp12_h_l_23')
// (12, 14, 'sp12_v_t_23')
// (12, 15, 'sp12_v_b_23')
// (12, 16, 'sp12_v_b_20')
// (12, 17, 'sp12_v_b_19')
// (12, 18, 'sp12_v_b_16')
// (12, 19, 'sp12_v_b_15')
// (12, 20, 'sp12_v_b_12')
// (12, 21, 'sp12_v_b_11')
// (12, 22, 'sp12_v_b_8')
// (12, 23, 'sp12_v_b_7')
// (12, 24, 'sp12_v_b_4')
// (12, 25, 'sp12_v_b_3')
// (12, 26, 'sp12_h_l_23')
// (12, 26, 'sp12_v_b_0')

wire read_clk;
// (0, 15, 'span4_vert_t_12')
// (0, 16, 'span4_vert_b_12')
// (0, 17, 'io_0/D_IN_0')
// (0, 17, 'io_0/PAD')
// (0, 17, 'span4_vert_b_8')
// (0, 18, 'span4_vert_b_4')
// (0, 19, 'span4_horz_1')
// (0, 19, 'span4_vert_b_0')
// (1, 16, 'neigh_op_tnl_0')
// (1, 16, 'neigh_op_tnl_4')
// (1, 17, 'neigh_op_lft_0')
// (1, 17, 'neigh_op_lft_4')
// (1, 18, 'neigh_op_bnl_0')
// (1, 18, 'neigh_op_bnl_4')
// (1, 19, 'sp4_h_r_12')
// (2, 19, 'sp4_h_r_25')
// (3, 19, 'sp4_h_r_36')
// (4, 19, 'sp4_h_l_36')
// (4, 19, 'sp4_h_r_1')
// (5, 19, 'sp4_h_r_12')
// (6, 19, 'sp4_h_r_25')
// (7, 19, 'sp4_h_r_36')
// (7, 20, 'sp4_r_v_b_36')
// (7, 21, 'sp4_r_v_b_25')
// (7, 22, 'sp4_r_v_b_12')
// (7, 23, 'sp4_r_v_b_1')
// (7, 24, 'sp4_r_v_b_36')
// (7, 25, 'sp4_r_v_b_25')
// (7, 26, 'sp4_r_v_b_12')
// (7, 27, 'sp4_r_v_b_1')
// (8, 19, 'sp4_h_l_36')
// (8, 19, 'sp4_v_t_36')
// (8, 20, 'sp4_v_b_36')
// (8, 21, 'sp4_v_b_25')
// (8, 22, 'sp4_v_b_12')
// (8, 23, 'local_g1_1')
// (8, 23, 'ram/RCLK')
// (8, 23, 'sp4_v_b_1')
// (8, 23, 'sp4_v_t_36')
// (8, 24, 'sp4_v_b_36')
// (8, 25, 'local_g3_1')
// (8, 25, 'ram/RCLK')
// (8, 25, 'sp4_v_b_25')
// (8, 26, 'sp4_v_b_12')
// (8, 27, 'sp4_v_b_1')

wire \data_out[30] ;
// (0, 16, 'io_0/D_OUT_0')
// (0, 16, 'io_0/PAD')
// (0, 16, 'local_g0_0')
// (0, 16, 'span4_horz_0')
// (1, 16, 'sp4_h_r_13')
// (2, 16, 'sp4_h_r_24')
// (3, 16, 'sp4_h_r_37')
// (3, 17, 'sp4_r_v_b_43')
// (3, 18, 'sp4_r_v_b_30')
// (3, 19, 'sp4_r_v_b_19')
// (3, 20, 'sp4_r_v_b_6')
// (4, 16, 'sp4_h_l_37')
// (4, 16, 'sp4_v_t_43')
// (4, 17, 'sp4_v_b_43')
// (4, 18, 'sp4_v_b_30')
// (4, 19, 'sp4_v_b_19')
// (4, 20, 'sp4_h_r_1')
// (4, 20, 'sp4_v_b_6')
// (5, 20, 'sp4_h_r_12')
// (6, 20, 'sp4_h_r_25')
// (7, 20, 'sp4_h_r_36')
// (7, 21, 'sp4_r_v_b_42')
// (7, 22, 'neigh_op_tnr_1')
// (7, 22, 'sp4_r_v_b_31')
// (7, 23, 'neigh_op_rgt_1')
// (7, 23, 'sp4_r_v_b_18')
// (7, 24, 'neigh_op_bnr_1')
// (7, 24, 'sp4_r_v_b_7')
// (8, 20, 'sp4_h_l_36')
// (8, 20, 'sp4_v_t_42')
// (8, 21, 'sp4_v_b_42')
// (8, 22, 'neigh_op_top_1')
// (8, 22, 'sp4_v_b_31')
// (8, 23, 'ram/RDATA_14')
// (8, 23, 'sp4_v_b_18')
// (8, 24, 'neigh_op_bot_1')
// (8, 24, 'sp4_v_b_7')
// (9, 22, 'neigh_op_tnl_1')
// (9, 23, 'neigh_op_lft_1')
// (9, 24, 'neigh_op_bnl_1')

wire write_clk;
// (0, 16, 'io_1/D_IN_0')
// (0, 16, 'io_1/PAD')
// (0, 16, 'span12_horz_12')
// (1, 15, 'neigh_op_tnl_2')
// (1, 15, 'neigh_op_tnl_6')
// (1, 16, 'neigh_op_lft_2')
// (1, 16, 'neigh_op_lft_6')
// (1, 16, 'sp12_h_r_15')
// (1, 17, 'neigh_op_bnl_2')
// (1, 17, 'neigh_op_bnl_6')
// (2, 16, 'sp12_h_r_16')
// (3, 16, 'sp12_h_r_19')
// (4, 16, 'sp12_h_r_20')
// (5, 16, 'sp12_h_r_23')
// (5, 25, 'sp4_r_v_b_37')
// (5, 26, 'sp4_r_v_b_24')
// (5, 27, 'sp4_r_v_b_13')
// (5, 28, 'sp4_h_r_1')
// (5, 28, 'sp4_r_v_b_0')
// (6, 16, 'sp12_h_l_23')
// (6, 16, 'sp12_v_t_23')
// (6, 17, 'sp12_v_b_23')
// (6, 18, 'sp12_v_b_20')
// (6, 19, 'sp12_v_b_19')
// (6, 20, 'sp12_v_b_16')
// (6, 21, 'sp12_v_b_15')
// (6, 22, 'sp12_v_b_12')
// (6, 23, 'sp12_v_b_11')
// (6, 24, 'sp12_v_b_8')
// (6, 24, 'sp4_h_r_0')
// (6, 24, 'sp4_v_t_37')
// (6, 25, 'sp12_v_b_7')
// (6, 25, 'sp4_v_b_37')
// (6, 26, 'sp12_v_b_4')
// (6, 26, 'sp4_v_b_24')
// (6, 27, 'sp12_v_b_3')
// (6, 27, 'sp4_v_b_13')
// (6, 28, 'sp12_h_r_0')
// (6, 28, 'sp12_v_b_0')
// (6, 28, 'sp4_h_r_12')
// (6, 28, 'sp4_v_b_0')
// (7, 24, 'sp4_h_r_13')
// (7, 28, 'sp12_h_r_3')
// (7, 28, 'sp4_h_r_25')
// (8, 24, 'local_g2_0')
// (8, 24, 'ram/WCLK')
// (8, 24, 'sp4_h_r_24')
// (8, 25, 'sp4_r_v_b_36')
// (8, 26, 'local_g1_1')
// (8, 26, 'ram/WCLK')
// (8, 26, 'sp4_r_v_b_25')
// (8, 27, 'sp4_r_v_b_12')
// (8, 28, 'sp12_h_r_4')
// (8, 28, 'sp4_h_r_36')
// (8, 28, 'sp4_r_v_b_1')
// (9, 24, 'sp4_h_r_37')
// (9, 24, 'sp4_v_t_36')
// (9, 25, 'sp4_v_b_36')
// (9, 26, 'sp4_v_b_25')
// (9, 27, 'sp4_v_b_12')
// (9, 28, 'sp12_h_r_7')
// (9, 28, 'sp4_h_l_36')
// (9, 28, 'sp4_v_b_1')
// (10, 24, 'sp4_h_l_37')
// (10, 28, 'sp12_h_r_8')
// (11, 28, 'sp12_h_r_11')
// (12, 28, 'sp12_h_r_12')
// (13, 28, 'sp12_h_r_15')
// (14, 28, 'sp12_h_r_16')
// (15, 28, 'sp12_h_r_19')
// (16, 28, 'sp12_h_r_20')
// (17, 28, 'sp12_h_r_23')
// (18, 28, 'sp12_h_l_23')

wire \data_out[31] ;
// (0, 17, 'io_1/D_OUT_0')
// (0, 17, 'io_1/PAD')
// (0, 17, 'local_g0_1')
// (0, 17, 'span4_horz_1')
// (1, 17, 'sp4_h_r_12')
// (2, 17, 'sp4_h_r_25')
// (3, 17, 'sp4_h_r_36')
// (3, 18, 'sp4_r_v_b_36')
// (3, 19, 'sp4_r_v_b_25')
// (3, 20, 'sp4_r_v_b_12')
// (3, 21, 'sp4_r_v_b_1')
// (4, 17, 'sp4_h_l_36')
// (4, 17, 'sp4_v_t_36')
// (4, 18, 'sp4_v_b_36')
// (4, 19, 'sp4_v_b_25')
// (4, 20, 'sp4_v_b_12')
// (4, 21, 'sp4_h_r_8')
// (4, 21, 'sp4_v_b_1')
// (5, 21, 'sp4_h_r_21')
// (6, 21, 'sp4_h_r_32')
// (7, 21, 'sp4_h_r_45')
// (7, 22, 'neigh_op_tnr_0')
// (7, 22, 'sp4_r_v_b_45')
// (7, 23, 'neigh_op_rgt_0')
// (7, 23, 'sp4_r_v_b_32')
// (7, 24, 'neigh_op_bnr_0')
// (7, 24, 'sp4_r_v_b_21')
// (7, 25, 'sp4_r_v_b_8')
// (8, 21, 'sp4_h_l_45')
// (8, 21, 'sp4_v_t_45')
// (8, 22, 'neigh_op_top_0')
// (8, 22, 'sp4_v_b_45')
// (8, 23, 'ram/RDATA_15')
// (8, 23, 'sp4_v_b_32')
// (8, 24, 'neigh_op_bot_0')
// (8, 24, 'sp4_v_b_21')
// (8, 25, 'sp4_v_b_8')
// (9, 22, 'neigh_op_tnl_0')
// (9, 23, 'neigh_op_lft_0')
// (9, 24, 'neigh_op_bnl_0')

wire \data_out[4] ;
// (0, 18, 'io_0/D_OUT_0')
// (0, 18, 'io_0/PAD')
// (0, 18, 'local_g0_0')
// (0, 18, 'span4_horz_0')
// (1, 18, 'sp4_h_r_13')
// (2, 18, 'sp4_h_r_24')
// (3, 18, 'sp4_h_r_37')
// (3, 19, 'sp4_r_v_b_37')
// (3, 20, 'sp4_r_v_b_24')
// (3, 21, 'sp4_r_v_b_13')
// (3, 22, 'sp4_r_v_b_0')
// (4, 18, 'sp4_h_l_37')
// (4, 18, 'sp4_v_t_37')
// (4, 19, 'sp4_v_b_37')
// (4, 20, 'sp4_v_b_24')
// (4, 21, 'sp4_v_b_13')
// (4, 22, 'sp4_h_r_0')
// (4, 22, 'sp4_v_b_0')
// (5, 22, 'sp4_h_r_13')
// (6, 22, 'sp4_h_r_24')
// (7, 22, 'sp4_h_r_37')
// (7, 23, 'sp4_r_v_b_43')
// (7, 24, 'sp4_r_v_b_30')
// (7, 25, 'neigh_op_tnr_3')
// (7, 25, 'sp4_r_v_b_19')
// (7, 26, 'neigh_op_rgt_3')
// (7, 26, 'sp4_r_v_b_6')
// (7, 27, 'neigh_op_bnr_3')
// (8, 22, 'sp4_h_l_37')
// (8, 22, 'sp4_v_t_43')
// (8, 23, 'sp4_v_b_43')
// (8, 24, 'sp4_v_b_30')
// (8, 25, 'neigh_op_top_3')
// (8, 25, 'sp4_v_b_19')
// (8, 26, 'ram/RDATA_4')
// (8, 26, 'sp4_v_b_6')
// (8, 27, 'neigh_op_bot_3')
// (9, 25, 'neigh_op_tnl_3')
// (9, 26, 'neigh_op_lft_3')
// (9, 27, 'neigh_op_bnl_3')

wire \data_out[5] ;
// (0, 18, 'io_1/D_OUT_0')
// (0, 18, 'io_1/PAD')
// (0, 18, 'local_g0_1')
// (0, 18, 'span4_horz_1')
// (1, 18, 'sp4_h_r_12')
// (2, 18, 'sp4_h_r_25')
// (3, 18, 'sp4_h_r_36')
// (4, 18, 'sp4_h_l_36')
// (4, 18, 'sp4_h_r_1')
// (5, 18, 'sp4_h_r_12')
// (6, 18, 'sp4_h_r_25')
// (7, 18, 'sp4_h_r_36')
// (7, 19, 'sp4_r_v_b_42')
// (7, 20, 'sp4_r_v_b_31')
// (7, 21, 'sp4_r_v_b_18')
// (7, 22, 'sp4_r_v_b_7')
// (7, 23, 'sp4_r_v_b_41')
// (7, 24, 'sp4_r_v_b_28')
// (7, 25, 'neigh_op_tnr_2')
// (7, 25, 'sp4_r_v_b_17')
// (7, 26, 'neigh_op_rgt_2')
// (7, 26, 'sp4_r_v_b_4')
// (7, 27, 'neigh_op_bnr_2')
// (8, 18, 'sp4_h_l_36')
// (8, 18, 'sp4_v_t_42')
// (8, 19, 'sp4_v_b_42')
// (8, 20, 'sp4_v_b_31')
// (8, 21, 'sp4_v_b_18')
// (8, 22, 'sp4_v_b_7')
// (8, 22, 'sp4_v_t_41')
// (8, 23, 'sp4_v_b_41')
// (8, 24, 'sp4_v_b_28')
// (8, 25, 'neigh_op_top_2')
// (8, 25, 'sp4_v_b_17')
// (8, 26, 'ram/RDATA_5')
// (8, 26, 'sp4_v_b_4')
// (8, 27, 'neigh_op_bot_2')
// (9, 25, 'neigh_op_tnl_2')
// (9, 26, 'neigh_op_lft_2')
// (9, 27, 'neigh_op_bnl_2')

wire \data_out[9] ;
// (0, 18, 'span4_vert_t_13')
// (0, 19, 'span4_vert_b_13')
// (0, 20, 'io_1/D_OUT_0')
// (0, 20, 'io_1/PAD')
// (0, 20, 'local_g0_1')
// (0, 20, 'span4_vert_b_9')
// (0, 21, 'span4_vert_b_5')
// (0, 22, 'span4_horz_7')
// (0, 22, 'span4_vert_b_1')
// (1, 22, 'sp4_h_r_18')
// (2, 22, 'sp4_h_r_31')
// (3, 22, 'sp4_h_r_42')
// (4, 22, 'sp4_h_l_42')
// (4, 22, 'sp4_h_r_7')
// (5, 22, 'sp4_h_r_18')
// (6, 22, 'sp4_h_r_31')
// (7, 22, 'sp4_h_r_42')
// (7, 23, 'sp4_r_v_b_36')
// (7, 24, 'neigh_op_tnr_6')
// (7, 24, 'sp4_r_v_b_25')
// (7, 25, 'neigh_op_rgt_6')
// (7, 25, 'sp4_r_v_b_12')
// (7, 26, 'neigh_op_bnr_6')
// (7, 26, 'sp4_r_v_b_1')
// (8, 22, 'sp4_h_l_42')
// (8, 22, 'sp4_v_t_36')
// (8, 23, 'sp4_v_b_36')
// (8, 24, 'neigh_op_top_6')
// (8, 24, 'sp4_v_b_25')
// (8, 25, 'ram/RDATA_9')
// (8, 25, 'sp4_v_b_12')
// (8, 26, 'neigh_op_bot_6')
// (8, 26, 'sp4_v_b_1')
// (9, 24, 'neigh_op_tnl_6')
// (9, 25, 'neigh_op_lft_6')
// (9, 26, 'neigh_op_bnl_6')

wire \data_out[6] ;
// (0, 19, 'io_0/D_OUT_0')
// (0, 19, 'io_0/PAD')
// (0, 19, 'local_g0_0')
// (0, 19, 'span4_horz_16')
// (1, 19, 'sp4_h_r_29')
// (2, 19, 'sp4_h_r_40')
// (2, 20, 'sp4_r_v_b_40')
// (2, 21, 'sp4_r_v_b_29')
// (2, 22, 'sp4_r_v_b_16')
// (2, 23, 'sp4_r_v_b_5')
// (3, 14, 'sp12_v_t_22')
// (3, 15, 'sp12_v_b_22')
// (3, 16, 'sp12_v_b_21')
// (3, 17, 'sp12_v_b_18')
// (3, 18, 'sp12_v_b_17')
// (3, 19, 'sp12_v_b_14')
// (3, 19, 'sp4_h_l_40')
// (3, 19, 'sp4_v_t_40')
// (3, 20, 'sp12_v_b_13')
// (3, 20, 'sp4_v_b_40')
// (3, 21, 'sp12_v_b_10')
// (3, 21, 'sp4_v_b_29')
// (3, 22, 'sp12_v_b_9')
// (3, 22, 'sp4_v_b_16')
// (3, 23, 'sp12_v_b_6')
// (3, 23, 'sp4_v_b_5')
// (3, 24, 'sp12_v_b_5')
// (3, 25, 'sp12_v_b_2')
// (3, 26, 'sp12_h_r_1')
// (3, 26, 'sp12_v_b_1')
// (4, 26, 'sp12_h_r_2')
// (5, 26, 'sp12_h_r_5')
// (6, 26, 'sp12_h_r_6')
// (7, 25, 'neigh_op_tnr_1')
// (7, 26, 'neigh_op_rgt_1')
// (7, 26, 'sp12_h_r_9')
// (7, 27, 'neigh_op_bnr_1')
// (8, 25, 'neigh_op_top_1')
// (8, 26, 'ram/RDATA_6')
// (8, 26, 'sp12_h_r_10')
// (8, 27, 'neigh_op_bot_1')
// (9, 25, 'neigh_op_tnl_1')
// (9, 26, 'neigh_op_lft_1')
// (9, 26, 'sp12_h_r_13')
// (9, 27, 'neigh_op_bnl_1')
// (10, 26, 'sp12_h_r_14')
// (11, 26, 'sp12_h_r_17')
// (12, 26, 'sp12_h_r_18')
// (13, 26, 'sp12_h_r_21')
// (14, 26, 'sp12_h_r_22')
// (15, 26, 'sp12_h_l_22')

wire \data_out[7] ;
// (0, 19, 'io_1/D_OUT_0')
// (0, 19, 'io_1/PAD')
// (0, 19, 'local_g0_1')
// (0, 19, 'span4_horz_41')
// (1, 19, 'sp4_h_l_41')
// (1, 19, 'sp4_h_r_1')
// (2, 19, 'sp4_h_r_12')
// (3, 19, 'sp4_h_r_25')
// (4, 19, 'sp4_h_r_36')
// (5, 19, 'sp4_h_l_36')
// (5, 19, 'sp4_h_r_1')
// (6, 19, 'sp4_h_r_12')
// (7, 19, 'sp4_h_r_25')
// (7, 25, 'neigh_op_tnr_0')
// (7, 26, 'neigh_op_rgt_0')
// (7, 27, 'neigh_op_bnr_0')
// (8, 19, 'sp4_h_r_36')
// (8, 20, 'sp4_r_v_b_42')
// (8, 21, 'sp4_r_v_b_31')
// (8, 22, 'sp4_r_v_b_18')
// (8, 23, 'sp4_r_v_b_7')
// (8, 24, 'sp4_r_v_b_41')
// (8, 25, 'neigh_op_top_0')
// (8, 25, 'sp4_r_v_b_28')
// (8, 26, 'ram/RDATA_7')
// (8, 26, 'sp4_r_v_b_17')
// (8, 27, 'neigh_op_bot_0')
// (8, 27, 'sp4_r_v_b_4')
// (9, 19, 'sp4_h_l_36')
// (9, 19, 'sp4_v_t_42')
// (9, 20, 'sp4_v_b_42')
// (9, 21, 'sp4_v_b_31')
// (9, 22, 'sp4_v_b_18')
// (9, 23, 'sp4_v_b_7')
// (9, 23, 'sp4_v_t_41')
// (9, 24, 'sp4_v_b_41')
// (9, 25, 'neigh_op_tnl_0')
// (9, 25, 'sp4_v_b_28')
// (9, 26, 'neigh_op_lft_0')
// (9, 26, 'sp4_v_b_17')
// (9, 27, 'neigh_op_bnl_0')
// (9, 27, 'sp4_v_b_4')

wire \data_out[8] ;
// (0, 20, 'io_0/D_OUT_0')
// (0, 20, 'io_0/PAD')
// (0, 20, 'local_g1_1')
// (0, 20, 'span12_horz_9')
// (1, 20, 'sp12_h_r_10')
// (2, 20, 'sp12_h_r_13')
// (3, 20, 'sp12_h_r_14')
// (4, 20, 'sp12_h_r_17')
// (5, 20, 'sp12_h_r_18')
// (6, 20, 'sp12_h_r_21')
// (7, 20, 'sp12_h_r_22')
// (7, 24, 'neigh_op_tnr_7')
// (7, 25, 'neigh_op_rgt_7')
// (7, 26, 'neigh_op_bnr_7')
// (8, 20, 'sp12_h_l_22')
// (8, 20, 'sp12_v_t_22')
// (8, 21, 'sp12_v_b_22')
// (8, 22, 'sp12_v_b_21')
// (8, 23, 'sp12_v_b_18')
// (8, 24, 'neigh_op_top_7')
// (8, 24, 'sp12_v_b_17')
// (8, 25, 'ram/RDATA_8')
// (8, 25, 'sp12_v_b_14')
// (8, 26, 'neigh_op_bot_7')
// (8, 26, 'sp12_v_b_13')
// (8, 27, 'sp12_v_b_10')
// (8, 28, 'sp12_v_b_9')
// (8, 29, 'sp12_v_b_6')
// (8, 30, 'sp12_v_b_5')
// (8, 31, 'sp12_v_b_2')
// (8, 32, 'sp12_v_b_1')
// (9, 24, 'neigh_op_tnl_7')
// (9, 25, 'neigh_op_lft_7')
// (9, 26, 'neigh_op_bnl_7')

wire rd_en;
// (0, 21, 'io_1/D_IN_0')
// (0, 21, 'io_1/PAD')
// (0, 21, 'span12_horz_4')
// (1, 20, 'neigh_op_tnl_2')
// (1, 20, 'neigh_op_tnl_6')
// (1, 21, 'neigh_op_lft_2')
// (1, 21, 'neigh_op_lft_6')
// (1, 21, 'sp12_h_r_7')
// (1, 22, 'neigh_op_bnl_2')
// (1, 22, 'neigh_op_bnl_6')
// (2, 21, 'sp12_h_r_8')
// (3, 21, 'sp12_h_r_11')
// (4, 21, 'sp12_h_r_12')
// (5, 21, 'sp12_h_r_15')
// (5, 21, 'sp4_h_r_9')
// (5, 25, 'sp4_h_r_7')
// (6, 21, 'sp12_h_r_16')
// (6, 21, 'sp4_h_r_20')
// (6, 25, 'sp4_h_r_18')
// (7, 21, 'sp12_h_r_19')
// (7, 21, 'sp4_h_r_33')
// (7, 25, 'sp4_h_r_31')
// (8, 21, 'sp12_h_r_20')
// (8, 21, 'sp4_h_r_44')
// (8, 22, 'sp4_r_v_b_39')
// (8, 23, 'local_g0_2')
// (8, 23, 'ram/RCLKE')
// (8, 23, 'sp4_r_v_b_26')
// (8, 24, 'sp4_r_v_b_15')
// (8, 25, 'local_g2_2')
// (8, 25, 'ram/RCLKE')
// (8, 25, 'sp4_h_r_42')
// (8, 25, 'sp4_r_v_b_2')
// (9, 21, 'sp12_h_r_23')
// (9, 21, 'sp4_h_l_44')
// (9, 21, 'sp4_v_t_39')
// (9, 22, 'sp4_v_b_39')
// (9, 23, 'sp4_v_b_26')
// (9, 24, 'sp4_v_b_15')
// (9, 25, 'sp4_h_l_42')
// (9, 25, 'sp4_v_b_2')
// (10, 21, 'sp12_h_l_23')

wire \read_address[0] ;
// (0, 22, 'io_0/D_IN_0')
// (0, 22, 'io_0/PAD')
// (0, 22, 'span4_horz_0')
// (1, 21, 'neigh_op_tnl_0')
// (1, 21, 'neigh_op_tnl_4')
// (1, 22, 'neigh_op_lft_0')
// (1, 22, 'neigh_op_lft_4')
// (1, 22, 'sp4_h_r_13')
// (1, 23, 'neigh_op_bnl_0')
// (1, 23, 'neigh_op_bnl_4')
// (2, 22, 'sp4_h_r_24')
// (3, 22, 'sp4_h_r_37')
// (4, 22, 'sp4_h_l_37')
// (4, 22, 'sp4_h_r_3')
// (5, 22, 'sp4_h_r_14')
// (6, 22, 'sp4_h_r_27')
// (7, 22, 'sp4_h_r_38')
// (7, 23, 'sp4_r_v_b_45')
// (7, 24, 'sp4_r_v_b_32')
// (7, 25, 'sp4_r_v_b_21')
// (7, 26, 'sp4_r_v_b_8')
// (8, 22, 'sp4_h_l_38')
// (8, 22, 'sp4_v_t_45')
// (8, 23, 'local_g2_5')
// (8, 23, 'ram/RADDR_0')
// (8, 23, 'sp4_v_b_45')
// (8, 24, 'sp4_v_b_32')
// (8, 25, 'local_g0_5')
// (8, 25, 'ram/RADDR_0')
// (8, 25, 'sp4_v_b_21')
// (8, 26, 'sp4_v_b_8')

wire \read_address[1] ;
// (0, 22, 'io_1/D_IN_0')
// (0, 22, 'io_1/PAD')
// (0, 22, 'span4_horz_4')
// (1, 21, 'neigh_op_tnl_2')
// (1, 21, 'neigh_op_tnl_6')
// (1, 22, 'neigh_op_lft_2')
// (1, 22, 'neigh_op_lft_6')
// (1, 22, 'sp4_h_r_17')
// (1, 23, 'neigh_op_bnl_2')
// (1, 23, 'neigh_op_bnl_6')
// (2, 22, 'sp4_h_r_28')
// (3, 22, 'sp4_h_r_41')
// (4, 22, 'sp4_h_l_41')
// (4, 22, 'sp4_h_r_4')
// (5, 22, 'sp4_h_r_17')
// (6, 22, 'sp4_h_r_28')
// (7, 19, 'sp4_r_v_b_40')
// (7, 20, 'sp4_r_v_b_29')
// (7, 21, 'sp4_r_v_b_16')
// (7, 22, 'sp4_h_r_41')
// (7, 22, 'sp4_r_v_b_5')
// (7, 23, 'sp4_r_v_b_40')
// (7, 23, 'sp4_r_v_b_44')
// (7, 24, 'sp4_r_v_b_29')
// (7, 24, 'sp4_r_v_b_33')
// (7, 25, 'sp4_r_v_b_16')
// (7, 25, 'sp4_r_v_b_20')
// (7, 26, 'sp4_r_v_b_5')
// (7, 26, 'sp4_r_v_b_9')
// (8, 18, 'sp4_v_t_40')
// (8, 19, 'sp4_v_b_40')
// (8, 20, 'sp4_v_b_29')
// (8, 21, 'sp4_v_b_16')
// (8, 22, 'sp4_h_l_41')
// (8, 22, 'sp4_v_b_5')
// (8, 22, 'sp4_v_t_40')
// (8, 22, 'sp4_v_t_44')
// (8, 23, 'local_g2_0')
// (8, 23, 'ram/RADDR_1')
// (8, 23, 'sp4_v_b_40')
// (8, 23, 'sp4_v_b_44')
// (8, 24, 'sp4_v_b_29')
// (8, 24, 'sp4_v_b_33')
// (8, 25, 'local_g0_4')
// (8, 25, 'ram/RADDR_1')
// (8, 25, 'sp4_v_b_16')
// (8, 25, 'sp4_v_b_20')
// (8, 26, 'sp4_v_b_5')
// (8, 26, 'sp4_v_b_9')

wire \read_address[2] ;
// (0, 23, 'io_0/D_IN_0')
// (0, 23, 'io_0/PAD')
// (0, 23, 'span12_horz_0')
// (1, 22, 'neigh_op_tnl_0')
// (1, 22, 'neigh_op_tnl_4')
// (1, 23, 'neigh_op_lft_0')
// (1, 23, 'neigh_op_lft_4')
// (1, 23, 'sp12_h_r_3')
// (1, 23, 'sp4_h_r_3')
// (1, 24, 'neigh_op_bnl_0')
// (1, 24, 'neigh_op_bnl_4')
// (2, 23, 'sp12_h_r_4')
// (2, 23, 'sp4_h_r_14')
// (3, 23, 'sp12_h_r_7')
// (3, 23, 'sp4_h_r_27')
// (4, 23, 'sp12_h_r_8')
// (4, 23, 'sp4_h_r_38')
// (5, 23, 'sp12_h_r_11')
// (5, 23, 'sp4_h_l_38')
// (5, 23, 'sp4_h_r_3')
// (6, 23, 'sp12_h_r_12')
// (6, 23, 'sp4_h_r_14')
// (7, 23, 'sp12_h_r_15')
// (7, 23, 'sp4_h_r_27')
// (8, 23, 'local_g1_0')
// (8, 23, 'ram/RADDR_2')
// (8, 23, 'sp12_h_r_16')
// (8, 23, 'sp4_h_r_38')
// (8, 24, 'sp4_r_v_b_38')
// (8, 25, 'local_g0_3')
// (8, 25, 'ram/RADDR_2')
// (8, 25, 'sp4_r_v_b_27')
// (8, 26, 'sp4_r_v_b_14')
// (8, 27, 'sp4_r_v_b_3')
// (9, 23, 'sp12_h_r_19')
// (9, 23, 'sp4_h_l_38')
// (9, 23, 'sp4_v_t_38')
// (9, 24, 'sp4_v_b_38')
// (9, 25, 'sp4_v_b_27')
// (9, 26, 'sp4_v_b_14')
// (9, 27, 'sp4_v_b_3')
// (10, 23, 'sp12_h_r_20')
// (11, 23, 'sp12_h_r_23')
// (12, 23, 'sp12_h_l_23')

wire \read_address[3] ;
// (0, 23, 'io_1/D_IN_0')
// (0, 23, 'io_1/PAD')
// (0, 23, 'span12_horz_4')
// (1, 22, 'neigh_op_tnl_2')
// (1, 22, 'neigh_op_tnl_6')
// (1, 23, 'neigh_op_lft_2')
// (1, 23, 'neigh_op_lft_6')
// (1, 23, 'sp12_h_r_7')
// (1, 24, 'neigh_op_bnl_2')
// (1, 24, 'neigh_op_bnl_6')
// (2, 23, 'sp12_h_r_8')
// (3, 23, 'sp12_h_r_11')
// (4, 23, 'sp12_h_r_12')
// (5, 23, 'sp12_h_r_15')
// (5, 23, 'sp4_h_r_9')
// (6, 23, 'sp12_h_r_16')
// (6, 23, 'sp4_h_r_20')
// (7, 23, 'sp12_h_r_19')
// (7, 23, 'sp4_h_r_11')
// (7, 23, 'sp4_h_r_33')
// (8, 23, 'local_g0_6')
// (8, 23, 'ram/RADDR_3')
// (8, 23, 'sp12_h_r_20')
// (8, 23, 'sp4_h_r_22')
// (8, 23, 'sp4_h_r_44')
// (8, 24, 'sp4_r_v_b_39')
// (8, 25, 'local_g0_2')
// (8, 25, 'ram/RADDR_3')
// (8, 25, 'sp4_r_v_b_26')
// (8, 26, 'sp4_r_v_b_15')
// (8, 27, 'sp4_r_v_b_2')
// (9, 23, 'sp12_h_r_23')
// (9, 23, 'sp4_h_l_44')
// (9, 23, 'sp4_h_r_35')
// (9, 23, 'sp4_v_t_39')
// (9, 24, 'sp4_v_b_39')
// (9, 25, 'sp4_v_b_26')
// (9, 26, 'sp4_v_b_15')
// (9, 27, 'sp4_v_b_2')
// (10, 23, 'sp12_h_l_23')
// (10, 23, 'sp4_h_r_46')
// (11, 23, 'sp4_h_l_46')

wire \read_address[4] ;
// (0, 24, 'io_0/D_IN_0')
// (0, 24, 'io_0/PAD')
// (0, 24, 'span12_horz_8')
// (1, 23, 'neigh_op_tnl_0')
// (1, 23, 'neigh_op_tnl_4')
// (1, 24, 'neigh_op_lft_0')
// (1, 24, 'neigh_op_lft_4')
// (1, 24, 'sp12_h_r_11')
// (1, 25, 'neigh_op_bnl_0')
// (1, 25, 'neigh_op_bnl_4')
// (2, 24, 'sp12_h_r_12')
// (3, 24, 'sp12_h_r_15')
// (4, 24, 'sp12_h_r_16')
// (5, 24, 'sp12_h_r_19')
// (6, 24, 'sp12_h_r_20')
// (7, 21, 'sp4_r_v_b_41')
// (7, 22, 'sp4_r_v_b_28')
// (7, 23, 'sp4_r_v_b_17')
// (7, 24, 'sp12_h_r_23')
// (7, 24, 'sp4_r_v_b_4')
// (7, 25, 'sp4_r_v_b_45')
// (7, 26, 'sp4_r_v_b_32')
// (7, 27, 'sp4_r_v_b_21')
// (7, 28, 'sp4_r_v_b_8')
// (8, 20, 'sp4_v_t_41')
// (8, 21, 'sp4_v_b_41')
// (8, 22, 'sp4_v_b_28')
// (8, 23, 'local_g0_1')
// (8, 23, 'ram/RADDR_4')
// (8, 23, 'sp4_v_b_17')
// (8, 24, 'sp12_h_l_23')
// (8, 24, 'sp12_v_t_23')
// (8, 24, 'sp4_v_b_4')
// (8, 24, 'sp4_v_t_45')
// (8, 25, 'local_g2_7')
// (8, 25, 'ram/RADDR_4')
// (8, 25, 'sp12_v_b_23')
// (8, 25, 'sp4_v_b_45')
// (8, 26, 'sp12_v_b_20')
// (8, 26, 'sp4_v_b_32')
// (8, 27, 'sp12_v_b_19')
// (8, 27, 'sp4_v_b_21')
// (8, 28, 'sp12_v_b_16')
// (8, 28, 'sp4_v_b_8')
// (8, 29, 'sp12_v_b_15')
// (8, 30, 'sp12_v_b_12')
// (8, 31, 'sp12_v_b_11')
// (8, 32, 'sp12_v_b_8')
// (8, 33, 'span12_vert_7')

wire \read_address[5] ;
// (0, 24, 'io_1/D_IN_0')
// (0, 24, 'io_1/PAD')
// (0, 24, 'span4_horz_4')
// (1, 23, 'neigh_op_tnl_2')
// (1, 23, 'neigh_op_tnl_6')
// (1, 24, 'neigh_op_lft_2')
// (1, 24, 'neigh_op_lft_6')
// (1, 24, 'sp4_h_r_17')
// (1, 25, 'neigh_op_bnl_2')
// (1, 25, 'neigh_op_bnl_6')
// (2, 24, 'sp4_h_r_28')
// (3, 24, 'sp4_h_r_41')
// (4, 24, 'sp4_h_l_41')
// (4, 24, 'sp4_h_r_0')
// (5, 24, 'sp4_h_r_13')
// (6, 24, 'sp4_h_r_24')
// (7, 21, 'sp4_r_v_b_37')
// (7, 22, 'sp4_r_v_b_24')
// (7, 23, 'sp4_r_v_b_13')
// (7, 24, 'sp4_h_r_37')
// (7, 24, 'sp4_r_v_b_0')
// (7, 25, 'sp4_r_v_b_38')
// (7, 26, 'sp4_r_v_b_27')
// (7, 27, 'sp4_r_v_b_14')
// (7, 28, 'sp4_r_v_b_3')
// (8, 20, 'sp4_v_t_37')
// (8, 21, 'sp4_v_b_37')
// (8, 22, 'sp4_v_b_24')
// (8, 23, 'local_g1_5')
// (8, 23, 'ram/RADDR_5')
// (8, 23, 'sp4_v_b_13')
// (8, 24, 'sp4_h_l_37')
// (8, 24, 'sp4_v_b_0')
// (8, 24, 'sp4_v_t_38')
// (8, 25, 'local_g2_6')
// (8, 25, 'ram/RADDR_5')
// (8, 25, 'sp4_v_b_38')
// (8, 26, 'sp4_v_b_27')
// (8, 27, 'sp4_v_b_14')
// (8, 28, 'sp4_v_b_3')

wire wr_en;
// (0, 27, 'io_0/D_IN_0')
// (0, 27, 'io_0/PAD')
// (0, 27, 'span12_horz_0')
// (0, 27, 'span4_horz_0')
// (1, 26, 'neigh_op_tnl_0')
// (1, 26, 'neigh_op_tnl_4')
// (1, 27, 'neigh_op_lft_0')
// (1, 27, 'neigh_op_lft_4')
// (1, 27, 'sp12_h_r_3')
// (1, 27, 'sp4_h_r_13')
// (1, 28, 'neigh_op_bnl_0')
// (1, 28, 'neigh_op_bnl_4')
// (2, 27, 'sp12_h_r_4')
// (2, 27, 'sp4_h_r_24')
// (3, 27, 'sp12_h_r_7')
// (3, 27, 'sp4_h_r_37')
// (4, 27, 'sp12_h_r_8')
// (4, 27, 'sp4_h_l_37')
// (4, 27, 'sp4_h_r_0')
// (5, 27, 'sp12_h_r_11')
// (5, 27, 'sp4_h_r_13')
// (5, 27, 'sp4_h_r_7')
// (6, 27, 'sp12_h_r_12')
// (6, 27, 'sp4_h_r_18')
// (6, 27, 'sp4_h_r_24')
// (7, 24, 'sp4_r_v_b_43')
// (7, 25, 'sp4_r_v_b_30')
// (7, 26, 'sp4_r_v_b_19')
// (7, 27, 'sp12_h_r_15')
// (7, 27, 'sp4_h_r_31')
// (7, 27, 'sp4_h_r_37')
// (7, 27, 'sp4_r_v_b_6')
// (8, 23, 'sp4_v_t_43')
// (8, 24, 'local_g3_3')
// (8, 24, 'ram/WCLKE')
// (8, 24, 'sp4_r_v_b_42')
// (8, 24, 'sp4_v_b_43')
// (8, 25, 'sp4_r_v_b_31')
// (8, 25, 'sp4_v_b_30')
// (8, 26, 'local_g1_3')
// (8, 26, 'ram/WCLKE')
// (8, 26, 'sp4_r_v_b_18')
// (8, 26, 'sp4_v_b_19')
// (8, 27, 'sp12_h_r_16')
// (8, 27, 'sp4_h_l_37')
// (8, 27, 'sp4_h_r_42')
// (8, 27, 'sp4_r_v_b_7')
// (8, 27, 'sp4_v_b_6')
// (9, 23, 'sp4_v_t_42')
// (9, 24, 'local_g3_2')
// (9, 24, 'lutff_7/in_0')
// (9, 24, 'sp4_v_b_42')
// (9, 25, 'sp4_v_b_31')
// (9, 26, 'sp4_v_b_18')
// (9, 27, 'sp12_h_r_19')
// (9, 27, 'sp4_h_l_42')
// (9, 27, 'sp4_v_b_7')
// (10, 27, 'sp12_h_r_20')
// (11, 27, 'sp12_h_r_23')
// (12, 27, 'sp12_h_l_23')

wire \write_address[0] ;
// (0, 27, 'io_1/D_IN_0')
// (0, 27, 'io_1/PAD')
// (0, 27, 'span4_horz_4')
// (1, 26, 'neigh_op_tnl_2')
// (1, 26, 'neigh_op_tnl_6')
// (1, 27, 'neigh_op_lft_2')
// (1, 27, 'neigh_op_lft_6')
// (1, 27, 'sp4_h_r_17')
// (1, 28, 'neigh_op_bnl_2')
// (1, 28, 'neigh_op_bnl_6')
// (2, 27, 'sp4_h_r_28')
// (3, 27, 'sp4_h_r_41')
// (4, 27, 'sp4_h_l_41')
// (4, 27, 'sp4_h_r_4')
// (5, 27, 'sp4_h_r_17')
// (6, 27, 'sp4_h_r_28')
// (7, 24, 'sp4_r_v_b_41')
// (7, 24, 'sp4_r_v_b_47')
// (7, 25, 'sp4_r_v_b_28')
// (7, 25, 'sp4_r_v_b_34')
// (7, 26, 'sp4_r_v_b_17')
// (7, 26, 'sp4_r_v_b_23')
// (7, 27, 'sp4_h_r_41')
// (7, 27, 'sp4_r_v_b_10')
// (7, 27, 'sp4_r_v_b_4')
// (8, 23, 'sp4_v_t_41')
// (8, 23, 'sp4_v_t_47')
// (8, 24, 'local_g2_1')
// (8, 24, 'ram/WADDR_0')
// (8, 24, 'sp4_v_b_41')
// (8, 24, 'sp4_v_b_47')
// (8, 25, 'sp4_v_b_28')
// (8, 25, 'sp4_v_b_34')
// (8, 26, 'local_g0_7')
// (8, 26, 'ram/WADDR_0')
// (8, 26, 'sp4_v_b_17')
// (8, 26, 'sp4_v_b_23')
// (8, 27, 'sp4_h_l_41')
// (8, 27, 'sp4_v_b_10')
// (8, 27, 'sp4_v_b_4')

wire \write_address[1] ;
// (0, 28, 'io_0/D_IN_0')
// (0, 28, 'io_0/PAD')
// (0, 28, 'span12_horz_0')
// (1, 27, 'neigh_op_tnl_0')
// (1, 27, 'neigh_op_tnl_4')
// (1, 28, 'neigh_op_lft_0')
// (1, 28, 'neigh_op_lft_4')
// (1, 28, 'sp12_h_r_3')
// (1, 29, 'neigh_op_bnl_0')
// (1, 29, 'neigh_op_bnl_4')
// (2, 28, 'sp12_h_r_4')
// (3, 28, 'sp12_h_r_7')
// (4, 28, 'sp12_h_r_8')
// (5, 28, 'sp12_h_r_11')
// (6, 28, 'sp12_h_r_12')
// (7, 28, 'sp12_h_r_15')
// (8, 21, 'sp4_r_v_b_42')
// (8, 22, 'sp4_r_v_b_31')
// (8, 23, 'sp4_r_v_b_18')
// (8, 24, 'local_g1_7')
// (8, 24, 'ram/WADDR_1')
// (8, 24, 'sp4_r_v_b_7')
// (8, 25, 'sp4_r_v_b_41')
// (8, 26, 'local_g0_4')
// (8, 26, 'ram/WADDR_1')
// (8, 26, 'sp4_r_v_b_28')
// (8, 27, 'sp4_r_v_b_17')
// (8, 28, 'sp12_h_r_16')
// (8, 28, 'sp4_r_v_b_4')
// (9, 20, 'sp4_v_t_42')
// (9, 21, 'sp4_v_b_42')
// (9, 22, 'sp4_v_b_31')
// (9, 23, 'sp4_v_b_18')
// (9, 24, 'sp4_v_b_7')
// (9, 24, 'sp4_v_t_41')
// (9, 25, 'sp4_v_b_41')
// (9, 26, 'sp4_v_b_28')
// (9, 27, 'sp4_v_b_17')
// (9, 28, 'sp12_h_r_19')
// (9, 28, 'sp4_h_r_11')
// (9, 28, 'sp4_v_b_4')
// (10, 28, 'sp12_h_r_20')
// (10, 28, 'sp4_h_r_22')
// (11, 28, 'sp12_h_r_23')
// (11, 28, 'sp4_h_r_35')
// (12, 28, 'sp12_h_l_23')
// (12, 28, 'sp4_h_r_46')
// (13, 28, 'sp4_h_l_46')

wire \write_address[2] ;
// (0, 28, 'io_1/D_IN_0')
// (0, 28, 'io_1/PAD')
// (0, 28, 'span12_horz_4')
// (1, 27, 'neigh_op_tnl_2')
// (1, 27, 'neigh_op_tnl_6')
// (1, 28, 'neigh_op_lft_2')
// (1, 28, 'neigh_op_lft_6')
// (1, 28, 'sp12_h_r_7')
// (1, 29, 'neigh_op_bnl_2')
// (1, 29, 'neigh_op_bnl_6')
// (2, 28, 'sp12_h_r_8')
// (3, 28, 'sp12_h_r_11')
// (4, 28, 'sp12_h_r_12')
// (5, 28, 'sp12_h_r_15')
// (5, 28, 'sp4_h_r_9')
// (6, 28, 'sp12_h_r_16')
// (6, 28, 'sp4_h_r_20')
// (7, 28, 'sp12_h_r_19')
// (7, 28, 'sp4_h_r_33')
// (8, 21, 'sp4_r_v_b_43')
// (8, 22, 'sp4_r_v_b_30')
// (8, 23, 'sp4_r_v_b_19')
// (8, 24, 'local_g1_6')
// (8, 24, 'ram/WADDR_2')
// (8, 24, 'sp4_r_v_b_6')
// (8, 25, 'sp4_r_v_b_38')
// (8, 26, 'local_g0_3')
// (8, 26, 'ram/WADDR_2')
// (8, 26, 'sp4_r_v_b_27')
// (8, 27, 'sp4_r_v_b_14')
// (8, 28, 'sp12_h_r_20')
// (8, 28, 'sp4_h_r_44')
// (8, 28, 'sp4_r_v_b_3')
// (9, 20, 'sp4_v_t_43')
// (9, 21, 'sp4_v_b_43')
// (9, 22, 'sp4_v_b_30')
// (9, 23, 'sp4_v_b_19')
// (9, 24, 'sp4_v_b_6')
// (9, 24, 'sp4_v_t_38')
// (9, 25, 'sp4_v_b_38')
// (9, 26, 'sp4_v_b_27')
// (9, 27, 'sp4_v_b_14')
// (9, 28, 'sp12_h_r_23')
// (9, 28, 'sp4_h_l_44')
// (9, 28, 'sp4_v_b_3')
// (10, 28, 'sp12_h_l_23')

wire \write_address[3] ;
// (0, 30, 'io_0/D_IN_0')
// (0, 30, 'io_0/PAD')
// (0, 30, 'span12_horz_0')
// (1, 29, 'neigh_op_tnl_0')
// (1, 29, 'neigh_op_tnl_4')
// (1, 30, 'neigh_op_lft_0')
// (1, 30, 'neigh_op_lft_4')
// (1, 30, 'sp12_h_r_3')
// (1, 31, 'neigh_op_bnl_0')
// (1, 31, 'neigh_op_bnl_4')
// (2, 30, 'sp12_h_r_4')
// (3, 30, 'sp12_h_r_7')
// (4, 30, 'sp12_h_r_8')
// (5, 30, 'sp12_h_r_11')
// (6, 30, 'sp12_h_r_12')
// (7, 30, 'sp12_h_r_15')
// (8, 24, 'local_g0_6')
// (8, 24, 'ram/WADDR_3')
// (8, 24, 'sp4_h_r_6')
// (8, 26, 'local_g0_6')
// (8, 26, 'ram/WADDR_3')
// (8, 26, 'sp4_h_r_6')
// (8, 30, 'sp12_h_r_16')
// (9, 24, 'sp4_h_r_19')
// (9, 26, 'sp4_h_r_19')
// (9, 30, 'sp12_h_r_19')
// (10, 24, 'sp4_h_r_30')
// (10, 26, 'sp4_h_r_30')
// (10, 30, 'sp12_h_r_20')
// (11, 21, 'sp4_r_v_b_43')
// (11, 22, 'sp4_r_v_b_30')
// (11, 23, 'sp4_r_v_b_19')
// (11, 24, 'sp4_h_r_43')
// (11, 24, 'sp4_r_v_b_6')
// (11, 26, 'sp4_h_r_43')
// (11, 27, 'sp4_r_v_b_37')
// (11, 28, 'sp4_r_v_b_24')
// (11, 29, 'sp4_r_v_b_13')
// (11, 30, 'sp12_h_r_23')
// (11, 30, 'sp4_r_v_b_0')
// (12, 18, 'sp12_v_t_23')
// (12, 19, 'sp12_v_b_23')
// (12, 20, 'sp12_v_b_20')
// (12, 20, 'sp4_v_t_43')
// (12, 21, 'sp12_v_b_19')
// (12, 21, 'sp4_v_b_43')
// (12, 22, 'sp12_v_b_16')
// (12, 22, 'sp4_v_b_30')
// (12, 23, 'sp12_v_b_15')
// (12, 23, 'sp4_v_b_19')
// (12, 24, 'sp12_v_b_12')
// (12, 24, 'sp4_h_l_43')
// (12, 24, 'sp4_v_b_6')
// (12, 25, 'sp12_v_b_11')
// (12, 26, 'sp12_v_b_8')
// (12, 26, 'sp4_h_l_43')
// (12, 26, 'sp4_v_t_37')
// (12, 27, 'sp12_v_b_7')
// (12, 27, 'sp4_v_b_37')
// (12, 28, 'sp12_v_b_4')
// (12, 28, 'sp4_v_b_24')
// (12, 29, 'sp12_v_b_3')
// (12, 29, 'sp4_v_b_13')
// (12, 30, 'sp12_h_l_23')
// (12, 30, 'sp12_v_b_0')
// (12, 30, 'sp4_v_b_0')

wire \write_address[4] ;
// (0, 30, 'io_1/D_IN_0')
// (0, 30, 'io_1/PAD')
// (0, 30, 'span12_horz_4')
// (1, 29, 'neigh_op_tnl_2')
// (1, 29, 'neigh_op_tnl_6')
// (1, 30, 'neigh_op_lft_2')
// (1, 30, 'neigh_op_lft_6')
// (1, 30, 'sp12_h_r_7')
// (1, 31, 'neigh_op_bnl_2')
// (1, 31, 'neigh_op_bnl_6')
// (2, 30, 'sp12_h_r_8')
// (3, 30, 'sp12_h_r_11')
// (4, 30, 'sp12_h_r_12')
// (5, 30, 'sp12_h_r_15')
// (5, 30, 'sp4_h_r_9')
// (6, 30, 'sp12_h_r_16')
// (6, 30, 'sp4_h_r_20')
// (7, 30, 'sp12_h_r_19')
// (7, 30, 'sp4_h_r_33')
// (8, 23, 'sp4_r_v_b_40')
// (8, 23, 'sp4_r_v_b_44')
// (8, 24, 'local_g0_5')
// (8, 24, 'ram/WADDR_4')
// (8, 24, 'sp4_r_v_b_29')
// (8, 24, 'sp4_r_v_b_33')
// (8, 25, 'sp4_r_v_b_16')
// (8, 25, 'sp4_r_v_b_20')
// (8, 26, 'local_g2_1')
// (8, 26, 'ram/WADDR_4')
// (8, 26, 'sp4_r_v_b_5')
// (8, 26, 'sp4_r_v_b_9')
// (8, 27, 'sp4_r_v_b_44')
// (8, 28, 'sp4_r_v_b_33')
// (8, 29, 'sp4_r_v_b_20')
// (8, 30, 'sp12_h_r_20')
// (8, 30, 'sp4_h_r_44')
// (8, 30, 'sp4_r_v_b_9')
// (9, 22, 'sp4_v_t_40')
// (9, 22, 'sp4_v_t_44')
// (9, 23, 'sp4_v_b_40')
// (9, 23, 'sp4_v_b_44')
// (9, 24, 'sp4_v_b_29')
// (9, 24, 'sp4_v_b_33')
// (9, 25, 'sp4_v_b_16')
// (9, 25, 'sp4_v_b_20')
// (9, 26, 'sp4_v_b_5')
// (9, 26, 'sp4_v_b_9')
// (9, 26, 'sp4_v_t_44')
// (9, 27, 'sp4_v_b_44')
// (9, 28, 'sp4_v_b_33')
// (9, 29, 'sp4_v_b_20')
// (9, 30, 'sp12_h_r_23')
// (9, 30, 'sp4_h_l_44')
// (9, 30, 'sp4_v_b_9')
// (10, 30, 'sp12_h_l_23')

wire \write_address[5] ;
// (0, 31, 'io_0/D_IN_0')
// (0, 31, 'io_0/PAD')
// (0, 31, 'span12_horz_8')
// (1, 30, 'neigh_op_tnl_0')
// (1, 30, 'neigh_op_tnl_4')
// (1, 31, 'neigh_op_lft_0')
// (1, 31, 'neigh_op_lft_4')
// (1, 31, 'sp12_h_r_11')
// (1, 32, 'neigh_op_bnl_0')
// (1, 32, 'neigh_op_bnl_4')
// (2, 31, 'sp12_h_r_12')
// (3, 31, 'sp12_h_r_15')
// (4, 31, 'sp12_h_r_16')
// (5, 31, 'sp12_h_r_19')
// (6, 31, 'sp12_h_r_20')
// (7, 24, 'sp4_r_v_b_38')
// (7, 25, 'sp4_r_v_b_27')
// (7, 26, 'sp4_r_v_b_14')
// (7, 27, 'sp4_r_v_b_3')
// (7, 28, 'sp4_r_v_b_37')
// (7, 29, 'sp4_r_v_b_24')
// (7, 30, 'sp4_r_v_b_13')
// (7, 31, 'sp12_h_r_23')
// (7, 31, 'sp4_r_v_b_0')
// (8, 19, 'sp12_v_t_23')
// (8, 20, 'sp12_v_b_23')
// (8, 21, 'sp12_v_b_20')
// (8, 22, 'sp12_v_b_19')
// (8, 23, 'sp12_v_b_16')
// (8, 23, 'sp4_v_t_38')
// (8, 24, 'local_g2_6')
// (8, 24, 'ram/WADDR_5')
// (8, 24, 'sp12_v_b_15')
// (8, 24, 'sp4_v_b_38')
// (8, 25, 'sp12_v_b_12')
// (8, 25, 'sp4_v_b_27')
// (8, 26, 'local_g3_3')
// (8, 26, 'ram/WADDR_5')
// (8, 26, 'sp12_v_b_11')
// (8, 26, 'sp4_v_b_14')
// (8, 27, 'sp12_v_b_8')
// (8, 27, 'sp4_v_b_3')
// (8, 27, 'sp4_v_t_37')
// (8, 28, 'sp12_v_b_7')
// (8, 28, 'sp4_v_b_37')
// (8, 29, 'sp12_v_b_4')
// (8, 29, 'sp4_v_b_24')
// (8, 30, 'sp12_v_b_3')
// (8, 30, 'sp4_v_b_13')
// (8, 31, 'sp12_h_l_23')
// (8, 31, 'sp12_v_b_0')
// (8, 31, 'sp4_v_b_0')

wire \data_in[20] ;
// (1, 21, 'sp12_h_r_0')
// (2, 21, 'sp12_h_r_3')
// (3, 21, 'sp12_h_r_4')
// (4, 21, 'sp12_h_r_7')
// (5, 21, 'sp12_h_r_8')
// (6, 21, 'sp12_h_r_11')
// (7, 21, 'sp12_h_r_12')
// (7, 22, 'sp4_r_v_b_44')
// (7, 23, 'sp4_r_v_b_33')
// (7, 24, 'sp4_r_v_b_20')
// (7, 25, 'sp4_r_v_b_9')
// (8, 21, 'sp12_h_r_15')
// (8, 21, 'sp4_h_r_9')
// (8, 21, 'sp4_v_t_44')
// (8, 22, 'sp4_v_b_44')
// (8, 23, 'sp4_v_b_33')
// (8, 24, 'local_g0_4')
// (8, 24, 'ram/WDATA_4')
// (8, 24, 'sp4_v_b_20')
// (8, 25, 'sp4_v_b_9')
// (9, 21, 'sp12_h_r_16')
// (9, 21, 'sp4_h_r_20')
// (10, 21, 'sp12_h_r_19')
// (10, 21, 'sp4_h_r_33')
// (11, 21, 'sp12_h_r_20')
// (11, 21, 'sp4_h_r_44')
// (12, 21, 'sp12_h_r_23')
// (12, 21, 'sp4_h_l_44')
// (12, 32, 'neigh_op_tnr_0')
// (12, 32, 'neigh_op_tnr_4')
// (13, 21, 'sp12_h_l_23')
// (13, 21, 'sp12_v_t_23')
// (13, 22, 'sp12_v_b_23')
// (13, 23, 'sp12_v_b_20')
// (13, 24, 'sp12_v_b_19')
// (13, 25, 'sp12_v_b_16')
// (13, 26, 'sp12_v_b_15')
// (13, 27, 'sp12_v_b_12')
// (13, 28, 'sp12_v_b_11')
// (13, 29, 'sp12_v_b_8')
// (13, 30, 'sp12_v_b_7')
// (13, 31, 'sp12_v_b_4')
// (13, 32, 'neigh_op_top_0')
// (13, 32, 'neigh_op_top_4')
// (13, 32, 'sp12_v_b_3')
// (13, 33, 'io_0/D_IN_0')
// (13, 33, 'io_0/PAD')
// (13, 33, 'span12_vert_0')
// (14, 32, 'neigh_op_tnl_0')
// (14, 32, 'neigh_op_tnl_4')

wire \data_in[0] ;
// (1, 23, 'sp12_h_r_0')
// (1, 23, 'sp12_v_t_23')
// (1, 24, 'sp12_v_b_23')
// (1, 25, 'sp12_v_b_20')
// (1, 26, 'sp12_v_b_19')
// (1, 27, 'sp12_v_b_16')
// (1, 28, 'sp12_v_b_15')
// (1, 29, 'sp12_v_b_12')
// (1, 30, 'sp12_v_b_11')
// (1, 31, 'sp12_v_b_8')
// (1, 32, 'neigh_op_top_2')
// (1, 32, 'neigh_op_top_6')
// (1, 32, 'sp12_v_b_7')
// (1, 33, 'io_1/D_IN_0')
// (1, 33, 'io_1/PAD')
// (1, 33, 'span12_vert_4')
// (2, 23, 'sp12_h_r_3')
// (2, 32, 'neigh_op_tnl_2')
// (2, 32, 'neigh_op_tnl_6')
// (3, 23, 'sp12_h_r_4')
// (4, 23, 'sp12_h_r_7')
// (4, 23, 'sp4_h_r_5')
// (5, 23, 'sp12_h_r_8')
// (5, 23, 'sp4_h_r_16')
// (6, 23, 'sp12_h_r_11')
// (6, 23, 'sp4_h_r_29')
// (7, 23, 'sp12_h_r_12')
// (7, 23, 'sp4_h_r_40')
// (7, 24, 'sp4_r_v_b_40')
// (7, 25, 'sp4_r_v_b_29')
// (7, 26, 'sp4_r_v_b_16')
// (7, 27, 'sp4_r_v_b_5')
// (8, 23, 'sp12_h_r_15')
// (8, 23, 'sp4_h_l_40')
// (8, 23, 'sp4_v_t_40')
// (8, 24, 'sp4_v_b_40')
// (8, 25, 'sp4_v_b_29')
// (8, 26, 'local_g0_0')
// (8, 26, 'ram/WDATA_0')
// (8, 26, 'sp4_v_b_16')
// (8, 27, 'sp4_v_b_5')
// (9, 23, 'sp12_h_r_16')
// (10, 23, 'sp12_h_r_19')
// (11, 23, 'sp12_h_r_20')
// (12, 23, 'sp12_h_r_23')
// (13, 23, 'sp12_h_l_23')

wire \data_in[9] ;
// (1, 32, 'neigh_op_tnr_0')
// (1, 32, 'neigh_op_tnr_4')
// (2, 25, 'sp12_h_r_0')
// (2, 25, 'sp12_v_t_23')
// (2, 26, 'sp12_v_b_23')
// (2, 27, 'sp12_v_b_20')
// (2, 28, 'sp12_v_b_19')
// (2, 29, 'sp12_v_b_16')
// (2, 30, 'sp12_v_b_15')
// (2, 31, 'sp12_v_b_12')
// (2, 32, 'neigh_op_top_0')
// (2, 32, 'neigh_op_top_4')
// (2, 32, 'sp12_v_b_11')
// (2, 33, 'io_0/D_IN_0')
// (2, 33, 'io_0/PAD')
// (2, 33, 'span12_vert_8')
// (3, 25, 'sp12_h_r_3')
// (3, 32, 'neigh_op_tnl_0')
// (3, 32, 'neigh_op_tnl_4')
// (4, 25, 'sp12_h_r_4')
// (5, 25, 'sp12_h_r_7')
// (6, 25, 'sp12_h_r_8')
// (7, 25, 'sp12_h_r_11')
// (8, 25, 'local_g1_4')
// (8, 25, 'ram/WDATA_9')
// (8, 25, 'sp12_h_r_12')
// (9, 25, 'sp12_h_r_15')
// (10, 25, 'sp12_h_r_16')
// (11, 25, 'sp12_h_r_19')
// (12, 25, 'sp12_h_r_20')
// (13, 25, 'sp12_h_r_23')
// (14, 25, 'sp12_h_l_23')

wire \data_in[8] ;
// (1, 32, 'neigh_op_tnr_2')
// (1, 32, 'neigh_op_tnr_6')
// (2, 27, 'sp12_h_r_0')
// (2, 27, 'sp12_v_t_23')
// (2, 28, 'sp12_v_b_23')
// (2, 29, 'sp12_v_b_20')
// (2, 30, 'sp12_v_b_19')
// (2, 31, 'sp12_v_b_16')
// (2, 32, 'neigh_op_top_2')
// (2, 32, 'neigh_op_top_6')
// (2, 32, 'sp12_v_b_15')
// (2, 33, 'io_1/D_IN_0')
// (2, 33, 'io_1/PAD')
// (2, 33, 'span12_vert_12')
// (3, 27, 'sp12_h_r_3')
// (3, 32, 'neigh_op_tnl_2')
// (3, 32, 'neigh_op_tnl_6')
// (4, 27, 'sp12_h_r_4')
// (5, 27, 'sp12_h_r_7')
// (5, 27, 'sp4_h_r_5')
// (6, 27, 'sp12_h_r_8')
// (6, 27, 'sp4_h_r_16')
// (7, 27, 'sp12_h_r_11')
// (7, 27, 'sp4_h_r_29')
// (8, 24, 'sp4_r_v_b_46')
// (8, 25, 'local_g0_0')
// (8, 25, 'ram/WDATA_8')
// (8, 25, 'sp4_r_v_b_35')
// (8, 26, 'sp4_r_v_b_22')
// (8, 27, 'sp12_h_r_12')
// (8, 27, 'sp4_h_r_40')
// (8, 27, 'sp4_r_v_b_11')
// (9, 23, 'sp4_v_t_46')
// (9, 24, 'sp4_v_b_46')
// (9, 25, 'sp4_v_b_35')
// (9, 26, 'sp4_v_b_22')
// (9, 27, 'sp12_h_r_15')
// (9, 27, 'sp4_h_l_40')
// (9, 27, 'sp4_v_b_11')
// (10, 27, 'sp12_h_r_16')
// (11, 27, 'sp12_h_r_19')
// (12, 27, 'sp12_h_r_20')
// (13, 27, 'sp12_h_r_23')
// (14, 27, 'sp12_h_l_23')

wire \data_in[21] ;
// (2, 23, 'sp12_h_r_0')
// (3, 23, 'sp12_h_r_3')
// (4, 23, 'sp12_h_r_4')
// (5, 23, 'sp12_h_r_7')
// (5, 23, 'sp4_h_r_5')
// (6, 23, 'sp12_h_r_8')
// (6, 23, 'sp4_h_r_16')
// (7, 23, 'sp12_h_r_11')
// (7, 23, 'sp4_h_r_29')
// (8, 23, 'sp12_h_r_12')
// (8, 23, 'sp4_h_r_40')
// (8, 24, 'local_g3_0')
// (8, 24, 'ram/WDATA_5')
// (8, 24, 'sp4_r_v_b_40')
// (8, 25, 'sp4_r_v_b_29')
// (8, 26, 'sp4_r_v_b_16')
// (8, 27, 'sp4_r_v_b_5')
// (9, 23, 'sp12_h_r_15')
// (9, 23, 'sp4_h_l_40')
// (9, 23, 'sp4_v_t_40')
// (9, 24, 'sp4_v_b_40')
// (9, 25, 'sp4_v_b_29')
// (9, 26, 'sp4_v_b_16')
// (9, 27, 'sp4_v_b_5')
// (10, 23, 'sp12_h_r_16')
// (11, 23, 'sp12_h_r_19')
// (12, 23, 'sp12_h_r_20')
// (13, 23, 'sp12_h_r_23')
// (13, 32, 'neigh_op_tnr_2')
// (13, 32, 'neigh_op_tnr_6')
// (14, 23, 'sp12_h_l_23')
// (14, 23, 'sp12_v_t_23')
// (14, 24, 'sp12_v_b_23')
// (14, 25, 'sp12_v_b_20')
// (14, 26, 'sp12_v_b_19')
// (14, 27, 'sp12_v_b_16')
// (14, 28, 'sp12_v_b_15')
// (14, 29, 'sp12_v_b_12')
// (14, 30, 'sp12_v_b_11')
// (14, 31, 'sp12_v_b_8')
// (14, 32, 'neigh_op_top_2')
// (14, 32, 'neigh_op_top_6')
// (14, 32, 'sp12_v_b_7')
// (14, 33, 'io_1/D_IN_0')
// (14, 33, 'io_1/PAD')
// (14, 33, 'span12_vert_4')
// (15, 32, 'neigh_op_tnl_2')
// (15, 32, 'neigh_op_tnl_6')

wire \data_in[7] ;
// (2, 27, 'sp4_r_v_b_36')
// (2, 28, 'sp4_r_v_b_25')
// (2, 29, 'sp4_r_v_b_12')
// (2, 30, 'sp4_r_v_b_1')
// (2, 31, 'sp4_r_v_b_40')
// (2, 32, 'neigh_op_tnr_0')
// (2, 32, 'neigh_op_tnr_4')
// (2, 32, 'sp4_r_v_b_29')
// (3, 26, 'sp4_h_r_1')
// (3, 26, 'sp4_v_t_36')
// (3, 27, 'sp4_v_b_36')
// (3, 28, 'sp4_v_b_25')
// (3, 29, 'sp4_v_b_12')
// (3, 30, 'sp4_v_b_1')
// (3, 30, 'sp4_v_t_40')
// (3, 31, 'sp4_v_b_40')
// (3, 32, 'neigh_op_top_0')
// (3, 32, 'neigh_op_top_4')
// (3, 32, 'sp4_v_b_29')
// (3, 33, 'io_0/D_IN_0')
// (3, 33, 'io_0/PAD')
// (3, 33, 'span4_vert_16')
// (4, 26, 'sp4_h_r_12')
// (4, 32, 'neigh_op_tnl_0')
// (4, 32, 'neigh_op_tnl_4')
// (5, 26, 'sp4_h_r_25')
// (6, 26, 'sp4_h_r_36')
// (7, 26, 'sp4_h_l_36')
// (7, 26, 'sp4_h_r_4')
// (8, 26, 'local_g0_1')
// (8, 26, 'ram/WDATA_7')
// (8, 26, 'sp4_h_r_17')
// (9, 26, 'sp4_h_r_28')
// (10, 26, 'sp4_h_r_41')
// (11, 26, 'sp4_h_l_41')

wire \data_in[6] ;
// (2, 32, 'neigh_op_tnr_2')
// (2, 32, 'neigh_op_tnr_6')
// (3, 23, 'sp12_h_r_0')
// (3, 23, 'sp12_v_t_23')
// (3, 24, 'sp12_v_b_23')
// (3, 25, 'sp12_v_b_20')
// (3, 26, 'sp12_v_b_19')
// (3, 27, 'sp12_v_b_16')
// (3, 28, 'sp12_v_b_15')
// (3, 29, 'sp12_v_b_12')
// (3, 30, 'sp12_v_b_11')
// (3, 31, 'sp12_v_b_8')
// (3, 32, 'neigh_op_top_2')
// (3, 32, 'neigh_op_top_6')
// (3, 32, 'sp12_v_b_7')
// (3, 33, 'io_1/D_IN_0')
// (3, 33, 'io_1/PAD')
// (3, 33, 'span12_vert_4')
// (4, 23, 'sp12_h_r_3')
// (4, 32, 'neigh_op_tnl_2')
// (4, 32, 'neigh_op_tnl_6')
// (5, 23, 'sp12_h_r_4')
// (6, 23, 'sp12_h_r_7')
// (7, 23, 'sp12_h_r_8')
// (7, 24, 'sp4_r_v_b_42')
// (7, 25, 'sp4_r_v_b_31')
// (7, 26, 'sp4_r_v_b_18')
// (7, 27, 'sp4_r_v_b_7')
// (8, 23, 'sp12_h_r_11')
// (8, 23, 'sp4_h_r_7')
// (8, 23, 'sp4_v_t_42')
// (8, 24, 'sp4_v_b_42')
// (8, 25, 'sp4_v_b_31')
// (8, 26, 'local_g0_2')
// (8, 26, 'ram/WDATA_6')
// (8, 26, 'sp4_v_b_18')
// (8, 27, 'sp4_v_b_7')
// (9, 23, 'sp12_h_r_12')
// (9, 23, 'sp4_h_r_18')
// (10, 23, 'sp12_h_r_15')
// (10, 23, 'sp4_h_r_31')
// (11, 23, 'sp12_h_r_16')
// (11, 23, 'sp4_h_r_42')
// (12, 23, 'sp12_h_r_19')
// (12, 23, 'sp4_h_l_42')
// (13, 23, 'sp12_h_r_20')
// (14, 23, 'sp12_h_r_23')
// (15, 23, 'sp12_h_l_23')

wire \data_in[4] ;
// (3, 30, 'sp4_r_v_b_41')
// (3, 31, 'sp4_r_v_b_28')
// (3, 32, 'neigh_op_tnr_2')
// (3, 32, 'neigh_op_tnr_6')
// (3, 32, 'sp4_r_v_b_17')
// (4, 29, 'sp4_h_r_9')
// (4, 29, 'sp4_v_t_41')
// (4, 30, 'sp4_v_b_41')
// (4, 31, 'sp4_v_b_28')
// (4, 32, 'neigh_op_top_2')
// (4, 32, 'neigh_op_top_6')
// (4, 32, 'sp4_v_b_17')
// (4, 33, 'io_1/D_IN_0')
// (4, 33, 'io_1/PAD')
// (4, 33, 'span4_vert_4')
// (5, 29, 'sp4_h_r_20')
// (5, 32, 'neigh_op_tnl_2')
// (5, 32, 'neigh_op_tnl_6')
// (6, 29, 'sp4_h_r_33')
// (7, 26, 'sp4_r_v_b_44')
// (7, 27, 'sp4_r_v_b_33')
// (7, 28, 'sp4_r_v_b_20')
// (7, 29, 'sp4_h_r_44')
// (7, 29, 'sp4_r_v_b_9')
// (8, 25, 'sp4_v_t_44')
// (8, 26, 'local_g2_4')
// (8, 26, 'ram/WDATA_4')
// (8, 26, 'sp4_v_b_44')
// (8, 27, 'sp4_v_b_33')
// (8, 28, 'sp4_v_b_20')
// (8, 29, 'sp4_h_l_44')
// (8, 29, 'sp4_v_b_9')

wire \data_in[5] ;
// (3, 30, 'sp4_r_v_b_45')
// (3, 31, 'sp4_r_v_b_32')
// (3, 32, 'neigh_op_tnr_0')
// (3, 32, 'neigh_op_tnr_4')
// (3, 32, 'sp4_r_v_b_21')
// (4, 29, 'sp4_h_r_8')
// (4, 29, 'sp4_v_t_45')
// (4, 30, 'sp4_v_b_45')
// (4, 31, 'sp4_v_b_32')
// (4, 32, 'neigh_op_top_0')
// (4, 32, 'neigh_op_top_4')
// (4, 32, 'sp4_v_b_21')
// (4, 33, 'io_0/D_IN_0')
// (4, 33, 'io_0/PAD')
// (4, 33, 'span4_vert_8')
// (5, 29, 'sp4_h_r_21')
// (5, 32, 'neigh_op_tnl_0')
// (5, 32, 'neigh_op_tnl_4')
// (6, 29, 'sp4_h_r_32')
// (7, 26, 'sp4_r_v_b_39')
// (7, 27, 'sp4_r_v_b_26')
// (7, 28, 'sp4_r_v_b_15')
// (7, 29, 'sp4_h_r_45')
// (7, 29, 'sp4_r_v_b_2')
// (8, 25, 'sp4_v_t_39')
// (8, 26, 'local_g2_7')
// (8, 26, 'ram/WDATA_5')
// (8, 26, 'sp4_v_b_39')
// (8, 27, 'sp4_v_b_26')
// (8, 28, 'sp4_v_b_15')
// (8, 29, 'sp4_h_l_45')
// (8, 29, 'sp4_v_b_2')

wire \data_in[22] ;
// (4, 21, 'sp12_h_r_0')
// (5, 21, 'sp12_h_r_3')
// (6, 21, 'sp12_h_r_4')
// (7, 21, 'sp12_h_r_7')
// (8, 21, 'sp12_h_r_8')
// (8, 22, 'sp4_r_v_b_36')
// (8, 23, 'sp4_r_v_b_25')
// (8, 24, 'local_g2_4')
// (8, 24, 'ram/WDATA_6')
// (8, 24, 'sp4_r_v_b_12')
// (8, 25, 'sp4_r_v_b_1')
// (9, 21, 'sp12_h_r_11')
// (9, 21, 'sp4_h_r_7')
// (9, 21, 'sp4_v_t_36')
// (9, 22, 'sp4_v_b_36')
// (9, 23, 'sp4_v_b_25')
// (9, 24, 'sp4_v_b_12')
// (9, 25, 'sp4_v_b_1')
// (10, 21, 'sp12_h_r_12')
// (10, 21, 'sp4_h_r_18')
// (11, 21, 'sp12_h_r_15')
// (11, 21, 'sp4_h_r_31')
// (12, 21, 'sp12_h_r_16')
// (12, 21, 'sp4_h_r_42')
// (13, 21, 'sp12_h_r_19')
// (13, 21, 'sp4_h_l_42')
// (14, 21, 'sp12_h_r_20')
// (15, 21, 'sp12_h_r_23')
// (15, 32, 'neigh_op_tnr_0')
// (15, 32, 'neigh_op_tnr_4')
// (16, 21, 'sp12_h_l_23')
// (16, 21, 'sp12_v_t_23')
// (16, 22, 'sp12_v_b_23')
// (16, 23, 'sp12_v_b_20')
// (16, 24, 'sp12_v_b_19')
// (16, 25, 'sp12_v_b_16')
// (16, 26, 'sp12_v_b_15')
// (16, 27, 'sp12_v_b_12')
// (16, 28, 'sp12_v_b_11')
// (16, 29, 'sp12_v_b_8')
// (16, 30, 'sp12_v_b_7')
// (16, 31, 'sp12_v_b_4')
// (16, 32, 'neigh_op_top_0')
// (16, 32, 'neigh_op_top_4')
// (16, 32, 'sp12_v_b_3')
// (16, 33, 'io_0/D_IN_0')
// (16, 33, 'io_0/PAD')
// (16, 33, 'span12_vert_0')
// (17, 32, 'neigh_op_tnl_0')
// (17, 32, 'neigh_op_tnl_4')

wire \data_in[23] ;
// (4, 27, 'sp12_h_r_0')
// (5, 27, 'sp12_h_r_3')
// (6, 27, 'sp12_h_r_4')
// (7, 27, 'sp12_h_r_7')
// (8, 24, 'local_g2_5')
// (8, 24, 'ram/WDATA_7')
// (8, 24, 'sp4_r_v_b_37')
// (8, 25, 'sp4_r_v_b_24')
// (8, 26, 'sp4_r_v_b_13')
// (8, 27, 'sp12_h_r_8')
// (8, 27, 'sp4_r_v_b_0')
// (9, 23, 'sp4_v_t_37')
// (9, 24, 'sp4_v_b_37')
// (9, 25, 'sp4_v_b_24')
// (9, 26, 'sp4_v_b_13')
// (9, 27, 'sp12_h_r_11')
// (9, 27, 'sp4_h_r_7')
// (9, 27, 'sp4_v_b_0')
// (10, 27, 'sp12_h_r_12')
// (10, 27, 'sp4_h_r_18')
// (11, 27, 'sp12_h_r_15')
// (11, 27, 'sp4_h_r_31')
// (12, 27, 'sp12_h_r_16')
// (12, 27, 'sp4_h_r_42')
// (13, 27, 'sp12_h_r_19')
// (13, 27, 'sp4_h_l_42')
// (14, 27, 'sp12_h_r_20')
// (15, 27, 'sp12_h_r_23')
// (15, 32, 'neigh_op_tnr_2')
// (15, 32, 'neigh_op_tnr_6')
// (16, 27, 'sp12_h_l_23')
// (16, 27, 'sp12_v_t_23')
// (16, 28, 'sp12_v_b_23')
// (16, 29, 'sp12_v_b_20')
// (16, 30, 'sp12_v_b_19')
// (16, 31, 'sp12_v_b_16')
// (16, 32, 'neigh_op_top_2')
// (16, 32, 'neigh_op_top_6')
// (16, 32, 'sp12_v_b_15')
// (16, 33, 'io_1/D_IN_0')
// (16, 33, 'io_1/PAD')
// (16, 33, 'span12_vert_12')
// (17, 32, 'neigh_op_tnl_2')
// (17, 32, 'neigh_op_tnl_6')

wire \data_in[3] ;
// (4, 27, 'sp4_r_v_b_36')
// (4, 28, 'sp4_r_v_b_25')
// (4, 29, 'sp4_r_v_b_12')
// (4, 30, 'sp4_r_v_b_1')
// (4, 31, 'sp4_r_v_b_40')
// (4, 32, 'neigh_op_tnr_0')
// (4, 32, 'neigh_op_tnr_4')
// (4, 32, 'sp4_r_v_b_29')
// (5, 26, 'sp4_h_r_6')
// (5, 26, 'sp4_v_t_36')
// (5, 27, 'sp4_v_b_36')
// (5, 28, 'sp4_v_b_25')
// (5, 29, 'sp4_v_b_12')
// (5, 30, 'sp4_v_b_1')
// (5, 30, 'sp4_v_t_40')
// (5, 31, 'sp4_v_b_40')
// (5, 32, 'neigh_op_top_0')
// (5, 32, 'neigh_op_top_4')
// (5, 32, 'sp4_v_b_29')
// (5, 33, 'io_0/D_IN_0')
// (5, 33, 'io_0/PAD')
// (5, 33, 'span4_vert_16')
// (6, 26, 'sp4_h_r_19')
// (6, 32, 'neigh_op_tnl_0')
// (6, 32, 'neigh_op_tnl_4')
// (7, 26, 'sp4_h_r_30')
// (8, 26, 'local_g2_3')
// (8, 26, 'ram/WDATA_3')
// (8, 26, 'sp4_h_r_43')
// (9, 26, 'sp4_h_l_43')

wire \data_in[2] ;
// (4, 27, 'sp4_r_v_b_37')
// (4, 28, 'sp4_r_v_b_24')
// (4, 29, 'sp4_r_v_b_13')
// (4, 30, 'sp4_r_v_b_0')
// (4, 31, 'sp4_r_v_b_44')
// (4, 32, 'neigh_op_tnr_2')
// (4, 32, 'neigh_op_tnr_6')
// (4, 32, 'sp4_r_v_b_33')
// (5, 26, 'sp4_h_r_5')
// (5, 26, 'sp4_v_t_37')
// (5, 27, 'sp4_v_b_37')
// (5, 28, 'sp4_v_b_24')
// (5, 29, 'sp4_v_b_13')
// (5, 30, 'sp4_v_b_0')
// (5, 30, 'sp4_v_t_44')
// (5, 31, 'sp4_v_b_44')
// (5, 32, 'neigh_op_top_2')
// (5, 32, 'neigh_op_top_6')
// (5, 32, 'sp4_v_b_33')
// (5, 33, 'io_1/D_IN_0')
// (5, 33, 'io_1/PAD')
// (5, 33, 'span4_vert_20')
// (6, 26, 'sp4_h_r_16')
// (6, 32, 'neigh_op_tnl_2')
// (6, 32, 'neigh_op_tnl_6')
// (7, 26, 'sp4_h_r_29')
// (8, 26, 'local_g2_0')
// (8, 26, 'ram/WDATA_2')
// (8, 26, 'sp4_h_r_40')
// (9, 26, 'sp4_h_l_40')

wire \data_in[25] ;
// (5, 23, 'sp12_h_r_0')
// (6, 23, 'sp12_h_r_3')
// (7, 23, 'sp12_h_r_4')
// (8, 23, 'local_g0_7')
// (8, 23, 'ram/WDATA_9')
// (8, 23, 'sp12_h_r_7')
// (9, 23, 'sp12_h_r_8')
// (10, 23, 'sp12_h_r_11')
// (11, 23, 'sp12_h_r_12')
// (12, 23, 'sp12_h_r_15')
// (13, 23, 'sp12_h_r_16')
// (14, 23, 'sp12_h_r_19')
// (15, 23, 'sp12_h_r_20')
// (16, 23, 'sp12_h_r_23')
// (16, 32, 'neigh_op_tnr_2')
// (16, 32, 'neigh_op_tnr_6')
// (17, 23, 'sp12_h_l_23')
// (17, 23, 'sp12_v_t_23')
// (17, 24, 'sp12_v_b_23')
// (17, 25, 'sp12_v_b_20')
// (17, 26, 'sp12_v_b_19')
// (17, 27, 'sp12_v_b_16')
// (17, 28, 'sp12_v_b_15')
// (17, 29, 'sp12_v_b_12')
// (17, 30, 'sp12_v_b_11')
// (17, 31, 'sp12_v_b_8')
// (17, 32, 'neigh_op_top_2')
// (17, 32, 'neigh_op_top_6')
// (17, 32, 'sp12_v_b_7')
// (17, 33, 'io_1/D_IN_0')
// (17, 33, 'io_1/PAD')
// (17, 33, 'span12_vert_4')
// (18, 32, 'neigh_op_tnl_2')
// (18, 32, 'neigh_op_tnl_6')

wire \data_in[24] ;
// (5, 25, 'sp12_h_r_0')
// (6, 25, 'sp12_h_r_3')
// (7, 22, 'sp4_r_v_b_47')
// (7, 23, 'sp4_r_v_b_34')
// (7, 24, 'sp4_r_v_b_23')
// (7, 25, 'sp12_h_r_4')
// (7, 25, 'sp4_r_v_b_10')
// (8, 21, 'sp4_v_t_47')
// (8, 22, 'sp4_v_b_47')
// (8, 23, 'local_g2_2')
// (8, 23, 'ram/WDATA_8')
// (8, 23, 'sp4_v_b_34')
// (8, 24, 'sp4_v_b_23')
// (8, 25, 'sp12_h_r_7')
// (8, 25, 'sp4_h_r_5')
// (8, 25, 'sp4_v_b_10')
// (9, 25, 'sp12_h_r_8')
// (9, 25, 'sp4_h_r_16')
// (10, 25, 'sp12_h_r_11')
// (10, 25, 'sp4_h_r_29')
// (11, 25, 'sp12_h_r_12')
// (11, 25, 'sp4_h_r_40')
// (12, 25, 'sp12_h_r_15')
// (12, 25, 'sp4_h_l_40')
// (13, 25, 'sp12_h_r_16')
// (14, 25, 'sp12_h_r_19')
// (15, 25, 'sp12_h_r_20')
// (16, 25, 'sp12_h_r_23')
// (16, 32, 'neigh_op_tnr_0')
// (16, 32, 'neigh_op_tnr_4')
// (17, 25, 'sp12_h_l_23')
// (17, 25, 'sp12_v_t_23')
// (17, 26, 'sp12_v_b_23')
// (17, 27, 'sp12_v_b_20')
// (17, 28, 'sp12_v_b_19')
// (17, 29, 'sp12_v_b_16')
// (17, 30, 'sp12_v_b_15')
// (17, 31, 'sp12_v_b_12')
// (17, 32, 'neigh_op_top_0')
// (17, 32, 'neigh_op_top_4')
// (17, 32, 'sp12_v_b_11')
// (17, 33, 'io_0/D_IN_0')
// (17, 33, 'io_0/PAD')
// (17, 33, 'span12_vert_8')
// (18, 32, 'neigh_op_tnl_0')
// (18, 32, 'neigh_op_tnl_4')

wire n64;
// (5, 26, 'sp4_h_r_11')
// (6, 26, 'sp4_h_r_22')
// (7, 26, 'sp4_h_r_35')
// (8, 23, 'local_g2_7')
// (8, 23, 'local_g3_7')
// (8, 23, 'neigh_op_tnr_7')
// (8, 23, 'ram/MASK_10')
// (8, 23, 'ram/MASK_11')
// (8, 23, 'ram/MASK_12')
// (8, 23, 'ram/MASK_13')
// (8, 23, 'ram/MASK_14')
// (8, 23, 'ram/MASK_15')
// (8, 23, 'ram/MASK_8')
// (8, 23, 'ram/MASK_9')
// (8, 23, 'sp4_r_v_b_43')
// (8, 24, 'local_g2_7')
// (8, 24, 'local_g3_7')
// (8, 24, 'neigh_op_rgt_7')
// (8, 24, 'ram/MASK_0')
// (8, 24, 'ram/MASK_1')
// (8, 24, 'ram/MASK_2')
// (8, 24, 'ram/MASK_3')
// (8, 24, 'ram/MASK_4')
// (8, 24, 'ram/MASK_5')
// (8, 24, 'ram/MASK_6')
// (8, 24, 'ram/MASK_7')
// (8, 24, 'sp4_r_v_b_30')
// (8, 25, 'local_g0_7')
// (8, 25, 'local_g1_7')
// (8, 25, 'neigh_op_bnr_7')
// (8, 25, 'ram/MASK_10')
// (8, 25, 'ram/MASK_11')
// (8, 25, 'ram/MASK_12')
// (8, 25, 'ram/MASK_13')
// (8, 25, 'ram/MASK_14')
// (8, 25, 'ram/MASK_15')
// (8, 25, 'ram/MASK_8')
// (8, 25, 'ram/MASK_9')
// (8, 25, 'sp4_r_v_b_19')
// (8, 26, 'local_g1_6')
// (8, 26, 'local_g2_6')
// (8, 26, 'ram/MASK_0')
// (8, 26, 'ram/MASK_1')
// (8, 26, 'ram/MASK_2')
// (8, 26, 'ram/MASK_3')
// (8, 26, 'ram/MASK_4')
// (8, 26, 'ram/MASK_5')
// (8, 26, 'ram/MASK_6')
// (8, 26, 'ram/MASK_7')
// (8, 26, 'sp4_h_r_46')
// (8, 26, 'sp4_r_v_b_6')
// (9, 22, 'sp4_v_t_43')
// (9, 23, 'neigh_op_top_7')
// (9, 23, 'sp4_v_b_43')
// (9, 24, 'lutff_7/out')
// (9, 24, 'sp4_v_b_30')
// (9, 25, 'neigh_op_bot_7')
// (9, 25, 'sp4_v_b_19')
// (9, 26, 'sp4_h_l_46')
// (9, 26, 'sp4_v_b_6')
// (10, 23, 'neigh_op_tnl_7')
// (10, 24, 'neigh_op_lft_7')
// (10, 25, 'neigh_op_bnl_7')

wire \data_in[15] ;
// (5, 26, 'sp4_r_v_b_41')
// (5, 27, 'sp4_r_v_b_28')
// (5, 28, 'sp4_r_v_b_17')
// (5, 29, 'sp4_r_v_b_4')
// (5, 30, 'sp4_r_v_b_41')
// (5, 31, 'sp4_r_v_b_28')
// (5, 32, 'neigh_op_tnr_2')
// (5, 32, 'neigh_op_tnr_6')
// (5, 32, 'sp4_r_v_b_17')
// (6, 25, 'sp4_h_r_9')
// (6, 25, 'sp4_v_t_41')
// (6, 26, 'sp4_v_b_41')
// (6, 27, 'sp4_v_b_28')
// (6, 28, 'sp4_v_b_17')
// (6, 29, 'sp4_v_b_4')
// (6, 29, 'sp4_v_t_41')
// (6, 30, 'sp4_v_b_41')
// (6, 31, 'sp4_v_b_28')
// (6, 32, 'neigh_op_top_2')
// (6, 32, 'neigh_op_top_6')
// (6, 32, 'sp4_v_b_17')
// (6, 33, 'io_1/D_IN_0')
// (6, 33, 'io_1/PAD')
// (6, 33, 'span4_vert_4')
// (7, 25, 'sp4_h_r_20')
// (7, 32, 'neigh_op_tnl_2')
// (7, 32, 'neigh_op_tnl_6')
// (8, 25, 'local_g2_1')
// (8, 25, 'ram/WDATA_15')
// (8, 25, 'sp4_h_r_33')
// (9, 25, 'sp4_h_r_44')
// (10, 25, 'sp4_h_l_44')

wire \data_in[13] ;
// (6, 22, 'sp4_r_v_b_47')
// (6, 23, 'sp4_r_v_b_34')
// (6, 24, 'sp4_r_v_b_23')
// (6, 25, 'sp4_r_v_b_10')
// (6, 32, 'neigh_op_tnr_2')
// (6, 32, 'neigh_op_tnr_6')
// (7, 21, 'sp4_v_t_47')
// (7, 22, 'sp4_v_b_47')
// (7, 23, 'sp12_v_t_23')
// (7, 23, 'sp4_v_b_34')
// (7, 24, 'sp12_v_b_23')
// (7, 24, 'sp4_v_b_23')
// (7, 25, 'sp12_v_b_20')
// (7, 25, 'sp4_h_r_4')
// (7, 25, 'sp4_v_b_10')
// (7, 26, 'sp12_v_b_19')
// (7, 27, 'sp12_v_b_16')
// (7, 28, 'sp12_v_b_15')
// (7, 29, 'sp12_v_b_12')
// (7, 30, 'sp12_v_b_11')
// (7, 31, 'sp12_v_b_8')
// (7, 32, 'neigh_op_top_2')
// (7, 32, 'neigh_op_top_6')
// (7, 32, 'sp12_v_b_7')
// (7, 33, 'io_1/D_IN_0')
// (7, 33, 'io_1/PAD')
// (7, 33, 'span12_vert_4')
// (8, 25, 'local_g0_1')
// (8, 25, 'ram/WDATA_13')
// (8, 25, 'sp4_h_r_17')
// (8, 32, 'neigh_op_tnl_2')
// (8, 32, 'neigh_op_tnl_6')
// (9, 25, 'sp4_h_r_28')
// (10, 25, 'sp4_h_r_41')
// (11, 25, 'sp4_h_l_41')

wire \data_in[26] ;
// (6, 23, 'sp12_h_r_0')
// (7, 23, 'sp12_h_r_3')
// (8, 23, 'local_g0_4')
// (8, 23, 'ram/WDATA_10')
// (8, 23, 'sp12_h_r_4')
// (9, 23, 'sp12_h_r_7')
// (10, 23, 'sp12_h_r_8')
// (11, 23, 'sp12_h_r_11')
// (12, 23, 'sp12_h_r_12')
// (13, 23, 'sp12_h_r_15')
// (14, 23, 'sp12_h_r_16')
// (15, 23, 'sp12_h_r_19')
// (16, 23, 'sp12_h_r_20')
// (17, 23, 'sp12_h_r_23')
// (17, 32, 'neigh_op_tnr_2')
// (17, 32, 'neigh_op_tnr_6')
// (18, 23, 'sp12_h_l_23')
// (18, 23, 'sp12_v_t_23')
// (18, 24, 'sp12_v_b_23')
// (18, 25, 'sp12_v_b_20')
// (18, 26, 'sp12_v_b_19')
// (18, 27, 'sp12_v_b_16')
// (18, 28, 'sp12_v_b_15')
// (18, 29, 'sp12_v_b_12')
// (18, 30, 'sp12_v_b_11')
// (18, 31, 'sp12_v_b_8')
// (18, 32, 'neigh_op_top_2')
// (18, 32, 'neigh_op_top_6')
// (18, 32, 'sp12_v_b_7')
// (18, 33, 'io_1/D_IN_0')
// (18, 33, 'io_1/PAD')
// (18, 33, 'span12_vert_4')
// (19, 32, 'neigh_op_tnl_2')
// (19, 32, 'neigh_op_tnl_6')

wire \data_in[14] ;
// (6, 32, 'neigh_op_tnr_0')
// (6, 32, 'neigh_op_tnr_4')
// (7, 25, 'sp12_h_r_0')
// (7, 25, 'sp12_v_t_23')
// (7, 26, 'sp12_v_b_23')
// (7, 27, 'sp12_v_b_20')
// (7, 28, 'sp12_v_b_19')
// (7, 29, 'sp12_v_b_16')
// (7, 30, 'sp12_v_b_15')
// (7, 31, 'sp12_v_b_12')
// (7, 32, 'neigh_op_top_0')
// (7, 32, 'neigh_op_top_4')
// (7, 32, 'sp12_v_b_11')
// (7, 33, 'io_0/D_IN_0')
// (7, 33, 'io_0/PAD')
// (7, 33, 'span12_vert_8')
// (8, 25, 'local_g1_3')
// (8, 25, 'ram/WDATA_14')
// (8, 25, 'sp12_h_r_3')
// (8, 32, 'neigh_op_tnl_0')
// (8, 32, 'neigh_op_tnl_4')
// (9, 25, 'sp12_h_r_4')
// (10, 25, 'sp12_h_r_7')
// (11, 25, 'sp12_h_r_8')
// (12, 25, 'sp12_h_r_11')
// (13, 25, 'sp12_h_r_12')
// (14, 25, 'sp12_h_r_15')
// (15, 25, 'sp12_h_r_16')
// (16, 25, 'sp12_h_r_19')
// (17, 25, 'sp12_h_r_20')
// (18, 25, 'sp12_h_r_23')
// (19, 25, 'sp12_h_l_23')

wire \data_in[27] ;
// (7, 21, 'sp12_h_r_0')
// (7, 22, 'sp4_r_v_b_38')
// (7, 23, 'sp4_r_v_b_27')
// (7, 24, 'sp4_r_v_b_14')
// (7, 25, 'sp4_r_v_b_3')
// (8, 21, 'sp12_h_r_3')
// (8, 21, 'sp4_h_r_3')
// (8, 21, 'sp4_v_t_38')
// (8, 22, 'sp4_v_b_38')
// (8, 23, 'local_g2_3')
// (8, 23, 'ram/WDATA_11')
// (8, 23, 'sp4_v_b_27')
// (8, 24, 'sp4_v_b_14')
// (8, 25, 'sp4_v_b_3')
// (9, 21, 'sp12_h_r_4')
// (9, 21, 'sp4_h_r_14')
// (10, 21, 'sp12_h_r_7')
// (10, 21, 'sp4_h_r_27')
// (11, 21, 'sp12_h_r_8')
// (11, 21, 'sp4_h_r_38')
// (12, 21, 'sp12_h_r_11')
// (12, 21, 'sp4_h_l_38')
// (13, 21, 'sp12_h_r_12')
// (14, 21, 'sp12_h_r_15')
// (15, 21, 'sp12_h_r_16')
// (16, 21, 'sp12_h_r_19')
// (17, 21, 'sp12_h_r_20')
// (18, 21, 'sp12_h_r_23')
// (18, 32, 'neigh_op_tnr_0')
// (18, 32, 'neigh_op_tnr_4')
// (19, 21, 'sp12_h_l_23')
// (19, 21, 'sp12_v_t_23')
// (19, 22, 'sp12_v_b_23')
// (19, 23, 'sp12_v_b_20')
// (19, 24, 'sp12_v_b_19')
// (19, 25, 'sp12_v_b_16')
// (19, 26, 'sp12_v_b_15')
// (19, 27, 'sp12_v_b_12')
// (19, 28, 'sp12_v_b_11')
// (19, 29, 'sp12_v_b_8')
// (19, 30, 'sp12_v_b_7')
// (19, 31, 'sp12_v_b_4')
// (19, 32, 'neigh_op_top_0')
// (19, 32, 'neigh_op_top_4')
// (19, 32, 'sp12_v_b_3')
// (19, 33, 'io_0/D_IN_0')
// (19, 33, 'io_0/PAD')
// (19, 33, 'span12_vert_0')
// (20, 32, 'neigh_op_tnl_0')
// (20, 32, 'neigh_op_tnl_4')

wire \data_in[17] ;
// (7, 22, 'sp4_r_v_b_41')
// (7, 23, 'sp4_r_v_b_28')
// (7, 24, 'sp4_r_v_b_17')
// (7, 25, 'sp4_r_v_b_4')
// (7, 26, 'sp4_r_v_b_36')
// (7, 27, 'sp4_r_v_b_25')
// (7, 28, 'sp4_r_v_b_12')
// (7, 29, 'sp4_r_v_b_1')
// (7, 30, 'sp4_r_v_b_36')
// (7, 31, 'sp4_r_v_b_25')
// (7, 32, 'sp4_r_v_b_12')
// (8, 21, 'sp4_v_t_41')
// (8, 22, 'sp4_v_b_41')
// (8, 23, 'sp4_v_b_28')
// (8, 24, 'local_g0_1')
// (8, 24, 'ram/WDATA_1')
// (8, 24, 'sp4_v_b_17')
// (8, 25, 'sp4_v_b_4')
// (8, 25, 'sp4_v_t_36')
// (8, 26, 'sp4_v_b_36')
// (8, 27, 'sp4_v_b_25')
// (8, 28, 'sp4_v_b_12')
// (8, 29, 'sp4_v_b_1')
// (8, 29, 'sp4_v_t_36')
// (8, 30, 'sp4_v_b_36')
// (8, 31, 'sp4_v_b_25')
// (8, 32, 'sp4_v_b_12')
// (8, 33, 'span4_horz_r_0')
// (8, 33, 'span4_vert_1')
// (9, 33, 'span4_horz_r_4')
// (10, 32, 'neigh_op_tnr_0')
// (10, 32, 'neigh_op_tnr_4')
// (10, 33, 'span4_horz_r_8')
// (11, 32, 'neigh_op_top_0')
// (11, 32, 'neigh_op_top_4')
// (11, 33, 'io_0/D_IN_0')
// (11, 33, 'io_0/PAD')
// (11, 33, 'span4_horz_r_12')
// (12, 32, 'neigh_op_tnl_0')
// (12, 32, 'neigh_op_tnl_4')
// (12, 33, 'span4_horz_l_12')

wire \data_in[19] ;
// (7, 22, 'sp4_r_v_b_43')
// (7, 23, 'sp4_r_v_b_30')
// (7, 24, 'sp4_r_v_b_19')
// (7, 25, 'sp4_r_v_b_6')
// (7, 26, 'sp4_r_v_b_43')
// (7, 27, 'sp4_r_v_b_30')
// (7, 28, 'sp4_r_v_b_19')
// (7, 29, 'sp4_r_v_b_6')
// (8, 21, 'sp4_v_t_43')
// (8, 22, 'sp4_v_b_43')
// (8, 23, 'sp4_v_b_30')
// (8, 24, 'local_g0_3')
// (8, 24, 'ram/WDATA_3')
// (8, 24, 'sp4_v_b_19')
// (8, 25, 'sp4_v_b_6')
// (8, 25, 'sp4_v_t_43')
// (8, 26, 'sp4_v_b_43')
// (8, 27, 'sp4_v_b_30')
// (8, 28, 'sp4_v_b_19')
// (8, 29, 'sp4_h_r_6')
// (8, 29, 'sp4_v_b_6')
// (9, 29, 'sp4_h_r_19')
// (10, 29, 'sp4_h_r_30')
// (11, 29, 'sp4_h_r_43')
// (11, 30, 'sp4_r_v_b_37')
// (11, 31, 'sp4_r_v_b_24')
// (11, 32, 'neigh_op_tnr_0')
// (11, 32, 'neigh_op_tnr_4')
// (11, 32, 'sp4_r_v_b_13')
// (12, 29, 'sp4_h_l_43')
// (12, 29, 'sp4_v_t_37')
// (12, 30, 'sp4_v_b_37')
// (12, 31, 'sp4_v_b_24')
// (12, 32, 'neigh_op_top_0')
// (12, 32, 'neigh_op_top_4')
// (12, 32, 'sp4_v_b_13')
// (12, 33, 'io_0/D_IN_0')
// (12, 33, 'io_0/PAD')
// (12, 33, 'span4_vert_0')
// (13, 32, 'neigh_op_tnl_0')
// (13, 32, 'neigh_op_tnl_4')

wire \data_in[28] ;
// (7, 23, 'sp12_h_r_0')
// (8, 23, 'local_g1_3')
// (8, 23, 'ram/WDATA_12')
// (8, 23, 'sp12_h_r_3')
// (9, 23, 'sp12_h_r_4')
// (10, 23, 'sp12_h_r_7')
// (11, 23, 'sp12_h_r_8')
// (12, 23, 'sp12_h_r_11')
// (13, 23, 'sp12_h_r_12')
// (14, 23, 'sp12_h_r_15')
// (15, 23, 'sp12_h_r_16')
// (16, 23, 'sp12_h_r_19')
// (17, 23, 'sp12_h_r_20')
// (18, 23, 'sp12_h_r_23')
// (18, 32, 'neigh_op_tnr_2')
// (18, 32, 'neigh_op_tnr_6')
// (19, 23, 'sp12_h_l_23')
// (19, 23, 'sp12_v_t_23')
// (19, 24, 'sp12_v_b_23')
// (19, 25, 'sp12_v_b_20')
// (19, 26, 'sp12_v_b_19')
// (19, 27, 'sp12_v_b_16')
// (19, 28, 'sp12_v_b_15')
// (19, 29, 'sp12_v_b_12')
// (19, 30, 'sp12_v_b_11')
// (19, 31, 'sp12_v_b_8')
// (19, 32, 'neigh_op_top_2')
// (19, 32, 'neigh_op_top_6')
// (19, 32, 'sp12_v_b_7')
// (19, 33, 'io_1/D_IN_0')
// (19, 33, 'io_1/PAD')
// (19, 33, 'span12_vert_4')
// (20, 32, 'neigh_op_tnl_2')
// (20, 32, 'neigh_op_tnl_6')

wire \data_in[18] ;
// (7, 24, 'sp4_h_r_7')
// (8, 24, 'local_g0_2')
// (8, 24, 'ram/WDATA_2')
// (8, 24, 'sp4_h_r_18')
// (9, 24, 'sp4_h_r_31')
// (10, 24, 'sp4_h_r_42')
// (10, 25, 'sp4_r_v_b_36')
// (10, 26, 'sp4_r_v_b_25')
// (10, 27, 'sp4_r_v_b_12')
// (10, 28, 'sp4_r_v_b_1')
// (10, 29, 'sp4_r_v_b_36')
// (10, 30, 'sp4_r_v_b_25')
// (10, 31, 'sp4_r_v_b_12')
// (10, 32, 'neigh_op_tnr_2')
// (10, 32, 'neigh_op_tnr_6')
// (10, 32, 'sp4_r_v_b_1')
// (11, 24, 'sp4_h_l_42')
// (11, 24, 'sp4_v_t_36')
// (11, 25, 'sp4_v_b_36')
// (11, 26, 'sp4_v_b_25')
// (11, 27, 'sp4_v_b_12')
// (11, 28, 'sp4_v_b_1')
// (11, 28, 'sp4_v_t_36')
// (11, 29, 'sp4_v_b_36')
// (11, 30, 'sp4_v_b_25')
// (11, 31, 'sp4_v_b_12')
// (11, 32, 'neigh_op_top_2')
// (11, 32, 'neigh_op_top_6')
// (11, 32, 'sp4_v_b_1')
// (11, 32, 'sp4_v_t_36')
// (11, 33, 'io_1/D_IN_0')
// (11, 33, 'io_1/PAD')
// (11, 33, 'span4_vert_36')
// (12, 32, 'neigh_op_tnl_2')
// (12, 32, 'neigh_op_tnl_6')

wire \data_in[12] ;
// (7, 32, 'neigh_op_tnr_0')
// (7, 32, 'neigh_op_tnr_4')
// (8, 21, 'sp12_v_t_23')
// (8, 22, 'sp12_v_b_23')
// (8, 23, 'sp12_v_b_20')
// (8, 24, 'sp12_v_b_19')
// (8, 25, 'local_g2_0')
// (8, 25, 'ram/WDATA_12')
// (8, 25, 'sp12_v_b_16')
// (8, 26, 'sp12_v_b_15')
// (8, 27, 'sp12_v_b_12')
// (8, 28, 'sp12_v_b_11')
// (8, 29, 'sp12_v_b_8')
// (8, 30, 'sp12_v_b_7')
// (8, 31, 'sp12_v_b_4')
// (8, 32, 'neigh_op_top_0')
// (8, 32, 'neigh_op_top_4')
// (8, 32, 'sp12_v_b_3')
// (8, 33, 'io_0/D_IN_0')
// (8, 33, 'io_0/PAD')
// (8, 33, 'span12_vert_0')
// (9, 32, 'neigh_op_tnl_0')
// (9, 32, 'neigh_op_tnl_4')

wire \data_in[11] ;
// (7, 32, 'neigh_op_tnr_2')
// (7, 32, 'neigh_op_tnr_6')
// (8, 23, 'sp12_v_t_23')
// (8, 24, 'sp12_v_b_23')
// (8, 25, 'local_g3_4')
// (8, 25, 'ram/WDATA_11')
// (8, 25, 'sp12_v_b_20')
// (8, 26, 'sp12_v_b_19')
// (8, 27, 'sp12_v_b_16')
// (8, 28, 'sp12_v_b_15')
// (8, 29, 'sp12_v_b_12')
// (8, 30, 'sp12_v_b_11')
// (8, 31, 'sp12_v_b_8')
// (8, 32, 'neigh_op_top_2')
// (8, 32, 'neigh_op_top_6')
// (8, 32, 'sp12_v_b_7')
// (8, 33, 'io_1/D_IN_0')
// (8, 33, 'io_1/PAD')
// (8, 33, 'span12_vert_4')
// (9, 32, 'neigh_op_tnl_2')
// (9, 32, 'neigh_op_tnl_6')

wire \data_in[29] ;
// (8, 13, 'sp12_v_t_23')
// (8, 14, 'sp12_v_b_23')
// (8, 15, 'sp12_v_b_20')
// (8, 16, 'sp12_v_b_19')
// (8, 17, 'sp12_v_b_16')
// (8, 18, 'sp12_v_b_15')
// (8, 19, 'sp12_v_b_12')
// (8, 20, 'sp12_v_b_11')
// (8, 21, 'sp12_v_b_8')
// (8, 22, 'sp12_v_b_7')
// (8, 23, 'local_g3_4')
// (8, 23, 'ram/WDATA_13')
// (8, 23, 'sp12_v_b_4')
// (8, 24, 'sp12_v_b_3')
// (8, 25, 'sp12_h_r_0')
// (8, 25, 'sp12_v_b_0')
// (9, 25, 'sp12_h_r_3')
// (10, 25, 'sp12_h_r_4')
// (11, 25, 'sp12_h_r_7')
// (12, 25, 'sp12_h_r_8')
// (13, 25, 'sp12_h_r_11')
// (14, 25, 'sp12_h_r_12')
// (15, 25, 'sp12_h_r_15')
// (16, 25, 'sp12_h_r_16')
// (17, 25, 'sp12_h_r_19')
// (18, 25, 'sp12_h_r_20')
// (19, 25, 'sp12_h_r_23')
// (19, 32, 'neigh_op_tnr_0')
// (19, 32, 'neigh_op_tnr_4')
// (20, 25, 'sp12_h_l_23')
// (20, 25, 'sp12_v_t_23')
// (20, 26, 'sp12_v_b_23')
// (20, 27, 'sp12_v_b_20')
// (20, 28, 'sp12_v_b_19')
// (20, 29, 'sp12_v_b_16')
// (20, 30, 'sp12_v_b_15')
// (20, 31, 'sp12_v_b_12')
// (20, 32, 'neigh_op_top_0')
// (20, 32, 'neigh_op_top_4')
// (20, 32, 'sp12_v_b_11')
// (20, 33, 'io_0/D_IN_0')
// (20, 33, 'io_0/PAD')
// (20, 33, 'span12_vert_8')
// (21, 32, 'neigh_op_tnl_0')
// (21, 32, 'neigh_op_tnl_4')

wire n77;
// (8, 17, 'sp4_r_v_b_36')
// (8, 18, 'sp4_r_v_b_25')
// (8, 19, 'sp4_r_v_b_12')
// (8, 20, 'sp4_r_v_b_1')
// (8, 21, 'sp4_r_v_b_36')
// (8, 21, 'sp4_r_v_b_40')
// (8, 22, 'sp4_r_v_b_25')
// (8, 22, 'sp4_r_v_b_29')
// (8, 23, 'local_g2_4')
// (8, 23, 'ram/RE')
// (8, 23, 'sp4_r_v_b_12')
// (8, 23, 'sp4_r_v_b_16')
// (8, 24, 'local_g1_5')
// (8, 24, 'ram/WE')
// (8, 24, 'sp4_r_v_b_1')
// (8, 24, 'sp4_r_v_b_5')
// (8, 25, 'local_g3_5')
// (8, 25, 'neigh_op_tnr_5')
// (8, 25, 'ram/RE')
// (8, 25, 'sp4_r_v_b_39')
// (8, 26, 'local_g3_5')
// (8, 26, 'neigh_op_rgt_5')
// (8, 26, 'ram/WE')
// (8, 26, 'sp4_r_v_b_26')
// (8, 27, 'neigh_op_bnr_5')
// (8, 27, 'sp4_r_v_b_15')
// (8, 28, 'sp4_r_v_b_2')
// (9, 16, 'sp4_v_t_36')
// (9, 17, 'sp4_v_b_36')
// (9, 18, 'sp4_v_b_25')
// (9, 19, 'sp4_v_b_12')
// (9, 20, 'sp4_v_b_1')
// (9, 20, 'sp4_v_t_36')
// (9, 20, 'sp4_v_t_40')
// (9, 21, 'sp4_v_b_36')
// (9, 21, 'sp4_v_b_40')
// (9, 22, 'sp4_v_b_25')
// (9, 22, 'sp4_v_b_29')
// (9, 23, 'sp4_v_b_12')
// (9, 23, 'sp4_v_b_16')
// (9, 24, 'sp4_v_b_1')
// (9, 24, 'sp4_v_b_5')
// (9, 24, 'sp4_v_t_39')
// (9, 25, 'neigh_op_top_5')
// (9, 25, 'sp4_v_b_39')
// (9, 26, 'lutff_5/out')
// (9, 26, 'sp4_v_b_26')
// (9, 27, 'neigh_op_bot_5')
// (9, 27, 'sp4_v_b_15')
// (9, 28, 'sp4_v_b_2')
// (10, 25, 'neigh_op_tnl_5')
// (10, 26, 'neigh_op_lft_5')
// (10, 27, 'neigh_op_bnl_5')

wire \data_in[31] ;
// (8, 22, 'sp4_r_v_b_43')
// (8, 23, 'local_g1_6')
// (8, 23, 'ram/WDATA_15')
// (8, 23, 'sp4_r_v_b_30')
// (8, 24, 'sp4_r_v_b_19')
// (8, 25, 'sp4_r_v_b_6')
// (9, 21, 'sp4_v_t_43')
// (9, 22, 'sp4_v_b_43')
// (9, 23, 'sp4_v_b_30')
// (9, 24, 'sp4_v_b_19')
// (9, 25, 'sp4_h_r_1')
// (9, 25, 'sp4_v_b_6')
// (10, 25, 'sp12_h_r_0')
// (10, 25, 'sp4_h_r_12')
// (11, 25, 'sp12_h_r_3')
// (11, 25, 'sp4_h_r_25')
// (12, 25, 'sp12_h_r_4')
// (12, 25, 'sp4_h_r_36')
// (13, 25, 'sp12_h_r_7')
// (13, 25, 'sp4_h_l_36')
// (14, 25, 'sp12_h_r_8')
// (15, 25, 'sp12_h_r_11')
// (16, 25, 'sp12_h_r_12')
// (17, 25, 'sp12_h_r_15')
// (18, 25, 'sp12_h_r_16')
// (19, 25, 'sp12_h_r_19')
// (20, 25, 'sp12_h_r_20')
// (21, 25, 'sp12_h_r_23')
// (21, 32, 'neigh_op_tnr_0')
// (21, 32, 'neigh_op_tnr_4')
// (22, 25, 'sp12_h_l_23')
// (22, 25, 'sp12_v_t_23')
// (22, 26, 'sp12_v_b_23')
// (22, 27, 'sp12_v_b_20')
// (22, 28, 'sp12_v_b_19')
// (22, 29, 'sp12_v_b_16')
// (22, 30, 'sp12_v_b_15')
// (22, 31, 'sp12_v_b_12')
// (22, 32, 'neigh_op_top_0')
// (22, 32, 'neigh_op_top_4')
// (22, 32, 'sp12_v_b_11')
// (22, 33, 'io_0/D_IN_0')
// (22, 33, 'io_0/PAD')
// (22, 33, 'span12_vert_8')
// (23, 32, 'neigh_op_tnl_0')
// (23, 32, 'neigh_op_tnl_4')

wire \data_in[30] ;
// (8, 23, 'local_g0_0')
// (8, 23, 'ram/WDATA_14')
// (8, 23, 'sp12_h_r_0')
// (9, 23, 'sp12_h_r_3')
// (10, 23, 'sp12_h_r_4')
// (11, 23, 'sp12_h_r_7')
// (12, 23, 'sp12_h_r_8')
// (13, 23, 'sp12_h_r_11')
// (14, 23, 'sp12_h_r_12')
// (15, 23, 'sp12_h_r_15')
// (16, 23, 'sp12_h_r_16')
// (17, 23, 'sp12_h_r_19')
// (18, 23, 'sp12_h_r_20')
// (19, 23, 'sp12_h_r_23')
// (19, 32, 'neigh_op_tnr_2')
// (19, 32, 'neigh_op_tnr_6')
// (20, 23, 'sp12_h_l_23')
// (20, 23, 'sp12_v_t_23')
// (20, 24, 'sp12_v_b_23')
// (20, 25, 'sp12_v_b_20')
// (20, 26, 'sp12_v_b_19')
// (20, 27, 'sp12_v_b_16')
// (20, 28, 'sp12_v_b_15')
// (20, 29, 'sp12_v_b_12')
// (20, 30, 'sp12_v_b_11')
// (20, 31, 'sp12_v_b_8')
// (20, 32, 'neigh_op_top_2')
// (20, 32, 'neigh_op_top_6')
// (20, 32, 'sp12_v_b_7')
// (20, 33, 'io_1/D_IN_0')
// (20, 33, 'io_1/PAD')
// (20, 33, 'span12_vert_4')
// (21, 32, 'neigh_op_tnl_2')
// (21, 32, 'neigh_op_tnl_6')

wire \data_in[16] ;
// (8, 23, 'sp4_r_v_b_37')
// (8, 24, 'local_g0_0')
// (8, 24, 'ram/WDATA_0')
// (8, 24, 'sp4_r_v_b_24')
// (8, 25, 'sp4_r_v_b_13')
// (8, 26, 'sp4_r_v_b_0')
// (8, 27, 'sp4_r_v_b_37')
// (8, 28, 'sp4_r_v_b_24')
// (8, 29, 'sp4_r_v_b_13')
// (8, 30, 'sp4_r_v_b_0')
// (8, 31, 'sp4_r_v_b_37')
// (8, 32, 'sp4_r_v_b_24')
// (9, 22, 'sp4_v_t_37')
// (9, 23, 'sp4_v_b_37')
// (9, 24, 'sp4_v_b_24')
// (9, 25, 'sp4_v_b_13')
// (9, 26, 'sp4_v_b_0')
// (9, 26, 'sp4_v_t_37')
// (9, 27, 'sp4_v_b_37')
// (9, 28, 'sp4_v_b_24')
// (9, 29, 'sp4_v_b_13')
// (9, 30, 'sp4_v_b_0')
// (9, 30, 'sp4_v_t_37')
// (9, 31, 'sp4_v_b_37')
// (9, 32, 'neigh_op_tnr_2')
// (9, 32, 'neigh_op_tnr_6')
// (9, 32, 'sp4_v_b_24')
// (9, 33, 'span4_horz_r_2')
// (9, 33, 'span4_vert_13')
// (10, 32, 'neigh_op_top_2')
// (10, 32, 'neigh_op_top_6')
// (10, 33, 'io_1/D_IN_0')
// (10, 33, 'io_1/PAD')
// (10, 33, 'span4_horz_r_6')
// (11, 32, 'neigh_op_tnl_2')
// (11, 32, 'neigh_op_tnl_6')
// (11, 33, 'span4_horz_r_10')
// (12, 33, 'span4_horz_r_14')
// (13, 33, 'span4_horz_l_14')

wire \data_in[10] ;
// (8, 24, 'sp4_r_v_b_43')
// (8, 25, 'local_g0_6')
// (8, 25, 'ram/WDATA_10')
// (8, 25, 'sp4_r_v_b_30')
// (8, 26, 'sp4_r_v_b_19')
// (8, 27, 'sp4_r_v_b_6')
// (8, 32, 'neigh_op_tnr_0')
// (8, 32, 'neigh_op_tnr_4')
// (9, 21, 'sp12_v_t_23')
// (9, 22, 'sp12_v_b_23')
// (9, 23, 'sp12_v_b_20')
// (9, 23, 'sp4_v_t_43')
// (9, 24, 'sp12_v_b_19')
// (9, 24, 'sp4_v_b_43')
// (9, 25, 'sp12_v_b_16')
// (9, 25, 'sp4_v_b_30')
// (9, 26, 'sp12_v_b_15')
// (9, 26, 'sp4_v_b_19')
// (9, 27, 'sp12_v_b_12')
// (9, 27, 'sp4_v_b_6')
// (9, 28, 'sp12_v_b_11')
// (9, 29, 'sp12_v_b_8')
// (9, 30, 'sp12_v_b_7')
// (9, 31, 'sp12_v_b_4')
// (9, 32, 'neigh_op_top_0')
// (9, 32, 'neigh_op_top_4')
// (9, 32, 'sp12_v_b_3')
// (9, 33, 'io_0/D_IN_0')
// (9, 33, 'io_0/PAD')
// (9, 33, 'span12_vert_0')
// (10, 32, 'neigh_op_tnl_0')
// (10, 32, 'neigh_op_tnl_4')

wire \data_in[1] ;
// (8, 26, 'local_g2_5')
// (8, 26, 'ram/WDATA_1')
// (8, 26, 'sp4_r_v_b_37')
// (8, 27, 'sp4_r_v_b_24')
// (8, 28, 'sp4_r_v_b_13')
// (8, 29, 'sp4_r_v_b_0')
// (8, 30, 'sp4_r_v_b_41')
// (8, 31, 'sp4_r_v_b_28')
// (8, 32, 'neigh_op_tnr_2')
// (8, 32, 'neigh_op_tnr_6')
// (8, 32, 'sp4_r_v_b_17')
// (9, 25, 'sp4_v_t_37')
// (9, 26, 'sp4_v_b_37')
// (9, 27, 'sp4_v_b_24')
// (9, 28, 'sp4_v_b_13')
// (9, 29, 'sp4_v_b_0')
// (9, 29, 'sp4_v_t_41')
// (9, 30, 'sp4_v_b_41')
// (9, 31, 'sp4_v_b_28')
// (9, 32, 'neigh_op_top_2')
// (9, 32, 'neigh_op_top_6')
// (9, 32, 'sp4_v_b_17')
// (9, 33, 'io_1/D_IN_0')
// (9, 33, 'io_1/PAD')
// (9, 33, 'span4_vert_4')
// (10, 32, 'neigh_op_tnl_2')
// (10, 32, 'neigh_op_tnl_6')

wire open_0;
wire open_1;
wire open_2;
wire open_3;
wire open_4;
wire open_5;
wire open_6;
wire open_7;
wire open_8;
wire open_9;
wire open_10;
wire open_11;
wire open_12;
wire open_13;
wire open_14;
wire open_15;
wire n83;
// (9, 24, 'lutff_7/lout')

wire n84;
// (9, 26, 'lutff_5/lout')

// RAM TILE 8 25
SB_RAM40_4K #(
  .READ_MODE(0),
  .WRITE_MODE(0),
  .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
) ram40_8_25 (
  .WADDR({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \write_address[5] , \write_address[4] , \write_address[3] , \write_address[2] , \write_address[1] , \write_address[0] }),
  .RADDR({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \read_address[5] , \read_address[4] , \read_address[3] , \read_address[2] , \read_address[1] , \read_address[0] }),
  .MASK({n64, n64, n64, n64, n64, n64, n64, n64, n64, n64, n64, n64, n64, n64, n64, n64}),
  .WDATA({\data_in[15] , \data_in[14] , \data_in[13] , \data_in[12] , \data_in[11] , \data_in[10] , \data_in[9] , \data_in[8] , \data_in[7] , \data_in[6] , \data_in[5] , \data_in[4] , \data_in[3] , \data_in[2] , \data_in[1] , \data_in[0] }),
  .RDATA({\data_out[15] , \data_out[14] , \data_out[13] , \data_out[12] , \data_out[11] , \data_out[10] , \data_out[9] , \data_out[8] , \data_out[7] , \data_out[6] , \data_out[5] , \data_out[4] , \data_out[3] , \data_out[2] , \data_out[1] , \data_out[0] }),
  .WE(n77),
  .WCLKE(wr_en),
  .WCLK(write_clk),
  .RE(n77),
  .RCLKE(rd_en),
  .RCLK(read_clk)
);

// RAM TILE 8 23
SB_RAM40_4K #(
  .READ_MODE(0),
  .WRITE_MODE(0),
  .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
) ram40_8_23 (
  .WADDR({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \write_address[5] , \write_address[4] , \write_address[3] , \write_address[2] , \write_address[1] , \write_address[0] }),
  .RADDR({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \read_address[5] , \read_address[4] , \read_address[3] , \read_address[2] , \read_address[1] , \read_address[0] }),
  .MASK({n64, n64, n64, n64, n64, n64, n64, n64, n64, n64, n64, n64, n64, n64, n64, n64}),
  .WDATA({\data_in[31] , \data_in[30] , \data_in[29] , \data_in[28] , \data_in[27] , \data_in[26] , \data_in[25] , \data_in[24] , \data_in[23] , \data_in[22] , \data_in[21] , \data_in[20] , \data_in[19] , \data_in[18] , \data_in[17] , \data_in[16] }),
  .RDATA({\data_out[31] , \data_out[30] , \data_out[29] , \data_out[28] , \data_out[27] , \data_out[26] , \data_out[25] , \data_out[24] , \data_out[23] , \data_out[22] , \data_out[21] , \data_out[20] , \data_out[19] , \data_out[18] , \data_out[17] , \data_out[16] }),
  .WE(n77),
  .WCLKE(wr_en),
  .WCLK(write_clk),
  .RE(n77),
  .RCLKE(rd_en),
  .RCLK(read_clk)
);

assign n83 = /* LUT    9 24  7 */ !wr_en;
assign n84 = /* LUT    9 26  5 */ 1'b1;
/* FF  9 24  7 */ assign n64 = n83;
/* FF  9 26  5 */ assign n77 = n84;

// Warning: unmatched port '\write_address[6] '
// Warning: unmatched port '\read_address[6] '
// Warning: unmatched port '\write_address[7] '
// Warning: unmatched port '\read_address[7] '

endmodule

