module top(
  input clk,
  input down1,
  input down2,
  input rst,
  input up1,
  input up2,
  output b,
  output g,
  output hs,
  output r,
  output vs
  );
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRL0;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRL1;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRL10;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRL11;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRL12;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRL13;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRL14;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRL15;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRL2;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRL3;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRL4;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRL5;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRL6;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRL7;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRL8;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRL9;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRU0;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRU1;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRU10;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRU11;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRU12;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRU13;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRU14;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRU2;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRU3;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRU4;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRU5;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRU6;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRU7;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRU8;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRU9;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRL0;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRL1;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRL10;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRL11;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRL12;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRL13;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRL14;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRL15;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRL2;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRL3;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRL4;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRL5;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRL6;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRL7;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRL8;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRL9;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRU0;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRU1;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRU10;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRU11;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRU12;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRU13;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRU14;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRU2;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRU3;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRU4;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRU5;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRU6;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRU7;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRU8;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRU9;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_CLKARDCLKL;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_CLKARDCLKU;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_CLKBWRCLKL;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_CLKBWRCLKU;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIADI0;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIADI1;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIADI10;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIADI11;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIADI12;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIADI13;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIADI14;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIADI15;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIADI16;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIADI17;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIADI18;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIADI19;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIADI2;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIADI20;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIADI21;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIADI22;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIADI23;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIADI24;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIADI25;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIADI26;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIADI27;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIADI28;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIADI29;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIADI3;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIADI30;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIADI31;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIADI4;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIADI5;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIADI6;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIADI7;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIADI8;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIADI9;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI0;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI1;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI10;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI11;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI12;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI13;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI14;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI15;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI16;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI17;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI18;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI19;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI2;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI20;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI21;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI22;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI23;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI24;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI25;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI26;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI27;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI28;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI29;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI3;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI30;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI31;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI4;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI5;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI6;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI7;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI8;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI9;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIPADIP0;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIPADIP1;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIPADIP2;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIPADIP3;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIPBDIP0;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIPBDIP1;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIPBDIP2;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DIPBDIP3;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOADO0;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOADO1;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOADO10;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOADO11;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOADO12;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOADO13;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOADO14;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOADO15;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOADO16;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOADO17;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOADO18;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOADO19;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOADO2;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOADO20;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOADO21;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOADO22;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOADO23;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOADO24;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOADO25;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOADO26;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOADO27;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOADO28;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOADO29;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOADO3;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOADO30;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOADO31;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOADO4;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOADO5;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOADO6;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOADO7;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOADO8;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOADO9;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO0;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO1;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO10;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO11;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO12;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO13;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO14;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO15;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO16;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO17;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO18;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO19;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO2;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO20;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO21;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO22;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO23;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO24;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO25;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO26;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO27;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO28;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO29;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO3;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO30;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO31;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO4;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO5;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO6;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO7;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO8;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO9;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOPADOP0;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOPADOP1;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOPADOP2;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOPADOP3;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOPBDOP0;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOPBDOP1;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOPBDOP2;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_DOPBDOP3;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ENARDENL;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ENARDENU;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ENBWRENL;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_ENBWRENU;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_REGCEAREGCEL;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_REGCEAREGCEU;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_REGCEBL;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_REGCEBU;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_REGCLKARDRCLKL;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_REGCLKARDRCLKU;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_REGCLKBL;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_REGCLKBU;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_RSTRAMARSTRAMLRST;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_RSTRAMARSTRAMU;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_RSTRAMBL;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_RSTRAMBU;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_RSTREGARSTREGL;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_RSTREGARSTREGU;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_RSTREGBL;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_RSTREGBU;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_WEAL0;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_WEAL1;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_WEAL2;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_WEAL3;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_WEAU0;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_WEAU1;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_WEAU2;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_WEAU3;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_WEBWEL0;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_WEBWEL1;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_WEBWEL2;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_WEBWEL3;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_WEBWEL4;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_WEBWEL5;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_WEBWEL6;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_WEBWEL7;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_WEBWEU0;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_WEBWEU1;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_WEBWEU2;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_WEBWEU3;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_WEBWEU4;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_WEBWEU5;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_WEBWEU6;
  wire [0:0] BRAM_L_X6Y90_RAMB36_X0Y18_WEBWEU7;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRL0;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRL1;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRL10;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRL11;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRL12;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRL13;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRL14;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRL15;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRL2;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRL3;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRL4;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRL5;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRL6;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRL7;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRL8;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRL9;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRU0;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRU1;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRU10;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRU11;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRU12;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRU13;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRU14;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRU2;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRU3;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRU4;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRU5;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRU6;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRU7;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRU8;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRU9;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRL0;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRL1;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRL10;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRL11;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRL12;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRL13;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRL14;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRL15;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRL2;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRL3;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRL4;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRL5;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRL6;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRL7;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRL8;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRL9;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRU0;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRU1;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRU10;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRU11;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRU12;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRU13;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRU14;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRU2;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRU3;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRU4;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRU5;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRU6;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRU7;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRU8;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRU9;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_CLKARDCLKL;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_CLKARDCLKU;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_CLKBWRCLKL;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_CLKBWRCLKU;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIADI0;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIADI1;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIADI10;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIADI11;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIADI12;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIADI13;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIADI14;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIADI15;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIADI16;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIADI17;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIADI18;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIADI19;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIADI2;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIADI20;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIADI21;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIADI22;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIADI23;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIADI24;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIADI25;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIADI26;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIADI27;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIADI28;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIADI29;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIADI3;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIADI30;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIADI31;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIADI4;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIADI5;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIADI6;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIADI7;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIADI8;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIADI9;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI0;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI1;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI10;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI11;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI12;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI13;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI14;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI15;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI16;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI17;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI18;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI19;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI2;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI20;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI21;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI22;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI23;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI24;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI25;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI26;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI27;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI28;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI29;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI3;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI30;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI31;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI4;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI5;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI6;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI7;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI8;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI9;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIPADIP0;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIPADIP1;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIPADIP2;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIPADIP3;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIPBDIP0;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIPBDIP1;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIPBDIP2;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DIPBDIP3;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOADO0;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOADO1;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOADO10;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOADO11;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOADO12;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOADO13;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOADO14;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOADO15;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOADO16;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOADO17;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOADO18;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOADO19;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOADO2;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOADO20;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOADO21;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOADO22;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOADO23;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOADO24;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOADO25;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOADO26;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOADO27;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOADO28;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOADO29;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOADO3;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOADO30;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOADO31;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOADO4;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOADO5;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOADO6;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOADO7;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOADO8;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOADO9;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO0;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO1;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO10;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO11;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO12;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO13;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO14;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO15;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO16;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO17;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO18;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO19;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO2;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO20;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO21;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO22;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO23;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO24;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO25;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO26;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO27;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO28;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO29;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO3;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO30;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO31;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO4;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO5;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO6;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO7;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO8;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO9;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOPADOP0;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOPADOP1;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOPADOP2;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOPADOP3;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOPBDOP0;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOPBDOP1;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOPBDOP2;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_DOPBDOP3;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ENARDENL;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ENARDENU;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ENBWRENL;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_ENBWRENU;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_REGCEAREGCEL;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_REGCEAREGCEU;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_REGCEBL;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_REGCEBU;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_REGCLKARDRCLKL;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_REGCLKARDRCLKU;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_REGCLKBL;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_REGCLKBU;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_RSTRAMARSTRAMLRST;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_RSTRAMARSTRAMU;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_RSTRAMBL;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_RSTRAMBU;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_RSTREGARSTREGL;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_RSTREGARSTREGU;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_RSTREGBL;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_RSTREGBU;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_WEAL0;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_WEAL1;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_WEAL2;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_WEAL3;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_WEAU0;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_WEAU1;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_WEAU2;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_WEAU3;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_WEBWEL0;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_WEBWEL1;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_WEBWEL2;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_WEBWEL3;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_WEBWEL4;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_WEBWEL5;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_WEBWEL6;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_WEBWEL7;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_WEBWEU0;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_WEBWEU1;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_WEBWEU2;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_WEBWEU3;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_WEBWEU4;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_WEBWEU5;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_WEBWEU6;
  wire [0:0] BRAM_L_X6Y95_RAMB36_X0Y19_WEBWEU7;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_A;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_A1;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_A2;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_A3;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_A4;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_A5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_A6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_AO5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_AO6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_AQ;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_AX;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_A_CY;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_A_XOR;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_B;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_B1;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_B2;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_B3;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_B4;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_B5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_B6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_BO5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_BO6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_B_CY;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_B_XOR;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_C;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_C1;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_C2;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_C3;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_C4;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_C5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_C6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_CLK;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_CO5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_CO6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_C_CY;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_C_XOR;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_D;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_D1;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_D2;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_D3;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_D4;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_D5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_D6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_DO5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_DO6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_D_CY;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_D_XOR;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_SR;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_A;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_A1;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_A2;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_A3;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_A4;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_A5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_A6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_AO5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_AO6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_A_CY;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_A_XOR;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_B;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_B1;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_B2;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_B3;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_B4;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_B5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_B6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_BO5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_BO6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_B_CY;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_B_XOR;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_C;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_C1;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_C2;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_C3;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_C4;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_C5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_C6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_CO5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_CO6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_C_CY;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_C_XOR;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_D;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_D1;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_D2;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_D3;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_D4;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_D5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_D6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_DO5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_DO6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_D_CY;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_D_XOR;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_A;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_A1;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_A2;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_A3;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_A4;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_A5;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_A6;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_AO5;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_AO6;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_A_CY;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_A_XOR;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_B;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_B1;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_B2;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_B3;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_B4;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_B5;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_B6;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_BO5;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_BO6;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_B_CY;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_B_XOR;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_C;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_C1;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_C2;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_C3;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_C4;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_C5;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_C6;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_CO5;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_CO6;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_C_CY;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_C_XOR;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_D;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_D1;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_D2;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_D3;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_D4;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_D5;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_D6;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_DO5;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_DO6;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_D_CY;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X0Y90_D_XOR;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_A;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_A1;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_A2;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_A3;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_A4;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_A5;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_A6;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_AO5;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_AO6;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_AQ;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_AX;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_A_CY;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_A_XOR;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_B;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_B1;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_B2;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_B3;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_B4;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_B5;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_B6;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_BO5;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_BO6;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_B_CY;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_B_XOR;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_C;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_C1;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_C2;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_C3;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_C4;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_C5;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_C6;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_CE;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_CLK;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_CO5;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_CO6;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_C_CY;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_C_XOR;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_D;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_D1;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_D2;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_D3;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_D4;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_D5;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_D6;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_DO5;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_DO6;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_D_CY;
  wire [0:0] CLBLL_L_X2Y90_SLICE_X1Y90_D_XOR;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_A;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_A1;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_A2;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_A3;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_A4;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_A5;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_A6;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_AO5;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_AO6;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_AQ;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_AX;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_A_CY;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_A_XOR;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_B;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_B1;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_B2;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_B3;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_B4;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_B5;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_B6;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_BO5;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_BO6;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_B_CY;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_B_XOR;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_C;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_C1;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_C2;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_C3;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_C4;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_C5;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_C6;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_CE;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_CLK;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_CO5;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_CO6;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_C_CY;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_C_XOR;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_D;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_D1;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_D2;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_D3;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_D4;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_D5;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_D6;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_DO5;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_DO6;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_D_CY;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X0Y91_D_XOR;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_A;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_A1;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_A2;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_A3;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_A4;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_A5;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_A6;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_AO5;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_AO6;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_AQ;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_AX;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_A_CY;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_A_XOR;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_B;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_B1;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_B2;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_B3;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_B4;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_B5;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_B6;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_BO5;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_BO6;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_BQ;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_BX;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_B_CY;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_B_XOR;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_C;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_C1;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_C2;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_C3;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_C4;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_C5;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_C6;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_CE;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_CLK;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_CO5;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_CO6;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_CQ;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_CX;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_C_CY;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_C_XOR;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_D;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_D1;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_D2;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_D3;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_D4;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_D5;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_D6;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_DO5;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_DO6;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_D_CY;
  wire [0:0] CLBLL_L_X2Y91_SLICE_X1Y91_D_XOR;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_A;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_A1;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_A2;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_A3;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_A4;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_A5;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_A6;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_AO5;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_AO6;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_AQ;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_AX;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_A_CY;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_A_XOR;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_B;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_B1;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_B2;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_B3;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_B4;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_B5;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_B6;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_BO5;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_BO6;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_B_CY;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_B_XOR;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_C;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_C1;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_C2;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_C3;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_C4;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_C5;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_C6;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_CE;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_CLK;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_CO5;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_CO6;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_C_CY;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_C_XOR;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_D;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_D1;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_D2;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_D3;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_D4;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_D5;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_D6;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_DO5;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_DO6;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_D_CY;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X0Y92_D_XOR;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_A;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_A1;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_A2;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_A3;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_A4;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_A5;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_A6;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_AO5;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_AO6;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_AQ;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_AX;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_A_CY;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_A_XOR;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_B;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_B1;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_B2;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_B3;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_B4;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_B5;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_B6;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_BO5;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_BO6;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_BQ;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_BX;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_B_CY;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_B_XOR;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_C;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_C1;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_C2;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_C3;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_C4;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_C5;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_C6;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_CE;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_CLK;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_CO5;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_CO6;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_CQ;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_CX;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_C_CY;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_C_XOR;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_D;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_D1;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_D2;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_D3;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_D4;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_D5;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_D6;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_DO5;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_DO6;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_D_CY;
  wire [0:0] CLBLL_L_X2Y92_SLICE_X1Y92_D_XOR;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_A;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_A1;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_A2;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_A3;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_A4;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_A5;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_A6;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_AMUX;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_AO5;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_AO6;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_AX;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_A_CY;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_A_XOR;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_B;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_B1;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_B2;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_B3;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_B4;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_B5;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_B6;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_BO5;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_BO6;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_BQ;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_BX;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_B_CY;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_B_XOR;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_C;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_C1;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_C2;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_C3;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_C4;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_C5;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_C6;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_CE;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_CLK;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_CMUX;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_CO5;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_CO6;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_CQ;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_CX;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_C_CY;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_C_XOR;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_D;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_D1;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_D2;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_D3;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_D4;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_D5;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_D6;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_DMUX;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_DO5;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_DO6;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_D_CY;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_D_XOR;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X0Y93_F7AMUX_O;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_A;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_A1;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_A2;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_A3;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_A4;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_A5;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_A6;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_AMUX;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_AO5;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_AO6;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_AX;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_A_CY;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_A_XOR;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_B;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_B1;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_B2;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_B3;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_B4;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_B5;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_B6;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_BO5;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_BO6;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_BQ;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_BX;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_B_CY;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_B_XOR;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_C;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_C1;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_C2;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_C3;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_C4;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_C5;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_C6;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_CE;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_CLK;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_CO5;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_CO6;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_C_CY;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_C_XOR;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_D;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_D1;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_D2;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_D3;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_D4;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_D5;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_D6;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_DMUX;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_DO5;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_DO6;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_D_CY;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_D_XOR;
  wire [0:0] CLBLL_L_X2Y93_SLICE_X1Y93_F7AMUX_O;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_A;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_A1;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_A2;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_A3;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_A4;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_A5;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_A6;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_AO5;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_AO6;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_A_CY;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_A_XOR;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_B;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_B1;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_B2;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_B3;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_B4;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_B5;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_B6;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_BO5;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_BO6;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_B_CY;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_B_XOR;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_C;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_C1;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_C2;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_C3;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_C4;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_C5;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_C6;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_CMUX;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_CO5;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_CO6;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_C_CY;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_C_XOR;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_D;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_D1;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_D2;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_D3;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_D4;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_D5;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_D6;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_DMUX;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_DO5;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_DO6;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_D_CY;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X0Y94_D_XOR;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_A;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_A1;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_A2;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_A3;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_A4;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_A5;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_A6;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_AMUX;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_AO5;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_AO6;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_AX;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_A_CY;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_A_XOR;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_B;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_B1;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_B2;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_B3;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_B4;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_B5;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_B6;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_BMUX;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_BO5;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_BO6;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_BQ;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_BX;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_B_CY;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_B_XOR;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_C;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_C1;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_C2;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_C3;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_C4;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_C5;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_C6;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_CE;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_CLK;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_CMUX;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_CO5;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_CO6;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_COUT;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_CQ;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_CX;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_C_CY;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_C_XOR;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_D;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_D1;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_D2;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_D3;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_D4;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_D5;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_D6;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_DMUX;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_DO5;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_DO6;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_DQ;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_DX;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_D_CY;
  wire [0:0] CLBLL_L_X2Y94_SLICE_X1Y94_D_XOR;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_A;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_A1;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_A2;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_A3;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_A4;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_A5;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_A6;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_AO5;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_AO6;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_A_CY;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_A_XOR;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_B;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_B1;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_B2;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_B3;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_B4;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_B5;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_B6;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_BO5;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_BO6;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_B_CY;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_B_XOR;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_C;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_C1;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_C2;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_C3;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_C4;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_C5;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_C6;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_CO5;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_CO6;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_COUT;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_C_CY;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_C_XOR;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_D;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_D1;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_D2;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_D3;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_D4;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_D5;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_D6;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_DMUX;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_DO5;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_DO6;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_D_CY;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X0Y95_D_XOR;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_A;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_A1;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_A2;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_A3;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_A4;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_A5;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_A6;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_AMUX;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_AO5;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_AO6;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_AX;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_A_CY;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_A_XOR;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_B;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_B1;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_B2;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_B3;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_B4;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_B5;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_B6;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_BMUX;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_BO5;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_BO6;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_BX;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_B_CY;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_B_XOR;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_C;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_C1;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_C2;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_C3;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_C4;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_C5;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_C6;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_CIN;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_CMUX;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_CO5;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_CO6;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_COUT;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_CX;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_C_CY;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_C_XOR;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_D;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_D1;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_D2;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_D3;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_D4;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_D5;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_D6;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_DMUX;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_DO5;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_DO6;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_DX;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_D_CY;
  wire [0:0] CLBLL_L_X2Y95_SLICE_X1Y95_D_XOR;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_A;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_A1;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_A2;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_A3;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_A4;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_A5;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_A6;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_AO5;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_AO6;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_A_CY;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_A_XOR;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_B;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_B1;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_B2;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_B3;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_B4;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_B5;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_B6;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_BMUX;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_BO5;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_BO6;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_B_CY;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_B_XOR;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_C;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_C1;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_C2;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_C3;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_C4;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_C5;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_C6;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_CO5;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_CO6;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_C_CY;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_C_XOR;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_D;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_D1;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_D2;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_D3;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_D4;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_D5;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_D6;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_DO5;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_DO6;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_D_CY;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X0Y96_D_XOR;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_A;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_A1;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_A2;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_A3;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_A4;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_A5;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_A6;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_AMUX;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_AO5;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_AO6;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_A_CY;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_A_XOR;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_B;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_B1;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_B2;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_B3;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_B4;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_B5;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_B6;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_BO5;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_BO6;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_B_CY;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_B_XOR;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_C;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_C1;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_C2;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_C3;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_C4;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_C5;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_C6;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_CO5;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_CO6;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_C_CY;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_C_XOR;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_D;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_D1;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_D2;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_D3;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_D4;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_D5;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_D6;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_DMUX;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_DO5;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_DO6;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_D_CY;
  wire [0:0] CLBLL_L_X2Y96_SLICE_X1Y96_D_XOR;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_A;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_A1;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_A2;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_A3;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_A4;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_A5;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_A6;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_AMUX;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_AO5;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_AO6;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_A_CY;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_A_XOR;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_B;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_B1;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_B2;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_B3;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_B4;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_B5;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_B6;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_BO5;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_BO6;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_B_CY;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_B_XOR;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_C;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_C1;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_C2;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_C3;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_C4;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_C5;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_C6;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_CO5;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_CO6;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_C_CY;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_C_XOR;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_D;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_D1;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_D2;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_D3;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_D4;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_D5;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_D6;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_DMUX;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_DO5;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_DO6;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_D_CY;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X0Y97_D_XOR;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_A;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_A1;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_A2;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_A3;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_A4;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_A5;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_A6;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_AO5;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_AO6;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_A_CY;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_A_XOR;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_B;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_B1;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_B2;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_B3;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_B4;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_B5;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_B6;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_BO5;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_BO6;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_B_CY;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_B_XOR;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_C;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_C1;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_C2;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_C3;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_C4;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_C5;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_C6;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_CO5;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_CO6;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_C_CY;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_C_XOR;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_D;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_D1;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_D2;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_D3;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_D4;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_D5;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_D6;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_DO5;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_DO6;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_D_CY;
  wire [0:0] CLBLL_L_X2Y97_SLICE_X1Y97_D_XOR;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_A;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_A1;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_A2;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_A3;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_A4;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_A5;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_A6;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_AO5;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_AO6;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_AQ;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_AX;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_A_CY;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_A_XOR;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_B;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_B1;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_B2;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_B3;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_B4;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_B5;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_B6;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_BO5;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_BO6;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_B_CY;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_B_XOR;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_C;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_C1;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_C2;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_C3;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_C4;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_C5;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_C6;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_CE;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_CLK;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_CO5;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_CO6;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_C_CY;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_C_XOR;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_D;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_D1;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_D2;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_D3;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_D4;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_D5;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_D6;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_DO5;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_DO6;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_D_CY;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_D_XOR;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_SR;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_A;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_A1;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_A2;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_A3;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_A4;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_A5;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_A6;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_AO5;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_AO6;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_AQ;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_A_CY;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_A_XOR;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_B;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_B1;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_B2;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_B3;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_B4;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_B5;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_B6;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_BO5;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_BO6;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_B_CY;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_B_XOR;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_C;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_C1;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_C2;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_C3;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_C4;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_C5;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_C6;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_CLK;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_CO5;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_CO6;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_C_CY;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_C_XOR;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_D;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_D1;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_D2;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_D3;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_D4;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_D5;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_D6;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_DO5;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_DO6;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_D_CY;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_D_XOR;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_SR;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_A;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_A1;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_A2;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_A3;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_A4;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_A5;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_A6;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_AO5;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_AO6;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_AQ;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_AX;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_A_CY;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_A_XOR;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_B;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_B1;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_B2;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_B3;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_B4;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_B5;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_B6;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_BO5;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_BO6;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_B_CY;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_B_XOR;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_C;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_C1;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_C2;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_C3;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_C4;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_C5;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_C6;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_CE;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_CLK;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_CO5;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_CO6;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_C_CY;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_C_XOR;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_D;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_D1;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_D2;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_D3;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_D4;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_D5;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_D6;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_DO5;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_DO6;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_D_CY;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_D_XOR;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X0Y99_SR;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_A;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_A1;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_A2;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_A3;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_A4;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_A5;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_A6;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_AO5;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_AO6;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_AQ;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_AX;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_A_CY;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_A_XOR;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_B;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_B1;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_B2;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_B3;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_B4;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_B5;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_B6;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_BO5;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_BO6;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_B_CY;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_B_XOR;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_C;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_C1;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_C2;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_C3;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_C4;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_C5;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_C6;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_CE;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_CLK;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_CO5;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_CO6;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_C_CY;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_C_XOR;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_D;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_D1;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_D2;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_D3;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_D4;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_D5;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_D6;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_DO5;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_DO6;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_D_CY;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_D_XOR;
  wire [0:0] CLBLL_L_X2Y99_SLICE_X1Y99_SR;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_A;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_A1;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_A2;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_A3;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_A4;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_A5;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_A6;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_AO5;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_AO6;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_A_CY;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_A_XOR;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_B;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_B1;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_B2;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_B3;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_B4;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_B5;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_B6;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_BO5;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_BO6;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_B_CY;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_B_XOR;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_C;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_C1;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_C2;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_C3;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_C4;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_C5;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_C6;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_CO5;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_CO6;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_C_CY;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_C_XOR;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_D;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_D1;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_D2;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_D3;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_D4;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_D5;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_D6;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_DO5;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_DO6;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_D_CY;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X4Y90_D_XOR;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_A;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_A1;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_A2;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_A3;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_A4;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_A5;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_A6;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_AO5;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_AO6;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_AQ;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_AX;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_A_CY;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_A_XOR;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_B;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_B1;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_B2;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_B3;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_B4;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_B5;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_B6;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_BO5;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_BO6;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_B_CY;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_B_XOR;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_C;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_C1;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_C2;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_C3;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_C4;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_C5;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_C6;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_CLK;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_CO5;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_CO6;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_C_CY;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_C_XOR;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_D;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_D1;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_D2;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_D3;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_D4;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_D5;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_D6;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_DO5;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_DO6;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_D_CY;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_D_XOR;
  wire [0:0] CLBLL_L_X4Y90_SLICE_X5Y90_SR;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_A;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_A1;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_A2;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_A3;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_A4;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_A5;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_A6;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_AMUX;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_AO5;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_AO6;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_AQ;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_AX;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_A_CY;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_A_XOR;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_B;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_B1;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_B2;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_B3;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_B4;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_B5;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_B6;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_BO5;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_BO6;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_BQ;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_BX;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_B_CY;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_B_XOR;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_C;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_C1;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_C2;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_C3;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_C4;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_C5;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_C6;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_CE;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_CLK;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_CO5;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_CO6;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_C_CY;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_C_XOR;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_D;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_D1;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_D2;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_D3;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_D4;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_D5;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_D6;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_DO5;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_DO6;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_D_CY;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X4Y91_D_XOR;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_A;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_A1;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_A2;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_A3;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_A4;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_A5;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_A6;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_AMUX;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_AO5;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_AO6;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_AX;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_A_CY;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_A_XOR;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_B;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_B1;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_B2;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_B3;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_B4;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_B5;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_B6;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_BO5;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_BO6;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_BQ;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_BX;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_B_CY;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_B_XOR;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_C;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_C1;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_C2;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_C3;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_C4;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_C5;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_C6;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_CE;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_CLK;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_CO5;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_CO6;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_C_CY;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_C_XOR;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_D;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_D1;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_D2;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_D3;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_D4;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_D5;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_D6;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_DO5;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_DO6;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_D_CY;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_D_XOR;
  wire [0:0] CLBLL_L_X4Y91_SLICE_X5Y91_F7AMUX_O;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_A;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_A1;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_A2;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_A3;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_A4;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_A5;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_A6;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_AMUX;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_AO5;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_AO6;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_AQ;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_AX;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_A_CY;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_A_XOR;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_B;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_B1;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_B2;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_B3;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_B4;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_B5;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_B5Q;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_B6;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_BMUX;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_BO5;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_BO6;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_BQ;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_BX;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_B_CY;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_B_XOR;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_C;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_C1;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_C2;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_C3;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_C4;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_C5;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_C6;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_CE;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_CLK;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_CO5;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_CO6;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_CQ;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_CX;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_C_CY;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_C_XOR;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_D;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_D1;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_D2;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_D3;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_D4;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_D5;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_D6;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_DO5;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_DO6;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_DQ;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_DX;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_D_CY;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X4Y92_D_XOR;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_A;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_A1;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_A2;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_A3;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_A4;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_A5;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_A6;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_AMUX;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_AO5;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_AO6;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_AX;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_A_CY;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_A_XOR;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_B;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_B1;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_B2;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_B3;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_B4;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_B5;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_B6;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_BO5;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_BO6;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_BQ;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_BX;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_B_CY;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_B_XOR;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_C;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_C1;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_C2;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_C3;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_C4;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_C5;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_C6;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_CE;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_CLK;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_CO5;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_CO6;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_CQ;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_CX;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_C_CY;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_C_XOR;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_D;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_D1;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_D2;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_D3;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_D4;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_D5;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_D6;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_DO5;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_DO6;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_D_CY;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_D_XOR;
  wire [0:0] CLBLL_L_X4Y92_SLICE_X5Y92_F7AMUX_O;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_A;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_A1;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_A2;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_A3;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_A4;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_A5;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_A6;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_AMUX;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_AO5;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_AO6;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_AX;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_A_CY;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_A_XOR;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_B;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_B1;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_B2;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_B3;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_B4;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_B5;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_B6;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_BO5;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_BO6;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_BQ;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_BX;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_B_CY;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_B_XOR;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_C;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_C1;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_C2;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_C3;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_C4;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_C5;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_C6;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_CE;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_CLK;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_CMUX;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_CO5;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_CO6;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_CQ;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_C_CY;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_C_XOR;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_D;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_D1;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_D2;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_D3;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_D4;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_D5;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_D6;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_DO5;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_DO6;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_DQ;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_DX;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_D_CY;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_D_XOR;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X4Y93_F7AMUX_O;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_A;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_A1;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_A2;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_A3;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_A4;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_A5;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_A6;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_AMUX;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_AO5;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_AO6;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_AX;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_A_CY;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_A_XOR;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_B;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_B1;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_B2;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_B3;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_B4;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_B5;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_B6;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_BO5;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_BO6;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_BQ;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_BX;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_B_CY;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_B_XOR;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_C;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_C1;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_C2;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_C3;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_C4;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_C5;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_C6;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_CE;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_CLK;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_CO5;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_CO6;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_CQ;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_CX;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_C_CY;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_C_XOR;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_D;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_D1;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_D2;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_D3;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_D4;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_D5;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_D6;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_DO5;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_DO6;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_DQ;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_DX;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_D_CY;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_D_XOR;
  wire [0:0] CLBLL_L_X4Y93_SLICE_X5Y93_F7AMUX_O;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_A;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_A1;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_A2;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_A3;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_A4;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_A5;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_A6;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_AO5;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_AO6;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_AQ;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_A_CY;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_A_XOR;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_B;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_B1;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_B2;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_B3;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_B4;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_B5;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_B6;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_BO5;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_BO6;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_BQ;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_B_CY;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_B_XOR;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_C;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_C1;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_C2;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_C3;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_C4;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_C5;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_C6;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_CLK;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_CMUX;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_CO5;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_CO6;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_C_CY;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_C_XOR;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_D;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_D1;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_D2;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_D3;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_D4;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_D5;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_D6;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_DO5;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_DO6;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_D_CY;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_D_XOR;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X4Y94_SR;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_A;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_A1;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_A2;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_A3;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_A4;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_A5;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_A6;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_AMUX;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_AO5;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_AO6;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_AX;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_A_CY;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_A_XOR;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_B;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_B1;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_B2;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_B3;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_B4;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_B5;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_B6;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_BO5;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_BO6;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_BQ;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_BX;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_B_CY;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_B_XOR;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_C;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_C1;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_C2;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_C3;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_C4;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_C5;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_C6;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_CE;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_CLK;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_CO5;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_CO6;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_CQ;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_CX;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_C_CY;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_C_XOR;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_D;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_D1;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_D2;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_D3;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_D4;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_D5;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_D6;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_DO5;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_DO6;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_DQ;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_DX;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_D_CY;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_D_XOR;
  wire [0:0] CLBLL_L_X4Y94_SLICE_X5Y94_F7AMUX_O;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_A;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_A1;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_A2;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_A3;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_A4;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_A5;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_A6;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_AO5;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_AO6;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_AQ;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_AX;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_A_CY;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_A_XOR;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_B;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_B1;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_B2;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_B3;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_B4;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_B5;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_B6;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_BO5;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_BO6;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_B_CY;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_B_XOR;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_C;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_C1;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_C2;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_C3;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_C4;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_C5;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_C6;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_CE;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_CLK;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_CO5;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_CO6;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_C_CY;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_C_XOR;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_D;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_D1;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_D2;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_D3;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_D4;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_D5;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_D6;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_DO5;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_DO6;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_D_CY;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X4Y95_D_XOR;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_A;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_A1;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_A2;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_A3;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_A4;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_A5;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_A6;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_AMUX;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_AO5;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_AO6;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_AX;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_A_CY;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_A_XOR;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_B;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_B1;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_B2;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_B3;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_B4;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_B5;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_B6;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_BO5;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_BO6;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_B_CY;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_B_XOR;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_C;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_C1;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_C2;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_C3;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_C4;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_C5;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_C6;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_CO5;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_CO6;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_C_CY;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_C_XOR;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_D;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_D1;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_D2;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_D3;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_D4;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_D5;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_D6;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_DO5;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_DO6;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_D_CY;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_D_XOR;
  wire [0:0] CLBLL_L_X4Y95_SLICE_X5Y95_F7AMUX_O;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_A;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_A1;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_A2;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_A3;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_A4;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_A5;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_A6;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_AO5;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_AO6;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_A_CY;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_A_XOR;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_B;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_B1;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_B2;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_B3;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_B4;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_B5;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_B6;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_BO5;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_BO6;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_B_CY;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_B_XOR;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_C;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_C1;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_C2;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_C3;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_C4;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_C5;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_C6;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_CO5;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_CO6;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_C_CY;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_C_XOR;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_D;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_D1;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_D2;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_D3;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_D4;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_D5;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_D6;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_DO5;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_DO6;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_D_CY;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X4Y96_D_XOR;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_A;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_A1;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_A2;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_A3;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_A4;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_A5;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_A6;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_AO5;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_AO6;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_A_CY;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_A_XOR;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_B;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_B1;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_B2;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_B3;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_B4;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_B5;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_B6;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_BO5;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_BO6;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_B_CY;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_B_XOR;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_C;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_C1;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_C2;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_C3;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_C4;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_C5;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_C6;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_CO5;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_CO6;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_C_CY;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_C_XOR;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_D;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_D1;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_D2;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_D3;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_D4;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_D5;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_D6;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_DO5;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_DO6;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_D_CY;
  wire [0:0] CLBLL_L_X4Y96_SLICE_X5Y96_D_XOR;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_A;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_A1;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_A2;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_A3;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_A4;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_A5;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_A6;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_AMUX;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_AO5;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_AO6;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_A_CY;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_A_XOR;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_B;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_B1;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_B2;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_B3;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_B4;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_B5;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_B6;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_BO5;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_BO6;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_BQ;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_B_CY;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_B_XOR;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_C;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_C1;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_C2;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_C3;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_C4;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_C5;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_C6;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_CLK;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_CO5;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_CO6;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_C_CY;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_C_XOR;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_D;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_D1;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_D2;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_D3;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_D4;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_D5;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_D6;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_DO5;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_DO6;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_D_CY;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_D_XOR;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X4Y97_SR;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_A;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_A1;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_A2;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_A3;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_A4;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_A5;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_A6;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_AMUX;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_AO5;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_AO6;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_A_CY;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_A_XOR;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_B;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_B1;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_B2;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_B3;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_B4;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_B5;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_B6;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_BO5;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_BO6;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_B_CY;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_B_XOR;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_C;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_C1;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_C2;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_C3;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_C4;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_C5;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_C6;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_CO5;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_CO6;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_C_CY;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_C_XOR;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_D;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_D1;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_D2;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_D3;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_D4;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_D5;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_D6;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_DO5;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_DO6;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_D_CY;
  wire [0:0] CLBLL_L_X4Y97_SLICE_X5Y97_D_XOR;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_A;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_A1;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_A2;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_A3;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_A4;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_A5;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_A6;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_AMUX;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_AO5;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_AO6;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_A_CY;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_A_XOR;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_B;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_B1;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_B2;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_B3;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_B4;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_B5;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_B6;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_BO5;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_BO6;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_B_CY;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_B_XOR;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_C;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_C1;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_C2;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_C3;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_C4;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_C5;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_C6;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_CO5;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_CO6;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_C_CY;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_C_XOR;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_D;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_D1;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_D2;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_D3;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_D4;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_D5;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_D6;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_DO5;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_DO6;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_D_CY;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X4Y98_D_XOR;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_A;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_A1;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_A2;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_A3;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_A4;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_A5;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_A6;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_AO5;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_AO6;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_A_CY;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_A_XOR;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_B;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_B1;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_B2;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_B3;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_B4;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_B5;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_B6;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_BO5;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_BO6;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_B_CY;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_B_XOR;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_C;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_C1;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_C2;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_C3;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_C4;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_C5;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_C6;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_CO5;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_CO6;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_C_CY;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_C_XOR;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_D;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_D1;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_D2;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_D3;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_D4;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_D5;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_D6;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_DO5;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_DO6;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_D_CY;
  wire [0:0] CLBLL_L_X4Y98_SLICE_X5Y98_D_XOR;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_A;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_A1;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_A2;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_A3;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_A4;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_A5;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_A5Q;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_A6;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_AMUX;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_AO5;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_AO6;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_AQ;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_A_CY;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_A_XOR;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_B;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_B1;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_B2;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_B3;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_B4;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_B5;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_B6;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_BO5;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_BO6;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_BQ;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_B_CY;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_B_XOR;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_C;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_C1;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_C2;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_C3;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_C4;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_C5;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_C6;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_CE;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_CLK;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_CO5;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_CO6;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_CQ;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_C_CY;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_C_XOR;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_D;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_D1;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_D2;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_D3;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_D4;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_D5;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_D6;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_DO5;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_DO6;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_D_CY;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_D_XOR;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X10Y89_SR;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_A;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_A1;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_A2;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_A3;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_A4;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_A5;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_A6;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_AO5;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_AO6;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_A_CY;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_A_XOR;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_B;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_B1;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_B2;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_B3;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_B4;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_B5;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_B6;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_BO5;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_BO6;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_B_CY;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_B_XOR;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_C;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_C1;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_C2;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_C3;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_C4;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_C5;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_C6;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_CO5;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_CO6;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_C_CY;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_C_XOR;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_D;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_D1;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_D2;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_D3;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_D4;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_D5;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_D6;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_DO5;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_DO6;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_D_CY;
  wire [0:0] CLBLM_L_X8Y89_SLICE_X11Y89_D_XOR;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X10Y97_A;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X10Y97_A1;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X10Y97_A2;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X10Y97_A3;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X10Y97_A4;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X10Y97_A5;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X10Y97_A6;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X10Y97_AO5;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X10Y97_AO6;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X10Y97_AX;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X10Y97_B;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X10Y97_B1;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X10Y97_B2;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X10Y97_B3;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X10Y97_B4;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X10Y97_B5;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X10Y97_B6;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X10Y97_BO5;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X10Y97_BO6;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X10Y97_BX;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X10Y97_C;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X10Y97_C1;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X10Y97_C2;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X10Y97_C3;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X10Y97_C4;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X10Y97_C5;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X10Y97_C6;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X10Y97_CE;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X10Y97_CLK;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X10Y97_CO5;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X10Y97_CO6;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X10Y97_D;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X10Y97_D1;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X10Y97_D2;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X10Y97_D3;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X10Y97_D4;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X10Y97_D5;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X10Y97_DI;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X10Y97_DO5;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X10Y97_DO6;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X10Y97_DX;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_A;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_A1;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_A2;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_A3;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_A4;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_A5;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_A6;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_AO5;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_AO6;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_AQ;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_AX;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_A_CY;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_A_XOR;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_B;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_B1;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_B2;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_B3;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_B4;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_B5;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_B6;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_BO5;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_BO6;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_B_CY;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_B_XOR;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_C;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_C1;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_C2;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_C3;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_C4;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_C5;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_C6;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_CLK;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_CO5;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_CO6;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_C_CY;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_C_XOR;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_D;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_D1;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_D2;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_D3;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_D4;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_D5;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_D6;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_DO5;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_DO6;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_D_CY;
  wire [0:0] CLBLM_L_X8Y97_SLICE_X11Y97_D_XOR;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_A;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_A1;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_A2;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_A3;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_A4;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_A5;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_A6;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_AMUX;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_AO5;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_AO6;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_A_CY;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_A_XOR;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_B;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_B1;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_B2;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_B3;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_B4;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_B5;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_B6;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_BO5;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_BO6;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_B_CY;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_B_XOR;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_C;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_C1;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_C2;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_C3;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_C4;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_C5;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_C6;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_CO5;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_CO6;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_C_CY;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_C_XOR;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_D;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_D1;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_D2;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_D3;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_D4;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_D5;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_D6;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_DO5;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_DO6;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_D_CY;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X10Y98_D_XOR;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_A;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_A1;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_A2;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_A3;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_A4;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_A5;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_A6;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_AO5;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_AO6;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_A_CY;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_A_XOR;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_B;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_B1;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_B2;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_B3;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_B4;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_B5;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_B6;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_BO5;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_BO6;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_B_CY;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_B_XOR;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_C;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_C1;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_C2;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_C3;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_C4;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_C5;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_C6;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_CO5;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_CO6;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_C_CY;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_C_XOR;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_D;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_D1;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_D2;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_D3;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_D4;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_D5;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_D6;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_DO5;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_DO6;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_D_CY;
  wire [0:0] CLBLM_L_X8Y98_SLICE_X11Y98_D_XOR;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_A;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_A1;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_A2;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_A3;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_A4;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_A5;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_A6;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_AO5;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_AO6;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_AQ;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_AX;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_A_CY;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_A_XOR;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_B;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_B1;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_B2;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_B3;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_B4;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_B5;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_B6;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_BO5;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_BO6;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_B_CY;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_B_XOR;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_C;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_C1;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_C2;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_C3;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_C4;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_C5;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_C6;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_CE;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_CLK;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_CO5;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_CO6;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_C_CY;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_C_XOR;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_D;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_D1;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_D2;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_D3;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_D4;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_D5;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_D6;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_DO5;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_DO6;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_D_CY;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X2Y90_D_XOR;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_A;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_A1;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_A2;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_A3;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_A4;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_A5;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_A6;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_AO5;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_AO6;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_AQ;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_AX;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_A_CY;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_A_XOR;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_B;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_B1;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_B2;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_B3;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_B4;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_B5;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_B6;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_BO5;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_BO6;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_B_CY;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_B_XOR;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_C;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_C1;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_C2;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_C3;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_C4;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_C5;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_C6;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_CE;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_CLK;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_CO5;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_CO6;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_C_CY;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_C_XOR;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_D;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_D1;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_D2;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_D3;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_D4;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_D5;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_D6;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_DO5;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_DO6;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_D_CY;
  wire [0:0] CLBLM_R_X3Y90_SLICE_X3Y90_D_XOR;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_A;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_A1;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_A2;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_A3;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_A4;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_A5;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_A6;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_AMUX;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_AO5;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_AO6;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_AX;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_A_CY;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_A_XOR;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_B;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_B1;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_B2;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_B3;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_B4;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_B5;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_B6;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_BO5;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_BO6;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_BQ;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_BX;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_B_CY;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_B_XOR;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_C;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_C1;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_C2;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_C3;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_C4;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_C5;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_C6;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_CE;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_CLK;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_CMUX;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_CO5;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_CO6;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_CX;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_C_CY;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_C_XOR;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_D;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_D1;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_D2;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_D3;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_D4;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_D5;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_D6;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_DO5;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_DO6;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_DQ;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_DX;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_D_CY;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_D_XOR;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_F7AMUX_O;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X2Y91_F7BMUX_O;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_A;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_A1;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_A2;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_A3;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_A4;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_A5;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_A6;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_AMUX;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_AO5;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_AO6;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_AX;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_A_CY;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_A_XOR;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_B;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_B1;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_B2;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_B3;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_B4;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_B5;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_B6;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_BO5;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_BO6;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_BQ;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_BX;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_B_CY;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_B_XOR;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_C;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_C1;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_C2;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_C3;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_C4;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_C5;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_C6;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_CE;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_CLK;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_CMUX;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_CO5;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_CO6;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_CX;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_C_CY;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_C_XOR;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_D;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_D1;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_D2;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_D3;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_D4;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_D5;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_D6;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_DO5;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_DO6;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_DQ;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_DX;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_D_CY;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_D_XOR;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_F7AMUX_O;
  wire [0:0] CLBLM_R_X3Y91_SLICE_X3Y91_F7BMUX_O;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_A;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_A1;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_A2;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_A3;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_A4;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_A5;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_A6;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_AMUX;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_AO5;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_AO6;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_AX;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_A_CY;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_A_XOR;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_B;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_B1;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_B2;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_B3;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_B4;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_B5;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_B6;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_BO5;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_BO6;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_BQ;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_BX;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_B_CY;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_B_XOR;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_C;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_C1;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_C2;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_C3;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_C4;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_C5;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_C6;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_CE;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_CLK;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_CMUX;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_CO5;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_CO6;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_CX;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_C_CY;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_C_XOR;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_D;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_D1;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_D2;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_D3;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_D4;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_D5;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_D6;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_DO5;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_DO6;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_DQ;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_DX;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_D_CY;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_D_XOR;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_F7AMUX_O;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X2Y92_F7BMUX_O;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_A;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_A1;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_A2;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_A3;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_A4;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_A5;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_A6;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_AO5;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_AO6;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_AQ;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_AX;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_A_CY;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_A_XOR;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_B;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_B1;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_B2;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_B3;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_B4;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_B5;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_B6;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_BO5;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_BO6;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_BQ;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_BX;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_B_CY;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_B_XOR;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_C;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_C1;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_C2;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_C3;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_C4;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_C5;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_C6;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_CE;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_CLK;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_CO5;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_CO6;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_CQ;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_CX;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_C_CY;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_C_XOR;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_D;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_D1;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_D2;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_D3;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_D4;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_D5;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_D6;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_DO5;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_DO6;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_D_CY;
  wire [0:0] CLBLM_R_X3Y92_SLICE_X3Y92_D_XOR;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_A;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_A1;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_A2;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_A3;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_A4;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_A5;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_A6;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_AMUX;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_AO5;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_AO6;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_AX;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_A_CY;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_A_XOR;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_B;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_B1;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_B2;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_B3;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_B4;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_B5;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_B6;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_BO5;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_BO6;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_BQ;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_BX;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_B_CY;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_B_XOR;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_C;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_C1;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_C2;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_C3;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_C4;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_C5;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_C6;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_CE;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_CLK;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_CMUX;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_CO5;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_CO6;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_CQ;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_CX;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_C_CY;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_C_XOR;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_D;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_D1;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_D2;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_D3;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_D4;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_D5;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_D6;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_DO5;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_DO6;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_D_CY;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_D_XOR;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X2Y93_F7AMUX_O;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_A;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_A1;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_A2;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_A3;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_A4;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_A5;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_A6;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_AMUX;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_AO5;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_AO6;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_AQ;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_AX;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_A_CY;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_A_XOR;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_B;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_B1;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_B2;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_B3;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_B4;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_B5;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_B6;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_BO5;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_BO6;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_BQ;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_BX;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_B_CY;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_B_XOR;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_C;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_C1;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_C2;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_C3;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_C4;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_C5;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_C6;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_CE;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_CLK;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_CO5;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_CO6;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_CQ;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_CX;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_C_CY;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_C_XOR;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_D;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_D1;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_D2;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_D3;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_D4;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_D5;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_D6;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_DO5;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_DO6;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_DQ;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_DX;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_D_CY;
  wire [0:0] CLBLM_R_X3Y93_SLICE_X3Y93_D_XOR;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_A;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_A1;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_A2;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_A3;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_A4;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_A5;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_A6;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_AO5;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_AO6;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_AQ;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_A_CY;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_A_XOR;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_B;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_B1;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_B2;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_B3;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_B4;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_B5;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_B6;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_BO5;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_BO6;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_BQ;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_B_CY;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_B_XOR;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_C;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_C1;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_C2;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_C3;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_C4;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_C5;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_C6;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_CLK;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_CO5;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_CO6;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_CQ;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_C_CY;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_C_XOR;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_D;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_D1;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_D2;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_D3;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_D4;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_D5;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_D6;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_DMUX;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_DO5;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_DO6;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_D_CY;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_D_XOR;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X2Y94_SR;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_A;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_A1;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_A2;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_A3;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_A4;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_A5;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_A6;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_AMUX;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_AO5;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_AO6;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_AX;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_A_CY;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_A_XOR;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_B;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_B1;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_B2;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_B3;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_B4;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_B5;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_B6;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_BO5;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_BO6;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_BQ;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_BX;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_B_CY;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_B_XOR;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_C;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_C1;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_C2;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_C3;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_C4;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_C5;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_C6;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_CE;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_CLK;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_CMUX;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_CO5;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_CO6;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_CX;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_C_CY;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_C_XOR;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_D;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_D1;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_D2;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_D3;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_D4;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_D5;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_D6;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_DO5;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_DO6;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_D_CY;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_D_XOR;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_F7AMUX_O;
  wire [0:0] CLBLM_R_X3Y94_SLICE_X3Y94_F7BMUX_O;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_A;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_A1;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_A2;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_A3;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_A4;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_A5;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_A6;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_AO5;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_AO6;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_A_CY;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_A_XOR;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_B;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_B1;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_B2;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_B3;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_B4;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_B5;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_B6;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_BO5;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_BO6;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_B_CY;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_B_XOR;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_C;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_C1;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_C2;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_C3;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_C4;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_C5;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_C6;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_CO5;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_CO6;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_C_CY;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_C_XOR;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_D;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_D1;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_D2;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_D3;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_D4;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_D5;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_D6;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_DO5;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_DO6;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_D_CY;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X2Y95_D_XOR;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_A;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_A1;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_A2;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_A3;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_A4;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_A5;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_A6;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_AO5;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_AO6;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_A_CY;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_A_XOR;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_B;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_B1;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_B2;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_B3;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_B4;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_B5;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_B6;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_BO5;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_BO6;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_B_CY;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_B_XOR;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_C;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_C1;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_C2;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_C3;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_C4;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_C5;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_C6;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_CO5;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_CO6;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_C_CY;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_C_XOR;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_D;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_D1;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_D2;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_D3;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_D4;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_D5;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_D6;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_DO5;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_DO6;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_D_CY;
  wire [0:0] CLBLM_R_X3Y95_SLICE_X3Y95_D_XOR;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_A;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_A1;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_A2;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_A3;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_A4;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_A5;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_A6;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_AO5;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_AO6;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_AX;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_B;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_B1;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_B2;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_B3;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_B4;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_B5;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_B6;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_BO5;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_BO6;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_BX;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_C;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_C1;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_C2;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_C3;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_C4;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_C5;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_C6;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_CE;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_CLK;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_CO5;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_CO6;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_CX;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_D;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_D1;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_D2;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_D3;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_D4;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_D5;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_D6;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_DI;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_DO5;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_DO6;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X2Y96_DX;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_A;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_A1;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_A2;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_A3;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_A4;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_A5;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_A6;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_AMUX;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_AO5;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_AO6;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_A_CY;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_A_XOR;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_B;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_B1;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_B2;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_B3;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_B4;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_B5;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_B6;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_BMUX;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_BO5;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_BO6;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_B_CY;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_B_XOR;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_C;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_C1;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_C2;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_C3;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_C4;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_C5;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_C6;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_CO5;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_CO6;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_C_CY;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_C_XOR;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_D;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_D1;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_D2;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_D3;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_D4;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_D5;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_D6;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_DO5;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_DO6;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_D_CY;
  wire [0:0] CLBLM_R_X3Y96_SLICE_X3Y96_D_XOR;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_A;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_A1;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_A2;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_A3;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_A4;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_A5;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_A6;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_AO5;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_AO6;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_AX;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_B;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_B1;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_B2;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_B3;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_B4;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_B5;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_B6;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_BO5;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_BO6;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_BX;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_C;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_C1;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_C2;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_C3;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_C4;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_C5;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_C6;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_CE;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_CLK;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_CO5;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_CO6;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_CX;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_D;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_D1;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_D2;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_D3;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_D4;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_D5;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_D6;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_DI;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_DO5;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_DO6;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X2Y97_DX;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_A;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_A1;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_A2;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_A3;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_A4;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_A5;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_A6;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_AO5;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_AO6;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_A_CY;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_A_XOR;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_B;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_B1;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_B2;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_B3;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_B4;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_B5;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_B6;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_BO5;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_BO6;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_B_CY;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_B_XOR;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_C;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_C1;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_C2;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_C3;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_C4;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_C5;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_C6;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_CO5;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_CO6;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_C_CY;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_C_XOR;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_D;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_D1;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_D2;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_D3;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_D4;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_D5;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_D6;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_DMUX;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_DO5;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_DO6;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_D_CY;
  wire [0:0] CLBLM_R_X3Y97_SLICE_X3Y97_D_XOR;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_A;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_A1;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_A2;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_A3;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_A4;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_A5;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_A6;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_AO5;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_AO6;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_A_CY;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_A_XOR;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_B;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_B1;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_B2;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_B3;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_B4;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_B5;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_B6;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_BO5;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_BO6;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_B_CY;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_B_XOR;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_C;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_C1;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_C2;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_C3;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_C4;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_C5;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_C6;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_CO5;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_CO6;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_C_CY;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_C_XOR;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_D;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_D1;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_D2;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_D3;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_D4;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_D5;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_D6;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_DMUX;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_DO5;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_DO6;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_D_CY;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X2Y98_D_XOR;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_A;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_A1;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_A2;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_A3;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_A4;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_A5;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_A6;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_AMUX;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_AO5;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_AO6;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_A_CY;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_A_XOR;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_B;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_B1;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_B2;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_B3;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_B4;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_B5;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_B6;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_BO5;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_BO6;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_B_CY;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_B_XOR;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_C;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_C1;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_C2;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_C3;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_C4;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_C5;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_C6;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_CO5;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_CO6;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_C_CY;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_C_XOR;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_D;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_D1;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_D2;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_D3;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_D4;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_D5;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_D6;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_DMUX;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_DO5;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_DO6;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_D_CY;
  wire [0:0] CLBLM_R_X3Y98_SLICE_X3Y98_D_XOR;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_A;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_A1;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_A2;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_A3;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_A4;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_A5;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_A6;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_AMUX;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_AO5;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_AO6;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_AQ;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_AX;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_A_CY;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_A_XOR;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_B;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_B1;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_B2;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_B3;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_B4;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_B5;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_B6;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_BO5;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_BO6;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_B_CY;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_B_XOR;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_C;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_C1;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_C2;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_C3;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_C4;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_C5;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_C6;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_CE;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_CLK;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_CO5;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_CO6;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_C_CY;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_C_XOR;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_D;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_D1;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_D2;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_D3;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_D4;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_D5;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_D6;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_DO5;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_DO6;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_D_CY;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_D_XOR;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X2Y99_SR;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_A;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_A1;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_A2;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_A3;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_A4;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_A5;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_A6;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_AO5;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_AO6;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_A_CY;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_A_XOR;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_B;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_B1;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_B2;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_B3;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_B4;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_B5;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_B6;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_BO5;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_BO6;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_B_CY;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_B_XOR;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_C;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_C1;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_C2;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_C3;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_C4;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_C5;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_C6;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_CO5;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_CO6;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_C_CY;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_C_XOR;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_D;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_D1;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_D2;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_D3;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_D4;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_D5;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_D6;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_DO5;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_DO6;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_D_CY;
  wire [0:0] CLBLM_R_X3Y99_SLICE_X3Y99_D_XOR;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_A;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_A1;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_A2;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_A3;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_A4;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_A5;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_A5Q;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_A6;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_AMUX;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_AO5;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_AO6;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_AQ;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_AX;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_A_CY;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_A_XOR;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_B;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_B1;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_B2;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_B3;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_B4;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_B5;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_B5Q;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_B6;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_BMUX;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_BO5;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_BO6;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_BQ;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_BX;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_B_CY;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_B_XOR;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_C;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_C1;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_C2;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_C3;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_C4;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_C5;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_C6;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_CE;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_CLK;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_CO5;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_CO6;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_CQ;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_CX;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_C_CY;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_C_XOR;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_D;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_D1;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_D2;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_D3;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_D4;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_D5;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_D6;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_DO5;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_DO6;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_DQ;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_DX;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_D_CY;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_D_XOR;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X6Y90_SR;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_A;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_A1;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_A2;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_A3;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_A4;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_A5;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_A5Q;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_A6;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_AMUX;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_AO5;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_AO6;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_AQ;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_AX;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_A_CY;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_A_XOR;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_B;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_B1;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_B2;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_B3;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_B4;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_B5;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_B5Q;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_B6;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_BMUX;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_BO5;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_BO6;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_BQ;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_BX;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_B_CY;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_B_XOR;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_C;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_C1;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_C2;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_C3;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_C4;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_C5;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_C5Q;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_C6;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_CE;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_CLK;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_CMUX;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_CO5;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_CO6;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_CQ;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_CX;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_C_CY;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_C_XOR;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_D;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_D1;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_D2;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_D3;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_D4;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_D5;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_D6;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_DO5;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_DO6;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_DQ;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_DX;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_D_CY;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_D_XOR;
  wire [0:0] CLBLM_R_X5Y90_SLICE_X7Y90_SR;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_A;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_A1;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_A2;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_A3;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_A4;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_A5;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_A6;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_AO5;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_AO6;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_AQ;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_A_CY;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_A_XOR;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_B;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_B1;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_B2;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_B3;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_B4;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_B5;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_B6;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_BO5;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_BO6;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_B_CY;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_B_XOR;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_C;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_C1;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_C2;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_C3;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_C4;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_C5;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_C6;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_CLK;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_CO5;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_CO6;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_C_CY;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_C_XOR;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_D;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_D1;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_D2;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_D3;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_D4;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_D5;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_D6;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_DO5;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_DO6;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_D_CY;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_D_XOR;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X6Y91_SR;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_A;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_A1;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_A2;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_A3;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_A4;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_A5;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_A6;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_AO5;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_AO6;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_A_CY;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_A_XOR;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_B;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_B1;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_B2;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_B3;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_B4;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_B5;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_B6;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_BO5;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_BO6;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_B_CY;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_B_XOR;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_C;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_C1;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_C2;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_C3;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_C4;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_C5;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_C6;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_CO5;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_CO6;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_C_CY;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_C_XOR;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_D;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_D1;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_D2;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_D3;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_D4;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_D5;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_D6;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_DO5;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_DO6;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_D_CY;
  wire [0:0] CLBLM_R_X5Y91_SLICE_X7Y91_D_XOR;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_A;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_A1;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_A2;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_A3;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_A4;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_A5;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_A6;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_AO5;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_AO6;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_AQ;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_A_CY;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_A_XOR;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_B;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_B1;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_B2;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_B3;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_B4;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_B5;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_B6;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_BO5;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_BO6;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_BQ;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_B_CY;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_B_XOR;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_C;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_C1;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_C2;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_C3;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_C4;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_C5;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_C6;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_CLK;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_CO5;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_CO6;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_CQ;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_C_CY;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_C_XOR;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_D;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_D1;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_D2;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_D3;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_D4;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_D5;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_D6;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_DO5;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_DO6;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_D_CY;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_D_XOR;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X6Y92_SR;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_A;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_A1;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_A2;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_A3;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_A4;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_A5;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_A6;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_AO5;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_AO6;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_A_CY;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_A_XOR;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_B;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_B1;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_B2;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_B3;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_B4;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_B5;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_B6;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_BO5;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_BO6;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_B_CY;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_B_XOR;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_C;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_C1;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_C2;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_C3;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_C4;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_C5;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_C6;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_CO5;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_CO6;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_C_CY;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_C_XOR;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_D;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_D1;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_D2;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_D3;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_D4;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_D5;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_D6;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_DO5;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_DO6;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_D_CY;
  wire [0:0] CLBLM_R_X5Y92_SLICE_X7Y92_D_XOR;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_A;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_A1;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_A2;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_A3;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_A4;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_A5;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_A6;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_AMUX;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_AO5;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_AO6;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_AX;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_A_CY;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_A_XOR;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_B;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_B1;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_B2;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_B3;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_B4;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_B5;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_B6;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_BO5;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_BO6;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_BQ;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_BX;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_B_CY;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_B_XOR;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_C;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_C1;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_C2;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_C3;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_C4;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_C5;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_C6;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_CE;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_CLK;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_CO5;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_CO6;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_C_CY;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_C_XOR;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_D;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_D1;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_D2;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_D3;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_D4;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_D5;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_D6;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_DO5;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_DO6;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_D_CY;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_D_XOR;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X6Y93_F7AMUX_O;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_A;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_A1;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_A2;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_A3;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_A4;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_A5;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_A6;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_AO5;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_AO6;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_AQ;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_A_CY;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_A_XOR;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_B;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_B1;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_B2;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_B3;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_B4;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_B5;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_B6;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_BO5;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_BO6;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_BQ;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_B_CY;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_B_XOR;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_C;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_C1;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_C2;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_C3;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_C4;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_C5;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_C6;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_CLK;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_CO5;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_CO6;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_CQ;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_C_CY;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_C_XOR;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_D;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_D1;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_D2;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_D3;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_D4;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_D5;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_D6;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_DO5;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_DO6;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_D_CY;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_D_XOR;
  wire [0:0] CLBLM_R_X5Y93_SLICE_X7Y93_SR;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_A;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_A1;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_A2;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_A3;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_A4;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_A5;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_A6;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_AMUX;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_AO5;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_AO6;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_AQ;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_AX;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_A_CY;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_A_XOR;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_B;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_B1;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_B2;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_B3;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_B4;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_B5;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_B6;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_BO5;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_BO6;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_BQ;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_BX;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_B_CY;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_B_XOR;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_C;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_C1;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_C2;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_C3;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_C4;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_C5;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_C6;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_CE;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_CLK;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_CO5;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_CO6;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_C_CY;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_C_XOR;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_D;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_D1;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_D2;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_D3;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_D4;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_D5;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_D6;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_DO5;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_DO6;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_D_CY;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X6Y94_D_XOR;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_A;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_A1;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_A2;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_A3;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_A4;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_A5;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_A6;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_AMUX;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_AO5;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_AO6;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_A_CY;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_A_XOR;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_B;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_B1;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_B2;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_B3;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_B4;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_B5;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_B6;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_BO5;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_BO6;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_B_CY;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_B_XOR;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_C;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_C1;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_C2;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_C3;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_C4;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_C5;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_C6;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_CO5;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_CO6;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_C_CY;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_C_XOR;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_D;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_D1;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_D2;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_D3;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_D4;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_D5;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_D6;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_DO5;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_DO6;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_D_CY;
  wire [0:0] CLBLM_R_X5Y94_SLICE_X7Y94_D_XOR;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_A;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_A1;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_A2;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_A3;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_A4;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_A5;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_A6;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_AO5;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_AO6;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_AQ;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_A_CY;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_A_XOR;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_B;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_B1;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_B2;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_B3;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_B4;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_B5;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_B6;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_BMUX;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_BO5;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_BO6;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_B_CY;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_B_XOR;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_C;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_C1;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_C2;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_C3;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_C4;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_C5;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_C6;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_CLK;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_CO5;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_CO6;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_C_CY;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_C_XOR;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_D;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_D1;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_D2;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_D3;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_D4;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_D5;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_D6;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_DO5;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_DO6;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_D_CY;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_D_XOR;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X6Y95_SR;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_A;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_A1;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_A2;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_A3;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_A4;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_A5;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_A6;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_AO5;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_AO6;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_A_CY;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_A_XOR;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_B;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_B1;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_B2;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_B3;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_B4;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_B5;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_B6;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_BO5;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_BO6;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_B_CY;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_B_XOR;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_C;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_C1;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_C2;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_C3;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_C4;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_C5;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_C6;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_CO5;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_CO6;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_C_CY;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_C_XOR;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_D;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_D1;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_D2;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_D3;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_D4;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_D5;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_D6;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_DO5;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_DO6;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_D_CY;
  wire [0:0] CLBLM_R_X5Y95_SLICE_X7Y95_D_XOR;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_A;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_A1;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_A2;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_A3;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_A4;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_A5;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_A6;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_AO5;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_AO6;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_AQ;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_A_CY;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_A_XOR;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_B;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_B1;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_B2;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_B3;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_B4;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_B5;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_B6;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_BO5;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_BO6;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_B_CY;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_B_XOR;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_C;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_C1;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_C2;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_C3;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_C4;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_C5;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_C6;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_CE;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_CLK;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_CO5;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_CO6;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_C_CY;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_C_XOR;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_D;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_D1;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_D2;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_D3;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_D4;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_D5;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_D6;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_DO5;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_DO6;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_D_CY;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_D_XOR;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X6Y96_SR;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_A;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_A1;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_A2;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_A3;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_A4;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_A5;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_A6;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_AO5;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_AO6;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_AQ;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_A_CY;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_A_XOR;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_B;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_B1;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_B2;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_B3;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_B4;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_B5;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_B6;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_BO5;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_BO6;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_BQ;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_B_CY;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_B_XOR;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_C;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_C1;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_C2;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_C3;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_C4;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_C5;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_C6;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_CE;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_CLK;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_CMUX;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_CO5;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_CO6;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_C_CY;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_C_XOR;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_D;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_D1;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_D2;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_D3;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_D4;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_D5;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_D6;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_DO5;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_DO6;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_D_CY;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_D_XOR;
  wire [0:0] CLBLM_R_X5Y96_SLICE_X7Y96_SR;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_A;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_A1;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_A2;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_A3;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_A4;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_A5;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_A6;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_AMUX;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_AO5;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_AO6;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_AX;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_B;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_B1;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_B2;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_B3;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_B4;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_B5;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_B6;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_BMUX;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_BO5;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_BO6;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_BX;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_C;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_C1;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_C2;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_C3;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_C4;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_C5;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_C6;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_CE;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_CLK;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_CO5;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_CO6;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_CX;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_D;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_D1;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_D2;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_D3;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_D4;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_D5;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_D6;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_DI;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_DO5;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_DO6;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X6Y97_DX;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_A;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_A1;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_A2;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_A3;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_A4;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_A5;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_A6;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_AMUX;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_AO5;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_AO6;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_A_CY;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_A_XOR;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_B;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_B1;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_B2;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_B3;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_B4;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_B5;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_B6;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_BO5;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_BO6;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_B_CY;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_B_XOR;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_C;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_C1;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_C2;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_C3;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_C4;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_C5;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_C6;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_CO5;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_CO6;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_C_CY;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_C_XOR;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_D;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_D1;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_D2;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_D3;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_D4;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_D5;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_D6;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_DO5;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_DO6;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_D_CY;
  wire [0:0] CLBLM_R_X5Y97_SLICE_X7Y97_D_XOR;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_A;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_A1;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_A2;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_A3;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_A4;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_A5;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_A6;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_AO5;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_AO6;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_AX;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_B;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_B1;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_B2;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_B3;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_B4;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_B5;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_B6;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_BO5;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_BO6;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_BX;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_C;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_C1;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_C2;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_C3;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_C4;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_C5;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_C6;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_CE;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_CLK;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_CMUX;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_CO5;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_CO6;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_CX;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_D;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_D1;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_D2;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_D3;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_D4;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_D5;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_D6;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_DI;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_DMUX;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_DO5;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_DO6;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X6Y98_DX;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_A;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_A1;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_A2;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_A3;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_A4;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_A5;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_A6;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_AMUX;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_AO5;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_AO6;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_A_CY;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_A_XOR;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_B;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_B1;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_B2;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_B3;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_B4;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_B5;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_B6;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_BO5;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_BO6;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_B_CY;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_B_XOR;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_C;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_C1;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_C2;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_C3;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_C4;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_C5;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_C6;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_CO5;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_CO6;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_C_CY;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_C_XOR;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_D;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_D1;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_D2;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_D3;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_D4;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_D5;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_D6;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_DO5;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_DO6;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_D_CY;
  wire [0:0] CLBLM_R_X5Y98_SLICE_X7Y98_D_XOR;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_A;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_A1;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_A2;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_A3;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_A4;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_A5;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_A6;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_AO5;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_AO6;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_AQ;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_A_CY;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_A_XOR;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_B;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_B1;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_B2;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_B3;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_B4;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_B5;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_B6;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_BO5;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_BO6;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_B_CY;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_B_XOR;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_C;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_C1;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_C2;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_C3;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_C4;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_C5;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_C6;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_CE;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_CLK;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_CO5;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_CO6;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_C_CY;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_C_XOR;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_D;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_D1;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_D2;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_D3;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_D4;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_D5;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_D6;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_DO5;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_DO6;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_D_CY;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_D_XOR;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X6Y99_SR;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_A;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_A1;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_A2;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_A3;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_A4;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_A5;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_A6;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_AO5;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_AO6;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_AQ;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_A_CY;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_A_XOR;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_B;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_B1;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_B2;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_B3;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_B4;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_B5;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_B6;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_BMUX;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_BO5;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_BO6;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_B_CY;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_B_XOR;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_C;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_C1;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_C2;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_C3;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_C4;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_C5;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_C6;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_CE;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_CLK;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_CO5;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_CO6;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_C_CY;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_C_XOR;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_D;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_D1;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_D2;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_D3;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_D4;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_D5;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_D6;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_DO5;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_DO6;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_D_CY;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_D_XOR;
  wire [0:0] CLBLM_R_X5Y99_SLICE_X7Y99_SR;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_A;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_A1;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_A2;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_A3;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_A4;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_A5;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_A6;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_AO5;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_AO6;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_AQ;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_A_CY;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_A_XOR;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_B;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_B1;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_B2;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_B3;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_B4;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_B5;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_B6;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_BO5;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_BO6;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_BQ;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_B_CY;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_B_XOR;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_C;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_C1;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_C2;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_C3;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_C4;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_C5;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_C6;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_CLK;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_CO5;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_CO6;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_C_CY;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_C_XOR;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_D;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_D1;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_D2;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_D3;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_D4;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_D5;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_D6;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_DO5;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_DO6;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_D_CY;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_D_XOR;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X8Y87_SR;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_A;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_A1;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_A2;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_A3;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_A4;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_A5;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_A6;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_AO5;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_AO6;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_A_CY;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_A_XOR;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_B;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_B1;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_B2;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_B3;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_B4;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_B5;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_B6;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_BO5;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_BO6;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_B_CY;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_B_XOR;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_C;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_C1;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_C2;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_C3;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_C4;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_C5;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_C6;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_CO5;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_CO6;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_C_CY;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_C_XOR;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_D;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_D1;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_D2;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_D3;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_D4;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_D5;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_D6;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_DO5;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_DO6;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_D_CY;
  wire [0:0] CLBLM_R_X7Y87_SLICE_X9Y87_D_XOR;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_A;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_A1;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_A2;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_A3;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_A4;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_A5;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_A6;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_AO5;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_AO6;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_AQ;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_A_CY;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_A_XOR;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_B;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_B1;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_B2;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_B3;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_B4;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_B5;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_B6;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_BO5;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_BO6;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_B_CY;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_B_XOR;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_C;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_C1;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_C2;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_C3;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_C4;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_C5;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_C6;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_CLK;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_CO5;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_CO6;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_C_CY;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_C_XOR;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_D;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_D1;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_D2;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_D3;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_D4;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_D5;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_D6;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_DO5;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_DO6;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_D_CY;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_D_XOR;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X8Y88_SR;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_A;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_A1;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_A2;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_A3;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_A4;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_A5;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_A6;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_AO5;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_AO6;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_A_CY;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_A_XOR;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_B;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_B1;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_B2;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_B3;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_B4;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_B5;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_B6;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_BO5;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_BO6;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_B_CY;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_B_XOR;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_C;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_C1;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_C2;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_C3;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_C4;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_C5;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_C6;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_CO5;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_CO6;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_C_CY;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_C_XOR;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_D;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_D1;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_D2;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_D3;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_D4;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_D5;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_D6;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_DO5;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_DO6;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_D_CY;
  wire [0:0] CLBLM_R_X7Y88_SLICE_X9Y88_D_XOR;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_A;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_A1;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_A2;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_A3;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_A4;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_A5;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_A6;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_AO5;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_AO6;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_AQ;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_A_CY;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_A_XOR;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_B;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_B1;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_B2;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_B3;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_B4;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_B5;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_B5Q;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_B6;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_BMUX;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_BO5;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_BO6;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_BQ;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_B_CY;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_B_XOR;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_C;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_C1;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_C2;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_C3;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_C4;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_C5;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_C6;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_CE;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_CLK;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_CO5;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_CO6;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_C_CY;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_C_XOR;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_D;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_D1;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_D2;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_D3;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_D4;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_D5;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_D6;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_DO5;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_DO6;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_D_CY;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_D_XOR;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X8Y89_SR;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_A;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_A1;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_A2;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_A3;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_A4;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_A5;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_A6;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_AMUX;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_AO5;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_AO6;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_AQ;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_A_CY;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_A_XOR;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_B;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_B1;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_B2;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_B3;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_B4;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_B5;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_B6;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_BO5;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_BO6;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_BQ;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_B_CY;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_B_XOR;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_C;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_C1;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_C2;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_C3;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_C4;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_C5;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_C6;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_CE;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_CLK;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_CO5;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_CO6;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_C_CY;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_C_XOR;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_D;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_D1;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_D2;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_D3;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_D4;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_D5;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_D6;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_DO5;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_DO6;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_D_CY;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_D_XOR;
  wire [0:0] CLBLM_R_X7Y89_SLICE_X9Y89_SR;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_A;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_A1;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_A2;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_A3;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_A4;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_A5;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_A6;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_AO5;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_AO6;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_AQ;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_A_CY;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_A_XOR;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_B;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_B1;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_B2;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_B3;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_B4;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_B5;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_B6;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_BO5;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_BO6;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_BQ;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_B_CY;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_B_XOR;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_C;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_C1;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_C2;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_C3;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_C4;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_C5;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_C6;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_CLK;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_CO5;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_CO6;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_C_CY;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_C_XOR;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_D;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_D1;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_D2;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_D3;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_D4;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_D5;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_D6;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_DO5;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_DO6;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_D_CY;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_D_XOR;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X8Y90_SR;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_A;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_A1;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_A2;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_A3;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_A4;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_A5;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_A5Q;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_A6;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_AMUX;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_AO5;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_AO6;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_AQ;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_A_CY;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_A_XOR;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_B;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_B1;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_B2;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_B3;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_B4;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_B5;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_B6;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_BO5;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_BO6;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_BQ;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_B_CY;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_B_XOR;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_C;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_C1;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_C2;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_C3;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_C4;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_C5;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_C6;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_CLK;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_CO5;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_CO6;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_CQ;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_C_CY;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_C_XOR;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_D;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_D1;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_D2;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_D3;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_D4;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_D5;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_D6;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_DO5;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_DO6;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_D_CY;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_D_XOR;
  wire [0:0] CLBLM_R_X7Y90_SLICE_X9Y90_SR;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_A;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_A1;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_A2;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_A3;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_A4;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_A5;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_A6;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_AO5;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_AO6;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_AQ;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_A_CY;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_A_XOR;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_B;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_B1;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_B2;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_B3;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_B4;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_B5;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_B6;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_BO5;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_BO6;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_B_CY;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_B_XOR;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_C;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_C1;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_C2;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_C3;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_C4;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_C5;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_C6;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_CLK;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_CO5;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_CO6;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_C_CY;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_C_XOR;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_D;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_D1;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_D2;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_D3;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_D4;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_D5;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_D6;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_DO5;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_DO6;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_D_CY;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_D_XOR;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X8Y91_SR;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_A;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_A1;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_A2;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_A3;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_A4;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_A5;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_A6;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_AO5;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_AO6;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_AQ;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_A_CY;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_A_XOR;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_B;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_B1;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_B2;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_B3;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_B4;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_B5;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_B6;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_BO5;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_BO6;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_BQ;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_B_CY;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_B_XOR;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_C;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_C1;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_C2;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_C3;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_C4;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_C5;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_C6;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_CLK;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_CO5;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_CO6;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_CQ;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_C_CY;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_C_XOR;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_D;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_D1;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_D2;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_D3;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_D4;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_D5;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_D6;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_DO5;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_DO6;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_D_CY;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_D_XOR;
  wire [0:0] CLBLM_R_X7Y91_SLICE_X9Y91_SR;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_A;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_A1;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_A2;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_A3;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_A4;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_A5;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_A6;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_AO5;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_AO6;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_A_CY;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_A_XOR;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_B;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_B1;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_B2;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_B3;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_B4;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_B5;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_B6;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_BO5;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_BO6;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_B_CY;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_B_XOR;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_C;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_C1;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_C2;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_C3;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_C4;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_C5;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_C6;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_CE;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_CLK;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_CO5;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_CO6;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_C_CY;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_C_XOR;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_D;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_D1;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_D2;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_D3;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_D4;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_D5;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_D6;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_DO5;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_DO6;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_D_CY;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_D_XOR;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X8Y93_SR;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_A;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_A1;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_A2;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_A3;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_A4;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_A5;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_A6;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_AO5;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_AO6;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_A_CY;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_A_XOR;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_B;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_B1;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_B2;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_B3;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_B4;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_B5;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_B6;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_BO5;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_BO6;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_B_CY;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_B_XOR;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_C;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_C1;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_C2;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_C3;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_C4;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_C5;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_C6;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_CO5;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_CO6;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_C_CY;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_C_XOR;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_D;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_D1;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_D2;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_D3;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_D4;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_D5;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_D6;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_DO5;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_DO6;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_D_CY;
  wire [0:0] CLBLM_R_X7Y93_SLICE_X9Y93_D_XOR;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_A;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_A1;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_A2;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_A3;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_A4;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_A5;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_A6;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_AO5;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_AO6;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_A_CY;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_A_XOR;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_B;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_B1;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_B2;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_B3;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_B4;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_B5;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_B6;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_BO5;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_BO6;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_B_CY;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_B_XOR;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_C;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_C1;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_C2;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_C3;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_C4;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_C5;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_C6;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_CE;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_CLK;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_CO5;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_CO6;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_C_CY;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_C_XOR;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_D;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_D1;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_D2;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_D3;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_D4;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_D5;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_D6;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_DO5;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_DO6;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_D_CY;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_D_XOR;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X8Y94_SR;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_A;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_A1;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_A2;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_A3;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_A4;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_A5;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_A6;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_AO5;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_AO6;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_A_CY;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_A_XOR;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_B;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_B1;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_B2;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_B3;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_B4;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_B5;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_B6;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_BO5;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_BO6;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_B_CY;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_B_XOR;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_C;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_C1;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_C2;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_C3;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_C4;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_C5;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_C6;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_CE;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_CLK;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_CO5;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_CO6;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_C_CY;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_C_XOR;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_D;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_D1;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_D2;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_D3;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_D4;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_D5;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_D6;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_DO5;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_DO6;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_D_CY;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_D_XOR;
  wire [0:0] CLBLM_R_X7Y94_SLICE_X9Y94_SR;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_A;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_A1;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_A2;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_A3;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_A4;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_A5;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_A6;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_AO5;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_AO6;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_AQ;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_A_CY;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_A_XOR;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_B;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_B1;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_B2;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_B3;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_B4;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_B5;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_B6;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_BMUX;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_BO5;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_BO6;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_B_CY;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_B_XOR;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_C;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_C1;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_C2;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_C3;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_C4;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_C5;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_C6;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_CE;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_CLK;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_CMUX;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_CO5;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_CO6;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_C_CY;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_C_XOR;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_D;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_D1;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_D2;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_D3;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_D4;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_D5;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_D6;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_DO5;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_DO6;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_D_CY;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_D_XOR;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X8Y96_SR;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_A;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_A1;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_A2;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_A3;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_A4;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_A5;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_A6;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_AO5;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_AO6;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_AQ;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_A_CY;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_A_XOR;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_B;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_B1;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_B2;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_B3;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_B4;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_B5;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_B6;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_BO5;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_BO6;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_B_CY;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_B_XOR;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_C;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_C1;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_C2;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_C3;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_C4;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_C5;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_C6;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_CE;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_CLK;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_CO5;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_CO6;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_C_CY;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_C_XOR;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_D;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_D1;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_D2;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_D3;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_D4;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_D5;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_D6;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_DO5;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_DO6;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_D_CY;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_D_XOR;
  wire [0:0] CLBLM_R_X7Y96_SLICE_X9Y96_SR;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_A;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_A1;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_A2;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_A3;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_A4;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_A5;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_A6;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_AO5;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_AO6;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_AQ;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_A_CY;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_A_XOR;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_B;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_B1;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_B2;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_B3;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_B4;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_B5;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_B6;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_BMUX;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_BO5;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_BO6;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_B_CY;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_B_XOR;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_C;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_C1;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_C2;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_C3;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_C4;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_C5;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_C6;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_CE;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_CLK;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_CO5;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_CO6;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_C_CY;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_C_XOR;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_D;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_D1;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_D2;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_D3;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_D4;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_D5;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_D6;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_DMUX;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_DO5;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_DO6;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_D_CY;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_D_XOR;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X8Y97_SR;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_A;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_A1;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_A2;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_A3;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_A4;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_A5;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_A5Q;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_A6;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_AMUX;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_AO5;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_AO6;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_AQ;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_A_CY;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_A_XOR;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_B;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_B1;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_B2;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_B3;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_B4;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_B5;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_B5Q;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_B6;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_BMUX;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_BO5;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_BO6;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_BQ;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_B_CY;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_B_XOR;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_C;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_C1;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_C2;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_C3;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_C4;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_C5;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_C6;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_CE;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_CLK;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_CMUX;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_CO5;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_CO6;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_C_CY;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_C_XOR;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_D;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_D1;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_D2;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_D3;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_D4;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_D5;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_D6;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_DO5;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_DO6;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_D_CY;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_D_XOR;
  wire [0:0] CLBLM_R_X7Y97_SLICE_X9Y97_SR;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_A;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_A1;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_A2;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_A3;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_A4;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_A5;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_A6;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_AMUX;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_AO5;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_AO6;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_AX;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_A_CY;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_A_XOR;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_B;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_B1;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_B2;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_B3;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_B4;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_B5;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_B6;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_BO5;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_BO6;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_B_CY;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_B_XOR;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_C;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_C1;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_C2;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_C3;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_C4;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_C5;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_C6;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_CO5;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_CO6;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_C_CY;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_C_XOR;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_D;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_D1;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_D2;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_D3;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_D4;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_D5;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_D6;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_DO5;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_DO6;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_D_CY;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_D_XOR;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X8Y98_F7AMUX_O;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_A;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_A1;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_A2;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_A3;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_A4;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_A5;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_A6;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_AO5;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_AO6;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_AQ;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_A_CY;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_A_XOR;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_B;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_B1;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_B2;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_B3;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_B4;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_B5;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_B6;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_BO5;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_BO6;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_B_CY;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_B_XOR;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_C;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_C1;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_C2;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_C3;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_C4;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_C5;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_C6;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_CE;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_CLK;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_CO5;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_CO6;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_C_CY;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_C_XOR;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_D;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_D1;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_D2;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_D3;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_D4;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_D5;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_D6;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_DO5;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_DO6;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_D_CY;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_D_XOR;
  wire [0:0] CLBLM_R_X7Y98_SLICE_X9Y98_SR;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_A;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_A1;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_A2;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_A3;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_A4;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_A5;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_A6;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_AO5;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_AO6;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_AQ;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_A_CY;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_A_XOR;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_B;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_B1;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_B2;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_B3;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_B4;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_B5;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_B6;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_BO5;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_BO6;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_B_CY;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_B_XOR;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_C;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_C1;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_C2;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_C3;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_C4;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_C5;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_C6;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_CE;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_CLK;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_CO5;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_CO6;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_C_CY;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_C_XOR;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_D;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_D1;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_D2;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_D3;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_D4;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_D5;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_D6;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_DO5;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_DO6;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_D_CY;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_D_XOR;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X8Y99_SR;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_A;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_A1;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_A2;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_A3;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_A4;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_A5;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_A6;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_AO5;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_AO6;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_AQ;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_A_CY;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_A_XOR;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_B;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_B1;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_B2;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_B3;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_B4;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_B5;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_B6;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_BO5;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_BO6;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_B_CY;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_B_XOR;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_C;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_C1;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_C2;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_C3;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_C4;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_C5;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_C6;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_CE;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_CLK;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_CO5;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_CO6;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_C_CY;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_C_XOR;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_D;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_D1;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_D2;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_D3;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_D4;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_D5;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_D6;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_DO5;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_DO6;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_D_CY;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_D_XOR;
  wire [0:0] CLBLM_R_X7Y99_SLICE_X9Y99_SR;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_O;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_O;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_I;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_I;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_TQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_TQ;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_O;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_D;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_O;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y128_D;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y128_O;


  (* KEEP, DONT_TOUCH, BEL = "RAMB36E1" *)
  RAMB36E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_40(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_41(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_42(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_43(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_44(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_45(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_46(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_47(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_48(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_49(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_50(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_51(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_52(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_53(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_54(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_55(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_56(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_59(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_61(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_62(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_63(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_64(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_65(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_66(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_67(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_68(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_69(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_70(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(36'h000000000),
    .INIT_B(36'h000000000),
    .IS_CLKARDCLK_INVERTED(0),
    .IS_CLKBWRCLK_INVERTED(0),
    .IS_ENARDEN_INVERTED(0),
    .IS_ENBWREN_INVERTED(0),
    .IS_RSTRAMARSTRAM_INVERTED(1),
    .IS_RSTRAMB_INVERTED(1),
    .IS_RSTREGARSTREG_INVERTED(1),
    .IS_RSTREGB_INVERTED(1),
    .RAM_MODE("TDP"),
    .READ_WIDTH_A(4),
    .READ_WIDTH_B(4),
    .SRVAL_A(36'h000000000),
    .SRVAL_B(36'h000000000),
    .WRITE_MODE_A("READ_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(4),
    .WRITE_WIDTH_B(4)
  ) BRAM_L_X6Y90_RAMB36_X0Y18_RAMB36E1 (
.ADDRARDADDR({1'b1, CLBLM_R_X5Y90_SLICE_X6Y90_B5Q, CLBLM_R_X5Y90_SLICE_X6Y90_A5Q, CLBLM_R_X5Y90_SLICE_X6Y90_DQ, CLBLM_R_X5Y90_SLICE_X6Y90_CQ, CLBLM_R_X5Y90_SLICE_X6Y90_BQ, CLBLM_R_X5Y90_SLICE_X6Y90_AQ, CLBLM_R_X5Y90_SLICE_X7Y90_C5Q, CLBLM_R_X5Y90_SLICE_X7Y90_B5Q, CLBLM_R_X5Y90_SLICE_X7Y90_A5Q, CLBLM_R_X5Y90_SLICE_X7Y90_DQ, CLBLM_R_X5Y90_SLICE_X7Y90_CQ, CLBLM_R_X5Y90_SLICE_X7Y90_BQ, CLBLM_R_X5Y90_SLICE_X7Y90_AQ, 1'b1, 1'b1}),
.ADDRBWRADDR({1'b1, CLBLM_R_X7Y89_SLICE_X8Y89_B5Q, CLBLM_R_X7Y89_SLICE_X8Y89_BQ, CLBLM_R_X7Y89_SLICE_X8Y89_AQ, CLBLM_R_X7Y89_SLICE_X9Y89_BQ, CLBLM_R_X7Y89_SLICE_X9Y89_AQ, CLBLM_L_X8Y89_SLICE_X10Y89_A5Q, CLBLM_R_X7Y87_SLICE_X8Y87_AQ, CLBLM_R_X7Y91_SLICE_X8Y91_AQ, CLBLM_R_X7Y87_SLICE_X8Y87_BQ, CLBLM_R_X7Y91_SLICE_X9Y91_AQ, CLBLM_R_X7Y90_SLICE_X9Y90_CQ, CLBLM_R_X7Y90_SLICE_X9Y90_BQ, CLBLM_R_X7Y90_SLICE_X9Y90_A5Q, 1'b1, 1'b1}),
.CLKARDCLK(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CLKBWRCLK(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.DIADI({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, CLBLM_R_X5Y91_SLICE_X6Y91_AQ, CLBLM_R_X5Y93_SLICE_X7Y93_AQ, CLBLM_R_X5Y93_SLICE_X7Y93_BQ}),
.DIBDI({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1}),
.DIPADIP({1'b0, 1'b0, 1'b1, 1'b1}),
.DIPBDIP({1'b0, 1'b0, 1'b1, 1'b1}),
.DOADO({BRAM_L_X6Y90_RAMB36_X0Y18_DOADO31, BRAM_L_X6Y90_RAMB36_X0Y18_DOADO30, BRAM_L_X6Y90_RAMB36_X0Y18_DOADO29, BRAM_L_X6Y90_RAMB36_X0Y18_DOADO28, BRAM_L_X6Y90_RAMB36_X0Y18_DOADO27, BRAM_L_X6Y90_RAMB36_X0Y18_DOADO26, BRAM_L_X6Y90_RAMB36_X0Y18_DOADO25, BRAM_L_X6Y90_RAMB36_X0Y18_DOADO24, BRAM_L_X6Y90_RAMB36_X0Y18_DOADO23, BRAM_L_X6Y90_RAMB36_X0Y18_DOADO22, BRAM_L_X6Y90_RAMB36_X0Y18_DOADO21, BRAM_L_X6Y90_RAMB36_X0Y18_DOADO20, BRAM_L_X6Y90_RAMB36_X0Y18_DOADO19, BRAM_L_X6Y90_RAMB36_X0Y18_DOADO18, BRAM_L_X6Y90_RAMB36_X0Y18_DOADO17, BRAM_L_X6Y90_RAMB36_X0Y18_DOADO16, BRAM_L_X6Y90_RAMB36_X0Y18_DOADO15, BRAM_L_X6Y90_RAMB36_X0Y18_DOADO14, BRAM_L_X6Y90_RAMB36_X0Y18_DOADO13, BRAM_L_X6Y90_RAMB36_X0Y18_DOADO12, BRAM_L_X6Y90_RAMB36_X0Y18_DOADO11, BRAM_L_X6Y90_RAMB36_X0Y18_DOADO10, BRAM_L_X6Y90_RAMB36_X0Y18_DOADO9, BRAM_L_X6Y90_RAMB36_X0Y18_DOADO8, BRAM_L_X6Y90_RAMB36_X0Y18_DOADO7, BRAM_L_X6Y90_RAMB36_X0Y18_DOADO6, BRAM_L_X6Y90_RAMB36_X0Y18_DOADO5, BRAM_L_X6Y90_RAMB36_X0Y18_DOADO4, BRAM_L_X6Y90_RAMB36_X0Y18_DOADO3, BRAM_L_X6Y90_RAMB36_X0Y18_DOADO2, BRAM_L_X6Y90_RAMB36_X0Y18_DOADO1, BRAM_L_X6Y90_RAMB36_X0Y18_DOADO0}),
.DOBDO({BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO31, BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO30, BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO29, BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO28, BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO27, BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO26, BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO25, BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO24, BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO23, BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO22, BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO21, BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO20, BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO19, BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO18, BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO17, BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO16, BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO15, BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO14, BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO13, BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO12, BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO11, BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO10, BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO9, BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO8, BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO7, BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO6, BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO5, BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO4, BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO3, BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO2, BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO1, BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO0}),
.DOPADOP({BRAM_L_X6Y90_RAMB36_X0Y18_DOPADOP3, BRAM_L_X6Y90_RAMB36_X0Y18_DOPADOP2, BRAM_L_X6Y90_RAMB36_X0Y18_DOPADOP1, BRAM_L_X6Y90_RAMB36_X0Y18_DOPADOP0}),
.DOPBDOP({BRAM_L_X6Y90_RAMB36_X0Y18_DOPBDOP3, BRAM_L_X6Y90_RAMB36_X0Y18_DOPBDOP2, BRAM_L_X6Y90_RAMB36_X0Y18_DOPBDOP1, BRAM_L_X6Y90_RAMB36_X0Y18_DOPBDOP0}),
.ENARDEN(CLBLM_R_X5Y93_SLICE_X7Y93_CQ),
.ENBWREN(1'b1),
.REGCEAREGCE(1'b0),
.REGCEB(1'b0),
.RSTRAMARSTRAM(1'b1),
.RSTRAMB(1'b1),
.RSTREGARSTREG(1'b1),
.RSTREGB(1'b1),
.WEA({1'b1, 1'b1, 1'b1, 1'b1}),
.WEBWE({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0})
  );


  (* KEEP, DONT_TOUCH, BEL = "RAMB36E1" *)
  RAMB36E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h210A112821092008110120062005210C114B210B110521162115111980F61000),
    .INIT_01(256'h810F810F810F810F810F810F810F810F810F810F810F810F810F810F2114111E),
    .INIT_02(256'h16041D201A16221580C0CF0047A0170246A016011D201A1580CE80F680D880CE),
    .INIT_03(256'h80EB14071A15190B80628074221680C0CF00CF00CF0047A01708CE00CE0046A0),
    .INIT_04(256'h13FF120011005820208027801701804D804D804D804D805A80EB14071A16190C),
    .INIT_05(256'h24602240212014071A14190A88005850120091015852920160562A6060592960),
    .INIT_06(256'h5871910168702CA09201586C3AA0606B2BA015011C091B081A14190A8800810A),
    .INIT_07(256'h26091601260696011E06688129E01702143A134E1A14190A88002214210A39A0),
    .INIT_08(256'h1B0B2008688F2A8026081601688C2AE0580E2009260596011E0568882960580E),
    .INIT_09(256'h940160A52A80940160A52A80940160A52A80940160A52A8068A7296093011C15),
    .INIT_0A(256'h940160BE2A8068BF29603CC01C1616011B0C2609160168A72A80940160A52A80),
    .INIT_0B(256'h8800200968BF2A80940160BE2A80940160BE2A80940160BE2A80940160BE2A80),
    .INIT_0C(256'h11131D05880032A060CD2A8068CD2F603AA060CD2A6068C82E60150214371301),
    .INIT_0D(256'h14041A16190C68E2296013061A0619058800815A120511391D06815A14061205),
    .INIT_0E(256'h224078F52A6033401305880058E980EB14041A15190B68EA2A60130658E180EB),
    .INIT_0F(256'h234061032C2014001300123C1150206027A01701880058ED9201810A24602120),
    .INIT_10(256'h804D880027A0170027A01701880020A058FD930161082B40140058FD94012420),
    .INIT_11(256'h61262960332013038800805A80EB14021A16190C80EB14021A15190B804D804D),
    .INIT_12(256'h24602120224061332A6033401303880039601303591E9101810A246021202240),
    .INIT_13(256'h31E01702880039E01702812931E017028800811C88003A601303592B9201810A),
    .INIT_14(256'h170281299202170288003AE01704811C9204170488003AE039E01702812932E0),
    .INIT_15(256'h61612DE0170461612DE0170188003AE01702811C920217028800812988003AE0),
    .INIT_16(256'h170461762DE01701813E616C2DE01702813861682DE0170661682DE017058136),
    .INIT_17(256'h170861822DE0170661822DE0170261822DE01700814661762DE0170761762DE0),
    .INIT_18(256'h815261902DE0170761902DE0170361902DE0170261902DE01701814C69832DE0),
    .INIT_19(256'h000000000000000000000000000000008800815461972DE0170161972DE01700),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_40(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_41(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_42(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_43(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_44(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_45(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_46(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_47(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_48(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_49(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_50(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_51(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_52(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_53(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_54(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_55(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_56(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_59(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_61(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_62(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_63(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_64(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_65(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_66(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_67(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_68(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_69(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_70(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(36'h000000000),
    .INIT_B(36'h000000000),
    .IS_CLKARDCLK_INVERTED(0),
    .IS_CLKBWRCLK_INVERTED(1),
    .IS_ENARDEN_INVERTED(0),
    .IS_ENBWREN_INVERTED(1),
    .IS_RSTRAMARSTRAM_INVERTED(1),
    .IS_RSTRAMB_INVERTED(1),
    .IS_RSTREGARSTREG_INVERTED(1),
    .IS_RSTREGB_INVERTED(1),
    .RAM_MODE("TDP"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(2),
    .SRVAL_A(36'h000000000),
    .SRVAL_B(36'h000000000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(2)
  ) BRAM_L_X6Y95_RAMB36_X0Y19_RAMB36E1 (
.ADDRARDADDR({1'b1, CLBLM_R_X7Y97_SLICE_X8Y97_AQ, CLBLM_R_X7Y99_SLICE_X9Y99_AQ, CLBLM_R_X7Y98_SLICE_X9Y98_AQ, CLBLM_R_X7Y96_SLICE_X9Y96_AQ, CLBLM_R_X7Y96_SLICE_X8Y96_AQ, CLBLM_R_X5Y96_SLICE_X6Y96_AQ, CLBLM_R_X5Y96_SLICE_X7Y96_BQ, CLBLM_R_X5Y96_SLICE_X7Y96_AQ, CLBLM_R_X5Y99_SLICE_X6Y99_AQ, CLBLM_R_X5Y99_SLICE_X7Y99_AQ, CLBLM_R_X7Y99_SLICE_X8Y99_AQ, 1'b0, 1'b0, 1'b0, 1'b0}),
.ADDRBWRADDR({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
.CLKARDCLK(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CLKBWRCLK(1'b1),
.DIADI({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
.DIBDI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
.DIPADIP({1'b0, 1'b0, 1'b0, 1'b0}),
.DIPBDIP({1'b1, 1'b1, 1'b1, 1'b1}),
.DOADO({BRAM_L_X6Y95_RAMB36_X0Y19_DOADO31, BRAM_L_X6Y95_RAMB36_X0Y19_DOADO30, BRAM_L_X6Y95_RAMB36_X0Y19_DOADO29, BRAM_L_X6Y95_RAMB36_X0Y19_DOADO28, BRAM_L_X6Y95_RAMB36_X0Y19_DOADO27, BRAM_L_X6Y95_RAMB36_X0Y19_DOADO26, BRAM_L_X6Y95_RAMB36_X0Y19_DOADO25, BRAM_L_X6Y95_RAMB36_X0Y19_DOADO24, BRAM_L_X6Y95_RAMB36_X0Y19_DOADO23, BRAM_L_X6Y95_RAMB36_X0Y19_DOADO22, BRAM_L_X6Y95_RAMB36_X0Y19_DOADO21, BRAM_L_X6Y95_RAMB36_X0Y19_DOADO20, BRAM_L_X6Y95_RAMB36_X0Y19_DOADO19, BRAM_L_X6Y95_RAMB36_X0Y19_DOADO18, BRAM_L_X6Y95_RAMB36_X0Y19_DOADO17, BRAM_L_X6Y95_RAMB36_X0Y19_DOADO16, BRAM_L_X6Y95_RAMB36_X0Y19_DOADO15, BRAM_L_X6Y95_RAMB36_X0Y19_DOADO14, BRAM_L_X6Y95_RAMB36_X0Y19_DOADO13, BRAM_L_X6Y95_RAMB36_X0Y19_DOADO12, BRAM_L_X6Y95_RAMB36_X0Y19_DOADO11, BRAM_L_X6Y95_RAMB36_X0Y19_DOADO10, BRAM_L_X6Y95_RAMB36_X0Y19_DOADO9, BRAM_L_X6Y95_RAMB36_X0Y19_DOADO8, BRAM_L_X6Y95_RAMB36_X0Y19_DOADO7, BRAM_L_X6Y95_RAMB36_X0Y19_DOADO6, BRAM_L_X6Y95_RAMB36_X0Y19_DOADO5, BRAM_L_X6Y95_RAMB36_X0Y19_DOADO4, BRAM_L_X6Y95_RAMB36_X0Y19_DOADO3, BRAM_L_X6Y95_RAMB36_X0Y19_DOADO2, BRAM_L_X6Y95_RAMB36_X0Y19_DOADO1, BRAM_L_X6Y95_RAMB36_X0Y19_DOADO0}),
.DOBDO({BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO31, BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO30, BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO29, BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO28, BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO27, BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO26, BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO25, BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO24, BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO23, BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO22, BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO21, BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO20, BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO19, BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO18, BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO17, BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO16, BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO15, BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO14, BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO13, BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO12, BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO11, BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO10, BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO9, BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO8, BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO7, BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO6, BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO5, BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO4, BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO3, BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO2, BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO1, BRAM_L_X6Y95_RAMB36_X0Y19_DOBDO0}),
.DOPADOP({BRAM_L_X6Y95_RAMB36_X0Y19_DOPADOP3, BRAM_L_X6Y95_RAMB36_X0Y19_DOPADOP2, BRAM_L_X6Y95_RAMB36_X0Y19_DOPADOP1, BRAM_L_X6Y95_RAMB36_X0Y19_DOPADOP0}),
.DOPBDOP({BRAM_L_X6Y95_RAMB36_X0Y19_DOPBDOP3, BRAM_L_X6Y95_RAMB36_X0Y19_DOPBDOP2, BRAM_L_X6Y95_RAMB36_X0Y19_DOPBDOP1, BRAM_L_X6Y95_RAMB36_X0Y19_DOPBDOP0}),
.ENARDEN(CLBLM_L_X8Y97_SLICE_X11Y97_CO6),
.ENBWREN(1'b1),
.REGCEAREGCE(1'b0),
.REGCEB(1'b0),
.RSTRAMARSTRAM(1'b1),
.RSTRAMB(1'b1),
.RSTREGARSTREG(1'b1),
.RSTREGB(1'b1),
.WEA({1'b0, 1'b0, 1'b0, 1'b0}),
.WEBWE({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y90_SLICE_X0Y90_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y90_SLICE_X0Y90_DO5),
.O6(CLBLL_L_X2Y90_SLICE_X0Y90_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y90_SLICE_X0Y90_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y90_SLICE_X0Y90_CO5),
.O6(CLBLL_L_X2Y90_SLICE_X0Y90_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y90_SLICE_X0Y90_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y90_SLICE_X0Y90_BO5),
.O6(CLBLL_L_X2Y90_SLICE_X0Y90_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y90_SLICE_X0Y90_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y90_SLICE_X0Y90_AO5),
.O6(CLBLL_L_X2Y90_SLICE_X0Y90_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y90_SLICE_X1Y90_A_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLL_L_X2Y92_SLICE_X1Y92_AO6),
.D(CLBLL_L_X4Y92_SLICE_X4Y92_AO6),
.Q(CLBLL_L_X2Y90_SLICE_X1Y90_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y90_SLICE_X1Y90_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y90_SLICE_X1Y90_DO5),
.O6(CLBLL_L_X2Y90_SLICE_X1Y90_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y90_SLICE_X1Y90_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y90_SLICE_X1Y90_CO5),
.O6(CLBLL_L_X2Y90_SLICE_X1Y90_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y90_SLICE_X1Y90_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y90_SLICE_X1Y90_BO5),
.O6(CLBLL_L_X2Y90_SLICE_X1Y90_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y90_SLICE_X1Y90_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y90_SLICE_X1Y90_AO5),
.O6(CLBLL_L_X2Y90_SLICE_X1Y90_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y91_SLICE_X0Y91_A_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLL_L_X2Y93_SLICE_X0Y93_DO6),
.D(CLBLL_L_X4Y92_SLICE_X4Y92_AO6),
.Q(CLBLL_L_X2Y91_SLICE_X0Y91_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y91_SLICE_X0Y91_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y91_SLICE_X0Y91_DO5),
.O6(CLBLL_L_X2Y91_SLICE_X0Y91_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y91_SLICE_X0Y91_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y91_SLICE_X0Y91_CO5),
.O6(CLBLL_L_X2Y91_SLICE_X0Y91_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y91_SLICE_X0Y91_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y91_SLICE_X0Y91_BO5),
.O6(CLBLL_L_X2Y91_SLICE_X0Y91_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y91_SLICE_X0Y91_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y91_SLICE_X0Y91_AO5),
.O6(CLBLL_L_X2Y91_SLICE_X0Y91_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y91_SLICE_X1Y91_A_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLL_L_X2Y93_SLICE_X1Y93_CO6),
.D(CLBLM_R_X3Y94_SLICE_X2Y94_DO6),
.Q(CLBLL_L_X2Y91_SLICE_X1Y91_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y91_SLICE_X1Y91_B_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLL_L_X2Y93_SLICE_X1Y93_CO6),
.D(CLBLL_L_X4Y92_SLICE_X4Y92_AO6),
.Q(CLBLL_L_X2Y91_SLICE_X1Y91_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y91_SLICE_X1Y91_C_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLL_L_X2Y93_SLICE_X1Y93_CO6),
.D(CLBLL_L_X4Y94_SLICE_X4Y94_CO5),
.Q(CLBLL_L_X2Y91_SLICE_X1Y91_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y91_SLICE_X1Y91_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y91_SLICE_X1Y91_DO5),
.O6(CLBLL_L_X2Y91_SLICE_X1Y91_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y91_SLICE_X1Y91_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y91_SLICE_X1Y91_CO5),
.O6(CLBLL_L_X2Y91_SLICE_X1Y91_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y91_SLICE_X1Y91_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y91_SLICE_X1Y91_BO5),
.O6(CLBLL_L_X2Y91_SLICE_X1Y91_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y91_SLICE_X1Y91_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y91_SLICE_X1Y91_AO5),
.O6(CLBLL_L_X2Y91_SLICE_X1Y91_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y92_SLICE_X0Y92_A_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLL_L_X2Y93_SLICE_X0Y93_DO6),
.D(CLBLL_L_X4Y94_SLICE_X4Y94_CO5),
.Q(CLBLL_L_X2Y92_SLICE_X0Y92_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y92_SLICE_X0Y92_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y92_SLICE_X0Y92_DO5),
.O6(CLBLL_L_X2Y92_SLICE_X0Y92_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y92_SLICE_X0Y92_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y92_SLICE_X0Y92_CO5),
.O6(CLBLL_L_X2Y92_SLICE_X0Y92_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y92_SLICE_X0Y92_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y92_SLICE_X0Y92_BO5),
.O6(CLBLL_L_X2Y92_SLICE_X0Y92_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y92_SLICE_X0Y92_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y92_SLICE_X0Y92_AO5),
.O6(CLBLL_L_X2Y92_SLICE_X0Y92_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y92_SLICE_X1Y92_A_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLL_L_X4Y92_SLICE_X4Y92_BO6),
.D(CLBLM_R_X3Y94_SLICE_X2Y94_DO6),
.Q(CLBLL_L_X2Y92_SLICE_X1Y92_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y92_SLICE_X1Y92_B_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLL_L_X4Y92_SLICE_X4Y92_BO6),
.D(CLBLL_L_X4Y92_SLICE_X4Y92_AO6),
.Q(CLBLL_L_X2Y92_SLICE_X1Y92_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y92_SLICE_X1Y92_C_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLL_L_X4Y92_SLICE_X4Y92_BO6),
.D(CLBLL_L_X4Y94_SLICE_X4Y94_CO5),
.Q(CLBLL_L_X2Y92_SLICE_X1Y92_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y92_SLICE_X1Y92_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y92_SLICE_X1Y92_DO5),
.O6(CLBLL_L_X2Y92_SLICE_X1Y92_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y92_SLICE_X1Y92_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y92_SLICE_X1Y92_CO5),
.O6(CLBLL_L_X2Y92_SLICE_X1Y92_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y92_SLICE_X1Y92_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y92_SLICE_X1Y92_BO5),
.O6(CLBLL_L_X2Y92_SLICE_X1Y92_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000550000000000)
  ) CLBLL_L_X2Y92_SLICE_X1Y92_ALUT (
.I0(CLBLM_R_X5Y94_SLICE_X7Y94_DO6),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X5Y94_SLICE_X6Y94_BO6),
.I4(CLBLL_L_X4Y94_SLICE_X5Y94_DO6),
.I5(CLBLL_L_X2Y93_SLICE_X0Y93_CO6),
.O5(CLBLL_L_X2Y92_SLICE_X1Y92_AO5),
.O6(CLBLL_L_X2Y92_SLICE_X1Y92_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y93_SLICE_X0Y93_B_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLL_L_X2Y93_SLICE_X0Y93_DO6),
.D(CLBLM_R_X3Y94_SLICE_X2Y94_DO6),
.Q(CLBLL_L_X2Y93_SLICE_X0Y93_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y93_SLICE_X0Y93_C_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLL_L_X2Y93_SLICE_X0Y93_DO6),
.D(CLBLM_R_X3Y94_SLICE_X2Y94_DO5),
.Q(CLBLL_L_X2Y93_SLICE_X0Y93_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3000000030000000)
  ) CLBLL_L_X2Y93_SLICE_X0Y93_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y94_SLICE_X7Y94_DO6),
.I2(CLBLL_L_X4Y94_SLICE_X5Y94_DO6),
.I3(CLBLL_L_X2Y93_SLICE_X0Y93_CO6),
.I4(CLBLM_R_X5Y94_SLICE_X6Y94_BO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y93_SLICE_X0Y93_DO5),
.O6(CLBLL_L_X2Y93_SLICE_X0Y93_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a740b5c7fdff7af)
  ) CLBLL_L_X2Y93_SLICE_X0Y93_CLUT (
.I0(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I1(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I2(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I3(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I4(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y93_SLICE_X0Y93_CO5),
.O6(CLBLL_L_X2Y93_SLICE_X0Y93_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0edc0ec00010000)
  ) CLBLL_L_X2Y93_SLICE_X0Y93_BLUT (
.I0(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I1(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I2(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I3(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I4(CLBLM_R_X3Y93_SLICE_X2Y93_DO6),
.I5(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO10),
.O5(CLBLL_L_X2Y93_SLICE_X0Y93_BO5),
.O6(CLBLL_L_X2Y93_SLICE_X0Y93_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f005f0000000f00)
  ) CLBLL_L_X2Y93_SLICE_X0Y93_ALUT (
.I0(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I3(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO10),
.I4(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I5(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.O5(CLBLL_L_X2Y93_SLICE_X0Y93_AO5),
.O6(CLBLL_L_X2Y93_SLICE_X0Y93_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_L_X2Y93_SLICE_X0Y93_MUXF7A (
.I0(CLBLL_L_X2Y93_SLICE_X0Y93_BO6),
.I1(CLBLL_L_X2Y93_SLICE_X0Y93_AO6),
.O(CLBLL_L_X2Y93_SLICE_X0Y93_F7AMUX_O),
.S(CLBLL_L_X4Y91_SLICE_X5Y91_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y93_SLICE_X1Y93_B_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLL_L_X2Y93_SLICE_X1Y93_DO6),
.D(CLBLM_R_X3Y94_SLICE_X2Y94_DO6),
.Q(CLBLL_L_X2Y93_SLICE_X1Y93_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0000000c0000000)
  ) CLBLL_L_X2Y93_SLICE_X1Y93_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X2Y93_SLICE_X0Y93_CO6),
.I2(CLBLM_R_X5Y94_SLICE_X6Y94_BO6),
.I3(CLBLM_R_X5Y94_SLICE_X7Y94_DO6),
.I4(CLBLL_L_X4Y94_SLICE_X5Y94_DO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y93_SLICE_X1Y93_DO5),
.O6(CLBLL_L_X2Y93_SLICE_X1Y93_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000c0000000c000)
  ) CLBLL_L_X2Y93_SLICE_X1Y93_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X2Y93_SLICE_X0Y93_CO6),
.I2(CLBLM_R_X5Y94_SLICE_X6Y94_BO6),
.I3(CLBLM_R_X5Y94_SLICE_X7Y94_DO6),
.I4(CLBLL_L_X4Y94_SLICE_X5Y94_DO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y93_SLICE_X1Y93_CO5),
.O6(CLBLL_L_X2Y93_SLICE_X1Y93_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e2e2e2ff33cc00)
  ) CLBLL_L_X2Y93_SLICE_X1Y93_BLUT (
.I0(CLBLL_L_X2Y94_SLICE_X1Y94_BQ),
.I1(CLBLL_L_X4Y91_SLICE_X5Y91_F7AMUX_O),
.I2(CLBLL_L_X2Y91_SLICE_X1Y91_AQ),
.I3(CLBLL_L_X2Y92_SLICE_X1Y92_AQ),
.I4(CLBLM_R_X3Y94_SLICE_X2Y94_AQ),
.I5(CLBLM_R_X5Y93_SLICE_X6Y93_F7AMUX_O),
.O5(CLBLL_L_X2Y93_SLICE_X1Y93_BO5),
.O6(CLBLL_L_X2Y93_SLICE_X1Y93_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfd58f85dad08a80)
  ) CLBLL_L_X2Y93_SLICE_X1Y93_ALUT (
.I0(CLBLM_R_X5Y93_SLICE_X6Y93_F7AMUX_O),
.I1(CLBLL_L_X2Y93_SLICE_X1Y93_BQ),
.I2(CLBLL_L_X4Y91_SLICE_X5Y91_F7AMUX_O),
.I3(CLBLL_L_X2Y93_SLICE_X0Y93_BQ),
.I4(CLBLM_R_X3Y92_SLICE_X2Y92_BQ),
.I5(CLBLM_R_X3Y93_SLICE_X2Y93_BQ),
.O5(CLBLL_L_X2Y93_SLICE_X1Y93_AO5),
.O6(CLBLL_L_X2Y93_SLICE_X1Y93_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_L_X2Y93_SLICE_X1Y93_MUXF7A (
.I0(CLBLL_L_X2Y93_SLICE_X1Y93_BO6),
.I1(CLBLL_L_X2Y93_SLICE_X1Y93_AO6),
.O(CLBLL_L_X2Y93_SLICE_X1Y93_F7AMUX_O),
.S(CLBLL_L_X2Y93_SLICE_X0Y93_F7AMUX_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0ffffffaffaff)
  ) CLBLL_L_X2Y94_SLICE_X0Y94_DLUT (
.I0(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I3(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I4(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I5(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.O5(CLBLL_L_X2Y94_SLICE_X0Y94_DO5),
.O6(CLBLL_L_X2Y94_SLICE_X0Y94_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5e4a2d5e4a0e691)
  ) CLBLL_L_X2Y94_SLICE_X0Y94_CLUT (
.I0(CLBLL_L_X2Y93_SLICE_X0Y93_CO5),
.I1(CLBLM_R_X3Y93_SLICE_X2Y93_CO5),
.I2(CLBLL_L_X2Y94_SLICE_X1Y94_B_XOR),
.I3(CLBLL_L_X2Y93_SLICE_X1Y93_F7AMUX_O),
.I4(CLBLL_L_X2Y97_SLICE_X0Y97_AO6),
.I5(CLBLL_L_X4Y95_SLICE_X4Y95_CO6),
.O5(CLBLL_L_X2Y94_SLICE_X0Y94_CO5),
.O6(CLBLL_L_X2Y94_SLICE_X0Y94_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff2f9fff9df)
  ) CLBLL_L_X2Y94_SLICE_X0Y94_BLUT (
.I0(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I1(CLBLL_L_X4Y95_SLICE_X4Y95_CO6),
.I2(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I3(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I4(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I5(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.O5(CLBLL_L_X2Y94_SLICE_X0Y94_BO5),
.O6(CLBLL_L_X2Y94_SLICE_X0Y94_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffedffedffffcef7)
  ) CLBLL_L_X2Y94_SLICE_X0Y94_ALUT (
.I0(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I1(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I2(CLBLL_L_X4Y95_SLICE_X4Y95_BO6),
.I3(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I4(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I5(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.O5(CLBLL_L_X2Y94_SLICE_X0Y94_AO5),
.O6(CLBLL_L_X2Y94_SLICE_X0Y94_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y94_SLICE_X1Y94_B_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLL_L_X2Y92_SLICE_X1Y92_AO6),
.D(CLBLL_L_X2Y94_SLICE_X1Y94_BO5),
.Q(CLBLL_L_X2Y94_SLICE_X1Y94_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y94_SLICE_X1Y94_C_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLL_L_X2Y92_SLICE_X1Y92_AO6),
.D(CLBLL_L_X2Y94_SLICE_X1Y94_CO5),
.Q(CLBLL_L_X2Y94_SLICE_X1Y94_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y94_SLICE_X1Y94_D_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLL_L_X2Y92_SLICE_X1Y92_AO6),
.D(CLBLL_L_X2Y94_SLICE_X1Y94_DO5),
.Q(CLBLL_L_X2Y94_SLICE_X1Y94_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_L_X2Y94_SLICE_X1Y94_CARRY4 (
.CI(1'b0),
.CO({CLBLL_L_X2Y94_SLICE_X1Y94_D_CY, CLBLL_L_X2Y94_SLICE_X1Y94_C_CY, CLBLL_L_X2Y94_SLICE_X1Y94_B_CY, CLBLL_L_X2Y94_SLICE_X1Y94_A_CY}),
.CYINIT(CLBLL_L_X4Y93_SLICE_X4Y93_DO6),
.DI({CLBLL_L_X2Y94_SLICE_X0Y94_AO6, CLBLM_R_X3Y93_SLICE_X3Y93_AO6, CLBLL_L_X2Y94_SLICE_X0Y94_BO6, CLBLL_L_X2Y94_SLICE_X1Y94_AO5}),
.O({CLBLL_L_X2Y94_SLICE_X1Y94_D_XOR, CLBLL_L_X2Y94_SLICE_X1Y94_C_XOR, CLBLL_L_X2Y94_SLICE_X1Y94_B_XOR, CLBLL_L_X2Y94_SLICE_X1Y94_A_XOR}),
.S({CLBLL_L_X2Y94_SLICE_X1Y94_DO6, CLBLL_L_X2Y94_SLICE_X1Y94_CO6, CLBLL_L_X2Y94_SLICE_X1Y94_BO6, CLBLL_L_X2Y94_SLICE_X1Y94_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc030cf3aaaaaaaa)
  ) CLBLL_L_X2Y94_SLICE_X1Y94_DLUT (
.I0(CLBLL_L_X4Y94_SLICE_X4Y94_CO5),
.I1(CLBLL_L_X2Y97_SLICE_X0Y97_AO6),
.I2(CLBLL_L_X4Y95_SLICE_X4Y95_BO6),
.I3(CLBLL_L_X4Y93_SLICE_X4Y93_F7AMUX_O),
.I4(CLBLM_R_X3Y93_SLICE_X2Y93_CO5),
.I5(1'b1),
.O5(CLBLL_L_X2Y94_SLICE_X1Y94_DO5),
.O6(CLBLL_L_X2Y94_SLICE_X1Y94_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccc33c33aaaaaaaa)
  ) CLBLL_L_X2Y94_SLICE_X1Y94_CLUT (
.I0(CLBLM_R_X3Y94_SLICE_X2Y94_DO5),
.I1(CLBLM_R_X3Y94_SLICE_X3Y94_F7AMUX_O),
.I2(CLBLM_R_X3Y95_SLICE_X3Y95_DO6),
.I3(CLBLL_L_X2Y97_SLICE_X0Y97_AO6),
.I4(CLBLM_R_X3Y93_SLICE_X2Y93_CO5),
.I5(1'b1),
.O5(CLBLL_L_X2Y94_SLICE_X1Y94_CO5),
.O6(CLBLL_L_X2Y94_SLICE_X1Y94_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0cc0f33aaaaaaaa)
  ) CLBLL_L_X2Y94_SLICE_X1Y94_BLUT (
.I0(CLBLM_R_X3Y94_SLICE_X2Y94_DO6),
.I1(CLBLL_L_X2Y97_SLICE_X0Y97_AO6),
.I2(CLBLM_R_X3Y93_SLICE_X2Y93_CO5),
.I3(CLBLL_L_X4Y95_SLICE_X4Y95_CO6),
.I4(CLBLL_L_X2Y93_SLICE_X1Y93_F7AMUX_O),
.I5(1'b1),
.O5(CLBLL_L_X2Y94_SLICE_X1Y94_BO5),
.O6(CLBLL_L_X2Y94_SLICE_X1Y94_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000cccccccc)
  ) CLBLL_L_X2Y94_SLICE_X1Y94_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X2Y94_SLICE_X0Y94_DO6),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X2Y96_SLICE_X0Y96_AO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y94_SLICE_X1Y94_AO5),
.O6(CLBLL_L_X2Y94_SLICE_X1Y94_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_L_X2Y95_SLICE_X0Y95_CARRY4 (
.CI(1'b0),
.CO({CLBLL_L_X2Y95_SLICE_X0Y95_D_CY, CLBLL_L_X2Y95_SLICE_X0Y95_C_CY, CLBLL_L_X2Y95_SLICE_X0Y95_B_CY, CLBLL_L_X2Y95_SLICE_X0Y95_A_CY}),
.CYINIT(1'b0),
.DI({CLBLL_L_X2Y95_SLICE_X0Y95_DO5, CLBLL_L_X2Y95_SLICE_X0Y95_CO5, CLBLL_L_X2Y95_SLICE_X0Y95_BO5, CLBLL_L_X2Y95_SLICE_X0Y95_AO5}),
.O({CLBLL_L_X2Y95_SLICE_X0Y95_D_XOR, CLBLL_L_X2Y95_SLICE_X0Y95_C_XOR, CLBLL_L_X2Y95_SLICE_X0Y95_B_XOR, CLBLL_L_X2Y95_SLICE_X0Y95_A_XOR}),
.S({CLBLL_L_X2Y95_SLICE_X0Y95_DO6, CLBLL_L_X2Y95_SLICE_X0Y95_CO6, CLBLL_L_X2Y95_SLICE_X0Y95_BO6, CLBLL_L_X2Y95_SLICE_X0Y95_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc00c300300c0ccfc)
  ) CLBLL_L_X2Y95_SLICE_X0Y95_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y95_SLICE_X3Y95_BO6),
.I2(CLBLL_L_X4Y95_SLICE_X5Y95_CO6),
.I3(CLBLL_L_X4Y94_SLICE_X5Y94_F7AMUX_O),
.I4(CLBLM_R_X3Y92_SLICE_X2Y92_F7AMUX_O),
.I5(1'b1),
.O5(CLBLL_L_X2Y95_SLICE_X0Y95_DO5),
.O6(CLBLL_L_X2Y95_SLICE_X0Y95_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h842184212b0a2b0a)
  ) CLBLL_L_X2Y95_SLICE_X0Y95_CLUT (
.I0(CLBLL_L_X4Y91_SLICE_X4Y91_BO6),
.I1(CLBLM_R_X3Y91_SLICE_X2Y91_F7AMUX_O),
.I2(CLBLM_R_X3Y91_SLICE_X3Y91_F7AMUX_O),
.I3(CLBLM_R_X3Y95_SLICE_X3Y95_AO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y95_SLICE_X0Y95_CO5),
.O6(CLBLL_L_X2Y95_SLICE_X0Y95_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9900009922ff0022)
  ) CLBLL_L_X2Y95_SLICE_X0Y95_BLUT (
.I0(CLBLM_R_X3Y95_SLICE_X3Y95_DO6),
.I1(CLBLM_R_X3Y94_SLICE_X3Y94_F7AMUX_O),
.I2(1'b1),
.I3(CLBLL_L_X4Y93_SLICE_X4Y93_F7AMUX_O),
.I4(CLBLL_L_X4Y95_SLICE_X4Y95_BO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y95_SLICE_X0Y95_BO5),
.O6(CLBLL_L_X2Y95_SLICE_X0Y95_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h882244113300bb22)
  ) CLBLL_L_X2Y95_SLICE_X0Y95_ALUT (
.I0(CLBLL_L_X4Y95_SLICE_X4Y95_DO6),
.I1(CLBLL_L_X2Y93_SLICE_X1Y93_F7AMUX_O),
.I2(1'b1),
.I3(CLBLL_L_X4Y95_SLICE_X4Y95_CO6),
.I4(CLBLL_L_X4Y93_SLICE_X4Y93_DO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y95_SLICE_X0Y95_AO5),
.O6(CLBLL_L_X2Y95_SLICE_X0Y95_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_L_X2Y95_SLICE_X1Y95_CARRY4 (
.CI(CLBLL_L_X2Y94_SLICE_X1Y94_D_CY),
.CO({CLBLL_L_X2Y95_SLICE_X1Y95_D_CY, CLBLL_L_X2Y95_SLICE_X1Y95_C_CY, CLBLL_L_X2Y95_SLICE_X1Y95_B_CY, CLBLL_L_X2Y95_SLICE_X1Y95_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, CLBLL_L_X4Y95_SLICE_X4Y95_AO6, CLBLM_R_X3Y95_SLICE_X2Y95_AO6, CLBLM_R_X3Y95_SLICE_X3Y95_CO6}),
.O({CLBLL_L_X2Y95_SLICE_X1Y95_D_XOR, CLBLL_L_X2Y95_SLICE_X1Y95_C_XOR, CLBLL_L_X2Y95_SLICE_X1Y95_B_XOR, CLBLL_L_X2Y95_SLICE_X1Y95_A_XOR}),
.S({CLBLL_L_X2Y95_SLICE_X1Y95_DO6, CLBLL_L_X2Y95_SLICE_X1Y95_CO6, CLBLL_L_X2Y95_SLICE_X1Y95_BO6, CLBLL_L_X2Y95_SLICE_X1Y95_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3c0f3c00c3f0c3f)
  ) CLBLL_L_X2Y95_SLICE_X1Y95_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y95_SLICE_X3Y95_BO6),
.I2(CLBLM_R_X3Y93_SLICE_X2Y93_CO5),
.I3(CLBLL_L_X2Y97_SLICE_X0Y97_AO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y92_SLICE_X2Y92_F7AMUX_O),
.O5(CLBLL_L_X2Y95_SLICE_X1Y95_DO5),
.O6(CLBLL_L_X2Y95_SLICE_X1Y95_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc399c399c399c399)
  ) CLBLL_L_X2Y95_SLICE_X1Y95_CLUT (
.I0(CLBLL_L_X2Y97_SLICE_X0Y97_AO6),
.I1(CLBLL_L_X4Y94_SLICE_X5Y94_F7AMUX_O),
.I2(CLBLM_R_X3Y93_SLICE_X2Y93_CO5),
.I3(CLBLL_L_X4Y95_SLICE_X5Y95_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y95_SLICE_X1Y95_CO5),
.O6(CLBLL_L_X2Y95_SLICE_X1Y95_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9a9a95959a9a9595)
  ) CLBLL_L_X2Y95_SLICE_X1Y95_BLUT (
.I0(CLBLM_R_X3Y91_SLICE_X3Y91_F7AMUX_O),
.I1(CLBLM_R_X3Y93_SLICE_X2Y93_CO5),
.I2(CLBLL_L_X4Y91_SLICE_X4Y91_BO6),
.I3(1'b1),
.I4(CLBLL_L_X2Y97_SLICE_X0Y97_AO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y95_SLICE_X1Y95_BO5),
.O6(CLBLL_L_X2Y95_SLICE_X1Y95_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcf30c03fcf30c03f)
  ) CLBLL_L_X2Y95_SLICE_X1Y95_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y93_SLICE_X2Y93_CO5),
.I2(CLBLM_R_X3Y95_SLICE_X3Y95_AO6),
.I3(CLBLM_R_X3Y91_SLICE_X2Y91_F7AMUX_O),
.I4(CLBLL_L_X2Y97_SLICE_X0Y97_AO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y95_SLICE_X1Y95_AO5),
.O6(CLBLL_L_X2Y95_SLICE_X1Y95_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbf80b58fca50c05)
  ) CLBLL_L_X2Y96_SLICE_X0Y96_DLUT (
.I0(CLBLL_L_X2Y97_SLICE_X0Y97_AO6),
.I1(CLBLM_R_X3Y95_SLICE_X3Y95_DO6),
.I2(CLBLL_L_X2Y93_SLICE_X0Y93_CO5),
.I3(CLBLM_R_X3Y93_SLICE_X2Y93_CO5),
.I4(CLBLL_L_X2Y94_SLICE_X1Y94_C_XOR),
.I5(CLBLM_R_X3Y94_SLICE_X3Y94_F7AMUX_O),
.O5(CLBLL_L_X2Y96_SLICE_X0Y96_DO5),
.O6(CLBLL_L_X2Y96_SLICE_X0Y96_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeecdec3322012c3)
  ) CLBLL_L_X2Y96_SLICE_X0Y96_CLUT (
.I0(CLBLL_L_X4Y95_SLICE_X4Y95_DO6),
.I1(CLBLL_L_X2Y93_SLICE_X0Y93_CO5),
.I2(CLBLL_L_X4Y93_SLICE_X4Y93_DO6),
.I3(CLBLM_R_X3Y93_SLICE_X2Y93_CO5),
.I4(CLBLL_L_X2Y97_SLICE_X0Y97_AO6),
.I5(CLBLL_L_X2Y94_SLICE_X1Y94_A_XOR),
.O5(CLBLL_L_X2Y96_SLICE_X0Y96_CO5),
.O6(CLBLL_L_X2Y96_SLICE_X0Y96_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfebe5414ea994099)
  ) CLBLL_L_X2Y96_SLICE_X0Y96_BLUT (
.I0(CLBLL_L_X2Y93_SLICE_X0Y93_CO5),
.I1(CLBLM_R_X3Y92_SLICE_X2Y92_F7AMUX_O),
.I2(CLBLM_R_X3Y95_SLICE_X3Y95_BO6),
.I3(CLBLL_L_X2Y97_SLICE_X0Y97_AO6),
.I4(CLBLL_L_X2Y95_SLICE_X1Y95_D_XOR),
.I5(CLBLM_R_X3Y93_SLICE_X2Y93_CO5),
.O5(CLBLL_L_X2Y96_SLICE_X0Y96_BO5),
.O6(CLBLL_L_X2Y96_SLICE_X0Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffcebfffffcff)
  ) CLBLL_L_X2Y96_SLICE_X0Y96_ALUT (
.I0(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I1(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I2(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I3(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I4(CLBLL_L_X4Y95_SLICE_X4Y95_DO6),
.I5(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.O5(CLBLL_L_X2Y96_SLICE_X0Y96_AO5),
.O6(CLBLL_L_X2Y96_SLICE_X0Y96_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd4d4d4d4aa882200)
  ) CLBLL_L_X2Y96_SLICE_X1Y96_DLUT (
.I0(CLBLM_R_X3Y96_SLICE_X3Y96_BO5),
.I1(CLBLM_R_X3Y96_SLICE_X3Y96_BO6),
.I2(CLBLL_L_X2Y96_SLICE_X0Y96_BO6),
.I3(CLBLL_L_X2Y96_SLICE_X1Y96_CO6),
.I4(CLBLL_L_X2Y96_SLICE_X0Y96_CO6),
.I5(CLBLL_L_X2Y97_SLICE_X0Y97_AO5),
.O5(CLBLL_L_X2Y96_SLICE_X1Y96_DO5),
.O6(CLBLL_L_X2Y96_SLICE_X1Y96_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf3ccafa0c00f)
  ) CLBLL_L_X2Y96_SLICE_X1Y96_CLUT (
.I0(CLBLL_L_X2Y95_SLICE_X1Y95_C_XOR),
.I1(CLBLL_L_X4Y95_SLICE_X5Y95_CO6),
.I2(CLBLL_L_X2Y97_SLICE_X0Y97_AO6),
.I3(CLBLL_L_X4Y94_SLICE_X5Y94_F7AMUX_O),
.I4(CLBLL_L_X2Y93_SLICE_X0Y93_CO5),
.I5(CLBLM_R_X3Y93_SLICE_X2Y93_CO5),
.O5(CLBLL_L_X2Y96_SLICE_X1Y96_CO5),
.O6(CLBLL_L_X2Y96_SLICE_X1Y96_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5ff5088a0005088)
  ) CLBLL_L_X2Y96_SLICE_X1Y96_BLUT (
.I0(CLBLM_R_X3Y96_SLICE_X3Y96_BO5),
.I1(CLBLM_R_X3Y95_SLICE_X2Y95_CO6),
.I2(CLBLM_R_X3Y95_SLICE_X2Y95_DO6),
.I3(CLBLL_L_X2Y97_SLICE_X0Y97_AO5),
.I4(CLBLM_R_X3Y96_SLICE_X3Y96_BO6),
.I5(CLBLL_L_X2Y96_SLICE_X1Y96_CO6),
.O5(CLBLL_L_X2Y96_SLICE_X1Y96_BO5),
.O6(CLBLL_L_X2Y96_SLICE_X1Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8f0f04444aa00)
  ) CLBLL_L_X2Y96_SLICE_X1Y96_ALUT (
.I0(CLBLM_R_X3Y96_SLICE_X3Y96_BO5),
.I1(CLBLM_R_X3Y95_SLICE_X2Y95_CO6),
.I2(CLBLM_R_X3Y95_SLICE_X2Y95_DO6),
.I3(CLBLM_R_X3Y95_SLICE_X2Y95_BO6),
.I4(CLBLL_L_X2Y97_SLICE_X0Y97_AO5),
.I5(CLBLM_R_X3Y96_SLICE_X3Y96_BO6),
.O5(CLBLL_L_X2Y96_SLICE_X1Y96_AO5),
.O6(CLBLL_L_X2Y96_SLICE_X1Y96_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffeeffee)
  ) CLBLL_L_X2Y97_SLICE_X0Y97_DLUT (
.I0(CLBLL_L_X2Y94_SLICE_X0Y94_CO6),
.I1(CLBLL_L_X2Y96_SLICE_X0Y96_CO6),
.I2(1'b1),
.I3(CLBLL_L_X2Y96_SLICE_X0Y96_DO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y95_SLICE_X2Y95_BO6),
.O5(CLBLL_L_X2Y97_SLICE_X0Y97_DO5),
.O6(CLBLL_L_X2Y97_SLICE_X0Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff5f4a40a0004a40)
  ) CLBLL_L_X2Y97_SLICE_X0Y97_CLUT (
.I0(CLBLL_L_X2Y97_SLICE_X0Y97_AO5),
.I1(CLBLL_L_X2Y94_SLICE_X0Y94_CO6),
.I2(CLBLM_R_X3Y96_SLICE_X3Y96_BO5),
.I3(CLBLL_L_X2Y96_SLICE_X0Y96_DO6),
.I4(CLBLM_R_X3Y96_SLICE_X3Y96_BO6),
.I5(CLBLM_R_X3Y95_SLICE_X2Y95_BO6),
.O5(CLBLL_L_X2Y97_SLICE_X0Y97_CO5),
.O6(CLBLL_L_X2Y97_SLICE_X0Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbe2e2f3c0c0c0)
  ) CLBLL_L_X2Y97_SLICE_X0Y97_BLUT (
.I0(CLBLL_L_X2Y96_SLICE_X0Y96_CO6),
.I1(CLBLM_R_X3Y96_SLICE_X3Y96_BO6),
.I2(CLBLL_L_X2Y94_SLICE_X0Y94_CO6),
.I3(CLBLL_L_X2Y96_SLICE_X0Y96_BO6),
.I4(CLBLM_R_X3Y96_SLICE_X3Y96_BO5),
.I5(CLBLL_L_X2Y97_SLICE_X0Y97_AO5),
.O5(CLBLL_L_X2Y97_SLICE_X0Y97_BO5),
.O6(CLBLL_L_X2Y97_SLICE_X0Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0001202873fbbfff)
  ) CLBLL_L_X2Y97_SLICE_X0Y97_ALUT (
.I0(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I1(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I2(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I3(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I4(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y97_SLICE_X0Y97_AO5),
.O6(CLBLL_L_X2Y97_SLICE_X0Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000300000003)
  ) CLBLL_L_X2Y97_SLICE_X1Y97_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y95_SLICE_X2Y95_CO6),
.I2(CLBLL_L_X2Y96_SLICE_X0Y96_BO6),
.I3(CLBLL_L_X2Y96_SLICE_X1Y96_CO6),
.I4(CLBLM_R_X3Y95_SLICE_X2Y95_DO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y97_SLICE_X1Y97_DO5),
.O6(CLBLL_L_X2Y97_SLICE_X1Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h88e488e4f5a0a0a0)
  ) CLBLL_L_X2Y97_SLICE_X1Y97_CLUT (
.I0(CLBLM_R_X3Y96_SLICE_X3Y96_BO6),
.I1(CLBLL_L_X2Y96_SLICE_X1Y96_CO6),
.I2(CLBLL_L_X2Y96_SLICE_X0Y96_BO6),
.I3(CLBLM_R_X3Y96_SLICE_X3Y96_BO5),
.I4(CLBLM_R_X3Y95_SLICE_X2Y95_DO6),
.I5(CLBLL_L_X2Y97_SLICE_X0Y97_AO5),
.O5(CLBLL_L_X2Y97_SLICE_X1Y97_CO5),
.O6(CLBLL_L_X2Y97_SLICE_X1Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa058585f000808)
  ) CLBLL_L_X2Y97_SLICE_X1Y97_BLUT (
.I0(CLBLM_R_X3Y96_SLICE_X3Y96_BO5),
.I1(CLBLL_L_X2Y96_SLICE_X0Y96_DO6),
.I2(CLBLL_L_X2Y97_SLICE_X0Y97_AO5),
.I3(CLBLM_R_X3Y95_SLICE_X2Y95_CO6),
.I4(CLBLM_R_X3Y96_SLICE_X3Y96_BO6),
.I5(CLBLM_R_X3Y95_SLICE_X2Y95_BO6),
.O5(CLBLL_L_X2Y97_SLICE_X1Y97_BO5),
.O6(CLBLL_L_X2Y97_SLICE_X1Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0a0c0accf0cc00)
  ) CLBLL_L_X2Y97_SLICE_X1Y97_ALUT (
.I0(CLBLL_L_X2Y96_SLICE_X0Y96_CO6),
.I1(CLBLL_L_X2Y96_SLICE_X0Y96_DO6),
.I2(CLBLL_L_X2Y97_SLICE_X0Y97_AO5),
.I3(CLBLM_R_X3Y96_SLICE_X3Y96_BO6),
.I4(CLBLL_L_X2Y94_SLICE_X0Y94_CO6),
.I5(CLBLM_R_X3Y96_SLICE_X3Y96_BO5),
.O5(CLBLL_L_X2Y97_SLICE_X1Y97_AO5),
.O6(CLBLL_L_X2Y97_SLICE_X1Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y98_SLICE_X0Y98_A_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(LIOB33_X0Y105_IOB_X0Y105_I),
.D(LIOB33_X0Y105_IOB_X0Y105_I),
.Q(CLBLL_L_X2Y98_SLICE_X0Y98_AQ),
.R(CLBLL_L_X2Y98_SLICE_X1Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y98_SLICE_X0Y98_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y98_SLICE_X0Y98_DO5),
.O6(CLBLL_L_X2Y98_SLICE_X0Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y98_SLICE_X0Y98_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y98_SLICE_X0Y98_CO5),
.O6(CLBLL_L_X2Y98_SLICE_X0Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y98_SLICE_X0Y98_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y98_SLICE_X0Y98_BO5),
.O6(CLBLL_L_X2Y98_SLICE_X0Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y98_SLICE_X0Y98_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y98_SLICE_X0Y98_AO5),
.O6(CLBLL_L_X2Y98_SLICE_X0Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y98_SLICE_X1Y98_A_FDCE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(1'b1),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLL_L_X2Y98_SLICE_X1Y98_AO6),
.Q(CLBLL_L_X2Y98_SLICE_X1Y98_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y98_SLICE_X1Y98_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y98_SLICE_X1Y98_DO5),
.O6(CLBLL_L_X2Y98_SLICE_X1Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y98_SLICE_X1Y98_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y98_SLICE_X1Y98_CO5),
.O6(CLBLL_L_X2Y98_SLICE_X1Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff0f0fffff0f0)
  ) CLBLL_L_X2Y98_SLICE_X1Y98_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X2Y98_SLICE_X1Y98_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y98_SLICE_X1Y98_BO5),
.O6(CLBLL_L_X2Y98_SLICE_X1Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0f0d8f0f0)
  ) CLBLL_L_X2Y98_SLICE_X1Y98_ALUT (
.I0(CLBLM_R_X3Y98_SLICE_X3Y98_AO6),
.I1(CLBLL_L_X2Y97_SLICE_X0Y97_BO6),
.I2(CLBLL_L_X2Y98_SLICE_X1Y98_AQ),
.I3(CLBLL_L_X4Y97_SLICE_X4Y97_CO6),
.I4(CLBLM_R_X5Y94_SLICE_X6Y94_CO6),
.I5(CLBLL_L_X4Y98_SLICE_X4Y98_AO6),
.O5(CLBLL_L_X2Y98_SLICE_X1Y98_AO5),
.O6(CLBLL_L_X2Y98_SLICE_X1Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y99_SLICE_X0Y99_A_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(LIOB33_X0Y107_IOB_X0Y108_I),
.D(LIOB33_X0Y107_IOB_X0Y108_I),
.Q(CLBLL_L_X2Y99_SLICE_X0Y99_AQ),
.R(CLBLL_L_X2Y98_SLICE_X1Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y99_SLICE_X0Y99_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y99_SLICE_X0Y99_DO5),
.O6(CLBLL_L_X2Y99_SLICE_X0Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y99_SLICE_X0Y99_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y99_SLICE_X0Y99_CO5),
.O6(CLBLL_L_X2Y99_SLICE_X0Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y99_SLICE_X0Y99_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y99_SLICE_X0Y99_BO5),
.O6(CLBLL_L_X2Y99_SLICE_X0Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y99_SLICE_X0Y99_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y99_SLICE_X0Y99_AO5),
.O6(CLBLL_L_X2Y99_SLICE_X0Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y99_SLICE_X1Y99_A_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLL_L_X2Y99_SLICE_X1Y99_AQ),
.R(CLBLL_L_X2Y98_SLICE_X1Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y99_SLICE_X1Y99_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y99_SLICE_X1Y99_DO5),
.O6(CLBLL_L_X2Y99_SLICE_X1Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y99_SLICE_X1Y99_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y99_SLICE_X1Y99_CO5),
.O6(CLBLL_L_X2Y99_SLICE_X1Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y99_SLICE_X1Y99_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y99_SLICE_X1Y99_BO5),
.O6(CLBLL_L_X2Y99_SLICE_X1Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y99_SLICE_X1Y99_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y99_SLICE_X1Y99_AO5),
.O6(CLBLL_L_X2Y99_SLICE_X1Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y102_SLICE_X0Y102_A_FDPE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(1'b1),
.D(CLBLM_R_X7Y90_SLICE_X8Y90_BQ),
.PRE(LIOB33_X0Y107_IOB_X0Y107_I),
.Q(CLBLL_L_X2Y102_SLICE_X0Y102_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y102_SLICE_X0Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y102_SLICE_X0Y102_DO5),
.O6(CLBLL_L_X2Y102_SLICE_X0Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y102_SLICE_X0Y102_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y102_SLICE_X0Y102_CO5),
.O6(CLBLL_L_X2Y102_SLICE_X0Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y102_SLICE_X0Y102_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y102_SLICE_X0Y102_BO5),
.O6(CLBLL_L_X2Y102_SLICE_X0Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y102_SLICE_X0Y102_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y102_SLICE_X0Y102_AO5),
.O6(CLBLL_L_X2Y102_SLICE_X0Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y102_SLICE_X1Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y102_SLICE_X1Y102_DO5),
.O6(CLBLL_L_X2Y102_SLICE_X1Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y102_SLICE_X1Y102_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y102_SLICE_X1Y102_CO5),
.O6(CLBLL_L_X2Y102_SLICE_X1Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y102_SLICE_X1Y102_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y102_SLICE_X1Y102_BO5),
.O6(CLBLL_L_X2Y102_SLICE_X1Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y102_SLICE_X1Y102_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y102_SLICE_X1Y102_AO5),
.O6(CLBLL_L_X2Y102_SLICE_X1Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y90_SLICE_X4Y90_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y90_SLICE_X4Y90_DO5),
.O6(CLBLL_L_X4Y90_SLICE_X4Y90_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y90_SLICE_X4Y90_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y90_SLICE_X4Y90_CO5),
.O6(CLBLL_L_X4Y90_SLICE_X4Y90_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y90_SLICE_X4Y90_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y90_SLICE_X4Y90_BO5),
.O6(CLBLL_L_X4Y90_SLICE_X4Y90_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y90_SLICE_X4Y90_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y90_SLICE_X4Y90_AO5),
.O6(CLBLL_L_X4Y90_SLICE_X4Y90_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y90_SLICE_X5Y90_A_FDPE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(1'b1),
.D(CLBLM_R_X7Y90_SLICE_X8Y90_AQ),
.PRE(LIOB33_X0Y107_IOB_X0Y107_I),
.Q(CLBLL_L_X4Y90_SLICE_X5Y90_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y90_SLICE_X5Y90_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y90_SLICE_X5Y90_DO5),
.O6(CLBLL_L_X4Y90_SLICE_X5Y90_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y90_SLICE_X5Y90_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y90_SLICE_X5Y90_CO5),
.O6(CLBLL_L_X4Y90_SLICE_X5Y90_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y90_SLICE_X5Y90_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y90_SLICE_X5Y90_BO5),
.O6(CLBLL_L_X4Y90_SLICE_X5Y90_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y90_SLICE_X5Y90_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y90_SLICE_X5Y90_AO5),
.O6(CLBLL_L_X4Y90_SLICE_X5Y90_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y91_SLICE_X4Y91_A_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLL_L_X2Y93_SLICE_X1Y93_CO6),
.D(CLBLL_L_X4Y93_SLICE_X4Y93_CO5),
.Q(CLBLL_L_X4Y91_SLICE_X4Y91_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y91_SLICE_X4Y91_B_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLL_L_X2Y93_SLICE_X1Y93_CO6),
.D(CLBLL_L_X4Y92_SLICE_X4Y92_AO5),
.Q(CLBLL_L_X4Y91_SLICE_X4Y91_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y91_SLICE_X4Y91_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y91_SLICE_X4Y91_DO5),
.O6(CLBLL_L_X4Y91_SLICE_X4Y91_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y91_SLICE_X4Y91_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y91_SLICE_X4Y91_CO5),
.O6(CLBLL_L_X4Y91_SLICE_X4Y91_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaaeaaa2aa)
  ) CLBLL_L_X4Y91_SLICE_X4Y91_BLUT (
.I0(CLBLM_R_X3Y91_SLICE_X3Y91_F7BMUX_O),
.I1(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I2(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I3(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I4(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO5),
.I5(CLBLL_L_X4Y91_SLICE_X4Y91_AO5),
.O5(CLBLL_L_X4Y91_SLICE_X4Y91_BO5),
.O6(CLBLL_L_X4Y91_SLICE_X4Y91_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00440008fafafafa)
  ) CLBLL_L_X4Y91_SLICE_X4Y91_ALUT (
.I0(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I1(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO5),
.I2(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I3(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I4(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y91_SLICE_X4Y91_AO5),
.O6(CLBLL_L_X4Y91_SLICE_X4Y91_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y91_SLICE_X5Y91_B_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLL_L_X2Y93_SLICE_X0Y93_DO6),
.D(CLBLL_L_X4Y92_SLICE_X4Y92_AO5),
.Q(CLBLL_L_X4Y91_SLICE_X5Y91_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y91_SLICE_X5Y91_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y91_SLICE_X5Y91_DO5),
.O6(CLBLL_L_X4Y91_SLICE_X5Y91_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff4400ffff4400)
  ) CLBLL_L_X4Y91_SLICE_X5Y91_CLUT (
.I0(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I1(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I4(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y91_SLICE_X5Y91_CO5),
.O6(CLBLL_L_X4Y91_SLICE_X5Y91_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f0303200000002)
  ) CLBLL_L_X4Y91_SLICE_X5Y91_BLUT (
.I0(CLBLL_L_X4Y94_SLICE_X5Y94_CO6),
.I1(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I2(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I3(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I4(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I5(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO8),
.O5(CLBLL_L_X4Y91_SLICE_X5Y91_BO5),
.O6(CLBLL_L_X4Y91_SLICE_X5Y91_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0044ccff00000000)
  ) CLBLL_L_X4Y91_SLICE_X5Y91_ALUT (
.I0(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I1(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I4(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I5(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO8),
.O5(CLBLL_L_X4Y91_SLICE_X5Y91_AO5),
.O6(CLBLL_L_X4Y91_SLICE_X5Y91_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_L_X4Y91_SLICE_X5Y91_MUXF7A (
.I0(CLBLL_L_X4Y91_SLICE_X5Y91_BO6),
.I1(CLBLL_L_X4Y91_SLICE_X5Y91_AO6),
.O(CLBLL_L_X4Y91_SLICE_X5Y91_F7AMUX_O),
.S(CLBLL_L_X4Y91_SLICE_X5Y91_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y92_SLICE_X4Y92_B5_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLL_L_X4Y92_SLICE_X4Y92_BO6),
.D(CLBLL_L_X4Y94_SLICE_X4Y94_CO6),
.Q(CLBLL_L_X4Y92_SLICE_X4Y92_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y92_SLICE_X4Y92_A_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLL_L_X4Y92_SLICE_X4Y92_BO6),
.D(CLBLL_L_X4Y93_SLICE_X4Y93_CO5),
.Q(CLBLL_L_X4Y92_SLICE_X4Y92_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y92_SLICE_X4Y92_B_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLL_L_X4Y92_SLICE_X4Y92_BO6),
.D(CLBLL_L_X4Y92_SLICE_X4Y92_BO5),
.Q(CLBLL_L_X4Y92_SLICE_X4Y92_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y92_SLICE_X4Y92_C_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLL_L_X4Y92_SLICE_X4Y92_BO6),
.D(CLBLL_L_X4Y93_SLICE_X4Y93_CO6),
.Q(CLBLL_L_X4Y92_SLICE_X4Y92_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y92_SLICE_X4Y92_D_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLL_L_X4Y92_SLICE_X4Y92_BO6),
.D(CLBLL_L_X4Y92_SLICE_X4Y92_AO5),
.Q(CLBLL_L_X4Y92_SLICE_X4Y92_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y92_SLICE_X4Y92_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y92_SLICE_X4Y92_DO5),
.O6(CLBLL_L_X4Y92_SLICE_X4Y92_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y92_SLICE_X4Y92_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y92_SLICE_X4Y92_CO5),
.O6(CLBLL_L_X4Y92_SLICE_X4Y92_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000808ff00ff00)
  ) CLBLL_L_X4Y92_SLICE_X4Y92_BLUT (
.I0(CLBLM_R_X5Y94_SLICE_X7Y94_DO6),
.I1(CLBLL_L_X2Y93_SLICE_X0Y93_CO6),
.I2(CLBLL_L_X4Y94_SLICE_X5Y94_DO6),
.I3(CLBLM_R_X3Y94_SLICE_X2Y94_DO5),
.I4(CLBLM_R_X5Y94_SLICE_X6Y94_BO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y92_SLICE_X4Y92_BO5),
.O6(CLBLL_L_X4Y92_SLICE_X4Y92_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8d8d8ffaa5500)
  ) CLBLL_L_X4Y92_SLICE_X4Y92_ALUT (
.I0(CLBLM_R_X3Y93_SLICE_X2Y93_CO6),
.I1(CLBLL_L_X2Y96_SLICE_X1Y96_AO6),
.I2(CLBLL_L_X4Y96_SLICE_X4Y96_AO6),
.I3(CLBLL_L_X4Y96_SLICE_X5Y96_AO6),
.I4(CLBLL_L_X2Y96_SLICE_X1Y96_BO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y92_SLICE_X4Y92_AO5),
.O6(CLBLL_L_X4Y92_SLICE_X4Y92_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y92_SLICE_X5Y92_B_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLL_L_X2Y93_SLICE_X0Y93_DO6),
.D(CLBLL_L_X4Y93_SLICE_X4Y93_CO5),
.Q(CLBLL_L_X4Y92_SLICE_X5Y92_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y92_SLICE_X5Y92_C_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLL_L_X2Y93_SLICE_X0Y93_DO6),
.D(CLBLL_L_X4Y94_SLICE_X4Y94_CO6),
.Q(CLBLL_L_X4Y92_SLICE_X5Y92_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbf80bf80aaaaff00)
  ) CLBLL_L_X4Y92_SLICE_X5Y92_DLUT (
.I0(CLBLL_L_X4Y92_SLICE_X4Y92_AQ),
.I1(CLBLM_R_X5Y94_SLICE_X7Y94_AO5),
.I2(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO8),
.I3(CLBLM_R_X5Y92_SLICE_X6Y92_CQ),
.I4(CLBLL_L_X4Y91_SLICE_X5Y91_BO6),
.I5(CLBLL_L_X4Y91_SLICE_X5Y91_CO6),
.O5(CLBLL_L_X4Y92_SLICE_X5Y92_DO5),
.O6(CLBLL_L_X4Y92_SLICE_X5Y92_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff2aff7fd5008000)
  ) CLBLL_L_X4Y92_SLICE_X5Y92_CLUT (
.I0(CLBLL_L_X4Y91_SLICE_X5Y91_CO6),
.I1(CLBLM_R_X5Y94_SLICE_X7Y94_AO5),
.I2(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO8),
.I3(CLBLL_L_X4Y93_SLICE_X5Y93_BQ),
.I4(CLBLL_L_X4Y91_SLICE_X5Y91_BO6),
.I5(CLBLL_L_X4Y92_SLICE_X5Y92_BQ),
.O5(CLBLL_L_X4Y92_SLICE_X5Y92_CO5),
.O6(CLBLL_L_X4Y92_SLICE_X5Y92_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000ccaaccaa)
  ) CLBLL_L_X4Y92_SLICE_X5Y92_BLUT (
.I0(CLBLM_R_X5Y92_SLICE_X6Y92_CQ),
.I1(CLBLM_R_X5Y94_SLICE_X6Y94_AQ),
.I2(CLBLL_L_X4Y91_SLICE_X4Y91_AQ),
.I3(CLBLM_R_X3Y96_SLICE_X3Y96_AO6),
.I4(CLBLL_L_X4Y92_SLICE_X4Y92_AQ),
.I5(CLBLL_L_X4Y91_SLICE_X4Y91_AO6),
.O5(CLBLL_L_X4Y92_SLICE_X5Y92_BO5),
.O6(CLBLL_L_X4Y92_SLICE_X5Y92_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0ccaa00f0ccaa)
  ) CLBLL_L_X4Y92_SLICE_X5Y92_ALUT (
.I0(CLBLM_R_X3Y93_SLICE_X3Y93_AQ),
.I1(CLBLL_L_X4Y92_SLICE_X5Y92_BQ),
.I2(CLBLL_L_X4Y94_SLICE_X5Y94_BQ),
.I3(CLBLM_R_X3Y96_SLICE_X3Y96_AO6),
.I4(CLBLL_L_X4Y91_SLICE_X4Y91_AO6),
.I5(CLBLL_L_X4Y93_SLICE_X5Y93_BQ),
.O5(CLBLL_L_X4Y92_SLICE_X5Y92_AO5),
.O6(CLBLL_L_X4Y92_SLICE_X5Y92_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_L_X4Y92_SLICE_X5Y92_MUXF7A (
.I0(CLBLL_L_X4Y92_SLICE_X5Y92_BO6),
.I1(CLBLL_L_X4Y92_SLICE_X5Y92_AO6),
.O(CLBLL_L_X4Y92_SLICE_X5Y92_F7AMUX_O),
.S(CLBLL_L_X4Y95_SLICE_X5Y95_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y93_SLICE_X4Y93_B_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLL_L_X2Y93_SLICE_X1Y93_CO6),
.D(CLBLM_R_X3Y94_SLICE_X2Y94_DO5),
.Q(CLBLL_L_X4Y93_SLICE_X4Y93_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y93_SLICE_X4Y93_C_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLL_L_X2Y93_SLICE_X1Y93_CO6),
.D(CLBLL_L_X4Y93_SLICE_X4Y93_CO6),
.Q(CLBLL_L_X4Y93_SLICE_X4Y93_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y93_SLICE_X4Y93_D_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLL_L_X2Y93_SLICE_X1Y93_CO6),
.D(CLBLL_L_X4Y94_SLICE_X4Y94_CO6),
.Q(CLBLL_L_X4Y93_SLICE_X4Y93_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44f5f5ee44a0a0)
  ) CLBLL_L_X4Y93_SLICE_X4Y93_DLUT (
.I0(CLBLM_R_X5Y93_SLICE_X6Y93_F7AMUX_O),
.I1(CLBLL_L_X4Y93_SLICE_X5Y93_CO6),
.I2(CLBLL_L_X4Y93_SLICE_X5Y93_DO6),
.I3(CLBLL_L_X4Y92_SLICE_X5Y92_CO6),
.I4(CLBLL_L_X2Y93_SLICE_X0Y93_F7AMUX_O),
.I5(CLBLL_L_X4Y92_SLICE_X5Y92_DO6),
.O5(CLBLL_L_X4Y93_SLICE_X4Y93_DO5),
.O6(CLBLL_L_X4Y93_SLICE_X4Y93_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0ccaaffaa00)
  ) CLBLL_L_X4Y93_SLICE_X4Y93_CLUT (
.I0(CLBLL_L_X2Y97_SLICE_X0Y97_BO6),
.I1(CLBLM_R_X3Y98_SLICE_X2Y98_CO6),
.I2(CLBLL_L_X2Y97_SLICE_X1Y97_BO6),
.I3(CLBLM_R_X3Y93_SLICE_X2Y93_CO6),
.I4(CLBLM_R_X3Y99_SLICE_X2Y99_CO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y93_SLICE_X4Y93_CO5),
.O6(CLBLL_L_X4Y93_SLICE_X4Y93_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50fa50dddd8888)
  ) CLBLL_L_X4Y93_SLICE_X4Y93_BLUT (
.I0(CLBLM_R_X5Y93_SLICE_X6Y93_F7AMUX_O),
.I1(CLBLL_L_X4Y95_SLICE_X4Y95_AQ),
.I2(CLBLL_L_X4Y92_SLICE_X4Y92_CQ),
.I3(CLBLL_L_X4Y93_SLICE_X4Y93_CQ),
.I4(CLBLL_L_X4Y94_SLICE_X4Y94_AQ),
.I5(CLBLL_L_X4Y91_SLICE_X5Y91_F7AMUX_O),
.O5(CLBLL_L_X4Y93_SLICE_X4Y93_BO5),
.O6(CLBLL_L_X4Y93_SLICE_X4Y93_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdf85d58ada80d08)
  ) CLBLL_L_X4Y93_SLICE_X4Y93_ALUT (
.I0(CLBLM_R_X5Y93_SLICE_X6Y93_F7AMUX_O),
.I1(CLBLM_R_X5Y93_SLICE_X6Y93_BQ),
.I2(CLBLL_L_X4Y91_SLICE_X5Y91_F7AMUX_O),
.I3(CLBLM_R_X3Y93_SLICE_X3Y93_CQ),
.I4(CLBLL_L_X4Y93_SLICE_X5Y93_CQ),
.I5(CLBLL_L_X4Y94_SLICE_X5Y94_CQ),
.O5(CLBLL_L_X4Y93_SLICE_X4Y93_AO5),
.O6(CLBLL_L_X4Y93_SLICE_X4Y93_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_L_X4Y93_SLICE_X4Y93_MUXF7A (
.I0(CLBLL_L_X4Y93_SLICE_X4Y93_BO6),
.I1(CLBLL_L_X4Y93_SLICE_X4Y93_AO6),
.O(CLBLL_L_X4Y93_SLICE_X4Y93_F7AMUX_O),
.S(CLBLL_L_X2Y93_SLICE_X0Y93_F7AMUX_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y93_SLICE_X5Y93_B_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLL_L_X2Y93_SLICE_X1Y93_DO6),
.D(CLBLL_L_X4Y93_SLICE_X4Y93_CO5),
.Q(CLBLL_L_X4Y93_SLICE_X5Y93_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y93_SLICE_X5Y93_C_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLL_L_X2Y93_SLICE_X1Y93_DO6),
.D(CLBLL_L_X4Y93_SLICE_X4Y93_CO6),
.Q(CLBLL_L_X4Y93_SLICE_X5Y93_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y93_SLICE_X5Y93_D_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLL_L_X2Y93_SLICE_X1Y93_DO6),
.D(CLBLL_L_X4Y94_SLICE_X4Y94_CO6),
.Q(CLBLL_L_X4Y93_SLICE_X5Y93_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haae2e2e2b8f0f0f0)
  ) CLBLL_L_X4Y93_SLICE_X5Y93_DLUT (
.I0(CLBLL_L_X4Y91_SLICE_X4Y91_AQ),
.I1(CLBLL_L_X4Y91_SLICE_X5Y91_CO6),
.I2(CLBLM_R_X5Y94_SLICE_X6Y94_AQ),
.I3(CLBLM_R_X5Y94_SLICE_X7Y94_AO5),
.I4(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO8),
.I5(CLBLL_L_X4Y91_SLICE_X5Y91_BO6),
.O5(CLBLL_L_X4Y93_SLICE_X5Y93_DO5),
.O6(CLBLL_L_X4Y93_SLICE_X5Y93_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfef2f2f210d0d0d0)
  ) CLBLL_L_X4Y93_SLICE_X5Y93_CLUT (
.I0(CLBLL_L_X4Y91_SLICE_X5Y91_BO6),
.I1(CLBLL_L_X4Y91_SLICE_X5Y91_CO6),
.I2(CLBLM_R_X3Y93_SLICE_X3Y93_AQ),
.I3(CLBLM_R_X5Y94_SLICE_X7Y94_AO5),
.I4(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO8),
.I5(CLBLL_L_X4Y94_SLICE_X5Y94_BQ),
.O5(CLBLL_L_X4Y93_SLICE_X5Y93_CO5),
.O6(CLBLL_L_X4Y93_SLICE_X5Y93_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88dd88fafa5050)
  ) CLBLL_L_X4Y93_SLICE_X5Y93_BLUT (
.I0(CLBLM_R_X3Y96_SLICE_X3Y96_AO6),
.I1(CLBLL_L_X4Y93_SLICE_X4Y93_CQ),
.I2(CLBLL_L_X4Y94_SLICE_X4Y94_AQ),
.I3(CLBLL_L_X4Y92_SLICE_X4Y92_CQ),
.I4(CLBLL_L_X4Y95_SLICE_X4Y95_AQ),
.I5(CLBLL_L_X4Y91_SLICE_X4Y91_AO6),
.O5(CLBLL_L_X4Y93_SLICE_X5Y93_BO5),
.O6(CLBLL_L_X4Y93_SLICE_X5Y93_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5ee44a0a0ee44)
  ) CLBLL_L_X4Y93_SLICE_X5Y93_ALUT (
.I0(CLBLM_R_X3Y96_SLICE_X3Y96_AO6),
.I1(CLBLM_R_X3Y93_SLICE_X3Y93_CQ),
.I2(CLBLL_L_X4Y93_SLICE_X5Y93_CQ),
.I3(CLBLM_R_X5Y93_SLICE_X6Y93_BQ),
.I4(CLBLL_L_X4Y91_SLICE_X4Y91_AO6),
.I5(CLBLL_L_X4Y94_SLICE_X5Y94_CQ),
.O5(CLBLL_L_X4Y93_SLICE_X5Y93_AO5),
.O6(CLBLL_L_X4Y93_SLICE_X5Y93_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_L_X4Y93_SLICE_X5Y93_MUXF7A (
.I0(CLBLL_L_X4Y93_SLICE_X5Y93_BO6),
.I1(CLBLL_L_X4Y93_SLICE_X5Y93_AO6),
.O(CLBLL_L_X4Y93_SLICE_X5Y93_F7AMUX_O),
.S(CLBLL_L_X4Y95_SLICE_X5Y95_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y94_SLICE_X4Y94_A_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(1'b1),
.D(CLBLL_L_X4Y94_SLICE_X4Y94_AO6),
.Q(CLBLL_L_X4Y94_SLICE_X4Y94_AQ),
.R(CLBLM_R_X5Y92_SLICE_X7Y92_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y94_SLICE_X4Y94_B_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(1'b1),
.D(CLBLL_L_X4Y94_SLICE_X4Y94_BO6),
.Q(CLBLL_L_X4Y94_SLICE_X4Y94_BQ),
.R(CLBLM_R_X5Y92_SLICE_X7Y92_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8088808880c580c0)
  ) CLBLL_L_X4Y94_SLICE_X4Y94_DLUT (
.I0(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I1(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO10),
.I2(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I3(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I4(CLBLL_L_X4Y96_SLICE_X4Y96_DO6),
.I5(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.O5(CLBLL_L_X4Y94_SLICE_X4Y94_DO5),
.O6(CLBLL_L_X4Y94_SLICE_X4Y94_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88dd88f5f5a0a0)
  ) CLBLL_L_X4Y94_SLICE_X4Y94_CLUT (
.I0(CLBLM_R_X3Y93_SLICE_X2Y93_CO6),
.I1(CLBLL_L_X2Y97_SLICE_X1Y97_CO6),
.I2(CLBLL_L_X2Y96_SLICE_X1Y96_DO6),
.I3(CLBLL_L_X4Y96_SLICE_X4Y96_CO6),
.I4(CLBLM_R_X3Y96_SLICE_X3Y96_DO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y94_SLICE_X4Y94_CO5),
.O6(CLBLL_L_X4Y94_SLICE_X4Y94_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000011011000)
  ) CLBLL_L_X4Y94_SLICE_X4Y94_BLUT (
.I0(CLBLM_R_X5Y94_SLICE_X7Y94_DO6),
.I1(CLBLL_L_X4Y94_SLICE_X5Y94_DO6),
.I2(CLBLM_R_X3Y93_SLICE_X2Y93_CO6),
.I3(CLBLL_L_X2Y97_SLICE_X1Y97_CO6),
.I4(CLBLL_L_X4Y96_SLICE_X4Y96_CO6),
.I5(CLBLM_R_X5Y94_SLICE_X6Y94_BO6),
.O5(CLBLL_L_X4Y94_SLICE_X4Y94_BO5),
.O6(CLBLL_L_X4Y94_SLICE_X4Y94_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000004040500)
  ) CLBLL_L_X4Y94_SLICE_X4Y94_ALUT (
.I0(CLBLM_R_X5Y94_SLICE_X7Y94_DO6),
.I1(CLBLL_L_X2Y97_SLICE_X1Y97_BO6),
.I2(CLBLL_L_X4Y94_SLICE_X5Y94_DO6),
.I3(CLBLM_R_X3Y98_SLICE_X2Y98_CO6),
.I4(CLBLM_R_X3Y93_SLICE_X2Y93_CO6),
.I5(CLBLM_R_X5Y94_SLICE_X6Y94_BO6),
.O5(CLBLL_L_X4Y94_SLICE_X4Y94_AO5),
.O6(CLBLL_L_X4Y94_SLICE_X4Y94_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y94_SLICE_X5Y94_B_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X3Y93_SLICE_X3Y93_CO6),
.D(CLBLL_L_X4Y93_SLICE_X4Y93_CO5),
.Q(CLBLL_L_X4Y94_SLICE_X5Y94_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y94_SLICE_X5Y94_C_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X3Y93_SLICE_X3Y93_CO6),
.D(CLBLL_L_X4Y93_SLICE_X4Y93_CO6),
.Q(CLBLL_L_X4Y94_SLICE_X5Y94_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y94_SLICE_X5Y94_D_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X3Y93_SLICE_X3Y93_CO6),
.D(CLBLL_L_X4Y94_SLICE_X4Y94_CO6),
.Q(CLBLL_L_X4Y94_SLICE_X5Y94_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff004400f4f0f4f0)
  ) CLBLL_L_X4Y94_SLICE_X5Y94_DLUT (
.I0(CLBLM_R_X5Y94_SLICE_X7Y94_AO6),
.I1(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I2(CLBLL_L_X4Y94_SLICE_X4Y94_DO6),
.I3(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO10),
.I4(CLBLM_R_X5Y94_SLICE_X7Y94_AO5),
.I5(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.O5(CLBLL_L_X4Y94_SLICE_X5Y94_DO5),
.O6(CLBLL_L_X4Y94_SLICE_X5Y94_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010000000000)
  ) CLBLL_L_X4Y94_SLICE_X5Y94_CLUT (
.I0(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO14),
.I1(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO11),
.I2(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO15),
.I3(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO13),
.I4(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO12),
.I5(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO8),
.O5(CLBLL_L_X4Y94_SLICE_X5Y94_CO5),
.O6(CLBLL_L_X4Y94_SLICE_X5Y94_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacafff0caca0f00)
  ) CLBLL_L_X4Y94_SLICE_X5Y94_BLUT (
.I0(CLBLL_L_X4Y92_SLICE_X4Y92_B5Q),
.I1(CLBLL_L_X4Y93_SLICE_X4Y93_DQ),
.I2(CLBLM_R_X5Y93_SLICE_X6Y93_F7AMUX_O),
.I3(CLBLL_L_X4Y94_SLICE_X4Y94_BQ),
.I4(CLBLL_L_X4Y91_SLICE_X5Y91_F7AMUX_O),
.I5(CLBLM_R_X5Y94_SLICE_X6Y94_BQ),
.O5(CLBLL_L_X4Y94_SLICE_X5Y94_BO5),
.O6(CLBLL_L_X4Y94_SLICE_X5Y94_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacfff0acac0f00)
  ) CLBLL_L_X4Y94_SLICE_X5Y94_ALUT (
.I0(CLBLL_L_X4Y93_SLICE_X5Y93_DQ),
.I1(CLBLL_L_X4Y94_SLICE_X5Y94_DQ),
.I2(CLBLM_R_X5Y93_SLICE_X6Y93_F7AMUX_O),
.I3(CLBLM_R_X3Y93_SLICE_X3Y93_DQ),
.I4(CLBLL_L_X4Y91_SLICE_X5Y91_F7AMUX_O),
.I5(CLBLL_L_X4Y92_SLICE_X5Y92_CQ),
.O5(CLBLL_L_X4Y94_SLICE_X5Y94_AO5),
.O6(CLBLL_L_X4Y94_SLICE_X5Y94_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_L_X4Y94_SLICE_X5Y94_MUXF7A (
.I0(CLBLL_L_X4Y94_SLICE_X5Y94_BO6),
.I1(CLBLL_L_X4Y94_SLICE_X5Y94_AO6),
.O(CLBLL_L_X4Y94_SLICE_X5Y94_F7AMUX_O),
.S(CLBLL_L_X2Y93_SLICE_X0Y93_F7AMUX_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y95_SLICE_X4Y95_A_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLL_L_X2Y92_SLICE_X1Y92_AO6),
.D(CLBLL_L_X4Y93_SLICE_X4Y93_CO6),
.Q(CLBLL_L_X4Y95_SLICE_X4Y95_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0f0f0f870)
  ) CLBLL_L_X4Y95_SLICE_X4Y95_DLUT (
.I0(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I1(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I2(CLBLL_L_X4Y92_SLICE_X5Y92_F7AMUX_O),
.I3(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO0),
.I4(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I5(CLBLL_L_X4Y91_SLICE_X4Y91_AO5),
.O5(CLBLL_L_X4Y95_SLICE_X4Y95_DO5),
.O6(CLBLL_L_X4Y95_SLICE_X4Y95_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0f0f8f070)
  ) CLBLL_L_X4Y95_SLICE_X4Y95_CLUT (
.I0(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I1(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I2(CLBLM_R_X3Y93_SLICE_X2Y93_F7AMUX_O),
.I3(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I4(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO1),
.I5(CLBLL_L_X4Y91_SLICE_X4Y91_AO5),
.O5(CLBLL_L_X4Y95_SLICE_X4Y95_CO5),
.O6(CLBLL_L_X4Y95_SLICE_X4Y95_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffbf00400000)
  ) CLBLL_L_X4Y95_SLICE_X4Y95_BLUT (
.I0(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I1(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I2(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I3(CLBLL_L_X4Y91_SLICE_X4Y91_AO5),
.I4(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO3),
.I5(CLBLL_L_X4Y93_SLICE_X5Y93_F7AMUX_O),
.O5(CLBLL_L_X4Y95_SLICE_X4Y95_BO5),
.O6(CLBLL_L_X4Y95_SLICE_X4Y95_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefefdfdffe7fff3)
  ) CLBLL_L_X4Y95_SLICE_X4Y95_ALUT (
.I0(CLBLL_L_X4Y95_SLICE_X5Y95_CO6),
.I1(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I2(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I3(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I4(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I5(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.O5(CLBLL_L_X4Y95_SLICE_X4Y95_AO5),
.O6(CLBLL_L_X4Y95_SLICE_X4Y95_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0040004010401040)
  ) CLBLL_L_X4Y95_SLICE_X5Y95_DLUT (
.I0(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I1(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I2(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO7),
.I3(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.O5(CLBLL_L_X4Y95_SLICE_X5Y95_DO5),
.O6(CLBLL_L_X4Y95_SLICE_X5Y95_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00fd20ff00)
  ) CLBLL_L_X4Y95_SLICE_X5Y95_CLUT (
.I0(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I1(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I2(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO6),
.I3(CLBLL_L_X4Y95_SLICE_X5Y95_F7AMUX_O),
.I4(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I5(CLBLL_L_X4Y91_SLICE_X4Y91_AO5),
.O5(CLBLL_L_X4Y95_SLICE_X5Y95_CO5),
.O6(CLBLL_L_X4Y95_SLICE_X5Y95_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haffca0fcaf0ca00c)
  ) CLBLL_L_X4Y95_SLICE_X5Y95_BLUT (
.I0(CLBLL_L_X4Y93_SLICE_X4Y93_DQ),
.I1(CLBLL_L_X4Y94_SLICE_X4Y94_BQ),
.I2(CLBLL_L_X4Y91_SLICE_X4Y91_AO6),
.I3(CLBLM_R_X3Y96_SLICE_X3Y96_AO6),
.I4(CLBLM_R_X5Y94_SLICE_X6Y94_BQ),
.I5(CLBLL_L_X4Y92_SLICE_X4Y92_B5Q),
.O5(CLBLL_L_X4Y95_SLICE_X5Y95_BO5),
.O6(CLBLL_L_X4Y95_SLICE_X5Y95_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafcfa0cfafc0a0c0)
  ) CLBLL_L_X4Y95_SLICE_X5Y95_ALUT (
.I0(CLBLL_L_X4Y93_SLICE_X5Y93_DQ),
.I1(CLBLL_L_X4Y94_SLICE_X5Y94_DQ),
.I2(CLBLL_L_X4Y91_SLICE_X4Y91_AO6),
.I3(CLBLM_R_X3Y96_SLICE_X3Y96_AO6),
.I4(CLBLL_L_X4Y92_SLICE_X5Y92_CQ),
.I5(CLBLM_R_X3Y93_SLICE_X3Y93_DQ),
.O5(CLBLL_L_X4Y95_SLICE_X5Y95_AO5),
.O6(CLBLL_L_X4Y95_SLICE_X5Y95_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_L_X4Y95_SLICE_X5Y95_MUXF7A (
.I0(CLBLL_L_X4Y95_SLICE_X5Y95_BO6),
.I1(CLBLL_L_X4Y95_SLICE_X5Y95_AO6),
.O(CLBLL_L_X4Y95_SLICE_X5Y95_F7AMUX_O),
.S(CLBLL_L_X4Y95_SLICE_X5Y95_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0004000000000000)
  ) CLBLL_L_X4Y96_SLICE_X4Y96_DLUT (
.I0(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO14),
.I1(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO10),
.I2(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO15),
.I3(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO13),
.I4(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO12),
.I5(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO11),
.O5(CLBLL_L_X4Y96_SLICE_X4Y96_DO5),
.O6(CLBLL_L_X4Y96_SLICE_X4Y96_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888888888d8)
  ) CLBLL_L_X4Y96_SLICE_X4Y96_CLUT (
.I0(CLBLL_L_X4Y97_SLICE_X4Y97_AO6),
.I1(CLBLL_L_X4Y96_SLICE_X5Y96_CO6),
.I2(CLBLM_R_X3Y96_SLICE_X2Y96_BO6),
.I3(CLBLL_L_X4Y98_SLICE_X4Y98_AO6),
.I4(CLBLL_L_X4Y97_SLICE_X4Y97_CO6),
.I5(CLBLM_R_X3Y98_SLICE_X3Y98_AO6),
.O5(CLBLL_L_X4Y96_SLICE_X4Y96_CO5),
.O6(CLBLL_L_X4Y96_SLICE_X4Y96_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000200000000)
  ) CLBLL_L_X4Y96_SLICE_X4Y96_BLUT (
.I0(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO4),
.I1(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I2(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I3(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I4(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I5(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.O5(CLBLL_L_X4Y96_SLICE_X4Y96_BO5),
.O6(CLBLL_L_X4Y96_SLICE_X4Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000101ff000000)
  ) CLBLL_L_X4Y96_SLICE_X4Y96_ALUT (
.I0(CLBLM_R_X3Y98_SLICE_X3Y98_AO6),
.I1(CLBLL_L_X4Y98_SLICE_X4Y98_AO6),
.I2(CLBLL_L_X4Y97_SLICE_X4Y97_CO6),
.I3(CLBLL_L_X4Y96_SLICE_X4Y96_BO6),
.I4(CLBLL_L_X4Y97_SLICE_X4Y97_AO6),
.I5(CLBLM_R_X3Y96_SLICE_X2Y96_DO6),
.O5(CLBLL_L_X4Y96_SLICE_X4Y96_AO5),
.O6(CLBLL_L_X4Y96_SLICE_X4Y96_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y96_SLICE_X5Y96_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y96_SLICE_X5Y96_DO5),
.O6(CLBLL_L_X4Y96_SLICE_X5Y96_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000040000)
  ) CLBLL_L_X4Y96_SLICE_X5Y96_CLUT (
.I0(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I1(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I2(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I3(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I4(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO6),
.I5(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.O5(CLBLL_L_X4Y96_SLICE_X5Y96_CO5),
.O6(CLBLL_L_X4Y96_SLICE_X5Y96_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000200)
  ) CLBLL_L_X4Y96_SLICE_X5Y96_BLUT (
.I0(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I1(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I2(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I3(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO5),
.I4(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I5(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.O5(CLBLL_L_X4Y96_SLICE_X5Y96_BO5),
.O6(CLBLL_L_X4Y96_SLICE_X5Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000f000f404)
  ) CLBLL_L_X4Y96_SLICE_X5Y96_ALUT (
.I0(CLBLL_L_X4Y98_SLICE_X4Y98_AO6),
.I1(CLBLM_R_X3Y96_SLICE_X2Y96_AO6),
.I2(CLBLL_L_X4Y97_SLICE_X4Y97_AO6),
.I3(CLBLL_L_X4Y96_SLICE_X5Y96_BO6),
.I4(CLBLL_L_X4Y97_SLICE_X4Y97_CO6),
.I5(CLBLM_R_X3Y98_SLICE_X3Y98_AO6),
.O5(CLBLL_L_X4Y96_SLICE_X5Y96_AO5),
.O6(CLBLL_L_X4Y96_SLICE_X5Y96_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y97_SLICE_X4Y97_B_FDCE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(1'b1),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLL_L_X4Y97_SLICE_X4Y97_BO6),
.Q(CLBLL_L_X4Y97_SLICE_X4Y97_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000002001000)
  ) CLBLL_L_X4Y97_SLICE_X4Y97_DLUT (
.I0(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO11),
.I1(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO15),
.I2(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO13),
.I3(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO6),
.I4(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO12),
.I5(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO14),
.O5(CLBLL_L_X4Y97_SLICE_X4Y97_DO5),
.O6(CLBLL_L_X4Y97_SLICE_X4Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0100010001010000)
  ) CLBLL_L_X4Y97_SLICE_X4Y97_CLUT (
.I0(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I1(CLBLL_L_X4Y97_SLICE_X5Y97_AO6),
.I2(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I3(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO6),
.I4(CLBLL_L_X4Y97_SLICE_X4Y97_DO6),
.I5(CLBLM_R_X3Y96_SLICE_X3Y96_AO5),
.O5(CLBLL_L_X4Y97_SLICE_X4Y97_CO5),
.O6(CLBLL_L_X4Y97_SLICE_X4Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa00aacccccccc)
  ) CLBLL_L_X4Y97_SLICE_X4Y97_BLUT (
.I0(CLBLL_L_X2Y97_SLICE_X1Y97_DO6),
.I1(CLBLL_L_X4Y97_SLICE_X4Y97_BQ),
.I2(1'b1),
.I3(CLBLL_L_X2Y97_SLICE_X0Y97_DO6),
.I4(1'b1),
.I5(CLBLL_L_X4Y97_SLICE_X4Y97_AO5),
.O5(CLBLL_L_X4Y97_SLICE_X4Y97_BO5),
.O6(CLBLL_L_X4Y97_SLICE_X4Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000200000010)
  ) CLBLL_L_X4Y97_SLICE_X4Y97_ALUT (
.I0(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I1(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I2(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I3(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I4(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y97_SLICE_X4Y97_AO5),
.O6(CLBLL_L_X4Y97_SLICE_X4Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0800600008006000)
  ) CLBLL_L_X4Y97_SLICE_X5Y97_DLUT (
.I0(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I1(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I2(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I3(CLBLL_L_X4Y97_SLICE_X5Y97_AO5),
.I4(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y97_SLICE_X5Y97_DO5),
.O6(CLBLL_L_X4Y97_SLICE_X5Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0b0e0104a1a40104)
  ) CLBLL_L_X4Y97_SLICE_X5Y97_CLUT (
.I0(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I1(CLBLM_R_X5Y97_SLICE_X7Y97_AO5),
.I2(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I3(CLBLM_R_X5Y97_SLICE_X6Y97_BO6),
.I4(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO5),
.I5(CLBLL_L_X4Y97_SLICE_X4Y97_BQ),
.O5(CLBLL_L_X4Y97_SLICE_X5Y97_CO5),
.O6(CLBLL_L_X4Y97_SLICE_X5Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0220ffff02200000)
  ) CLBLL_L_X4Y97_SLICE_X5Y97_BLUT (
.I0(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO5),
.I1(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I2(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I3(CLBLM_R_X5Y95_SLICE_X6Y95_AQ),
.I4(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I5(CLBLL_L_X4Y97_SLICE_X5Y97_CO6),
.O5(CLBLL_L_X4Y97_SLICE_X5Y97_BO5),
.O6(CLBLL_L_X4Y97_SLICE_X5Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff3030d2d20fd2)
  ) CLBLL_L_X4Y97_SLICE_X5Y97_ALUT (
.I0(CLBLM_R_X5Y95_SLICE_X6Y95_AQ),
.I1(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I2(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I3(CLBLL_L_X4Y97_SLICE_X4Y97_BQ),
.I4(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y97_SLICE_X5Y97_AO5),
.O6(CLBLL_L_X4Y97_SLICE_X5Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000050400000100)
  ) CLBLL_L_X4Y98_SLICE_X4Y98_DLUT (
.I0(CLBLL_L_X4Y97_SLICE_X5Y97_AO6),
.I1(CLBLM_R_X3Y96_SLICE_X3Y96_AO5),
.I2(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I3(CLBLL_L_X4Y98_SLICE_X4Y98_CO6),
.I4(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I5(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO1),
.O5(CLBLL_L_X4Y98_SLICE_X4Y98_DO5),
.O6(CLBLL_L_X4Y98_SLICE_X4Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0002000400000000)
  ) CLBLL_L_X4Y98_SLICE_X4Y98_CLUT (
.I0(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO12),
.I1(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO13),
.I2(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO15),
.I3(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO14),
.I4(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO11),
.I5(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO1),
.O5(CLBLL_L_X4Y98_SLICE_X4Y98_CO5),
.O6(CLBLL_L_X4Y98_SLICE_X4Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000004000200)
  ) CLBLL_L_X4Y98_SLICE_X4Y98_BLUT (
.I0(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO13),
.I1(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO11),
.I2(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO14),
.I3(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO5),
.I4(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO12),
.I5(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO15),
.O5(CLBLL_L_X4Y98_SLICE_X4Y98_BO5),
.O6(CLBLL_L_X4Y98_SLICE_X4Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000050400000100)
  ) CLBLL_L_X4Y98_SLICE_X4Y98_ALUT (
.I0(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I1(CLBLM_R_X3Y96_SLICE_X3Y96_AO5),
.I2(CLBLL_L_X4Y97_SLICE_X5Y97_AO6),
.I3(CLBLL_L_X4Y98_SLICE_X4Y98_BO6),
.I4(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I5(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO5),
.O5(CLBLL_L_X4Y98_SLICE_X4Y98_AO5),
.O6(CLBLL_L_X4Y98_SLICE_X4Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000005040100)
  ) CLBLL_L_X4Y98_SLICE_X5Y98_DLUT (
.I0(CLBLL_L_X4Y97_SLICE_X5Y97_AO6),
.I1(CLBLM_R_X3Y96_SLICE_X3Y96_AO5),
.I2(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I3(CLBLL_L_X4Y98_SLICE_X5Y98_CO6),
.I4(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO4),
.I5(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.O5(CLBLL_L_X4Y98_SLICE_X5Y98_DO5),
.O6(CLBLL_L_X4Y98_SLICE_X5Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0010000000001000)
  ) CLBLL_L_X4Y98_SLICE_X5Y98_CLUT (
.I0(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO14),
.I1(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO15),
.I2(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO4),
.I3(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO13),
.I4(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO12),
.I5(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO11),
.O5(CLBLL_L_X4Y98_SLICE_X5Y98_CO5),
.O6(CLBLL_L_X4Y98_SLICE_X5Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010000000000)
  ) CLBLL_L_X4Y98_SLICE_X5Y98_BLUT (
.I0(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I1(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I2(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I3(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO1),
.I4(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I5(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.O5(CLBLL_L_X4Y98_SLICE_X5Y98_BO5),
.O6(CLBLL_L_X4Y98_SLICE_X5Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h557d002855550000)
  ) CLBLL_L_X4Y98_SLICE_X5Y98_ALUT (
.I0(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I1(CLBLM_R_X5Y95_SLICE_X6Y95_AQ),
.I2(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I3(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I4(CLBLM_R_X5Y98_SLICE_X7Y98_BO6),
.I5(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO2),
.O5(CLBLL_L_X4Y98_SLICE_X5Y98_AO5),
.O6(CLBLL_L_X4Y98_SLICE_X5Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y89_SLICE_X10Y89_A5_FDCE (
.C(CLBLM_R_X7Y88_SLICE_X8Y88_AQ),
.CE(CLBLM_R_X7Y88_SLICE_X8Y88_BO6),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_L_X8Y89_SLICE_X10Y89_AO5),
.Q(CLBLM_L_X8Y89_SLICE_X10Y89_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y89_SLICE_X10Y89_A_FDCE (
.C(CLBLM_R_X7Y88_SLICE_X8Y88_AQ),
.CE(CLBLM_R_X7Y88_SLICE_X8Y88_BO6),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_L_X8Y89_SLICE_X10Y89_AO6),
.Q(CLBLM_L_X8Y89_SLICE_X10Y89_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y89_SLICE_X10Y89_B_FDCE (
.C(CLBLM_R_X7Y88_SLICE_X8Y88_AQ),
.CE(CLBLM_R_X7Y88_SLICE_X8Y88_BO6),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_L_X8Y89_SLICE_X10Y89_BO5),
.Q(CLBLM_L_X8Y89_SLICE_X10Y89_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y89_SLICE_X10Y89_C_FDCE (
.C(CLBLM_R_X7Y88_SLICE_X8Y88_AQ),
.CE(CLBLM_R_X7Y88_SLICE_X8Y88_BO6),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_L_X8Y89_SLICE_X10Y89_CO6),
.Q(CLBLM_L_X8Y89_SLICE_X10Y89_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y89_SLICE_X10Y89_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y89_SLICE_X10Y89_DO5),
.O6(CLBLM_L_X8Y89_SLICE_X10Y89_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333333333333)
  ) CLBLM_L_X8Y89_SLICE_X10Y89_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y89_SLICE_X10Y89_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y89_SLICE_X10Y89_CO5),
.O6(CLBLM_L_X8Y89_SLICE_X10Y89_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888888866666666)
  ) CLBLM_L_X8Y89_SLICE_X10Y89_BLUT (
.I0(CLBLM_L_X8Y89_SLICE_X10Y89_CQ),
.I1(CLBLM_L_X8Y89_SLICE_X10Y89_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y89_SLICE_X10Y89_BO5),
.O6(CLBLM_L_X8Y89_SLICE_X10Y89_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h787878787f7f8080)
  ) CLBLM_L_X8Y89_SLICE_X10Y89_ALUT (
.I0(CLBLM_L_X8Y89_SLICE_X10Y89_CQ),
.I1(CLBLM_L_X8Y89_SLICE_X10Y89_BQ),
.I2(CLBLM_L_X8Y89_SLICE_X10Y89_AQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y89_SLICE_X10Y89_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y89_SLICE_X10Y89_AO5),
.O6(CLBLM_L_X8Y89_SLICE_X10Y89_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y89_SLICE_X11Y89_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y89_SLICE_X11Y89_DO5),
.O6(CLBLM_L_X8Y89_SLICE_X11Y89_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y89_SLICE_X11Y89_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y89_SLICE_X11Y89_CO5),
.O6(CLBLM_L_X8Y89_SLICE_X11Y89_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y89_SLICE_X11Y89_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y89_SLICE_X11Y89_BO5),
.O6(CLBLM_L_X8Y89_SLICE_X11Y89_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y89_SLICE_X11Y89_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y89_SLICE_X11Y89_AO5),
.O6(CLBLM_L_X8Y89_SLICE_X11Y89_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a03a0030a0ca00c)
  ) CLBLM_L_X8Y97_SLICE_X10Y97_CLUT (
.I0(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO6),
.I1(CLBLM_R_X5Y97_SLICE_X7Y97_DO6),
.I2(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I3(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I4(CLBLL_L_X4Y97_SLICE_X4Y97_BQ),
.I5(CLBLM_R_X5Y97_SLICE_X6Y97_CO6),
.O5(CLBLM_L_X8Y97_SLICE_X10Y97_CO5),
.O6(CLBLM_L_X8Y97_SLICE_X10Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  RAM32X1S #(
    .INIT(32'h00000000)
  ) CLBLM_L_X8Y97_SLICE_X10Y97_RAM32X1S_D_0 (
.A0(CLBLM_R_X7Y97_SLICE_X9Y97_AQ),
.A1(CLBLM_R_X7Y97_SLICE_X9Y97_A5Q),
.A2(CLBLM_R_X7Y97_SLICE_X9Y97_BQ),
.A3(CLBLM_R_X7Y97_SLICE_X9Y97_B5Q),
.A4(1'b0),
.D(CLBLM_R_X7Y96_SLICE_X9Y96_AQ),
.O(CLBLM_L_X8Y97_SLICE_X10Y97_DO6),
.WCLK(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.WE(CLBLL_L_X4Y97_SLICE_X5Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5LUT" *)
  RAM32X1S #(
    .INIT(32'h00000000)
  ) CLBLM_L_X8Y97_SLICE_X10Y97_RAM32X1S_D_1 (
.A0(CLBLM_R_X7Y97_SLICE_X9Y97_AQ),
.A1(CLBLM_R_X7Y97_SLICE_X9Y97_A5Q),
.A2(CLBLM_R_X7Y97_SLICE_X9Y97_BQ),
.A3(CLBLM_R_X7Y97_SLICE_X9Y97_B5Q),
.A4(1'b0),
.D(1'b1),
.O(CLBLM_L_X8Y97_SLICE_X10Y97_DO5),
.WCLK(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.WE(CLBLL_L_X4Y97_SLICE_X5Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5LUT" *)
  RAM32X1D #(
    .INIT(32'h00000000)
  ) CLBLM_L_X8Y97_SLICE_X10Y97_RAM32X1D_B_1 (
.A0(CLBLM_R_X7Y97_SLICE_X9Y97_AQ),
.A1(CLBLM_R_X7Y97_SLICE_X9Y97_A5Q),
.A2(CLBLM_R_X7Y97_SLICE_X9Y97_BQ),
.A3(CLBLM_R_X7Y97_SLICE_X9Y97_B5Q),
.A4(1'b0),
.D(1'b1),
.DPO(CLBLM_L_X8Y97_SLICE_X10Y97_AO5),
.DPRA0(CLBLM_R_X7Y97_SLICE_X9Y97_AQ),
.DPRA1(CLBLM_R_X7Y97_SLICE_X9Y97_A5Q),
.DPRA2(CLBLM_R_X7Y97_SLICE_X9Y97_BQ),
.DPRA3(CLBLM_R_X7Y97_SLICE_X9Y97_B5Q),
.DPRA4(1'b0),
.SPO(CLBLM_L_X8Y97_SLICE_X10Y97_BO5),
.WCLK(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.WE(CLBLL_L_X4Y97_SLICE_X5Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  RAM32X1D #(
    .INIT(32'h00000000)
  ) CLBLM_L_X8Y97_SLICE_X10Y97_RAM32X1D_B_0 (
.A0(CLBLM_R_X7Y97_SLICE_X9Y97_AQ),
.A1(CLBLM_R_X7Y97_SLICE_X9Y97_A5Q),
.A2(CLBLM_R_X7Y97_SLICE_X9Y97_BQ),
.A3(CLBLM_R_X7Y97_SLICE_X9Y97_B5Q),
.A4(1'b0),
.D(CLBLM_R_X7Y99_SLICE_X9Y99_AQ),
.DPO(CLBLM_L_X8Y97_SLICE_X10Y97_AO6),
.DPRA0(CLBLM_R_X7Y97_SLICE_X9Y97_AQ),
.DPRA1(CLBLM_R_X7Y97_SLICE_X9Y97_A5Q),
.DPRA2(CLBLM_R_X7Y97_SLICE_X9Y97_BQ),
.DPRA3(CLBLM_R_X7Y97_SLICE_X9Y97_B5Q),
.DPRA4(1'b0),
.SPO(CLBLM_L_X8Y97_SLICE_X10Y97_BO6),
.WCLK(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.WE(CLBLL_L_X4Y97_SLICE_X5Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y97_SLICE_X11Y97_A_FDCE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(1'b1),
.CLR(1'b0),
.D(CLBLM_R_X7Y99_SLICE_X9Y99_DO6),
.Q(CLBLM_L_X8Y97_SLICE_X11Y97_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y97_SLICE_X11Y97_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y97_SLICE_X11Y97_DO5),
.O6(CLBLM_L_X8Y97_SLICE_X11Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff0f0fffff0f0)
  ) CLBLM_L_X8Y97_SLICE_X11Y97_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(1'b1),
.I4(CLBLM_L_X8Y97_SLICE_X11Y97_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y97_SLICE_X11Y97_CO5),
.O6(CLBLM_L_X8Y97_SLICE_X11Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00000000)
  ) CLBLM_L_X8Y97_SLICE_X11Y97_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y97_SLICE_X6Y97_CO6),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X5Y97_SLICE_X7Y97_DO6),
.O5(CLBLM_L_X8Y97_SLICE_X11Y97_BO5),
.O6(CLBLM_L_X8Y97_SLICE_X11Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h40404040808f8f80)
  ) CLBLM_L_X8Y97_SLICE_X11Y97_ALUT (
.I0(CLBLL_L_X4Y97_SLICE_X4Y97_BQ),
.I1(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO7),
.I2(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I3(CLBLM_L_X8Y97_SLICE_X11Y97_BO6),
.I4(CLBLM_L_X8Y97_SLICE_X10Y97_DO6),
.I5(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.O5(CLBLM_L_X8Y97_SLICE_X11Y97_AO5),
.O6(CLBLM_L_X8Y97_SLICE_X11Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff0006600000066)
  ) CLBLM_L_X8Y98_SLICE_X10Y98_DLUT (
.I0(CLBLM_L_X8Y98_SLICE_X10Y98_AO6),
.I1(CLBLM_L_X8Y97_SLICE_X10Y97_BO6),
.I2(CLBLL_L_X4Y97_SLICE_X4Y97_BQ),
.I3(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I4(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I5(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO9),
.O5(CLBLM_L_X8Y98_SLICE_X10Y98_DO5),
.O6(CLBLM_L_X8Y98_SLICE_X10Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c0000050a050a)
  ) CLBLM_L_X8Y98_SLICE_X10Y98_CLUT (
.I0(CLBLM_L_X8Y97_SLICE_X10Y97_AO6),
.I1(CLBLL_L_X4Y97_SLICE_X4Y97_BQ),
.I2(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I3(CLBLM_L_X8Y98_SLICE_X10Y98_AO5),
.I4(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO8),
.I5(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.O5(CLBLM_L_X8Y98_SLICE_X10Y98_CO5),
.O6(CLBLM_L_X8Y98_SLICE_X10Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6ccccccccccccccc)
  ) CLBLM_L_X8Y98_SLICE_X10Y98_BLUT (
.I0(CLBLM_R_X5Y97_SLICE_X6Y97_CO6),
.I1(CLBLM_R_X5Y98_SLICE_X6Y98_AO6),
.I2(CLBLM_L_X8Y97_SLICE_X10Y97_AO6),
.I3(CLBLM_L_X8Y97_SLICE_X10Y97_DO6),
.I4(CLBLM_L_X8Y97_SLICE_X10Y97_BO6),
.I5(CLBLM_R_X5Y97_SLICE_X7Y97_DO6),
.O5(CLBLM_L_X8Y98_SLICE_X10Y98_BO5),
.O6(CLBLM_L_X8Y98_SLICE_X10Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000800088008800)
  ) CLBLM_L_X8Y98_SLICE_X10Y98_ALUT (
.I0(CLBLM_R_X5Y97_SLICE_X7Y97_DO6),
.I1(CLBLM_R_X5Y97_SLICE_X6Y97_CO6),
.I2(CLBLM_L_X8Y97_SLICE_X10Y97_AO6),
.I3(CLBLM_L_X8Y97_SLICE_X10Y97_DO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y98_SLICE_X10Y98_AO5),
.O6(CLBLM_L_X8Y98_SLICE_X10Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y98_SLICE_X11Y98_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y98_SLICE_X11Y98_DO5),
.O6(CLBLM_L_X8Y98_SLICE_X11Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y98_SLICE_X11Y98_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y98_SLICE_X11Y98_CO5),
.O6(CLBLM_L_X8Y98_SLICE_X11Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y98_SLICE_X11Y98_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y98_SLICE_X11Y98_BO5),
.O6(CLBLM_L_X8Y98_SLICE_X11Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y98_SLICE_X11Y98_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y98_SLICE_X11Y98_AO5),
.O6(CLBLM_L_X8Y98_SLICE_X11Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y90_SLICE_X2Y90_A_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLL_L_X2Y93_SLICE_X1Y93_DO6),
.D(CLBLL_L_X4Y92_SLICE_X4Y92_AO6),
.Q(CLBLM_R_X3Y90_SLICE_X2Y90_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y90_SLICE_X2Y90_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y90_SLICE_X2Y90_DO5),
.O6(CLBLM_R_X3Y90_SLICE_X2Y90_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y90_SLICE_X2Y90_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y90_SLICE_X2Y90_CO5),
.O6(CLBLM_R_X3Y90_SLICE_X2Y90_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y90_SLICE_X2Y90_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y90_SLICE_X2Y90_BO5),
.O6(CLBLM_R_X3Y90_SLICE_X2Y90_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y90_SLICE_X2Y90_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y90_SLICE_X2Y90_AO5),
.O6(CLBLM_R_X3Y90_SLICE_X2Y90_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y90_SLICE_X3Y90_A_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLL_L_X2Y92_SLICE_X1Y92_AO6),
.D(CLBLL_L_X4Y92_SLICE_X4Y92_AO5),
.Q(CLBLM_R_X3Y90_SLICE_X3Y90_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y90_SLICE_X3Y90_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y90_SLICE_X3Y90_DO5),
.O6(CLBLM_R_X3Y90_SLICE_X3Y90_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y90_SLICE_X3Y90_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y90_SLICE_X3Y90_CO5),
.O6(CLBLM_R_X3Y90_SLICE_X3Y90_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y90_SLICE_X3Y90_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y90_SLICE_X3Y90_BO5),
.O6(CLBLM_R_X3Y90_SLICE_X3Y90_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y90_SLICE_X3Y90_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y90_SLICE_X3Y90_AO5),
.O6(CLBLM_R_X3Y90_SLICE_X3Y90_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y91_SLICE_X2Y91_B_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X3Y93_SLICE_X3Y93_BO6),
.D(CLBLL_L_X4Y92_SLICE_X4Y92_AO6),
.Q(CLBLM_R_X3Y91_SLICE_X2Y91_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y91_SLICE_X2Y91_D_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X3Y93_SLICE_X3Y93_BO6),
.D(CLBLL_L_X4Y92_SLICE_X4Y92_AO5),
.Q(CLBLM_R_X3Y91_SLICE_X2Y91_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbf3c08888f3c0)
  ) CLBLM_R_X3Y91_SLICE_X2Y91_DLUT (
.I0(CLBLL_L_X2Y91_SLICE_X1Y91_BQ),
.I1(CLBLM_R_X3Y96_SLICE_X3Y96_AO6),
.I2(CLBLL_L_X2Y90_SLICE_X1Y90_AQ),
.I3(CLBLM_R_X5Y92_SLICE_X6Y92_AQ),
.I4(CLBLL_L_X4Y91_SLICE_X4Y91_AO6),
.I5(CLBLL_L_X2Y92_SLICE_X1Y92_BQ),
.O5(CLBLM_R_X3Y91_SLICE_X2Y91_DO5),
.O6(CLBLM_R_X3Y91_SLICE_X2Y91_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfb73ea62d951c840)
  ) CLBLM_R_X3Y91_SLICE_X2Y91_CLUT (
.I0(CLBLL_L_X4Y91_SLICE_X4Y91_AO6),
.I1(CLBLM_R_X3Y96_SLICE_X3Y96_AO6),
.I2(CLBLL_L_X2Y91_SLICE_X0Y91_AQ),
.I3(CLBLM_R_X3Y90_SLICE_X2Y90_AQ),
.I4(CLBLM_R_X3Y91_SLICE_X2Y91_BQ),
.I5(CLBLM_R_X3Y91_SLICE_X3Y91_BQ),
.O5(CLBLM_R_X3Y91_SLICE_X2Y91_CO5),
.O6(CLBLM_R_X3Y91_SLICE_X2Y91_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbd97351eac86240)
  ) CLBLM_R_X3Y91_SLICE_X2Y91_BLUT (
.I0(CLBLL_L_X4Y91_SLICE_X5Y91_F7AMUX_O),
.I1(CLBLM_R_X5Y93_SLICE_X6Y93_F7AMUX_O),
.I2(CLBLL_L_X2Y90_SLICE_X1Y90_AQ),
.I3(CLBLL_L_X2Y92_SLICE_X1Y92_BQ),
.I4(CLBLL_L_X2Y91_SLICE_X1Y91_BQ),
.I5(CLBLM_R_X5Y92_SLICE_X6Y92_AQ),
.O5(CLBLM_R_X3Y91_SLICE_X2Y91_BO5),
.O6(CLBLM_R_X3Y91_SLICE_X2Y91_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0acac0f00acac)
  ) CLBLM_R_X3Y91_SLICE_X2Y91_ALUT (
.I0(CLBLL_L_X2Y91_SLICE_X0Y91_AQ),
.I1(CLBLM_R_X3Y91_SLICE_X2Y91_BQ),
.I2(CLBLM_R_X5Y93_SLICE_X6Y93_F7AMUX_O),
.I3(CLBLM_R_X3Y91_SLICE_X3Y91_BQ),
.I4(CLBLL_L_X4Y91_SLICE_X5Y91_F7AMUX_O),
.I5(CLBLM_R_X3Y90_SLICE_X2Y90_AQ),
.O5(CLBLM_R_X3Y91_SLICE_X2Y91_AO5),
.O6(CLBLM_R_X3Y91_SLICE_X2Y91_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_R_X3Y91_SLICE_X2Y91_MUXF7A (
.I0(CLBLM_R_X3Y91_SLICE_X2Y91_BO6),
.I1(CLBLM_R_X3Y91_SLICE_X2Y91_AO6),
.O(CLBLM_R_X3Y91_SLICE_X2Y91_F7AMUX_O),
.S(CLBLL_L_X2Y93_SLICE_X0Y93_F7AMUX_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_R_X3Y91_SLICE_X2Y91_MUXF7B (
.I0(CLBLM_R_X3Y91_SLICE_X2Y91_DO6),
.I1(CLBLM_R_X3Y91_SLICE_X2Y91_CO6),
.O(CLBLM_R_X3Y91_SLICE_X2Y91_F7BMUX_O),
.S(CLBLL_L_X4Y95_SLICE_X5Y95_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y91_SLICE_X3Y91_B_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X3Y93_SLICE_X3Y93_CO6),
.D(CLBLL_L_X4Y92_SLICE_X4Y92_AO6),
.Q(CLBLM_R_X3Y91_SLICE_X3Y91_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y91_SLICE_X3Y91_D_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X3Y93_SLICE_X3Y93_CO6),
.D(CLBLL_L_X4Y92_SLICE_X4Y92_AO5),
.Q(CLBLM_R_X3Y91_SLICE_X3Y91_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccf0aaffaa00)
  ) CLBLM_R_X3Y91_SLICE_X3Y91_DLUT (
.I0(CLBLM_R_X3Y90_SLICE_X3Y90_AQ),
.I1(CLBLL_L_X4Y91_SLICE_X4Y91_BQ),
.I2(CLBLL_L_X4Y92_SLICE_X4Y92_DQ),
.I3(CLBLM_R_X3Y96_SLICE_X3Y96_AO6),
.I4(CLBLM_R_X5Y92_SLICE_X6Y92_BQ),
.I5(CLBLL_L_X4Y91_SLICE_X4Y91_AO6),
.O5(CLBLM_R_X3Y91_SLICE_X3Y91_DO5),
.O6(CLBLM_R_X3Y91_SLICE_X3Y91_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcbbfc8830bb3088)
  ) CLBLM_R_X3Y91_SLICE_X3Y91_CLUT (
.I0(CLBLL_L_X4Y91_SLICE_X5Y91_BQ),
.I1(CLBLM_R_X3Y96_SLICE_X3Y96_AO6),
.I2(CLBLM_R_X3Y91_SLICE_X3Y91_DQ),
.I3(CLBLL_L_X4Y91_SLICE_X4Y91_AO6),
.I4(CLBLM_R_X3Y91_SLICE_X2Y91_DQ),
.I5(CLBLM_R_X3Y92_SLICE_X3Y92_BQ),
.O5(CLBLM_R_X3Y91_SLICE_X3Y91_CO5),
.O6(CLBLM_R_X3Y91_SLICE_X3Y91_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafadd885050dd88)
  ) CLBLM_R_X3Y91_SLICE_X3Y91_BLUT (
.I0(CLBLL_L_X4Y91_SLICE_X5Y91_F7AMUX_O),
.I1(CLBLL_L_X4Y92_SLICE_X4Y92_DQ),
.I2(CLBLM_R_X3Y90_SLICE_X3Y90_AQ),
.I3(CLBLM_R_X5Y92_SLICE_X6Y92_BQ),
.I4(CLBLM_R_X5Y93_SLICE_X6Y93_F7AMUX_O),
.I5(CLBLL_L_X4Y91_SLICE_X4Y91_BQ),
.O5(CLBLM_R_X3Y91_SLICE_X3Y91_BO5),
.O6(CLBLM_R_X3Y91_SLICE_X3Y91_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0fafacfc00a0a)
  ) CLBLM_R_X3Y91_SLICE_X3Y91_ALUT (
.I0(CLBLM_R_X3Y91_SLICE_X2Y91_DQ),
.I1(CLBLM_R_X3Y92_SLICE_X3Y92_BQ),
.I2(CLBLL_L_X4Y91_SLICE_X5Y91_F7AMUX_O),
.I3(CLBLL_L_X4Y91_SLICE_X5Y91_BQ),
.I4(CLBLM_R_X5Y93_SLICE_X6Y93_F7AMUX_O),
.I5(CLBLM_R_X3Y91_SLICE_X3Y91_DQ),
.O5(CLBLM_R_X3Y91_SLICE_X3Y91_AO5),
.O6(CLBLM_R_X3Y91_SLICE_X3Y91_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_R_X3Y91_SLICE_X3Y91_MUXF7A (
.I0(CLBLM_R_X3Y91_SLICE_X3Y91_BO6),
.I1(CLBLM_R_X3Y91_SLICE_X3Y91_AO6),
.O(CLBLM_R_X3Y91_SLICE_X3Y91_F7AMUX_O),
.S(CLBLL_L_X2Y93_SLICE_X0Y93_F7AMUX_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_R_X3Y91_SLICE_X3Y91_MUXF7B (
.I0(CLBLM_R_X3Y91_SLICE_X3Y91_DO6),
.I1(CLBLM_R_X3Y91_SLICE_X3Y91_CO6),
.O(CLBLM_R_X3Y91_SLICE_X3Y91_F7BMUX_O),
.S(CLBLL_L_X4Y95_SLICE_X5Y95_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y92_SLICE_X2Y92_B_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X3Y93_SLICE_X3Y93_CO6),
.D(CLBLM_R_X3Y94_SLICE_X2Y94_DO6),
.Q(CLBLM_R_X3Y92_SLICE_X2Y92_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y92_SLICE_X2Y92_D_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X3Y93_SLICE_X3Y93_CO6),
.D(CLBLL_L_X4Y94_SLICE_X4Y94_CO5),
.Q(CLBLM_R_X3Y92_SLICE_X2Y92_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdecb9a875643120)
  ) CLBLM_R_X3Y92_SLICE_X2Y92_DLUT (
.I0(CLBLL_L_X4Y91_SLICE_X4Y91_AO6),
.I1(CLBLM_R_X3Y96_SLICE_X3Y96_AO6),
.I2(CLBLL_L_X2Y92_SLICE_X1Y92_CQ),
.I3(CLBLM_R_X3Y94_SLICE_X2Y94_CQ),
.I4(CLBLL_L_X2Y94_SLICE_X1Y94_DQ),
.I5(CLBLL_L_X2Y91_SLICE_X1Y91_CQ),
.O5(CLBLM_R_X3Y92_SLICE_X2Y92_DO5),
.O6(CLBLM_R_X3Y92_SLICE_X2Y92_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc30fc30bbbb8888)
  ) CLBLM_R_X3Y92_SLICE_X2Y92_CLUT (
.I0(CLBLL_L_X2Y92_SLICE_X0Y92_AQ),
.I1(CLBLM_R_X3Y96_SLICE_X3Y96_AO6),
.I2(CLBLM_R_X3Y92_SLICE_X2Y92_DQ),
.I3(CLBLM_R_X3Y92_SLICE_X3Y92_CQ),
.I4(CLBLM_R_X3Y93_SLICE_X2Y93_CQ),
.I5(CLBLL_L_X4Y91_SLICE_X4Y91_AO6),
.O5(CLBLM_R_X3Y92_SLICE_X2Y92_CO5),
.O6(CLBLM_R_X3Y92_SLICE_X2Y92_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ccccaaaaf0f0)
  ) CLBLM_R_X3Y92_SLICE_X2Y92_BLUT (
.I0(CLBLL_L_X2Y94_SLICE_X1Y94_DQ),
.I1(CLBLL_L_X2Y92_SLICE_X1Y92_CQ),
.I2(CLBLM_R_X3Y94_SLICE_X2Y94_CQ),
.I3(CLBLL_L_X2Y91_SLICE_X1Y91_CQ),
.I4(CLBLM_R_X5Y93_SLICE_X6Y93_F7AMUX_O),
.I5(CLBLL_L_X4Y91_SLICE_X5Y91_F7AMUX_O),
.O5(CLBLM_R_X3Y92_SLICE_X2Y92_BO5),
.O6(CLBLM_R_X3Y92_SLICE_X2Y92_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfafc0a0cfa0c0a)
  ) CLBLM_R_X3Y92_SLICE_X2Y92_ALUT (
.I0(CLBLM_R_X3Y93_SLICE_X2Y93_CQ),
.I1(CLBLM_R_X3Y92_SLICE_X2Y92_DQ),
.I2(CLBLM_R_X5Y93_SLICE_X6Y93_F7AMUX_O),
.I3(CLBLL_L_X4Y91_SLICE_X5Y91_F7AMUX_O),
.I4(CLBLL_L_X2Y92_SLICE_X0Y92_AQ),
.I5(CLBLM_R_X3Y92_SLICE_X3Y92_CQ),
.O5(CLBLM_R_X3Y92_SLICE_X2Y92_AO5),
.O6(CLBLM_R_X3Y92_SLICE_X2Y92_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_R_X3Y92_SLICE_X2Y92_MUXF7A (
.I0(CLBLM_R_X3Y92_SLICE_X2Y92_BO6),
.I1(CLBLM_R_X3Y92_SLICE_X2Y92_AO6),
.O(CLBLM_R_X3Y92_SLICE_X2Y92_F7AMUX_O),
.S(CLBLL_L_X2Y93_SLICE_X0Y93_F7AMUX_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_R_X3Y92_SLICE_X2Y92_MUXF7B (
.I0(CLBLM_R_X3Y92_SLICE_X2Y92_DO6),
.I1(CLBLM_R_X3Y92_SLICE_X2Y92_CO6),
.O(CLBLM_R_X3Y92_SLICE_X2Y92_F7BMUX_O),
.S(CLBLL_L_X4Y95_SLICE_X5Y95_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y92_SLICE_X3Y92_A_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLL_L_X2Y93_SLICE_X1Y93_DO6),
.D(CLBLM_R_X3Y94_SLICE_X2Y94_DO5),
.Q(CLBLM_R_X3Y92_SLICE_X3Y92_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y92_SLICE_X3Y92_B_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLL_L_X2Y93_SLICE_X1Y93_DO6),
.D(CLBLL_L_X4Y92_SLICE_X4Y92_AO5),
.Q(CLBLM_R_X3Y92_SLICE_X3Y92_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y92_SLICE_X3Y92_C_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLL_L_X2Y93_SLICE_X1Y93_DO6),
.D(CLBLL_L_X4Y94_SLICE_X4Y94_CO5),
.Q(CLBLM_R_X3Y92_SLICE_X3Y92_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y92_SLICE_X3Y92_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y92_SLICE_X3Y92_DO5),
.O6(CLBLM_R_X3Y92_SLICE_X3Y92_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y92_SLICE_X3Y92_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y92_SLICE_X3Y92_CO5),
.O6(CLBLM_R_X3Y92_SLICE_X3Y92_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y92_SLICE_X3Y92_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y92_SLICE_X3Y92_BO5),
.O6(CLBLM_R_X3Y92_SLICE_X3Y92_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y92_SLICE_X3Y92_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y92_SLICE_X3Y92_AO5),
.O6(CLBLM_R_X3Y92_SLICE_X3Y92_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y93_SLICE_X2Y93_B_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X3Y93_SLICE_X3Y93_BO6),
.D(CLBLM_R_X3Y94_SLICE_X2Y94_DO6),
.Q(CLBLM_R_X3Y93_SLICE_X2Y93_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y93_SLICE_X2Y93_C_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X3Y93_SLICE_X3Y93_BO6),
.D(CLBLL_L_X4Y94_SLICE_X4Y94_CO5),
.Q(CLBLM_R_X3Y93_SLICE_X2Y93_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000400)
  ) CLBLM_R_X3Y93_SLICE_X2Y93_DLUT (
.I0(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO15),
.I1(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO10),
.I2(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO12),
.I3(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO13),
.I4(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO14),
.I5(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO11),
.O5(CLBLM_R_X3Y93_SLICE_X2Y93_DO5),
.O6(CLBLM_R_X3Y93_SLICE_X2Y93_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0d4db4a001010030)
  ) CLBLM_R_X3Y93_SLICE_X2Y93_CLUT (
.I0(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I1(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I2(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I3(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I4(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y93_SLICE_X2Y93_CO5),
.O6(CLBLM_R_X3Y93_SLICE_X2Y93_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbf388f3bbc088c0)
  ) CLBLM_R_X3Y93_SLICE_X2Y93_BLUT (
.I0(CLBLL_L_X2Y91_SLICE_X1Y91_AQ),
.I1(CLBLL_L_X4Y91_SLICE_X4Y91_AO6),
.I2(CLBLL_L_X2Y92_SLICE_X1Y92_AQ),
.I3(CLBLM_R_X3Y96_SLICE_X3Y96_AO6),
.I4(CLBLL_L_X2Y94_SLICE_X1Y94_BQ),
.I5(CLBLM_R_X3Y94_SLICE_X2Y94_AQ),
.O5(CLBLM_R_X3Y93_SLICE_X2Y93_BO5),
.O6(CLBLM_R_X3Y93_SLICE_X2Y93_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa00aaf0ccf0cc)
  ) CLBLM_R_X3Y93_SLICE_X2Y93_ALUT (
.I0(CLBLL_L_X2Y93_SLICE_X0Y93_BQ),
.I1(CLBLM_R_X3Y93_SLICE_X2Y93_BQ),
.I2(CLBLM_R_X3Y92_SLICE_X2Y92_BQ),
.I3(CLBLL_L_X4Y91_SLICE_X4Y91_AO6),
.I4(CLBLL_L_X2Y93_SLICE_X1Y93_BQ),
.I5(CLBLM_R_X3Y96_SLICE_X3Y96_AO6),
.O5(CLBLM_R_X3Y93_SLICE_X2Y93_AO5),
.O6(CLBLM_R_X3Y93_SLICE_X2Y93_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_R_X3Y93_SLICE_X2Y93_MUXF7A (
.I0(CLBLM_R_X3Y93_SLICE_X2Y93_BO6),
.I1(CLBLM_R_X3Y93_SLICE_X2Y93_AO6),
.O(CLBLM_R_X3Y93_SLICE_X2Y93_F7AMUX_O),
.S(CLBLL_L_X4Y95_SLICE_X5Y95_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y93_SLICE_X3Y93_A_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X3Y93_SLICE_X3Y93_BO6),
.D(CLBLL_L_X4Y93_SLICE_X4Y93_CO5),
.Q(CLBLM_R_X3Y93_SLICE_X3Y93_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y93_SLICE_X3Y93_B_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X3Y93_SLICE_X3Y93_BO6),
.D(CLBLM_R_X3Y94_SLICE_X2Y94_DO5),
.Q(CLBLM_R_X3Y93_SLICE_X3Y93_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y93_SLICE_X3Y93_C_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X3Y93_SLICE_X3Y93_BO6),
.D(CLBLL_L_X4Y93_SLICE_X4Y93_CO6),
.Q(CLBLM_R_X3Y93_SLICE_X3Y93_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y93_SLICE_X3Y93_D_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X3Y93_SLICE_X3Y93_BO6),
.D(CLBLL_L_X4Y94_SLICE_X4Y94_CO6),
.Q(CLBLM_R_X3Y93_SLICE_X3Y93_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y93_SLICE_X3Y93_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y93_SLICE_X3Y93_DO5),
.O6(CLBLM_R_X3Y93_SLICE_X3Y93_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000a000a000)
  ) CLBLM_R_X3Y93_SLICE_X3Y93_CLUT (
.I0(CLBLL_L_X2Y93_SLICE_X0Y93_CO6),
.I1(1'b1),
.I2(CLBLL_L_X4Y94_SLICE_X5Y94_DO6),
.I3(CLBLM_R_X5Y94_SLICE_X7Y94_DO6),
.I4(1'b1),
.I5(CLBLM_R_X5Y94_SLICE_X6Y94_BO6),
.O5(CLBLM_R_X3Y93_SLICE_X3Y93_CO5),
.O6(CLBLM_R_X3Y93_SLICE_X3Y93_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000000cc00)
  ) CLBLM_R_X3Y93_SLICE_X3Y93_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X2Y93_SLICE_X0Y93_CO6),
.I2(1'b1),
.I3(CLBLL_L_X4Y94_SLICE_X5Y94_DO6),
.I4(CLBLM_R_X5Y94_SLICE_X6Y94_BO6),
.I5(CLBLM_R_X5Y94_SLICE_X7Y94_DO6),
.O5(CLBLM_R_X3Y93_SLICE_X3Y93_BO5),
.O6(CLBLM_R_X3Y93_SLICE_X3Y93_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffedffedffffef73)
  ) CLBLM_R_X3Y93_SLICE_X3Y93_ALUT (
.I0(CLBLM_R_X3Y95_SLICE_X3Y95_DO6),
.I1(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I2(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I3(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I4(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I5(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.O5(CLBLM_R_X3Y93_SLICE_X3Y93_AO5),
.O6(CLBLM_R_X3Y93_SLICE_X3Y93_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y94_SLICE_X2Y94_A_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(1'b1),
.D(CLBLM_R_X3Y94_SLICE_X2Y94_AO6),
.Q(CLBLM_R_X3Y94_SLICE_X2Y94_AQ),
.R(CLBLM_R_X5Y92_SLICE_X7Y92_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y94_SLICE_X2Y94_B_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(1'b1),
.D(CLBLM_R_X3Y94_SLICE_X2Y94_BO6),
.Q(CLBLM_R_X3Y94_SLICE_X2Y94_BQ),
.R(CLBLM_R_X5Y92_SLICE_X7Y92_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y94_SLICE_X2Y94_C_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(1'b1),
.D(CLBLM_R_X3Y94_SLICE_X2Y94_CO6),
.Q(CLBLM_R_X3Y94_SLICE_X2Y94_CQ),
.R(CLBLM_R_X5Y92_SLICE_X7Y92_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa00ccf0ccf0)
  ) CLBLM_R_X3Y94_SLICE_X2Y94_DLUT (
.I0(CLBLL_L_X2Y97_SLICE_X1Y97_AO6),
.I1(CLBLL_L_X2Y97_SLICE_X0Y97_CO6),
.I2(CLBLM_R_X3Y99_SLICE_X2Y99_DO6),
.I3(CLBLM_R_X3Y93_SLICE_X2Y93_CO6),
.I4(CLBLM_R_X3Y98_SLICE_X2Y98_BO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y94_SLICE_X2Y94_DO5),
.O6(CLBLM_R_X3Y94_SLICE_X2Y94_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000010111000)
  ) CLBLM_R_X3Y94_SLICE_X2Y94_CLUT (
.I0(CLBLM_R_X5Y94_SLICE_X6Y94_BO6),
.I1(CLBLL_L_X4Y94_SLICE_X5Y94_DO6),
.I2(CLBLL_L_X2Y96_SLICE_X1Y96_DO6),
.I3(CLBLM_R_X3Y93_SLICE_X2Y93_CO6),
.I4(CLBLM_R_X3Y96_SLICE_X3Y96_DO6),
.I5(CLBLM_R_X5Y94_SLICE_X7Y94_DO6),
.O5(CLBLM_R_X3Y94_SLICE_X2Y94_CO5),
.O6(CLBLM_R_X3Y94_SLICE_X2Y94_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000003200000002)
  ) CLBLM_R_X3Y94_SLICE_X2Y94_BLUT (
.I0(CLBLM_R_X3Y99_SLICE_X2Y99_DO6),
.I1(CLBLL_L_X4Y94_SLICE_X5Y94_DO6),
.I2(CLBLM_R_X3Y93_SLICE_X2Y93_CO6),
.I3(CLBLM_R_X5Y94_SLICE_X7Y94_DO6),
.I4(CLBLM_R_X5Y94_SLICE_X6Y94_BO6),
.I5(CLBLL_L_X2Y97_SLICE_X0Y97_CO6),
.O5(CLBLM_R_X3Y94_SLICE_X2Y94_BO5),
.O6(CLBLM_R_X3Y94_SLICE_X2Y94_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000320002)
  ) CLBLM_R_X3Y94_SLICE_X2Y94_ALUT (
.I0(CLBLM_R_X3Y98_SLICE_X2Y98_BO6),
.I1(CLBLM_R_X5Y94_SLICE_X6Y94_BO6),
.I2(CLBLM_R_X3Y93_SLICE_X2Y93_CO6),
.I3(CLBLM_R_X5Y94_SLICE_X7Y94_DO6),
.I4(CLBLL_L_X2Y97_SLICE_X1Y97_AO6),
.I5(CLBLL_L_X4Y94_SLICE_X5Y94_DO6),
.O5(CLBLM_R_X3Y94_SLICE_X2Y94_AO5),
.O6(CLBLM_R_X3Y94_SLICE_X2Y94_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y94_SLICE_X3Y94_B_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X3Y93_SLICE_X3Y93_CO6),
.D(CLBLM_R_X3Y94_SLICE_X2Y94_DO5),
.Q(CLBLM_R_X3Y94_SLICE_X3Y94_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacff0facacf000)
  ) CLBLM_R_X3Y94_SLICE_X3Y94_DLUT (
.I0(CLBLL_L_X4Y93_SLICE_X4Y93_BQ),
.I1(CLBLL_L_X4Y92_SLICE_X4Y92_BQ),
.I2(CLBLM_R_X3Y96_SLICE_X3Y96_AO6),
.I3(CLBLL_L_X2Y94_SLICE_X1Y94_CQ),
.I4(CLBLL_L_X4Y91_SLICE_X4Y91_AO6),
.I5(CLBLM_R_X3Y94_SLICE_X2Y94_BQ),
.O5(CLBLM_R_X3Y94_SLICE_X3Y94_DO5),
.O6(CLBLM_R_X3Y94_SLICE_X3Y94_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfadd50ddfa885088)
  ) CLBLM_R_X3Y94_SLICE_X3Y94_CLUT (
.I0(CLBLM_R_X3Y96_SLICE_X3Y96_AO6),
.I1(CLBLL_L_X2Y93_SLICE_X0Y93_CQ),
.I2(CLBLM_R_X3Y94_SLICE_X3Y94_BQ),
.I3(CLBLL_L_X4Y91_SLICE_X4Y91_AO6),
.I4(CLBLM_R_X3Y92_SLICE_X3Y92_AQ),
.I5(CLBLM_R_X3Y93_SLICE_X3Y93_BQ),
.O5(CLBLM_R_X3Y94_SLICE_X3Y94_CO5),
.O6(CLBLM_R_X3Y94_SLICE_X3Y94_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdf85d58ada80d08)
  ) CLBLM_R_X3Y94_SLICE_X3Y94_BLUT (
.I0(CLBLM_R_X5Y93_SLICE_X6Y93_F7AMUX_O),
.I1(CLBLL_L_X2Y94_SLICE_X1Y94_CQ),
.I2(CLBLL_L_X4Y91_SLICE_X5Y91_F7AMUX_O),
.I3(CLBLM_R_X3Y94_SLICE_X2Y94_BQ),
.I4(CLBLL_L_X4Y93_SLICE_X4Y93_BQ),
.I5(CLBLL_L_X4Y92_SLICE_X4Y92_BQ),
.O5(CLBLM_R_X3Y94_SLICE_X3Y94_BO5),
.O6(CLBLM_R_X3Y94_SLICE_X3Y94_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hefea4f4ae5e04540)
  ) CLBLM_R_X3Y94_SLICE_X3Y94_ALUT (
.I0(CLBLM_R_X5Y93_SLICE_X6Y93_F7AMUX_O),
.I1(CLBLM_R_X3Y94_SLICE_X3Y94_BQ),
.I2(CLBLL_L_X4Y91_SLICE_X5Y91_F7AMUX_O),
.I3(CLBLM_R_X3Y93_SLICE_X3Y93_BQ),
.I4(CLBLM_R_X3Y92_SLICE_X3Y92_AQ),
.I5(CLBLL_L_X2Y93_SLICE_X0Y93_CQ),
.O5(CLBLM_R_X3Y94_SLICE_X3Y94_AO5),
.O6(CLBLM_R_X3Y94_SLICE_X3Y94_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_R_X3Y94_SLICE_X3Y94_MUXF7A (
.I0(CLBLM_R_X3Y94_SLICE_X3Y94_BO6),
.I1(CLBLM_R_X3Y94_SLICE_X3Y94_AO6),
.O(CLBLM_R_X3Y94_SLICE_X3Y94_F7AMUX_O),
.S(CLBLL_L_X2Y93_SLICE_X0Y93_F7AMUX_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_R_X3Y94_SLICE_X3Y94_MUXF7B (
.I0(CLBLM_R_X3Y94_SLICE_X3Y94_DO6),
.I1(CLBLM_R_X3Y94_SLICE_X3Y94_CO6),
.O(CLBLM_R_X3Y94_SLICE_X3Y94_F7BMUX_O),
.S(CLBLL_L_X4Y95_SLICE_X5Y95_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe0ef434f808cb0b)
  ) CLBLM_R_X3Y95_SLICE_X2Y95_DLUT (
.I0(CLBLL_L_X4Y91_SLICE_X4Y91_BO6),
.I1(CLBLM_R_X3Y93_SLICE_X2Y93_CO5),
.I2(CLBLL_L_X2Y93_SLICE_X0Y93_CO5),
.I3(CLBLL_L_X2Y95_SLICE_X1Y95_B_XOR),
.I4(CLBLL_L_X2Y97_SLICE_X0Y97_AO6),
.I5(CLBLM_R_X3Y91_SLICE_X3Y91_F7AMUX_O),
.O5(CLBLM_R_X3Y95_SLICE_X2Y95_DO5),
.O6(CLBLM_R_X3Y95_SLICE_X2Y95_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeae5426ead94051)
  ) CLBLM_R_X3Y95_SLICE_X2Y95_CLUT (
.I0(CLBLL_L_X2Y93_SLICE_X0Y93_CO5),
.I1(CLBLM_R_X3Y93_SLICE_X2Y93_CO5),
.I2(CLBLM_R_X3Y95_SLICE_X3Y95_AO6),
.I3(CLBLL_L_X2Y97_SLICE_X0Y97_AO6),
.I4(CLBLL_L_X2Y95_SLICE_X1Y95_A_XOR),
.I5(CLBLM_R_X3Y91_SLICE_X2Y91_F7AMUX_O),
.O5(CLBLM_R_X3Y95_SLICE_X2Y95_CO5),
.O6(CLBLM_R_X3Y95_SLICE_X2Y95_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfaa0dd880af5)
  ) CLBLM_R_X3Y95_SLICE_X2Y95_BLUT (
.I0(CLBLM_R_X3Y93_SLICE_X2Y93_CO5),
.I1(CLBLL_L_X2Y94_SLICE_X1Y94_D_XOR),
.I2(CLBLL_L_X4Y95_SLICE_X4Y95_BO6),
.I3(CLBLL_L_X4Y93_SLICE_X4Y93_F7AMUX_O),
.I4(CLBLL_L_X2Y93_SLICE_X0Y93_CO5),
.I5(CLBLL_L_X2Y97_SLICE_X0Y97_AO6),
.O5(CLBLM_R_X3Y95_SLICE_X2Y95_BO5),
.O6(CLBLM_R_X3Y95_SLICE_X2Y95_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffdffdfffb9efdb)
  ) CLBLM_R_X3Y95_SLICE_X2Y95_ALUT (
.I0(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I1(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I2(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I3(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I4(CLBLL_L_X4Y91_SLICE_X4Y91_BO6),
.I5(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.O5(CLBLM_R_X3Y95_SLICE_X2Y95_AO5),
.O6(CLBLM_R_X3Y95_SLICE_X2Y95_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0d8f0f0f0f0)
  ) CLBLM_R_X3Y95_SLICE_X3Y95_DLUT (
.I0(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I1(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO2),
.I2(CLBLM_R_X3Y94_SLICE_X3Y94_F7BMUX_O),
.I3(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I4(CLBLL_L_X4Y91_SLICE_X4Y91_AO5),
.I5(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.O5(CLBLM_R_X3Y95_SLICE_X3Y95_DO5),
.O6(CLBLM_R_X3Y95_SLICE_X3Y95_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffdcffa5efff)
  ) CLBLM_R_X3Y95_SLICE_X3Y95_CLUT (
.I0(CLBLM_R_X3Y95_SLICE_X3Y95_AO6),
.I1(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I2(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I3(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I4(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I5(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.O5(CLBLM_R_X3Y95_SLICE_X3Y95_CO5),
.O6(CLBLM_R_X3Y95_SLICE_X3Y95_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0e2f0f0f0)
  ) CLBLM_R_X3Y95_SLICE_X3Y95_BLUT (
.I0(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO7),
.I1(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I2(CLBLM_R_X3Y92_SLICE_X2Y92_F7BMUX_O),
.I3(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I4(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I5(CLBLL_L_X4Y91_SLICE_X4Y91_AO5),
.O5(CLBLM_R_X3Y95_SLICE_X3Y95_BO5),
.O6(CLBLM_R_X3Y95_SLICE_X3Y95_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1f0f0f0e0f0f0f0)
  ) CLBLM_R_X3Y95_SLICE_X3Y95_ALUT (
.I0(CLBLL_L_X4Y91_SLICE_X4Y91_AO5),
.I1(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I2(CLBLM_R_X3Y91_SLICE_X2Y91_F7BMUX_O),
.I3(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I4(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I5(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO4),
.O5(CLBLM_R_X3Y95_SLICE_X3Y95_AO5),
.O6(CLBLM_R_X3Y95_SLICE_X3Y95_AO6)
  );


  (* KEEP, DONT_TOUCH *)
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000)
  ) CLBLM_R_X3Y96_SLICE_X2Y96_RAM32M (
.ADDRA({CLBLL_L_X4Y98_SLICE_X5Y98_DO6, CLBLM_R_X3Y98_SLICE_X3Y98_DO6, CLBLM_R_X3Y97_SLICE_X3Y97_DO6, CLBLL_L_X4Y98_SLICE_X4Y98_DO6, CLBLM_R_X3Y97_SLICE_X3Y97_CO6}),
.ADDRB({CLBLL_L_X4Y98_SLICE_X5Y98_DO6, CLBLM_R_X3Y98_SLICE_X3Y98_DO6, CLBLM_R_X3Y97_SLICE_X3Y97_DO6, CLBLL_L_X4Y98_SLICE_X4Y98_DO6, CLBLM_R_X3Y97_SLICE_X3Y97_CO6}),
.ADDRC({CLBLL_L_X4Y98_SLICE_X5Y98_DO6, CLBLM_R_X3Y98_SLICE_X3Y98_DO6, CLBLM_R_X3Y97_SLICE_X3Y97_DO6, CLBLL_L_X4Y98_SLICE_X4Y98_DO6, CLBLM_R_X3Y97_SLICE_X3Y97_CO6}),
.ADDRD({CLBLL_L_X4Y98_SLICE_X5Y98_DO6, CLBLM_R_X3Y98_SLICE_X3Y98_DO6, CLBLM_R_X3Y97_SLICE_X3Y97_DO6, CLBLL_L_X4Y98_SLICE_X4Y98_DO6, CLBLM_R_X3Y97_SLICE_X3Y97_CO6}),
.DIA({CLBLL_L_X2Y96_SLICE_X1Y96_BO6, CLBLL_L_X4Y98_SLICE_X4Y98_DO6}),
.DIB({CLBLL_L_X2Y97_SLICE_X1Y97_CO6, CLBLL_L_X4Y98_SLICE_X4Y98_DO6}),
.DIC({CLBLL_L_X2Y96_SLICE_X1Y96_DO6, CLBLL_L_X4Y98_SLICE_X4Y98_DO6}),
.DID({CLBLL_L_X2Y96_SLICE_X1Y96_AO6, CLBLL_L_X4Y98_SLICE_X4Y98_DO6}),
.DOA({CLBLM_R_X3Y96_SLICE_X2Y96_AO6, CLBLM_R_X3Y96_SLICE_X2Y96_AO5}),
.DOB({CLBLM_R_X3Y96_SLICE_X2Y96_BO6, CLBLM_R_X3Y96_SLICE_X2Y96_BO5}),
.DOC({CLBLM_R_X3Y96_SLICE_X2Y96_CO6, CLBLM_R_X3Y96_SLICE_X2Y96_CO5}),
.DOD({CLBLM_R_X3Y96_SLICE_X2Y96_DO6, CLBLM_R_X3Y96_SLICE_X2Y96_DO5}),
.WCLK(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.WE(CLBLM_R_X5Y94_SLICE_X6Y94_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000f000f404)
  ) CLBLM_R_X3Y96_SLICE_X3Y96_DLUT (
.I0(CLBLM_R_X3Y98_SLICE_X3Y98_AO6),
.I1(CLBLM_R_X3Y96_SLICE_X2Y96_CO6),
.I2(CLBLL_L_X4Y97_SLICE_X4Y97_AO6),
.I3(CLBLM_R_X3Y96_SLICE_X3Y96_CO6),
.I4(CLBLL_L_X4Y97_SLICE_X4Y97_CO6),
.I5(CLBLL_L_X4Y98_SLICE_X4Y98_AO6),
.O5(CLBLM_R_X3Y96_SLICE_X3Y96_DO5),
.O6(CLBLM_R_X3Y96_SLICE_X3Y96_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0001000000000000)
  ) CLBLM_R_X3Y96_SLICE_X3Y96_CLUT (
.I0(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I1(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I2(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I3(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I4(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I5(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO7),
.O5(CLBLM_R_X3Y96_SLICE_X3Y96_CO5),
.O6(CLBLM_R_X3Y96_SLICE_X3Y96_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000080c02000c000)
  ) CLBLM_R_X3Y96_SLICE_X3Y96_BLUT (
.I0(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I1(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I2(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I3(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I4(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y96_SLICE_X3Y96_BO5),
.O6(CLBLM_R_X3Y96_SLICE_X3Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h02000208ffffff00)
  ) CLBLM_R_X3Y96_SLICE_X3Y96_ALUT (
.I0(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO6),
.I1(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I2(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I3(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I4(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y96_SLICE_X3Y96_AO5),
.O6(CLBLM_R_X3Y96_SLICE_X3Y96_AO6)
  );


  (* KEEP, DONT_TOUCH *)
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000)
  ) CLBLM_R_X3Y97_SLICE_X2Y97_RAM32M (
.ADDRA({CLBLL_L_X4Y98_SLICE_X5Y98_DO6, CLBLM_R_X3Y98_SLICE_X3Y98_DO6, CLBLM_R_X3Y97_SLICE_X3Y97_DO6, CLBLL_L_X4Y98_SLICE_X4Y98_DO6, CLBLM_R_X3Y97_SLICE_X3Y97_CO6}),
.ADDRB({CLBLL_L_X4Y98_SLICE_X5Y98_DO6, CLBLM_R_X3Y98_SLICE_X3Y98_DO6, CLBLM_R_X3Y97_SLICE_X3Y97_DO6, CLBLL_L_X4Y98_SLICE_X4Y98_DO6, CLBLM_R_X3Y97_SLICE_X3Y97_CO6}),
.ADDRC({CLBLL_L_X4Y98_SLICE_X5Y98_DO6, CLBLM_R_X3Y98_SLICE_X3Y98_DO6, CLBLM_R_X3Y97_SLICE_X3Y97_DO6, CLBLL_L_X4Y98_SLICE_X4Y98_DO6, CLBLM_R_X3Y97_SLICE_X3Y97_CO6}),
.ADDRD({CLBLL_L_X4Y98_SLICE_X5Y98_DO6, CLBLM_R_X3Y98_SLICE_X3Y98_DO6, CLBLM_R_X3Y97_SLICE_X3Y97_DO6, CLBLL_L_X4Y98_SLICE_X4Y98_DO6, CLBLM_R_X3Y97_SLICE_X3Y97_CO6}),
.DIA({CLBLL_L_X2Y97_SLICE_X1Y97_AO6, 1'b1}),
.DIB({CLBLL_L_X2Y97_SLICE_X0Y97_CO6, 1'b1}),
.DIC({CLBLL_L_X2Y97_SLICE_X1Y97_BO6, 1'b1}),
.DID({CLBLL_L_X2Y97_SLICE_X0Y97_BO6, 1'b1}),
.DOA({CLBLM_R_X3Y97_SLICE_X2Y97_AO6, CLBLM_R_X3Y97_SLICE_X2Y97_AO5}),
.DOB({CLBLM_R_X3Y97_SLICE_X2Y97_BO6, CLBLM_R_X3Y97_SLICE_X2Y97_BO5}),
.DOC({CLBLM_R_X3Y97_SLICE_X2Y97_CO6, CLBLM_R_X3Y97_SLICE_X2Y97_CO5}),
.DOD({CLBLM_R_X3Y97_SLICE_X2Y97_DO6, CLBLM_R_X3Y97_SLICE_X2Y97_DO5}),
.WCLK(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.WE(CLBLM_R_X5Y94_SLICE_X6Y94_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0011000100100000)
  ) CLBLM_R_X3Y97_SLICE_X3Y97_DLUT (
.I0(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I1(CLBLL_L_X4Y97_SLICE_X5Y97_AO6),
.I2(CLBLM_R_X3Y96_SLICE_X3Y96_AO5),
.I3(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I4(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO2),
.I5(CLBLM_R_X3Y97_SLICE_X3Y97_BO6),
.O5(CLBLM_R_X3Y97_SLICE_X3Y97_DO5),
.O6(CLBLM_R_X3Y97_SLICE_X3Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000003202)
  ) CLBLM_R_X3Y97_SLICE_X3Y97_CLUT (
.I0(CLBLM_R_X3Y97_SLICE_X3Y97_AO6),
.I1(CLBLL_L_X4Y97_SLICE_X5Y97_AO6),
.I2(CLBLM_R_X3Y96_SLICE_X3Y96_AO5),
.I3(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO0),
.I4(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I5(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.O5(CLBLM_R_X3Y97_SLICE_X3Y97_CO5),
.O6(CLBLM_R_X3Y97_SLICE_X3Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000100200000000)
  ) CLBLM_R_X3Y97_SLICE_X3Y97_BLUT (
.I0(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO13),
.I1(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO15),
.I2(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO12),
.I3(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO11),
.I4(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO14),
.I5(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO2),
.O5(CLBLM_R_X3Y97_SLICE_X3Y97_BO5),
.O6(CLBLM_R_X3Y97_SLICE_X3Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000100200000000)
  ) CLBLM_R_X3Y97_SLICE_X3Y97_ALUT (
.I0(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO13),
.I1(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO15),
.I2(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO12),
.I3(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO11),
.I4(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO14),
.I5(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO0),
.O5(CLBLM_R_X3Y97_SLICE_X3Y97_AO5),
.O6(CLBLM_R_X3Y97_SLICE_X3Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffcfcfcfc)
  ) CLBLM_R_X3Y98_SLICE_X2Y98_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y98_SLICE_X3Y98_AO6),
.I2(CLBLL_L_X4Y97_SLICE_X4Y97_CO6),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X4Y98_SLICE_X4Y98_AO6),
.O5(CLBLM_R_X3Y98_SLICE_X2Y98_DO5),
.O6(CLBLM_R_X3Y98_SLICE_X2Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf0f0aaaaff00)
  ) CLBLM_R_X3Y98_SLICE_X2Y98_CLUT (
.I0(CLBLM_R_X3Y98_SLICE_X2Y98_AO6),
.I1(1'b1),
.I2(CLBLL_L_X2Y99_SLICE_X1Y99_AQ),
.I3(CLBLM_R_X3Y97_SLICE_X2Y97_CO6),
.I4(CLBLL_L_X4Y97_SLICE_X4Y97_AO6),
.I5(CLBLM_R_X3Y98_SLICE_X2Y98_DO6),
.O5(CLBLM_R_X3Y98_SLICE_X2Y98_CO5),
.O6(CLBLM_R_X3Y98_SLICE_X2Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfa50ccccfa50)
  ) CLBLM_R_X3Y98_SLICE_X2Y98_BLUT (
.I0(CLBLM_R_X3Y98_SLICE_X2Y98_DO6),
.I1(CLBLL_L_X4Y98_SLICE_X5Y98_BO6),
.I2(CLBLM_R_X3Y97_SLICE_X2Y97_AO6),
.I3(CLBLL_L_X2Y98_SLICE_X0Y98_AQ),
.I4(CLBLL_L_X4Y97_SLICE_X4Y97_AO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y98_SLICE_X2Y98_BO5),
.O6(CLBLM_R_X3Y98_SLICE_X2Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000200)
  ) CLBLM_R_X3Y98_SLICE_X2Y98_ALUT (
.I0(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO3),
.I1(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I2(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I3(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I4(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I5(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.O5(CLBLM_R_X3Y98_SLICE_X2Y98_AO5),
.O6(CLBLM_R_X3Y98_SLICE_X2Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000010101100)
  ) CLBLM_R_X3Y98_SLICE_X3Y98_DLUT (
.I0(CLBLL_L_X4Y97_SLICE_X5Y97_AO6),
.I1(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I2(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO3),
.I3(CLBLM_R_X3Y98_SLICE_X3Y98_CO6),
.I4(CLBLM_R_X3Y96_SLICE_X3Y96_AO5),
.I5(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.O5(CLBLM_R_X3Y98_SLICE_X3Y98_DO5),
.O6(CLBLM_R_X3Y98_SLICE_X3Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000010000020)
  ) CLBLM_R_X3Y98_SLICE_X3Y98_CLUT (
.I0(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO13),
.I1(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO14),
.I2(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO3),
.I3(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO11),
.I4(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO12),
.I5(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO15),
.O5(CLBLM_R_X3Y98_SLICE_X3Y98_CO5),
.O6(CLBLM_R_X3Y98_SLICE_X3Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000040080)
  ) CLBLM_R_X3Y98_SLICE_X3Y98_BLUT (
.I0(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO12),
.I1(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO7),
.I2(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO11),
.I3(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO15),
.I4(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO13),
.I5(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO14),
.O5(CLBLM_R_X3Y98_SLICE_X3Y98_BO5),
.O6(CLBLM_R_X3Y98_SLICE_X3Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000d08)
  ) CLBLM_R_X3Y98_SLICE_X3Y98_ALUT (
.I0(CLBLM_R_X3Y96_SLICE_X3Y96_AO5),
.I1(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO7),
.I2(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I3(CLBLM_R_X3Y98_SLICE_X3Y98_BO6),
.I4(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I5(CLBLL_L_X4Y97_SLICE_X5Y97_AO6),
.O5(CLBLM_R_X3Y98_SLICE_X3Y98_AO5),
.O6(CLBLM_R_X3Y98_SLICE_X3Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y99_SLICE_X2Y99_A_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(LIOB33_X0Y109_IOB_X0Y109_I),
.D(LIOB33_X0Y109_IOB_X0Y109_I),
.Q(CLBLM_R_X3Y99_SLICE_X2Y99_AQ),
.R(CLBLL_L_X2Y98_SLICE_X1Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heefaeefa44504450)
  ) CLBLM_R_X3Y99_SLICE_X2Y99_DLUT (
.I0(CLBLL_L_X4Y97_SLICE_X4Y97_AO6),
.I1(CLBLM_R_X3Y99_SLICE_X2Y99_AQ),
.I2(CLBLM_R_X3Y97_SLICE_X2Y97_BO6),
.I3(CLBLM_R_X3Y98_SLICE_X2Y98_DO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y99_SLICE_X2Y99_BO6),
.O5(CLBLM_R_X3Y99_SLICE_X2Y99_DO5),
.O6(CLBLM_R_X3Y99_SLICE_X2Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55aa00fa50fa50)
  ) CLBLM_R_X3Y99_SLICE_X2Y99_CLUT (
.I0(CLBLL_L_X4Y97_SLICE_X4Y97_AO6),
.I1(1'b1),
.I2(CLBLM_R_X3Y97_SLICE_X2Y97_DO6),
.I3(CLBLM_R_X3Y99_SLICE_X2Y99_AO6),
.I4(CLBLL_L_X2Y99_SLICE_X0Y99_AQ),
.I5(CLBLM_R_X3Y98_SLICE_X2Y98_DO6),
.O5(CLBLM_R_X3Y99_SLICE_X2Y99_CO5),
.O6(CLBLM_R_X3Y99_SLICE_X2Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000001000000)
  ) CLBLM_R_X3Y99_SLICE_X2Y99_BLUT (
.I0(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I1(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I2(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I3(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I4(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO2),
.I5(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.O5(CLBLM_R_X3Y99_SLICE_X2Y99_BO5),
.O6(CLBLM_R_X3Y99_SLICE_X2Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0001000000000000)
  ) CLBLM_R_X3Y99_SLICE_X2Y99_ALUT (
.I0(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I1(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I2(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I3(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I4(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I5(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO0),
.O5(CLBLM_R_X3Y99_SLICE_X2Y99_AO5),
.O6(CLBLM_R_X3Y99_SLICE_X2Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y99_SLICE_X3Y99_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y99_SLICE_X3Y99_DO5),
.O6(CLBLM_R_X3Y99_SLICE_X3Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y99_SLICE_X3Y99_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y99_SLICE_X3Y99_CO5),
.O6(CLBLM_R_X3Y99_SLICE_X3Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y99_SLICE_X3Y99_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y99_SLICE_X3Y99_BO5),
.O6(CLBLM_R_X3Y99_SLICE_X3Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y99_SLICE_X3Y99_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y99_SLICE_X3Y99_AO5),
.O6(CLBLM_R_X3Y99_SLICE_X3Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y90_SLICE_X6Y90_A5_FDCE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X5Y90_SLICE_X6Y90_AO6),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLL_L_X2Y96_SLICE_X1Y96_AO6),
.Q(CLBLM_R_X5Y90_SLICE_X6Y90_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y90_SLICE_X6Y90_B5_FDCE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X5Y90_SLICE_X6Y90_AO6),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLL_L_X2Y96_SLICE_X1Y96_BO6),
.Q(CLBLM_R_X5Y90_SLICE_X6Y90_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y90_SLICE_X6Y90_A_FDCE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X5Y90_SLICE_X6Y90_AO6),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_R_X5Y90_SLICE_X6Y90_AO5),
.Q(CLBLM_R_X5Y90_SLICE_X6Y90_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y90_SLICE_X6Y90_B_FDCE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X5Y90_SLICE_X6Y90_AO6),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_R_X5Y90_SLICE_X6Y90_BO6),
.Q(CLBLM_R_X5Y90_SLICE_X6Y90_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y90_SLICE_X6Y90_C_FDCE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X5Y90_SLICE_X6Y90_AO6),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLL_L_X2Y97_SLICE_X0Y97_CO6),
.Q(CLBLM_R_X5Y90_SLICE_X6Y90_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y90_SLICE_X6Y90_D_FDCE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X5Y90_SLICE_X6Y90_AO6),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLL_L_X2Y97_SLICE_X1Y97_BO6),
.Q(CLBLM_R_X5Y90_SLICE_X6Y90_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y90_SLICE_X6Y90_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y90_SLICE_X6Y90_DO5),
.O6(CLBLM_R_X5Y90_SLICE_X6Y90_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y90_SLICE_X6Y90_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y90_SLICE_X6Y90_CO5),
.O6(CLBLM_R_X5Y90_SLICE_X6Y90_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X5Y90_SLICE_X6Y90_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X2Y97_SLICE_X1Y97_AO6),
.O5(CLBLM_R_X5Y90_SLICE_X6Y90_BO5),
.O6(CLBLM_R_X5Y90_SLICE_X6Y90_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00500000cccccccc)
  ) CLBLM_R_X5Y90_SLICE_X6Y90_ALUT (
.I0(CLBLM_R_X3Y98_SLICE_X3Y98_AO6),
.I1(CLBLL_L_X2Y97_SLICE_X0Y97_BO6),
.I2(CLBLL_L_X4Y97_SLICE_X4Y97_CO6),
.I3(CLBLL_L_X4Y98_SLICE_X4Y98_AO6),
.I4(CLBLM_R_X5Y94_SLICE_X6Y94_CO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y90_SLICE_X6Y90_AO5),
.O6(CLBLM_R_X5Y90_SLICE_X6Y90_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y90_SLICE_X7Y90_A5_FDCE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X5Y90_SLICE_X7Y90_AO6),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLL_L_X2Y96_SLICE_X1Y96_AO6),
.Q(CLBLM_R_X5Y90_SLICE_X7Y90_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y90_SLICE_X7Y90_B5_FDCE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X5Y90_SLICE_X7Y90_AO6),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLL_L_X2Y96_SLICE_X1Y96_BO6),
.Q(CLBLM_R_X5Y90_SLICE_X7Y90_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y90_SLICE_X7Y90_C5_FDCE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X5Y90_SLICE_X7Y90_AO6),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLL_L_X2Y97_SLICE_X1Y97_CO6),
.Q(CLBLM_R_X5Y90_SLICE_X7Y90_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y90_SLICE_X7Y90_A_FDCE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X5Y90_SLICE_X7Y90_AO6),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_R_X5Y90_SLICE_X7Y90_AO5),
.Q(CLBLM_R_X5Y90_SLICE_X7Y90_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y90_SLICE_X7Y90_B_FDCE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X5Y90_SLICE_X7Y90_AO6),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_R_X5Y90_SLICE_X7Y90_BO6),
.Q(CLBLM_R_X5Y90_SLICE_X7Y90_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y90_SLICE_X7Y90_C_FDCE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X5Y90_SLICE_X7Y90_AO6),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_R_X5Y90_SLICE_X7Y90_CO6),
.Q(CLBLM_R_X5Y90_SLICE_X7Y90_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y90_SLICE_X7Y90_D_FDCE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X5Y90_SLICE_X7Y90_AO6),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLL_L_X2Y97_SLICE_X1Y97_BO6),
.Q(CLBLM_R_X5Y90_SLICE_X7Y90_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y90_SLICE_X7Y90_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y90_SLICE_X7Y90_DO5),
.O6(CLBLM_R_X5Y90_SLICE_X7Y90_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X5Y90_SLICE_X7Y90_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X2Y97_SLICE_X0Y97_CO6),
.O5(CLBLM_R_X5Y90_SLICE_X7Y90_CO5),
.O6(CLBLM_R_X5Y90_SLICE_X7Y90_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X5Y90_SLICE_X7Y90_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X2Y97_SLICE_X1Y97_AO6),
.O5(CLBLM_R_X5Y90_SLICE_X7Y90_BO5),
.O6(CLBLM_R_X5Y90_SLICE_X7Y90_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00004040ff00ff00)
  ) CLBLM_R_X5Y90_SLICE_X7Y90_ALUT (
.I0(CLBLM_R_X3Y98_SLICE_X3Y98_AO6),
.I1(CLBLL_L_X4Y98_SLICE_X4Y98_AO6),
.I2(CLBLM_R_X5Y94_SLICE_X6Y94_CO6),
.I3(CLBLL_L_X2Y97_SLICE_X0Y97_BO6),
.I4(CLBLL_L_X4Y97_SLICE_X4Y97_CO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y90_SLICE_X7Y90_AO5),
.O6(CLBLM_R_X5Y90_SLICE_X7Y90_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y91_SLICE_X6Y91_A_FDCE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(1'b1),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_R_X5Y91_SLICE_X6Y91_AO6),
.Q(CLBLM_R_X5Y91_SLICE_X6Y91_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y91_SLICE_X6Y91_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y91_SLICE_X6Y91_DO5),
.O6(CLBLM_R_X5Y91_SLICE_X6Y91_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y91_SLICE_X6Y91_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y91_SLICE_X6Y91_CO5),
.O6(CLBLM_R_X5Y91_SLICE_X6Y91_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y91_SLICE_X6Y91_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y91_SLICE_X6Y91_BO5),
.O6(CLBLM_R_X5Y91_SLICE_X6Y91_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0f870f0f0)
  ) CLBLM_R_X5Y91_SLICE_X6Y91_ALUT (
.I0(CLBLM_R_X5Y94_SLICE_X6Y94_CO6),
.I1(CLBLL_L_X4Y98_SLICE_X4Y98_AO6),
.I2(CLBLM_R_X5Y91_SLICE_X6Y91_AQ),
.I3(CLBLL_L_X2Y97_SLICE_X0Y97_CO6),
.I4(CLBLL_L_X4Y97_SLICE_X4Y97_CO6),
.I5(CLBLM_R_X3Y98_SLICE_X3Y98_AO6),
.O5(CLBLM_R_X5Y91_SLICE_X6Y91_AO5),
.O6(CLBLM_R_X5Y91_SLICE_X6Y91_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y91_SLICE_X7Y91_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y91_SLICE_X7Y91_DO5),
.O6(CLBLM_R_X5Y91_SLICE_X7Y91_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y91_SLICE_X7Y91_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y91_SLICE_X7Y91_CO5),
.O6(CLBLM_R_X5Y91_SLICE_X7Y91_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y91_SLICE_X7Y91_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y91_SLICE_X7Y91_BO5),
.O6(CLBLM_R_X5Y91_SLICE_X7Y91_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y91_SLICE_X7Y91_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y91_SLICE_X7Y91_AO5),
.O6(CLBLM_R_X5Y91_SLICE_X7Y91_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y92_SLICE_X6Y92_A_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(1'b1),
.D(CLBLM_R_X5Y92_SLICE_X6Y92_AO6),
.Q(CLBLM_R_X5Y92_SLICE_X6Y92_AQ),
.R(CLBLM_R_X5Y92_SLICE_X7Y92_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y92_SLICE_X6Y92_B_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(1'b1),
.D(CLBLM_R_X5Y92_SLICE_X6Y92_BO6),
.Q(CLBLM_R_X5Y92_SLICE_X6Y92_BQ),
.R(CLBLM_R_X5Y92_SLICE_X7Y92_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y92_SLICE_X6Y92_C_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(1'b1),
.D(CLBLM_R_X5Y92_SLICE_X6Y92_CO6),
.Q(CLBLM_R_X5Y92_SLICE_X6Y92_CQ),
.R(CLBLM_R_X5Y92_SLICE_X7Y92_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y92_SLICE_X6Y92_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y92_SLICE_X6Y92_DO5),
.O6(CLBLM_R_X5Y92_SLICE_X6Y92_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000320010)
  ) CLBLM_R_X5Y92_SLICE_X6Y92_CLUT (
.I0(CLBLM_R_X3Y93_SLICE_X2Y93_CO6),
.I1(CLBLM_R_X5Y94_SLICE_X7Y94_DO6),
.I2(CLBLM_R_X3Y99_SLICE_X2Y99_CO6),
.I3(CLBLL_L_X4Y94_SLICE_X5Y94_DO6),
.I4(CLBLL_L_X2Y97_SLICE_X0Y97_BO6),
.I5(CLBLM_R_X5Y94_SLICE_X6Y94_BO6),
.O5(CLBLM_R_X5Y92_SLICE_X6Y92_CO5),
.O6(CLBLM_R_X5Y92_SLICE_X6Y92_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000440050)
  ) CLBLM_R_X5Y92_SLICE_X6Y92_BLUT (
.I0(CLBLM_R_X5Y94_SLICE_X7Y94_DO6),
.I1(CLBLL_L_X2Y96_SLICE_X1Y96_BO6),
.I2(CLBLL_L_X4Y96_SLICE_X5Y96_AO6),
.I3(CLBLL_L_X4Y94_SLICE_X5Y94_DO6),
.I4(CLBLM_R_X3Y93_SLICE_X2Y93_CO6),
.I5(CLBLM_R_X5Y94_SLICE_X6Y94_BO6),
.O5(CLBLM_R_X5Y92_SLICE_X6Y92_BO5),
.O6(CLBLM_R_X5Y92_SLICE_X6Y92_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0010001100100000)
  ) CLBLM_R_X5Y92_SLICE_X6Y92_ALUT (
.I0(CLBLM_R_X5Y94_SLICE_X7Y94_DO6),
.I1(CLBLL_L_X4Y94_SLICE_X5Y94_DO6),
.I2(CLBLL_L_X2Y96_SLICE_X1Y96_AO6),
.I3(CLBLM_R_X5Y94_SLICE_X6Y94_BO6),
.I4(CLBLM_R_X3Y93_SLICE_X2Y93_CO6),
.I5(CLBLL_L_X4Y96_SLICE_X4Y96_AO6),
.O5(CLBLM_R_X5Y92_SLICE_X6Y92_AO5),
.O6(CLBLM_R_X5Y92_SLICE_X6Y92_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y92_SLICE_X7Y92_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y92_SLICE_X7Y92_DO5),
.O6(CLBLM_R_X5Y92_SLICE_X7Y92_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y92_SLICE_X7Y92_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y92_SLICE_X7Y92_CO5),
.O6(CLBLM_R_X5Y92_SLICE_X7Y92_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y92_SLICE_X7Y92_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y92_SLICE_X7Y92_BO5),
.O6(CLBLM_R_X5Y92_SLICE_X7Y92_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haeae7070a7a76565)
  ) CLBLM_R_X5Y92_SLICE_X7Y92_ALUT (
.I0(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I1(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I2(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I5(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.O5(CLBLM_R_X5Y92_SLICE_X7Y92_AO5),
.O6(CLBLM_R_X5Y92_SLICE_X7Y92_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y93_SLICE_X6Y93_B_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLL_L_X2Y93_SLICE_X0Y93_DO6),
.D(CLBLL_L_X4Y93_SLICE_X4Y93_CO6),
.Q(CLBLM_R_X5Y93_SLICE_X6Y93_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y93_SLICE_X6Y93_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y93_SLICE_X6Y93_DO5),
.O6(CLBLM_R_X5Y93_SLICE_X6Y93_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000400)
  ) CLBLM_R_X5Y93_SLICE_X6Y93_CLUT (
.I0(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO12),
.I1(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO13),
.I2(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO15),
.I3(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO9),
.I4(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO14),
.I5(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO11),
.O5(CLBLM_R_X5Y93_SLICE_X6Y93_CO5),
.O6(CLBLM_R_X5Y93_SLICE_X6Y93_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcf000901cf000800)
  ) CLBLM_R_X5Y93_SLICE_X6Y93_BLUT (
.I0(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I1(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I2(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I3(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO9),
.I4(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I5(CLBLM_R_X5Y93_SLICE_X6Y93_CO6),
.O5(CLBLM_R_X5Y93_SLICE_X6Y93_BO5),
.O6(CLBLM_R_X5Y93_SLICE_X6Y93_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000f3003000f300)
  ) CLBLM_R_X5Y93_SLICE_X6Y93_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I2(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I3(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO9),
.I4(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I5(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.O5(CLBLM_R_X5Y93_SLICE_X6Y93_AO5),
.O6(CLBLM_R_X5Y93_SLICE_X6Y93_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_R_X5Y93_SLICE_X6Y93_MUXF7A (
.I0(CLBLM_R_X5Y93_SLICE_X6Y93_BO6),
.I1(CLBLM_R_X5Y93_SLICE_X6Y93_AO6),
.O(CLBLM_R_X5Y93_SLICE_X6Y93_F7AMUX_O),
.S(CLBLL_L_X4Y91_SLICE_X5Y91_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y93_SLICE_X7Y93_A_FDCE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(1'b1),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_R_X5Y93_SLICE_X7Y93_AO6),
.Q(CLBLM_R_X5Y93_SLICE_X7Y93_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y93_SLICE_X7Y93_B_FDCE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(1'b1),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_R_X5Y93_SLICE_X7Y93_BO6),
.Q(CLBLM_R_X5Y93_SLICE_X7Y93_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y93_SLICE_X7Y93_C_FDCE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(1'b1),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_R_X5Y93_SLICE_X7Y93_CO6),
.Q(CLBLM_R_X5Y93_SLICE_X7Y93_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y93_SLICE_X7Y93_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y93_SLICE_X7Y93_DO5),
.O6(CLBLM_R_X5Y93_SLICE_X7Y93_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff4000bfff0000)
  ) CLBLM_R_X5Y93_SLICE_X7Y93_CLUT (
.I0(CLBLL_L_X4Y97_SLICE_X4Y97_CO6),
.I1(CLBLM_R_X5Y94_SLICE_X6Y94_CO6),
.I2(CLBLL_L_X4Y98_SLICE_X4Y98_AO6),
.I3(CLBLM_R_X3Y98_SLICE_X3Y98_AO6),
.I4(CLBLM_R_X5Y93_SLICE_X7Y93_CQ),
.I5(CLBLL_L_X2Y97_SLICE_X0Y97_BO6),
.O5(CLBLM_R_X5Y93_SLICE_X7Y93_CO5),
.O6(CLBLM_R_X5Y93_SLICE_X7Y93_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccaccccccc)
  ) CLBLM_R_X5Y93_SLICE_X7Y93_BLUT (
.I0(CLBLL_L_X2Y97_SLICE_X0Y97_BO6),
.I1(CLBLM_R_X5Y93_SLICE_X7Y93_BQ),
.I2(CLBLM_R_X5Y94_SLICE_X6Y94_CO6),
.I3(CLBLL_L_X4Y98_SLICE_X4Y98_AO6),
.I4(CLBLL_L_X4Y97_SLICE_X4Y97_CO6),
.I5(CLBLM_R_X3Y98_SLICE_X3Y98_AO6),
.O5(CLBLM_R_X5Y93_SLICE_X7Y93_BO5),
.O6(CLBLM_R_X5Y93_SLICE_X7Y93_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaacaaaaaaa)
  ) CLBLM_R_X5Y93_SLICE_X7Y93_ALUT (
.I0(CLBLM_R_X5Y93_SLICE_X7Y93_AQ),
.I1(CLBLL_L_X2Y97_SLICE_X1Y97_AO6),
.I2(CLBLM_R_X5Y94_SLICE_X6Y94_CO6),
.I3(CLBLL_L_X4Y97_SLICE_X4Y97_CO6),
.I4(CLBLL_L_X4Y98_SLICE_X4Y98_AO6),
.I5(CLBLM_R_X3Y98_SLICE_X3Y98_AO6),
.O5(CLBLM_R_X5Y93_SLICE_X7Y93_AO5),
.O6(CLBLM_R_X5Y93_SLICE_X7Y93_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y94_SLICE_X6Y94_A_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLL_L_X2Y92_SLICE_X1Y92_AO6),
.D(CLBLL_L_X4Y93_SLICE_X4Y93_CO5),
.Q(CLBLM_R_X5Y94_SLICE_X6Y94_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y94_SLICE_X6Y94_B_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLL_L_X2Y92_SLICE_X1Y92_AO6),
.D(CLBLL_L_X4Y94_SLICE_X4Y94_CO6),
.Q(CLBLM_R_X5Y94_SLICE_X6Y94_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y94_SLICE_X6Y94_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y94_SLICE_X6Y94_DO5),
.O6(CLBLM_R_X5Y94_SLICE_X6Y94_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000004000400)
  ) CLBLM_R_X5Y94_SLICE_X6Y94_CLUT (
.I0(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I1(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I2(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I3(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.O5(CLBLM_R_X5Y94_SLICE_X6Y94_CO5),
.O6(CLBLM_R_X5Y94_SLICE_X6Y94_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haeff00ffae0c0000)
  ) CLBLM_R_X5Y94_SLICE_X6Y94_BLUT (
.I0(CLBLM_R_X5Y94_SLICE_X7Y94_AO5),
.I1(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I2(CLBLM_R_X5Y94_SLICE_X7Y94_AO6),
.I3(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I4(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO9),
.I5(CLBLM_R_X5Y94_SLICE_X6Y94_AO6),
.O5(CLBLM_R_X5Y94_SLICE_X6Y94_BO5),
.O6(CLBLM_R_X5Y94_SLICE_X6Y94_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0d0d000009180)
  ) CLBLM_R_X5Y94_SLICE_X6Y94_ALUT (
.I0(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I1(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I2(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO9),
.I3(CLBLM_R_X5Y95_SLICE_X6Y95_DO6),
.I4(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I5(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.O5(CLBLM_R_X5Y94_SLICE_X6Y94_AO5),
.O6(CLBLM_R_X5Y94_SLICE_X6Y94_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc4ffc0ffc444c000)
  ) CLBLM_R_X5Y94_SLICE_X7Y94_DLUT (
.I0(CLBLM_R_X5Y94_SLICE_X7Y94_AO6),
.I1(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO8),
.I2(CLBLM_R_X5Y94_SLICE_X7Y94_AO5),
.I3(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I4(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I5(CLBLM_R_X5Y94_SLICE_X7Y94_BO6),
.O5(CLBLM_R_X5Y94_SLICE_X7Y94_DO5),
.O6(CLBLM_R_X5Y94_SLICE_X7Y94_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000020000000000)
  ) CLBLM_R_X5Y94_SLICE_X7Y94_CLUT (
.I0(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO12),
.I1(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO14),
.I2(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO13),
.I3(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO8),
.I4(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO15),
.I5(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO11),
.O5(CLBLM_R_X5Y94_SLICE_X7Y94_CO5),
.O6(CLBLM_R_X5Y94_SLICE_X7Y94_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8a88000b8a880008)
  ) CLBLM_R_X5Y94_SLICE_X7Y94_BLUT (
.I0(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO8),
.I1(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I2(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I3(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I4(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I5(CLBLM_R_X5Y94_SLICE_X7Y94_CO6),
.O5(CLBLM_R_X5Y94_SLICE_X7Y94_BO5),
.O6(CLBLM_R_X5Y94_SLICE_X7Y94_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffcccc0030f3f3)
  ) CLBLM_R_X5Y94_SLICE_X7Y94_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I2(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I3(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I4(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y94_SLICE_X7Y94_AO5),
.O6(CLBLM_R_X5Y94_SLICE_X7Y94_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y95_SLICE_X6Y95_A_FDCE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(1'b1),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_R_X5Y95_SLICE_X6Y95_AO6),
.Q(CLBLM_R_X5Y95_SLICE_X6Y95_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0100000000000000)
  ) CLBLM_R_X5Y95_SLICE_X6Y95_DLUT (
.I0(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO13),
.I1(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO14),
.I2(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO15),
.I3(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO9),
.I4(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO12),
.I5(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO11),
.O5(CLBLM_R_X5Y95_SLICE_X6Y95_DO5),
.O6(CLBLM_R_X5Y95_SLICE_X6Y95_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffefffffffff)
  ) CLBLM_R_X5Y95_SLICE_X6Y95_CLUT (
.I0(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I1(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO13),
.I2(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO15),
.I3(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO14),
.I4(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO12),
.I5(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO11),
.O5(CLBLM_R_X5Y95_SLICE_X6Y95_CO5),
.O6(CLBLM_R_X5Y95_SLICE_X6Y95_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafafafa00000001)
  ) CLBLM_R_X5Y95_SLICE_X6Y95_BLUT (
.I0(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I1(CLBLM_R_X5Y95_SLICE_X6Y95_CO6),
.I2(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I3(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I4(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y95_SLICE_X6Y95_BO5),
.O6(CLBLM_R_X5Y95_SLICE_X6Y95_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f1f0f0f0e0f0f0)
  ) CLBLM_R_X5Y95_SLICE_X6Y95_ALUT (
.I0(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I1(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I2(CLBLM_R_X5Y95_SLICE_X6Y95_AQ),
.I3(CLBLM_R_X5Y95_SLICE_X6Y95_BO6),
.I4(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I5(CLBLL_L_X2Y95_SLICE_X0Y95_D_CY),
.O5(CLBLM_R_X5Y95_SLICE_X6Y95_AO5),
.O6(CLBLM_R_X5Y95_SLICE_X6Y95_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y95_SLICE_X7Y95_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y95_SLICE_X7Y95_DO5),
.O6(CLBLM_R_X5Y95_SLICE_X7Y95_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y95_SLICE_X7Y95_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y95_SLICE_X7Y95_CO5),
.O6(CLBLM_R_X5Y95_SLICE_X7Y95_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y95_SLICE_X7Y95_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y95_SLICE_X7Y95_BO5),
.O6(CLBLM_R_X5Y95_SLICE_X7Y95_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y95_SLICE_X7Y95_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y95_SLICE_X7Y95_AO5),
.O6(CLBLM_R_X5Y95_SLICE_X7Y95_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y96_SLICE_X6Y96_A_FDCE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X7Y99_SLICE_X9Y99_DO6),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_R_X5Y96_SLICE_X6Y96_AO6),
.Q(CLBLM_R_X5Y96_SLICE_X6Y96_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f80ff00ff00ff00)
  ) CLBLM_R_X5Y96_SLICE_X6Y96_DLUT (
.I0(CLBLM_R_X5Y96_SLICE_X7Y96_AQ),
.I1(CLBLM_R_X5Y96_SLICE_X7Y96_BQ),
.I2(CLBLM_R_X7Y99_SLICE_X8Y99_AQ),
.I3(CLBLM_R_X5Y96_SLICE_X6Y96_AQ),
.I4(CLBLM_R_X5Y99_SLICE_X7Y99_AQ),
.I5(CLBLM_R_X5Y99_SLICE_X6Y99_AQ),
.O5(CLBLM_R_X5Y96_SLICE_X6Y96_DO5),
.O6(CLBLM_R_X5Y96_SLICE_X6Y96_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb0f090d08000c040)
  ) CLBLM_R_X5Y96_SLICE_X6Y96_CLUT (
.I0(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I1(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I2(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO5),
.I3(CLBLM_R_X5Y95_SLICE_X6Y95_AQ),
.I4(CLBLL_L_X4Y97_SLICE_X4Y97_BQ),
.I5(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.O5(CLBLM_R_X5Y96_SLICE_X6Y96_CO5),
.O6(CLBLM_R_X5Y96_SLICE_X6Y96_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heac846ce00000000)
  ) CLBLM_R_X5Y96_SLICE_X6Y96_BLUT (
.I0(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I1(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I2(CLBLL_L_X4Y97_SLICE_X4Y97_BQ),
.I3(CLBLM_R_X5Y95_SLICE_X6Y95_AQ),
.I4(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I5(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO4),
.O5(CLBLM_R_X5Y96_SLICE_X6Y96_BO5),
.O6(CLBLM_R_X5Y96_SLICE_X6Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h2e2ee2222222e222)
  ) CLBLM_R_X5Y96_SLICE_X6Y96_ALUT (
.I0(CLBLM_R_X5Y96_SLICE_X6Y96_DO6),
.I1(CLBLM_R_X7Y98_SLICE_X8Y98_F7AMUX_O),
.I2(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I3(CLBLL_L_X4Y97_SLICE_X5Y97_BO6),
.I4(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I5(CLBLM_R_X5Y96_SLICE_X6Y96_CO6),
.O5(CLBLM_R_X5Y96_SLICE_X6Y96_AO5),
.O6(CLBLM_R_X5Y96_SLICE_X6Y96_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y96_SLICE_X7Y96_A_FDCE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X7Y99_SLICE_X9Y99_DO6),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_R_X5Y96_SLICE_X7Y96_AO6),
.Q(CLBLM_R_X5Y96_SLICE_X7Y96_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y96_SLICE_X7Y96_B_FDCE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X7Y99_SLICE_X9Y99_DO6),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_R_X5Y96_SLICE_X7Y96_BO6),
.Q(CLBLM_R_X5Y96_SLICE_X7Y96_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc844c8cc88080008)
  ) CLBLM_R_X5Y96_SLICE_X7Y96_DLUT (
.I0(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I1(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO3),
.I2(CLBLL_L_X4Y97_SLICE_X4Y97_BQ),
.I3(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I4(CLBLM_R_X5Y95_SLICE_X6Y95_AQ),
.I5(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.O5(CLBLM_R_X5Y96_SLICE_X7Y96_DO5),
.O6(CLBLM_R_X5Y96_SLICE_X7Y96_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f80ff007f7f8080)
  ) CLBLM_R_X5Y96_SLICE_X7Y96_CLUT (
.I0(CLBLM_R_X7Y99_SLICE_X8Y99_AQ),
.I1(CLBLM_R_X5Y99_SLICE_X6Y99_AQ),
.I2(CLBLM_R_X5Y99_SLICE_X7Y99_AQ),
.I3(CLBLM_R_X5Y96_SLICE_X7Y96_BQ),
.I4(CLBLM_R_X5Y96_SLICE_X7Y96_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y96_SLICE_X7Y96_CO5),
.O6(CLBLM_R_X5Y96_SLICE_X7Y96_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f55d5d50a008080)
  ) CLBLM_R_X5Y96_SLICE_X7Y96_BLUT (
.I0(CLBLM_R_X7Y98_SLICE_X8Y98_F7AMUX_O),
.I1(CLBLM_R_X5Y96_SLICE_X6Y96_BO6),
.I2(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I3(CLBLM_R_X5Y98_SLICE_X7Y98_DO6),
.I4(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I5(CLBLM_R_X5Y96_SLICE_X7Y96_CO6),
.O5(CLBLM_R_X5Y96_SLICE_X7Y96_BO5),
.O6(CLBLM_R_X5Y96_SLICE_X7Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h2c202c20ffff0000)
  ) CLBLM_R_X5Y96_SLICE_X7Y96_ALUT (
.I0(CLBLM_R_X5Y96_SLICE_X7Y96_DO6),
.I1(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I2(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I3(CLBLM_R_X5Y97_SLICE_X7Y97_BO6),
.I4(CLBLM_R_X5Y96_SLICE_X7Y96_CO5),
.I5(CLBLM_R_X7Y98_SLICE_X8Y98_F7AMUX_O),
.O5(CLBLM_R_X5Y96_SLICE_X7Y96_AO5),
.O6(CLBLM_R_X5Y96_SLICE_X7Y96_AO6)
  );


  (* KEEP, DONT_TOUCH *)
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000)
  ) CLBLM_R_X5Y97_SLICE_X6Y97_RAM32M (
.ADDRA({1'b0, CLBLM_R_X7Y97_SLICE_X9Y97_B5Q, CLBLM_R_X7Y97_SLICE_X9Y97_BQ, CLBLM_R_X7Y97_SLICE_X9Y97_A5Q, CLBLM_R_X7Y97_SLICE_X9Y97_AQ}),
.ADDRB({1'b0, CLBLM_R_X7Y97_SLICE_X9Y97_B5Q, CLBLM_R_X7Y97_SLICE_X9Y97_BQ, CLBLM_R_X7Y97_SLICE_X9Y97_A5Q, CLBLM_R_X7Y97_SLICE_X9Y97_AQ}),
.ADDRC({1'b0, CLBLM_R_X7Y97_SLICE_X9Y97_B5Q, CLBLM_R_X7Y97_SLICE_X9Y97_BQ, CLBLM_R_X7Y97_SLICE_X9Y97_A5Q, CLBLM_R_X7Y97_SLICE_X9Y97_AQ}),
.ADDRD({1'b0, CLBLM_R_X7Y97_SLICE_X9Y97_B5Q, CLBLM_R_X7Y97_SLICE_X9Y97_BQ, CLBLM_R_X7Y97_SLICE_X9Y97_A5Q, CLBLM_R_X7Y97_SLICE_X9Y97_AQ}),
.DIA({CLBLM_R_X5Y96_SLICE_X7Y96_BQ, CLBLM_R_X5Y98_SLICE_X6Y98_CO6}),
.DIB({CLBLM_R_X5Y96_SLICE_X6Y96_AQ, CLBLM_R_X5Y98_SLICE_X6Y98_CO6}),
.DIC({CLBLM_R_X7Y96_SLICE_X8Y96_AQ, CLBLM_R_X5Y98_SLICE_X6Y98_CO6}),
.DID({CLBLM_R_X5Y96_SLICE_X7Y96_AQ, CLBLM_R_X5Y98_SLICE_X6Y98_CO6}),
.DOA({CLBLM_R_X5Y97_SLICE_X6Y97_AO6, CLBLM_R_X5Y97_SLICE_X6Y97_AO5}),
.DOB({CLBLM_R_X5Y97_SLICE_X6Y97_BO6, CLBLM_R_X5Y97_SLICE_X6Y97_BO5}),
.DOC({CLBLM_R_X5Y97_SLICE_X6Y97_CO6, CLBLM_R_X5Y97_SLICE_X6Y97_CO5}),
.DOD({CLBLM_R_X5Y97_SLICE_X6Y97_DO6, CLBLM_R_X5Y97_SLICE_X6Y97_DO5}),
.WCLK(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.WE(CLBLL_L_X4Y97_SLICE_X5Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X5Y97_SLICE_X7Y97_DLUT (
.I0(CLBLM_R_X5Y97_SLICE_X6Y97_DO6),
.I1(CLBLM_R_X5Y97_SLICE_X6Y97_AO6),
.I2(CLBLM_R_X5Y97_SLICE_X6Y97_BO6),
.I3(CLBLM_R_X5Y98_SLICE_X6Y98_CO6),
.I4(CLBLM_R_X5Y98_SLICE_X6Y98_BO6),
.I5(CLBLM_R_X5Y98_SLICE_X6Y98_DO6),
.O5(CLBLM_R_X5Y97_SLICE_X7Y97_DO5),
.O6(CLBLM_R_X5Y97_SLICE_X7Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f0f60600000606)
  ) CLBLM_R_X5Y97_SLICE_X7Y97_CLUT (
.I0(CLBLM_R_X5Y97_SLICE_X7Y97_AO6),
.I1(CLBLM_R_X5Y97_SLICE_X6Y97_AO6),
.I2(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I3(CLBLL_L_X4Y97_SLICE_X4Y97_BQ),
.I4(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I5(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO4),
.O5(CLBLM_R_X5Y97_SLICE_X7Y97_CO5),
.O6(CLBLM_R_X5Y97_SLICE_X7Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5775555502200000)
  ) CLBLM_R_X5Y97_SLICE_X7Y97_BLUT (
.I0(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I1(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I2(CLBLM_R_X5Y95_SLICE_X6Y95_AQ),
.I3(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I4(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO3),
.I5(CLBLM_R_X5Y98_SLICE_X7Y98_CO6),
.O5(CLBLM_R_X5Y97_SLICE_X7Y97_BO5),
.O6(CLBLM_R_X5Y97_SLICE_X7Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8800000080000000)
  ) CLBLM_R_X5Y97_SLICE_X7Y97_ALUT (
.I0(CLBLM_R_X5Y98_SLICE_X6Y98_BO6),
.I1(CLBLM_R_X5Y98_SLICE_X6Y98_CO6),
.I2(CLBLM_R_X5Y97_SLICE_X6Y97_AO6),
.I3(CLBLM_R_X5Y98_SLICE_X6Y98_DO6),
.I4(CLBLM_R_X5Y97_SLICE_X6Y97_DO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y97_SLICE_X7Y97_AO5),
.O6(CLBLM_R_X5Y97_SLICE_X7Y97_AO6)
  );


  (* KEEP, DONT_TOUCH *)
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000)
  ) CLBLM_R_X5Y98_SLICE_X6Y98_RAM32M (
.ADDRA({1'b0, CLBLM_R_X7Y97_SLICE_X9Y97_B5Q, CLBLM_R_X7Y97_SLICE_X9Y97_BQ, CLBLM_R_X7Y97_SLICE_X9Y97_A5Q, CLBLM_R_X7Y97_SLICE_X9Y97_AQ}),
.ADDRB({1'b0, CLBLM_R_X7Y97_SLICE_X9Y97_B5Q, CLBLM_R_X7Y97_SLICE_X9Y97_BQ, CLBLM_R_X7Y97_SLICE_X9Y97_A5Q, CLBLM_R_X7Y97_SLICE_X9Y97_AQ}),
.ADDRC({1'b0, CLBLM_R_X7Y97_SLICE_X9Y97_B5Q, CLBLM_R_X7Y97_SLICE_X9Y97_BQ, CLBLM_R_X7Y97_SLICE_X9Y97_A5Q, CLBLM_R_X7Y97_SLICE_X9Y97_AQ}),
.ADDRD({1'b0, CLBLM_R_X7Y97_SLICE_X9Y97_B5Q, CLBLM_R_X7Y97_SLICE_X9Y97_BQ, CLBLM_R_X7Y97_SLICE_X9Y97_A5Q, CLBLM_R_X7Y97_SLICE_X9Y97_AQ}),
.DIA({CLBLM_R_X7Y97_SLICE_X8Y97_AQ, CLBLL_L_X4Y97_SLICE_X5Y97_DO6}),
.DIB({CLBLM_R_X5Y99_SLICE_X7Y99_AQ, CLBLL_L_X4Y97_SLICE_X5Y97_DO6}),
.DIC({CLBLM_R_X5Y99_SLICE_X6Y99_AQ, CLBLL_L_X4Y97_SLICE_X5Y97_DO6}),
.DID({CLBLM_R_X7Y99_SLICE_X8Y99_AQ, CLBLL_L_X4Y97_SLICE_X5Y97_DO6}),
.DOA({CLBLM_R_X5Y98_SLICE_X6Y98_AO6, CLBLM_R_X5Y98_SLICE_X6Y98_AO5}),
.DOB({CLBLM_R_X5Y98_SLICE_X6Y98_BO6, CLBLM_R_X5Y98_SLICE_X6Y98_BO5}),
.DOC({CLBLM_R_X5Y98_SLICE_X6Y98_CO6, CLBLM_R_X5Y98_SLICE_X6Y98_CO5}),
.DOD({CLBLM_R_X5Y98_SLICE_X6Y98_DO6, CLBLM_R_X5Y98_SLICE_X6Y98_DO5}),
.WCLK(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.WE(CLBLL_L_X4Y97_SLICE_X5Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0a0aca0aca0a0a)
  ) CLBLM_R_X5Y98_SLICE_X7Y98_DLUT (
.I0(CLBLM_R_X5Y97_SLICE_X7Y97_CO6),
.I1(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO4),
.I2(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I3(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I4(CLBLM_R_X5Y95_SLICE_X6Y95_AQ),
.I5(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.O5(CLBLM_R_X5Y98_SLICE_X7Y98_DO5),
.O6(CLBLM_R_X5Y98_SLICE_X7Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h50500000a0a033cc)
  ) CLBLM_R_X5Y98_SLICE_X7Y98_CLUT (
.I0(CLBLL_L_X4Y97_SLICE_X4Y97_BQ),
.I1(CLBLM_R_X5Y97_SLICE_X6Y97_DO6),
.I2(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO3),
.I3(CLBLM_R_X5Y98_SLICE_X7Y98_AO5),
.I4(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I5(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.O5(CLBLM_R_X5Y98_SLICE_X7Y98_CO5),
.O6(CLBLM_R_X5Y98_SLICE_X7Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2301321089019810)
  ) CLBLM_R_X5Y98_SLICE_X7Y98_BLUT (
.I0(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I1(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I2(CLBLM_R_X5Y98_SLICE_X6Y98_CO6),
.I3(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO2),
.I4(CLBLM_R_X5Y98_SLICE_X7Y98_AO6),
.I5(CLBLL_L_X4Y97_SLICE_X4Y97_BQ),
.O5(CLBLM_R_X5Y98_SLICE_X7Y98_BO5),
.O6(CLBLM_R_X5Y98_SLICE_X7Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00c000c000)
  ) CLBLM_R_X5Y98_SLICE_X7Y98_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y98_SLICE_X6Y98_BO6),
.I2(CLBLM_R_X5Y98_SLICE_X6Y98_CO6),
.I3(CLBLM_R_X5Y98_SLICE_X6Y98_DO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y98_SLICE_X7Y98_AO5),
.O6(CLBLM_R_X5Y98_SLICE_X7Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y99_SLICE_X6Y99_A_FDCE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X7Y99_SLICE_X9Y99_DO6),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_R_X5Y99_SLICE_X6Y99_AO6),
.Q(CLBLM_R_X5Y99_SLICE_X6Y99_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y99_SLICE_X6Y99_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y99_SLICE_X6Y99_DO5),
.O6(CLBLM_R_X5Y99_SLICE_X6Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c48c00cc048c00)
  ) CLBLM_R_X5Y99_SLICE_X6Y99_CLUT (
.I0(CLBLL_L_X4Y97_SLICE_X4Y97_BQ),
.I1(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO2),
.I2(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I3(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I4(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I5(CLBLM_R_X5Y95_SLICE_X6Y95_AQ),
.O5(CLBLM_R_X5Y99_SLICE_X6Y99_CO5),
.O6(CLBLM_R_X5Y99_SLICE_X6Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hab00c400cd00c400)
  ) CLBLM_R_X5Y99_SLICE_X6Y99_BLUT (
.I0(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I1(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I2(CLBLL_L_X4Y97_SLICE_X4Y97_BQ),
.I3(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO1),
.I4(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I5(CLBLM_R_X5Y95_SLICE_X6Y95_AQ),
.O5(CLBLM_R_X5Y99_SLICE_X6Y99_BO5),
.O6(CLBLM_R_X5Y99_SLICE_X6Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h50aacccc5000cccc)
  ) CLBLM_R_X5Y99_SLICE_X6Y99_ALUT (
.I0(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I1(CLBLM_R_X5Y99_SLICE_X7Y99_BO6),
.I2(CLBLL_L_X4Y98_SLICE_X5Y98_AO6),
.I3(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I4(CLBLM_R_X7Y98_SLICE_X8Y98_F7AMUX_O),
.I5(CLBLM_R_X5Y99_SLICE_X6Y99_CO6),
.O5(CLBLM_R_X5Y99_SLICE_X6Y99_AO5),
.O6(CLBLM_R_X5Y99_SLICE_X6Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y99_SLICE_X7Y99_A_FDCE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X7Y99_SLICE_X9Y99_DO6),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_R_X5Y99_SLICE_X7Y99_AO6),
.Q(CLBLM_R_X5Y99_SLICE_X7Y99_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4444888800000ff0)
  ) CLBLM_R_X5Y99_SLICE_X7Y99_DLUT (
.I0(CLBLL_L_X4Y97_SLICE_X4Y97_BQ),
.I1(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO1),
.I2(CLBLM_R_X5Y98_SLICE_X6Y98_DO6),
.I3(CLBLM_R_X5Y98_SLICE_X6Y98_BO6),
.I4(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I5(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.O5(CLBLM_R_X5Y99_SLICE_X7Y99_DO5),
.O6(CLBLM_R_X5Y99_SLICE_X7Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h04400440ffff0000)
  ) CLBLM_R_X5Y99_SLICE_X7Y99_CLUT (
.I0(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I1(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO1),
.I2(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I3(CLBLM_R_X5Y95_SLICE_X6Y95_AQ),
.I4(CLBLM_R_X5Y99_SLICE_X7Y99_DO6),
.I5(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.O5(CLBLM_R_X5Y99_SLICE_X7Y99_CO5),
.O6(CLBLM_R_X5Y99_SLICE_X7Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ffff0000ff00ff0)
  ) CLBLM_R_X5Y99_SLICE_X7Y99_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X5Y99_SLICE_X7Y99_AQ),
.I3(CLBLM_R_X7Y99_SLICE_X8Y99_AQ),
.I4(CLBLM_R_X5Y99_SLICE_X6Y99_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y99_SLICE_X7Y99_BO5),
.O6(CLBLM_R_X5Y99_SLICE_X7Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f8f50800f8f0080)
  ) CLBLM_R_X5Y99_SLICE_X7Y99_ALUT (
.I0(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I1(CLBLM_R_X5Y99_SLICE_X6Y99_BO6),
.I2(CLBLM_R_X7Y98_SLICE_X8Y98_F7AMUX_O),
.I3(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I4(CLBLM_R_X5Y99_SLICE_X7Y99_BO5),
.I5(CLBLM_R_X5Y99_SLICE_X7Y99_CO6),
.O5(CLBLM_R_X5Y99_SLICE_X7Y99_AO5),
.O6(CLBLM_R_X5Y99_SLICE_X7Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y87_SLICE_X8Y87_A_FDCE (
.C(CLBLM_R_X7Y88_SLICE_X8Y88_AQ),
.CE(1'b1),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_R_X7Y87_SLICE_X8Y87_AO6),
.Q(CLBLM_R_X7Y87_SLICE_X8Y87_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y87_SLICE_X8Y87_B_FDCE (
.C(CLBLM_R_X7Y88_SLICE_X8Y88_AQ),
.CE(1'b1),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_R_X7Y87_SLICE_X8Y87_BO6),
.Q(CLBLM_R_X7Y87_SLICE_X8Y87_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y87_SLICE_X8Y87_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y87_SLICE_X8Y87_DO5),
.O6(CLBLM_R_X7Y87_SLICE_X8Y87_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y87_SLICE_X8Y87_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y87_SLICE_X8Y87_CO5),
.O6(CLBLM_R_X7Y87_SLICE_X8Y87_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h03330ccc0ccc0ccc)
  ) CLBLM_R_X7Y87_SLICE_X8Y87_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y87_SLICE_X8Y87_BQ),
.I2(CLBLM_R_X7Y87_SLICE_X8Y87_AQ),
.I3(CLBLM_R_X7Y91_SLICE_X8Y91_AQ),
.I4(CLBLM_R_X7Y91_SLICE_X9Y91_AQ),
.I5(CLBLM_R_X7Y90_SLICE_X8Y90_CO6),
.O5(CLBLM_R_X7Y87_SLICE_X8Y87_BO5),
.O6(CLBLM_R_X7Y87_SLICE_X8Y87_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0cf010f000f010f0)
  ) CLBLM_R_X7Y87_SLICE_X8Y87_ALUT (
.I0(CLBLM_R_X7Y90_SLICE_X9Y90_CQ),
.I1(CLBLM_R_X7Y87_SLICE_X8Y87_BQ),
.I2(CLBLM_R_X7Y87_SLICE_X8Y87_AQ),
.I3(CLBLM_R_X7Y91_SLICE_X8Y91_AQ),
.I4(CLBLM_R_X7Y91_SLICE_X9Y91_AQ),
.I5(CLBLM_R_X7Y90_SLICE_X8Y90_CO6),
.O5(CLBLM_R_X7Y87_SLICE_X8Y87_AO5),
.O6(CLBLM_R_X7Y87_SLICE_X8Y87_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y87_SLICE_X9Y87_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y87_SLICE_X9Y87_DO5),
.O6(CLBLM_R_X7Y87_SLICE_X9Y87_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y87_SLICE_X9Y87_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y87_SLICE_X9Y87_CO5),
.O6(CLBLM_R_X7Y87_SLICE_X9Y87_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y87_SLICE_X9Y87_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y87_SLICE_X9Y87_BO5),
.O6(CLBLM_R_X7Y87_SLICE_X9Y87_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y87_SLICE_X9Y87_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y87_SLICE_X9Y87_AO5),
.O6(CLBLM_R_X7Y87_SLICE_X9Y87_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y88_SLICE_X8Y88_A_FDCE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(1'b1),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_R_X7Y88_SLICE_X8Y88_AO6),
.Q(CLBLM_R_X7Y88_SLICE_X8Y88_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y88_SLICE_X8Y88_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y88_SLICE_X8Y88_DO5),
.O6(CLBLM_R_X7Y88_SLICE_X8Y88_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y88_SLICE_X8Y88_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y88_SLICE_X8Y88_CO5),
.O6(CLBLM_R_X7Y88_SLICE_X8Y88_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000202)
  ) CLBLM_R_X7Y88_SLICE_X8Y88_BLUT (
.I0(CLBLM_R_X7Y90_SLICE_X8Y90_DO6),
.I1(CLBLM_R_X7Y87_SLICE_X8Y87_BQ),
.I2(CLBLM_R_X7Y87_SLICE_X8Y87_AQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y91_SLICE_X9Y91_AQ),
.I5(CLBLM_R_X7Y91_SLICE_X8Y91_AQ),
.O5(CLBLM_R_X7Y88_SLICE_X8Y88_BO5),
.O6(CLBLM_R_X7Y88_SLICE_X8Y88_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0f0f0f0f)
  ) CLBLM_R_X7Y88_SLICE_X8Y88_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X7Y88_SLICE_X8Y88_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y88_SLICE_X8Y88_AO5),
.O6(CLBLM_R_X7Y88_SLICE_X8Y88_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y88_SLICE_X9Y88_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y88_SLICE_X9Y88_DO5),
.O6(CLBLM_R_X7Y88_SLICE_X9Y88_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y88_SLICE_X9Y88_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y88_SLICE_X9Y88_CO5),
.O6(CLBLM_R_X7Y88_SLICE_X9Y88_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y88_SLICE_X9Y88_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y88_SLICE_X9Y88_BO5),
.O6(CLBLM_R_X7Y88_SLICE_X9Y88_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y88_SLICE_X9Y88_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y88_SLICE_X9Y88_AO5),
.O6(CLBLM_R_X7Y88_SLICE_X9Y88_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y89_SLICE_X8Y89_B5_FDCE (
.C(CLBLM_R_X7Y88_SLICE_X8Y88_AQ),
.CE(CLBLM_R_X7Y88_SLICE_X8Y88_BO6),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_R_X7Y89_SLICE_X8Y89_BO5),
.Q(CLBLM_R_X7Y89_SLICE_X8Y89_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y89_SLICE_X8Y89_A_FDCE (
.C(CLBLM_R_X7Y88_SLICE_X8Y88_AQ),
.CE(CLBLM_R_X7Y88_SLICE_X8Y88_BO6),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_R_X7Y89_SLICE_X8Y89_AO6),
.Q(CLBLM_R_X7Y89_SLICE_X8Y89_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y89_SLICE_X8Y89_B_FDCE (
.C(CLBLM_R_X7Y88_SLICE_X8Y88_AQ),
.CE(CLBLM_R_X7Y88_SLICE_X8Y88_BO6),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_R_X7Y89_SLICE_X8Y89_BO6),
.Q(CLBLM_R_X7Y89_SLICE_X8Y89_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y89_SLICE_X8Y89_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y89_SLICE_X8Y89_DO5),
.O6(CLBLM_R_X7Y89_SLICE_X8Y89_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888000000000000)
  ) CLBLM_R_X7Y89_SLICE_X8Y89_CLUT (
.I0(CLBLM_R_X7Y89_SLICE_X8Y89_BQ),
.I1(CLBLM_R_X7Y89_SLICE_X8Y89_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X7Y89_SLICE_X8Y89_B5Q),
.I5(CLBLM_R_X7Y89_SLICE_X9Y89_BQ),
.O5(CLBLM_R_X7Y89_SLICE_X8Y89_CO5),
.O6(CLBLM_R_X7Y89_SLICE_X8Y89_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3ccc3ccc6aaa6aaa)
  ) CLBLM_R_X7Y89_SLICE_X8Y89_BLUT (
.I0(CLBLM_R_X7Y89_SLICE_X8Y89_B5Q),
.I1(CLBLM_R_X7Y89_SLICE_X8Y89_BQ),
.I2(CLBLM_R_X7Y89_SLICE_X8Y89_AQ),
.I3(CLBLM_R_X7Y89_SLICE_X9Y89_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y89_SLICE_X8Y89_BO5),
.O6(CLBLM_R_X7Y89_SLICE_X8Y89_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h78f0f0f0f0f0f0f0)
  ) CLBLM_R_X7Y89_SLICE_X8Y89_ALUT (
.I0(CLBLM_R_X7Y89_SLICE_X9Y89_BQ),
.I1(CLBLM_R_X7Y89_SLICE_X9Y89_AQ),
.I2(CLBLM_R_X7Y89_SLICE_X8Y89_AQ),
.I3(CLBLM_L_X8Y89_SLICE_X10Y89_A5Q),
.I4(CLBLM_L_X8Y89_SLICE_X10Y89_AQ),
.I5(CLBLM_L_X8Y89_SLICE_X10Y89_BO6),
.O5(CLBLM_R_X7Y89_SLICE_X8Y89_AO5),
.O6(CLBLM_R_X7Y89_SLICE_X8Y89_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y89_SLICE_X9Y89_A_FDCE (
.C(CLBLM_R_X7Y88_SLICE_X8Y88_AQ),
.CE(CLBLM_R_X7Y88_SLICE_X8Y88_BO6),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_R_X7Y89_SLICE_X9Y89_AO6),
.Q(CLBLM_R_X7Y89_SLICE_X9Y89_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y89_SLICE_X9Y89_B_FDCE (
.C(CLBLM_R_X7Y88_SLICE_X8Y88_AQ),
.CE(CLBLM_R_X7Y88_SLICE_X8Y88_BO6),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_R_X7Y89_SLICE_X9Y89_BO6),
.Q(CLBLM_R_X7Y89_SLICE_X9Y89_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f1f3f3f3f3f3f)
  ) CLBLM_R_X7Y89_SLICE_X9Y89_DLUT (
.I0(CLBLM_L_X8Y89_SLICE_X10Y89_BQ),
.I1(CLBLM_R_X7Y89_SLICE_X9Y89_AQ),
.I2(CLBLM_R_X7Y89_SLICE_X8Y89_B5Q),
.I3(CLBLM_L_X8Y89_SLICE_X10Y89_CQ),
.I4(CLBLM_L_X8Y89_SLICE_X10Y89_AQ),
.I5(CLBLM_L_X8Y89_SLICE_X10Y89_A5Q),
.O5(CLBLM_R_X7Y89_SLICE_X9Y89_DO5),
.O6(CLBLM_R_X7Y89_SLICE_X9Y89_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X7Y89_SLICE_X9Y89_CLUT (
.I0(CLBLM_L_X8Y89_SLICE_X10Y89_BQ),
.I1(CLBLM_L_X8Y89_SLICE_X10Y89_A5Q),
.I2(CLBLM_L_X8Y89_SLICE_X10Y89_CQ),
.I3(CLBLM_R_X7Y89_SLICE_X9Y89_BQ),
.I4(CLBLM_L_X8Y89_SLICE_X10Y89_AQ),
.I5(CLBLM_R_X7Y89_SLICE_X9Y89_AQ),
.O5(CLBLM_R_X7Y89_SLICE_X9Y89_CO5),
.O6(CLBLM_R_X7Y89_SLICE_X9Y89_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffffff80000000)
  ) CLBLM_R_X7Y89_SLICE_X9Y89_BLUT (
.I0(CLBLM_L_X8Y89_SLICE_X10Y89_CQ),
.I1(CLBLM_L_X8Y89_SLICE_X10Y89_A5Q),
.I2(CLBLM_L_X8Y89_SLICE_X10Y89_AQ),
.I3(CLBLM_R_X7Y89_SLICE_X9Y89_AQ),
.I4(CLBLM_L_X8Y89_SLICE_X10Y89_BQ),
.I5(CLBLM_R_X7Y89_SLICE_X9Y89_BQ),
.O5(CLBLM_R_X7Y89_SLICE_X9Y89_BO5),
.O6(CLBLM_R_X7Y89_SLICE_X9Y89_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f80ff00003f007f)
  ) CLBLM_R_X7Y89_SLICE_X9Y89_ALUT (
.I0(CLBLM_L_X8Y89_SLICE_X10Y89_CQ),
.I1(CLBLM_L_X8Y89_SLICE_X10Y89_A5Q),
.I2(CLBLM_L_X8Y89_SLICE_X10Y89_AQ),
.I3(CLBLM_R_X7Y89_SLICE_X9Y89_AQ),
.I4(CLBLM_L_X8Y89_SLICE_X10Y89_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y89_SLICE_X9Y89_AO5),
.O6(CLBLM_R_X7Y89_SLICE_X9Y89_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y90_SLICE_X8Y90_A_FDPE (
.C(CLBLM_R_X7Y88_SLICE_X8Y88_AQ),
.CE(1'b1),
.D(CLBLM_R_X7Y90_SLICE_X8Y90_AO6),
.PRE(LIOB33_X0Y107_IOB_X0Y107_I),
.Q(CLBLM_R_X7Y90_SLICE_X8Y90_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y90_SLICE_X8Y90_B_FDPE (
.C(CLBLM_R_X7Y88_SLICE_X8Y88_AQ),
.CE(1'b1),
.D(CLBLM_R_X7Y90_SLICE_X8Y90_BO6),
.PRE(LIOB33_X0Y107_IOB_X0Y107_I),
.Q(CLBLM_R_X7Y90_SLICE_X8Y90_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_R_X7Y90_SLICE_X8Y90_DLUT (
.I0(CLBLM_R_X7Y91_SLICE_X9Y91_CQ),
.I1(CLBLM_R_X7Y90_SLICE_X9Y90_A5Q),
.I2(CLBLM_R_X7Y91_SLICE_X9Y91_BQ),
.I3(CLBLM_R_X7Y90_SLICE_X9Y90_CQ),
.I4(CLBLM_R_X7Y90_SLICE_X9Y90_AQ),
.I5(CLBLM_R_X7Y90_SLICE_X9Y90_BQ),
.O5(CLBLM_R_X7Y90_SLICE_X8Y90_DO5),
.O6(CLBLM_R_X7Y90_SLICE_X8Y90_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X7Y90_SLICE_X8Y90_CLUT (
.I0(CLBLM_R_X7Y91_SLICE_X9Y91_CQ),
.I1(CLBLM_R_X7Y90_SLICE_X9Y90_A5Q),
.I2(CLBLM_R_X7Y91_SLICE_X9Y91_BQ),
.I3(CLBLM_R_X7Y90_SLICE_X9Y90_CQ),
.I4(CLBLM_R_X7Y90_SLICE_X9Y90_AQ),
.I5(CLBLM_R_X7Y90_SLICE_X9Y90_BQ),
.O5(CLBLM_R_X7Y90_SLICE_X8Y90_CO5),
.O6(CLBLM_R_X7Y90_SLICE_X8Y90_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbfbfffffffbfffff)
  ) CLBLM_R_X7Y90_SLICE_X8Y90_BLUT (
.I0(CLBLM_R_X7Y89_SLICE_X9Y89_DO6),
.I1(CLBLM_R_X7Y89_SLICE_X9Y89_BQ),
.I2(CLBLM_R_X7Y89_SLICE_X8Y89_AQ),
.I3(CLBLM_R_X7Y89_SLICE_X8Y89_B5Q),
.I4(CLBLM_R_X7Y89_SLICE_X8Y89_BQ),
.I5(CLBLM_R_X7Y89_SLICE_X9Y89_AO5),
.O5(CLBLM_R_X7Y90_SLICE_X8Y90_BO5),
.O6(CLBLM_R_X7Y90_SLICE_X8Y90_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffdf5f5f7f)
  ) CLBLM_R_X7Y90_SLICE_X8Y90_ALUT (
.I0(CLBLM_R_X7Y87_SLICE_X8Y87_BQ),
.I1(CLBLM_R_X7Y91_SLICE_X9Y91_AQ),
.I2(CLBLM_R_X7Y87_SLICE_X8Y87_AQ),
.I3(CLBLM_R_X7Y90_SLICE_X9Y90_BQ),
.I4(CLBLM_R_X7Y90_SLICE_X9Y90_CQ),
.I5(CLBLM_R_X7Y91_SLICE_X8Y91_AQ),
.O5(CLBLM_R_X7Y90_SLICE_X8Y90_AO5),
.O6(CLBLM_R_X7Y90_SLICE_X8Y90_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y90_SLICE_X9Y90_A5_FDCE (
.C(CLBLM_R_X7Y88_SLICE_X8Y88_AQ),
.CE(1'b1),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_R_X7Y90_SLICE_X9Y90_AO5),
.Q(CLBLM_R_X7Y90_SLICE_X9Y90_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y90_SLICE_X9Y90_A_FDCE (
.C(CLBLM_R_X7Y88_SLICE_X8Y88_AQ),
.CE(1'b1),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_R_X7Y90_SLICE_X9Y90_AO6),
.Q(CLBLM_R_X7Y90_SLICE_X9Y90_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y90_SLICE_X9Y90_B_FDCE (
.C(CLBLM_R_X7Y88_SLICE_X8Y88_AQ),
.CE(1'b1),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_R_X7Y90_SLICE_X9Y90_BO6),
.Q(CLBLM_R_X7Y90_SLICE_X9Y90_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y90_SLICE_X9Y90_C_FDCE (
.C(CLBLM_R_X7Y88_SLICE_X8Y88_AQ),
.CE(1'b1),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_R_X7Y90_SLICE_X9Y90_CO6),
.Q(CLBLM_R_X7Y90_SLICE_X9Y90_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8800000000000000)
  ) CLBLM_R_X7Y90_SLICE_X9Y90_DLUT (
.I0(CLBLM_R_X7Y90_SLICE_X9Y90_BQ),
.I1(CLBLM_R_X7Y91_SLICE_X9Y91_CQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y90_SLICE_X9Y90_A5Q),
.I4(CLBLM_R_X7Y90_SLICE_X9Y90_AQ),
.I5(CLBLM_R_X7Y91_SLICE_X9Y91_BQ),
.O5(CLBLM_R_X7Y90_SLICE_X9Y90_DO5),
.O6(CLBLM_R_X7Y90_SLICE_X9Y90_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h03330ccc13330ccc)
  ) CLBLM_R_X7Y90_SLICE_X9Y90_CLUT (
.I0(CLBLM_R_X7Y91_SLICE_X9Y91_AQ),
.I1(CLBLM_R_X7Y90_SLICE_X9Y90_CQ),
.I2(CLBLM_R_X7Y91_SLICE_X8Y91_AQ),
.I3(CLBLM_R_X7Y87_SLICE_X8Y87_AQ),
.I4(CLBLM_R_X7Y90_SLICE_X9Y90_DO6),
.I5(CLBLM_R_X7Y87_SLICE_X8Y87_BQ),
.O5(CLBLM_R_X7Y90_SLICE_X9Y90_CO5),
.O6(CLBLM_R_X7Y90_SLICE_X9Y90_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1444444444444444)
  ) CLBLM_R_X7Y90_SLICE_X9Y90_BLUT (
.I0(CLBLM_R_X7Y91_SLICE_X9Y91_DO6),
.I1(CLBLM_R_X7Y90_SLICE_X9Y90_BQ),
.I2(CLBLM_R_X7Y90_SLICE_X9Y90_AQ),
.I3(CLBLM_R_X7Y91_SLICE_X9Y91_BQ),
.I4(CLBLM_R_X7Y90_SLICE_X9Y90_A5Q),
.I5(CLBLM_R_X7Y91_SLICE_X9Y91_CQ),
.O5(CLBLM_R_X7Y90_SLICE_X9Y90_BO5),
.O6(CLBLM_R_X7Y90_SLICE_X9Y90_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h1450145015554000)
  ) CLBLM_R_X7Y90_SLICE_X9Y90_ALUT (
.I0(CLBLM_R_X7Y91_SLICE_X9Y91_DO6),
.I1(CLBLM_R_X7Y91_SLICE_X9Y91_BQ),
.I2(CLBLM_R_X7Y90_SLICE_X9Y90_AQ),
.I3(CLBLM_R_X7Y91_SLICE_X9Y91_CQ),
.I4(CLBLM_R_X7Y90_SLICE_X9Y90_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y90_SLICE_X9Y90_AO5),
.O6(CLBLM_R_X7Y90_SLICE_X9Y90_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y91_SLICE_X8Y91_A_FDCE (
.C(CLBLM_R_X7Y88_SLICE_X8Y88_AQ),
.CE(1'b1),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_R_X7Y91_SLICE_X8Y91_AO6),
.Q(CLBLM_R_X7Y91_SLICE_X8Y91_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0010001000f000f0)
  ) CLBLM_R_X7Y91_SLICE_X8Y91_DLUT (
.I0(CLBLM_R_X7Y87_SLICE_X8Y87_BQ),
.I1(CLBLM_R_X7Y91_SLICE_X8Y91_AQ),
.I2(BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO2),
.I3(CLBLM_R_X7Y89_SLICE_X8Y89_CO6),
.I4(1'b1),
.I5(CLBLM_R_X7Y87_SLICE_X8Y87_AQ),
.O5(CLBLM_R_X7Y91_SLICE_X8Y91_DO5),
.O6(CLBLM_R_X7Y91_SLICE_X8Y91_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000010f010f0)
  ) CLBLM_R_X7Y91_SLICE_X8Y91_CLUT (
.I0(CLBLM_R_X7Y87_SLICE_X8Y87_BQ),
.I1(CLBLM_R_X7Y91_SLICE_X8Y91_AQ),
.I2(BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO1),
.I3(CLBLM_R_X7Y87_SLICE_X8Y87_AQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y89_SLICE_X8Y89_CO6),
.O5(CLBLM_R_X7Y91_SLICE_X8Y91_CO5),
.O6(CLBLM_R_X7Y91_SLICE_X8Y91_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0003000000ff0000)
  ) CLBLM_R_X7Y91_SLICE_X8Y91_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y87_SLICE_X8Y87_BQ),
.I2(CLBLM_R_X7Y91_SLICE_X8Y91_AQ),
.I3(CLBLM_R_X7Y89_SLICE_X8Y89_CO6),
.I4(BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO0),
.I5(CLBLM_R_X7Y87_SLICE_X8Y87_AQ),
.O5(CLBLM_R_X7Y91_SLICE_X8Y91_BO5),
.O6(CLBLM_R_X7Y91_SLICE_X8Y91_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0000305af0f0f0)
  ) CLBLM_R_X7Y91_SLICE_X8Y91_ALUT (
.I0(CLBLM_R_X7Y90_SLICE_X8Y90_CO6),
.I1(CLBLM_R_X7Y90_SLICE_X9Y90_CQ),
.I2(CLBLM_R_X7Y91_SLICE_X8Y91_AQ),
.I3(CLBLM_R_X7Y87_SLICE_X8Y87_BQ),
.I4(CLBLM_R_X7Y91_SLICE_X9Y91_AQ),
.I5(CLBLM_R_X7Y87_SLICE_X8Y87_AQ),
.O5(CLBLM_R_X7Y91_SLICE_X8Y91_AO5),
.O6(CLBLM_R_X7Y91_SLICE_X8Y91_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y91_SLICE_X9Y91_A_FDCE (
.C(CLBLM_R_X7Y88_SLICE_X8Y88_AQ),
.CE(1'b1),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_R_X7Y91_SLICE_X9Y91_AO6),
.Q(CLBLM_R_X7Y91_SLICE_X9Y91_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y91_SLICE_X9Y91_B_FDCE (
.C(CLBLM_R_X7Y88_SLICE_X8Y88_AQ),
.CE(1'b1),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_R_X7Y91_SLICE_X9Y91_BO6),
.Q(CLBLM_R_X7Y91_SLICE_X9Y91_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y91_SLICE_X9Y91_C_FDCE (
.C(CLBLM_R_X7Y88_SLICE_X8Y88_AQ),
.CE(1'b1),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_R_X7Y91_SLICE_X9Y91_CO6),
.Q(CLBLM_R_X7Y91_SLICE_X9Y91_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00cc008800)
  ) CLBLM_R_X7Y91_SLICE_X9Y91_DLUT (
.I0(CLBLM_R_X7Y90_SLICE_X9Y90_CQ),
.I1(CLBLM_R_X7Y87_SLICE_X8Y87_AQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y91_SLICE_X8Y91_AQ),
.I4(CLBLM_R_X7Y91_SLICE_X9Y91_AQ),
.I5(CLBLM_R_X7Y87_SLICE_X8Y87_BQ),
.O5(CLBLM_R_X7Y91_SLICE_X9Y91_DO5),
.O6(CLBLM_R_X7Y91_SLICE_X9Y91_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00003c3c00003c3c)
  ) CLBLM_R_X7Y91_SLICE_X9Y91_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y91_SLICE_X9Y91_CQ),
.I2(CLBLM_R_X7Y91_SLICE_X9Y91_BQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y91_SLICE_X9Y91_DO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y91_SLICE_X9Y91_CO5),
.O6(CLBLM_R_X7Y91_SLICE_X9Y91_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1111111333333333)
  ) CLBLM_R_X7Y91_SLICE_X9Y91_BLUT (
.I0(CLBLM_R_X7Y87_SLICE_X8Y87_AQ),
.I1(CLBLM_R_X7Y91_SLICE_X9Y91_BQ),
.I2(CLBLM_R_X7Y91_SLICE_X9Y91_AQ),
.I3(CLBLM_R_X7Y87_SLICE_X8Y87_BQ),
.I4(CLBLM_R_X7Y90_SLICE_X9Y90_CQ),
.I5(CLBLM_R_X7Y91_SLICE_X8Y91_AQ),
.O5(CLBLM_R_X7Y91_SLICE_X9Y91_BO5),
.O6(CLBLM_R_X7Y91_SLICE_X9Y91_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h12125a5a121a5a5a)
  ) CLBLM_R_X7Y91_SLICE_X9Y91_ALUT (
.I0(CLBLM_R_X7Y90_SLICE_X8Y90_CO6),
.I1(CLBLM_R_X7Y87_SLICE_X8Y87_AQ),
.I2(CLBLM_R_X7Y91_SLICE_X9Y91_AQ),
.I3(CLBLM_R_X7Y90_SLICE_X9Y90_CQ),
.I4(CLBLM_R_X7Y91_SLICE_X8Y91_AQ),
.I5(CLBLM_R_X7Y87_SLICE_X8Y87_BQ),
.O5(CLBLM_R_X7Y91_SLICE_X9Y91_AO5),
.O6(CLBLM_R_X7Y91_SLICE_X9Y91_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y93_SLICE_X8Y93_A_FDCE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X7Y94_SLICE_X8Y94_CO6),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_R_X7Y93_SLICE_X8Y93_AO6),
.Q(CLBLM_R_X7Y93_SLICE_X8Y93_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y93_SLICE_X8Y93_B_FDCE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X7Y94_SLICE_X8Y94_CO6),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_R_X7Y93_SLICE_X8Y93_BO6),
.Q(CLBLM_R_X7Y93_SLICE_X8Y93_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcfcfcfcfcfcef)
  ) CLBLM_R_X7Y93_SLICE_X8Y93_DLUT (
.I0(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO11),
.I1(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I2(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO15),
.I3(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO13),
.I4(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO12),
.I5(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO14),
.O5(CLBLM_R_X7Y93_SLICE_X8Y93_DO5),
.O6(CLBLM_R_X7Y93_SLICE_X8Y93_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf2fafafafafafaf8)
  ) CLBLM_R_X7Y93_SLICE_X8Y93_CLUT (
.I0(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO11),
.I1(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO15),
.I2(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I3(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO13),
.I4(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO12),
.I5(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO14),
.O5(CLBLM_R_X7Y93_SLICE_X8Y93_CO5),
.O6(CLBLM_R_X7Y93_SLICE_X8Y93_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000003)
  ) CLBLM_R_X7Y93_SLICE_X8Y93_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I2(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I3(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I4(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I5(CLBLM_R_X7Y93_SLICE_X8Y93_CO6),
.O5(CLBLM_R_X7Y93_SLICE_X8Y93_BO5),
.O6(CLBLM_R_X7Y93_SLICE_X8Y93_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fffffffffffffee)
  ) CLBLM_R_X7Y93_SLICE_X8Y93_ALUT (
.I0(CLBLM_R_X7Y93_SLICE_X8Y93_DO6),
.I1(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I2(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I3(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I4(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I5(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.O5(CLBLM_R_X7Y93_SLICE_X8Y93_AO5),
.O6(CLBLM_R_X7Y93_SLICE_X8Y93_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y93_SLICE_X9Y93_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y93_SLICE_X9Y93_DO5),
.O6(CLBLM_R_X7Y93_SLICE_X9Y93_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y93_SLICE_X9Y93_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y93_SLICE_X9Y93_CO5),
.O6(CLBLM_R_X7Y93_SLICE_X9Y93_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y93_SLICE_X9Y93_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y93_SLICE_X9Y93_BO5),
.O6(CLBLM_R_X7Y93_SLICE_X9Y93_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y93_SLICE_X9Y93_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y93_SLICE_X9Y93_AO5),
.O6(CLBLM_R_X7Y93_SLICE_X9Y93_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y94_SLICE_X8Y94_A_FDCE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X7Y94_SLICE_X8Y94_CO6),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_R_X7Y94_SLICE_X8Y94_AO6),
.Q(CLBLM_R_X7Y94_SLICE_X8Y94_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y94_SLICE_X8Y94_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y94_SLICE_X8Y94_DO5),
.O6(CLBLM_R_X7Y94_SLICE_X8Y94_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h77ffffffffffffff)
  ) CLBLM_R_X7Y94_SLICE_X8Y94_CLUT (
.I0(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I1(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I4(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I5(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.O5(CLBLM_R_X7Y94_SLICE_X8Y94_CO5),
.O6(CLBLM_R_X7Y94_SLICE_X8Y94_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcfcfcfcfcfdf3)
  ) CLBLM_R_X7Y94_SLICE_X8Y94_BLUT (
.I0(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO15),
.I1(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO14),
.I2(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I3(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO11),
.I4(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO12),
.I5(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO13),
.O5(CLBLM_R_X7Y94_SLICE_X8Y94_BO5),
.O6(CLBLM_R_X7Y94_SLICE_X8Y94_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f7fffff7f7fffee)
  ) CLBLM_R_X7Y94_SLICE_X8Y94_ALUT (
.I0(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I1(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I2(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I3(CLBLM_R_X7Y94_SLICE_X8Y94_BO6),
.I4(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I5(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.O5(CLBLM_R_X7Y94_SLICE_X8Y94_AO5),
.O6(CLBLM_R_X7Y94_SLICE_X8Y94_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y94_SLICE_X9Y94_A_FDCE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X7Y94_SLICE_X8Y94_CO6),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_R_X7Y94_SLICE_X9Y94_AO6),
.Q(CLBLM_R_X7Y94_SLICE_X9Y94_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y94_SLICE_X9Y94_B_FDCE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X7Y94_SLICE_X8Y94_CO6),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_R_X7Y94_SLICE_X9Y94_BO6),
.Q(CLBLM_R_X7Y94_SLICE_X9Y94_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaffabeebbeebb)
  ) CLBLM_R_X7Y94_SLICE_X9Y94_DLUT (
.I0(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I1(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO12),
.I2(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO15),
.I3(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO13),
.I4(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO14),
.I5(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO11),
.O5(CLBLM_R_X7Y94_SLICE_X9Y94_DO5),
.O6(CLBLM_R_X7Y94_SLICE_X9Y94_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haeeeeeeebbbbbbba)
  ) CLBLM_R_X7Y94_SLICE_X9Y94_CLUT (
.I0(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I1(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO11),
.I2(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO15),
.I3(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO13),
.I4(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO14),
.I5(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO12),
.O5(CLBLM_R_X7Y94_SLICE_X9Y94_CO5),
.O6(CLBLM_R_X7Y94_SLICE_X9Y94_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f7fffff7f7efffe)
  ) CLBLM_R_X7Y94_SLICE_X9Y94_BLUT (
.I0(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I1(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I2(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I3(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I4(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I5(CLBLM_R_X7Y94_SLICE_X9Y94_CO6),
.O5(CLBLM_R_X7Y94_SLICE_X9Y94_BO5),
.O6(CLBLM_R_X7Y94_SLICE_X9Y94_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3ffffffffefffe)
  ) CLBLM_R_X7Y94_SLICE_X9Y94_ALUT (
.I0(CLBLM_R_X7Y94_SLICE_X9Y94_DO6),
.I1(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I2(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I3(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I4(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I5(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.O5(CLBLM_R_X7Y94_SLICE_X9Y94_AO5),
.O6(CLBLM_R_X7Y94_SLICE_X9Y94_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y96_SLICE_X8Y96_A_FDCE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X7Y99_SLICE_X9Y99_DO6),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_R_X7Y96_SLICE_X8Y96_AO6),
.Q(CLBLM_R_X7Y96_SLICE_X8Y96_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa88a000220aaa00)
  ) CLBLM_R_X7Y96_SLICE_X8Y96_DLUT (
.I0(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO6),
.I1(CLBLM_R_X5Y95_SLICE_X6Y95_AQ),
.I2(CLBLL_L_X4Y97_SLICE_X4Y97_BQ),
.I3(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I4(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I5(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.O5(CLBLM_R_X7Y96_SLICE_X8Y96_DO5),
.O6(CLBLM_R_X7Y96_SLICE_X8Y96_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X7Y96_SLICE_X8Y96_CLUT (
.I0(CLBLM_R_X5Y96_SLICE_X6Y96_AQ),
.I1(CLBLM_R_X5Y99_SLICE_X7Y99_AQ),
.I2(CLBLM_R_X5Y96_SLICE_X7Y96_AQ),
.I3(CLBLM_R_X7Y99_SLICE_X8Y99_AQ),
.I4(CLBLM_R_X5Y99_SLICE_X6Y99_AQ),
.I5(CLBLM_R_X5Y96_SLICE_X7Y96_BQ),
.O5(CLBLM_R_X7Y96_SLICE_X8Y96_CO5),
.O6(CLBLM_R_X7Y96_SLICE_X8Y96_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0ff0f05a5aaaaa)
  ) CLBLM_R_X7Y96_SLICE_X8Y96_BLUT (
.I0(CLBLM_R_X7Y96_SLICE_X9Y96_AQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y96_SLICE_X8Y96_AQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y96_SLICE_X8Y96_CO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y96_SLICE_X8Y96_BO5),
.O6(CLBLM_R_X7Y96_SLICE_X8Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0ca0a0ff00ff00)
  ) CLBLM_R_X7Y96_SLICE_X8Y96_ALUT (
.I0(CLBLM_R_X7Y96_SLICE_X8Y96_DO6),
.I1(CLBLM_R_X7Y96_SLICE_X9Y96_BO6),
.I2(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I3(CLBLM_R_X7Y96_SLICE_X8Y96_BO6),
.I4(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I5(CLBLM_R_X7Y98_SLICE_X8Y98_F7AMUX_O),
.O5(CLBLM_R_X7Y96_SLICE_X8Y96_AO5),
.O6(CLBLM_R_X7Y96_SLICE_X8Y96_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y96_SLICE_X9Y96_A_FDCE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X7Y99_SLICE_X9Y99_DO6),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_R_X7Y96_SLICE_X9Y96_AO6),
.Q(CLBLM_R_X7Y96_SLICE_X9Y96_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa77880a00000000)
  ) CLBLM_R_X7Y96_SLICE_X9Y96_DLUT (
.I0(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I1(CLBLM_R_X5Y95_SLICE_X6Y95_AQ),
.I2(CLBLL_L_X4Y97_SLICE_X4Y97_BQ),
.I3(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I4(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I5(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO7),
.O5(CLBLM_R_X7Y96_SLICE_X9Y96_DO5),
.O6(CLBLM_R_X7Y96_SLICE_X9Y96_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h505050d85050d850)
  ) CLBLM_R_X7Y96_SLICE_X9Y96_CLUT (
.I0(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I1(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO7),
.I2(CLBLM_L_X8Y97_SLICE_X11Y97_AO6),
.I3(CLBLM_R_X5Y95_SLICE_X6Y95_AQ),
.I4(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I5(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.O5(CLBLM_R_X7Y96_SLICE_X9Y96_CO5),
.O6(CLBLM_R_X7Y96_SLICE_X9Y96_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a3a0a0a3a0a0a0a)
  ) CLBLM_R_X7Y96_SLICE_X9Y96_BLUT (
.I0(CLBLM_L_X8Y97_SLICE_X10Y97_CO6),
.I1(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I2(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I3(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I4(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO6),
.I5(CLBLM_R_X5Y95_SLICE_X6Y95_AQ),
.O5(CLBLM_R_X7Y96_SLICE_X9Y96_BO5),
.O6(CLBLM_R_X7Y96_SLICE_X9Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fa0cccc00a0cccc)
  ) CLBLM_R_X7Y96_SLICE_X9Y96_ALUT (
.I0(CLBLM_R_X7Y96_SLICE_X9Y96_DO6),
.I1(CLBLM_R_X7Y96_SLICE_X8Y96_BO5),
.I2(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I3(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I4(CLBLM_R_X7Y98_SLICE_X8Y98_F7AMUX_O),
.I5(CLBLM_R_X7Y96_SLICE_X9Y96_CO6),
.O5(CLBLM_R_X7Y96_SLICE_X9Y96_AO5),
.O6(CLBLM_R_X7Y96_SLICE_X9Y96_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y97_SLICE_X8Y97_A_FDCE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X7Y99_SLICE_X9Y99_DO6),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_R_X7Y97_SLICE_X8Y97_AO6),
.Q(CLBLM_R_X7Y97_SLICE_X8Y97_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6ccccccccccccccc)
  ) CLBLM_R_X7Y97_SLICE_X8Y97_DLUT (
.I0(CLBLM_R_X7Y99_SLICE_X9Y99_AQ),
.I1(CLBLM_R_X7Y97_SLICE_X8Y97_AQ),
.I2(CLBLM_R_X7Y96_SLICE_X8Y96_AQ),
.I3(CLBLM_R_X7Y96_SLICE_X8Y96_CO6),
.I4(CLBLM_R_X7Y96_SLICE_X9Y96_AQ),
.I5(CLBLM_R_X7Y98_SLICE_X9Y98_AQ),
.O5(CLBLM_R_X7Y97_SLICE_X8Y97_DO5),
.O6(CLBLM_R_X7Y97_SLICE_X8Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f07250f0f0d850)
  ) CLBLM_R_X7Y97_SLICE_X8Y97_CLUT (
.I0(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I1(CLBLM_R_X5Y95_SLICE_X6Y95_AQ),
.I2(CLBLM_R_X7Y98_SLICE_X8Y98_DO6),
.I3(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO10),
.I4(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I5(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.O5(CLBLM_R_X7Y97_SLICE_X8Y97_CO5),
.O6(CLBLM_R_X7Y97_SLICE_X8Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7788ff0078f0f0f0)
  ) CLBLM_R_X7Y97_SLICE_X8Y97_BLUT (
.I0(CLBLM_R_X7Y96_SLICE_X9Y96_AQ),
.I1(CLBLM_R_X7Y96_SLICE_X8Y96_CO6),
.I2(CLBLM_R_X7Y99_SLICE_X9Y99_AQ),
.I3(CLBLM_R_X7Y98_SLICE_X9Y98_AQ),
.I4(CLBLM_R_X7Y96_SLICE_X8Y96_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y97_SLICE_X8Y97_BO5),
.O6(CLBLM_R_X7Y97_SLICE_X8Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f0cb3803300b380)
  ) CLBLM_R_X7Y97_SLICE_X8Y97_ALUT (
.I0(CLBLM_R_X7Y98_SLICE_X8Y98_CO6),
.I1(CLBLM_R_X7Y98_SLICE_X8Y98_F7AMUX_O),
.I2(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I3(CLBLM_R_X7Y97_SLICE_X8Y97_DO6),
.I4(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I5(CLBLM_R_X7Y97_SLICE_X8Y97_CO6),
.O5(CLBLM_R_X7Y97_SLICE_X8Y97_AO5),
.O6(CLBLM_R_X7Y97_SLICE_X8Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y97_SLICE_X9Y97_A5_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X7Y97_SLICE_X9Y97_CO6),
.D(CLBLM_R_X7Y97_SLICE_X9Y97_AO5),
.Q(CLBLM_R_X7Y97_SLICE_X9Y97_A5Q),
.R(LIOB33_X0Y107_IOB_X0Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y97_SLICE_X9Y97_B5_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X7Y97_SLICE_X9Y97_CO6),
.D(CLBLM_R_X7Y97_SLICE_X9Y97_BO5),
.Q(CLBLM_R_X7Y97_SLICE_X9Y97_B5Q),
.R(LIOB33_X0Y107_IOB_X0Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y97_SLICE_X9Y97_A_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X7Y97_SLICE_X9Y97_CO6),
.D(CLBLM_R_X7Y97_SLICE_X9Y97_AO6),
.Q(CLBLM_R_X7Y97_SLICE_X9Y97_AQ),
.R(LIOB33_X0Y107_IOB_X0Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y97_SLICE_X9Y97_B_FDRE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X7Y97_SLICE_X9Y97_CO6),
.D(CLBLM_R_X7Y97_SLICE_X9Y97_BO6),
.Q(CLBLM_R_X7Y97_SLICE_X9Y97_BQ),
.R(LIOB33_X0Y107_IOB_X0Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00ff00fe00)
  ) CLBLM_R_X7Y97_SLICE_X9Y97_DLUT (
.I0(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I1(CLBLM_R_X5Y95_SLICE_X6Y95_CO6),
.I2(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I3(CLBLL_L_X4Y97_SLICE_X5Y97_DO6),
.I4(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I5(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.O5(CLBLM_R_X7Y97_SLICE_X9Y97_DO5),
.O6(CLBLM_R_X7Y97_SLICE_X9Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2666666666666664)
  ) CLBLM_R_X7Y97_SLICE_X9Y97_CLUT (
.I0(CLBLM_R_X5Y95_SLICE_X6Y95_BO5),
.I1(CLBLL_L_X4Y97_SLICE_X5Y97_DO6),
.I2(CLBLM_R_X7Y97_SLICE_X9Y97_BQ),
.I3(CLBLM_R_X7Y97_SLICE_X9Y97_A5Q),
.I4(CLBLM_R_X7Y97_SLICE_X9Y97_B5Q),
.I5(CLBLM_R_X7Y97_SLICE_X9Y97_AQ),
.O5(CLBLM_R_X7Y97_SLICE_X9Y97_CO5),
.O6(CLBLM_R_X7Y97_SLICE_X9Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hec6cc9c9ff80fe01)
  ) CLBLM_R_X7Y97_SLICE_X9Y97_BLUT (
.I0(CLBLM_R_X7Y97_SLICE_X9Y97_DO6),
.I1(CLBLM_R_X7Y97_SLICE_X9Y97_BQ),
.I2(CLBLM_R_X7Y97_SLICE_X9Y97_AQ),
.I3(CLBLM_R_X7Y97_SLICE_X9Y97_B5Q),
.I4(CLBLM_R_X7Y97_SLICE_X9Y97_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y97_SLICE_X9Y97_BO5),
.O6(CLBLM_R_X7Y97_SLICE_X9Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0fda5aa5a5)
  ) CLBLM_R_X7Y97_SLICE_X9Y97_ALUT (
.I0(CLBLM_R_X7Y97_SLICE_X9Y97_DO6),
.I1(CLBLM_R_X7Y97_SLICE_X9Y97_BQ),
.I2(CLBLM_R_X7Y97_SLICE_X9Y97_AQ),
.I3(CLBLM_R_X7Y97_SLICE_X9Y97_B5Q),
.I4(CLBLM_R_X7Y97_SLICE_X9Y97_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y97_SLICE_X9Y97_AO5),
.O6(CLBLM_R_X7Y97_SLICE_X9Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000404000008f80)
  ) CLBLM_R_X7Y98_SLICE_X8Y98_DLUT (
.I0(CLBLL_L_X4Y97_SLICE_X4Y97_BQ),
.I1(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO10),
.I2(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I3(CLBLM_L_X8Y98_SLICE_X10Y98_BO6),
.I4(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I5(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.O5(CLBLM_R_X7Y98_SLICE_X8Y98_DO5),
.O6(CLBLM_R_X7Y98_SLICE_X8Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccc0808004c4c0c0)
  ) CLBLM_R_X7Y98_SLICE_X8Y98_CLUT (
.I0(CLBLL_L_X4Y97_SLICE_X4Y97_BQ),
.I1(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO10),
.I2(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I3(CLBLM_R_X5Y95_SLICE_X6Y95_AQ),
.I4(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I5(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.O5(CLBLM_R_X7Y98_SLICE_X8Y98_CO5),
.O6(CLBLM_R_X7Y98_SLICE_X8Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1300190043004900)
  ) CLBLM_R_X7Y98_SLICE_X8Y98_BLUT (
.I0(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I1(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I2(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I3(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I4(CLBLL_L_X4Y97_SLICE_X4Y97_BQ),
.I5(CLBLM_R_X5Y95_SLICE_X6Y95_AQ),
.O5(CLBLM_R_X7Y98_SLICE_X8Y98_BO5),
.O6(CLBLM_R_X7Y98_SLICE_X8Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ca00d200aa00b2)
  ) CLBLM_R_X7Y98_SLICE_X8Y98_ALUT (
.I0(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I1(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I2(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I3(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I4(CLBLL_L_X4Y97_SLICE_X4Y97_BQ),
.I5(CLBLM_R_X5Y95_SLICE_X6Y95_AQ),
.O5(CLBLM_R_X7Y98_SLICE_X8Y98_AO5),
.O6(CLBLM_R_X7Y98_SLICE_X8Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_R_X7Y98_SLICE_X8Y98_MUXF7A (
.I0(CLBLM_R_X7Y98_SLICE_X8Y98_BO6),
.I1(CLBLM_R_X7Y98_SLICE_X8Y98_AO6),
.O(CLBLM_R_X7Y98_SLICE_X8Y98_F7AMUX_O),
.S(CLBLM_R_X7Y94_SLICE_X8Y94_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y98_SLICE_X9Y98_A_FDCE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X7Y99_SLICE_X9Y99_DO6),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_R_X7Y98_SLICE_X9Y98_AO6),
.Q(CLBLM_R_X7Y98_SLICE_X9Y98_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y98_SLICE_X9Y98_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y98_SLICE_X9Y98_DO5),
.O6(CLBLM_R_X7Y98_SLICE_X9Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hece0000034f40000)
  ) CLBLM_R_X7Y98_SLICE_X9Y98_CLUT (
.I0(CLBLL_L_X4Y97_SLICE_X4Y97_BQ),
.I1(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I2(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I3(CLBLM_R_X5Y95_SLICE_X6Y95_AQ),
.I4(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO8),
.I5(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.O5(CLBLM_R_X7Y98_SLICE_X9Y98_CO5),
.O6(CLBLM_R_X7Y98_SLICE_X9Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c5c5c0c0c0c0c0c)
  ) CLBLM_R_X7Y98_SLICE_X9Y98_BLUT (
.I0(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I1(CLBLM_L_X8Y98_SLICE_X10Y98_CO6),
.I2(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I3(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I4(CLBLM_R_X5Y95_SLICE_X6Y95_AQ),
.I5(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO8),
.O5(CLBLM_R_X7Y98_SLICE_X9Y98_BO5),
.O6(CLBLM_R_X7Y98_SLICE_X9Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6f2f60204f0f4000)
  ) CLBLM_R_X7Y98_SLICE_X9Y98_ALUT (
.I0(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I1(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I2(CLBLM_R_X7Y98_SLICE_X8Y98_F7AMUX_O),
.I3(CLBLM_R_X7Y98_SLICE_X9Y98_BO6),
.I4(CLBLM_R_X7Y97_SLICE_X8Y97_BO6),
.I5(CLBLM_R_X7Y98_SLICE_X9Y98_CO6),
.O5(CLBLM_R_X7Y98_SLICE_X9Y98_AO5),
.O6(CLBLM_R_X7Y98_SLICE_X9Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y99_SLICE_X8Y99_A_FDCE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X7Y99_SLICE_X9Y99_DO6),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_R_X7Y99_SLICE_X8Y99_AO6),
.Q(CLBLM_R_X7Y99_SLICE_X8Y99_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0020002020002303)
  ) CLBLM_R_X7Y99_SLICE_X8Y99_DLUT (
.I0(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO0),
.I1(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I2(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I3(CLBLL_L_X4Y97_SLICE_X4Y97_BQ),
.I4(CLBLM_R_X5Y98_SLICE_X6Y98_DO6),
.I5(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.O5(CLBLM_R_X7Y99_SLICE_X8Y99_DO5),
.O6(CLBLM_R_X7Y99_SLICE_X8Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaa080802a2a00a0)
  ) CLBLM_R_X7Y99_SLICE_X8Y99_CLUT (
.I0(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO0),
.I1(CLBLM_R_X5Y95_SLICE_X6Y95_AQ),
.I2(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I3(CLBLL_L_X4Y97_SLICE_X4Y97_BQ),
.I4(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I5(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.O5(CLBLM_R_X7Y99_SLICE_X8Y99_CO5),
.O6(CLBLM_R_X7Y99_SLICE_X8Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa30aaaaaac0aaaa)
  ) CLBLM_R_X7Y99_SLICE_X8Y99_BLUT (
.I0(CLBLM_R_X7Y99_SLICE_X8Y99_DO6),
.I1(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I2(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO0),
.I3(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I4(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I5(CLBLM_R_X5Y95_SLICE_X6Y95_AQ),
.O5(CLBLM_R_X7Y99_SLICE_X8Y99_BO5),
.O6(CLBLM_R_X7Y99_SLICE_X8Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h47038b8b47030303)
  ) CLBLM_R_X7Y99_SLICE_X8Y99_ALUT (
.I0(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I1(CLBLM_R_X7Y98_SLICE_X8Y98_F7AMUX_O),
.I2(CLBLM_R_X7Y99_SLICE_X8Y99_AQ),
.I3(CLBLM_R_X7Y99_SLICE_X8Y99_BO6),
.I4(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I5(CLBLM_R_X7Y99_SLICE_X8Y99_CO6),
.O5(CLBLM_R_X7Y99_SLICE_X8Y99_AO5),
.O6(CLBLM_R_X7Y99_SLICE_X8Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y99_SLICE_X9Y99_A_FDCE (
.C(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.CE(CLBLM_R_X7Y99_SLICE_X9Y99_DO6),
.CLR(LIOB33_X0Y107_IOB_X0Y107_I),
.D(CLBLM_R_X7Y99_SLICE_X9Y99_AO6),
.Q(CLBLM_R_X7Y99_SLICE_X9Y99_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ffffffffffffffa)
  ) CLBLM_R_X7Y99_SLICE_X9Y99_DLUT (
.I0(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I3(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I4(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I5(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.O5(CLBLM_R_X7Y99_SLICE_X9Y99_DO5),
.O6(CLBLM_R_X7Y99_SLICE_X9Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccc0808004c4c0c0)
  ) CLBLM_R_X7Y99_SLICE_X9Y99_CLUT (
.I0(CLBLL_L_X4Y97_SLICE_X4Y97_BQ),
.I1(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO9),
.I2(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I3(CLBLM_R_X5Y95_SLICE_X6Y95_AQ),
.I4(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I5(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.O5(CLBLM_R_X7Y99_SLICE_X9Y99_CO5),
.O6(CLBLM_R_X7Y99_SLICE_X9Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0044f0f04400f0f0)
  ) CLBLM_R_X7Y99_SLICE_X9Y99_BLUT (
.I0(CLBLM_R_X7Y94_SLICE_X9Y94_BQ),
.I1(BRAM_L_X6Y95_RAMB36_X0Y19_DOADO9),
.I2(CLBLM_L_X8Y98_SLICE_X10Y98_DO6),
.I3(CLBLM_R_X7Y93_SLICE_X8Y93_BQ),
.I4(CLBLM_R_X7Y94_SLICE_X9Y94_AQ),
.I5(CLBLM_R_X5Y95_SLICE_X6Y95_AQ),
.O5(CLBLM_R_X7Y99_SLICE_X9Y99_BO5),
.O6(CLBLM_R_X7Y99_SLICE_X9Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a0acccc5000cccc)
  ) CLBLM_R_X7Y99_SLICE_X9Y99_ALUT (
.I0(CLBLM_R_X7Y94_SLICE_X8Y94_AQ),
.I1(CLBLM_R_X7Y97_SLICE_X8Y97_BO5),
.I2(CLBLM_R_X7Y93_SLICE_X8Y93_AQ),
.I3(CLBLM_R_X7Y99_SLICE_X9Y99_BO6),
.I4(CLBLM_R_X7Y98_SLICE_X8Y98_F7AMUX_O),
.I5(CLBLM_R_X7Y99_SLICE_X9Y99_CO6),
.O5(CLBLM_R_X7Y99_SLICE_X9Y99_AO5),
.O6(CLBLM_R_X7Y99_SLICE_X9Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(LIOB33_X0Y127_IOB_X0Y128_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12.0"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y101_OBUF (
.I(CLBLM_R_X7Y91_SLICE_X8Y91_CO6),
.O(g)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12.0"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y102_OBUF (
.I(CLBLL_L_X4Y90_SLICE_X5Y90_AQ),
.O(hs)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12.0"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y103_OBUF (
.I(CLBLM_R_X7Y91_SLICE_X8Y91_DO6),
.O(r)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12.0"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y104_OBUF (
.I(CLBLL_L_X2Y102_SLICE_X0Y102_AQ),
.O(vs)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y105_IOB_X0Y105_IBUF (
.I(down1),
.O(LIOB33_X0Y105_IOB_X0Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y105_IOB_X0Y106_IBUF (
.I(down2),
.O(LIOB33_X0Y105_IOB_X0Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y107_IOB_X0Y107_IBUF (
.I(rst),
.O(LIOB33_X0Y107_IOB_X0Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y107_IOB_X0Y108_IBUF (
.I(up1),
.O(LIOB33_X0Y107_IOB_X0Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y109_IOB_X0Y109_IBUF (
.I(up2),
.O(LIOB33_X0Y109_IOB_X0Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y127_IOB_X0Y128_IBUF (
.I(clk),
.O(LIOB33_X0Y127_IOB_X0Y128_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12.0"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y100_IOB_X0Y100_OBUF (
.I(CLBLM_R_X7Y91_SLICE_X8Y91_BO6),
.O(b)
  );
  assign CLBLL_L_X2Y90_SLICE_X0Y90_COUT = CLBLL_L_X2Y90_SLICE_X0Y90_D_CY;
  assign CLBLL_L_X2Y90_SLICE_X0Y90_A = CLBLL_L_X2Y90_SLICE_X0Y90_AO6;
  assign CLBLL_L_X2Y90_SLICE_X0Y90_B = CLBLL_L_X2Y90_SLICE_X0Y90_BO6;
  assign CLBLL_L_X2Y90_SLICE_X0Y90_C = CLBLL_L_X2Y90_SLICE_X0Y90_CO6;
  assign CLBLL_L_X2Y90_SLICE_X0Y90_D = CLBLL_L_X2Y90_SLICE_X0Y90_DO6;
  assign CLBLL_L_X2Y90_SLICE_X1Y90_COUT = CLBLL_L_X2Y90_SLICE_X1Y90_D_CY;
  assign CLBLL_L_X2Y90_SLICE_X1Y90_A = CLBLL_L_X2Y90_SLICE_X1Y90_AO6;
  assign CLBLL_L_X2Y90_SLICE_X1Y90_B = CLBLL_L_X2Y90_SLICE_X1Y90_BO6;
  assign CLBLL_L_X2Y90_SLICE_X1Y90_C = CLBLL_L_X2Y90_SLICE_X1Y90_CO6;
  assign CLBLL_L_X2Y90_SLICE_X1Y90_D = CLBLL_L_X2Y90_SLICE_X1Y90_DO6;
  assign CLBLL_L_X2Y91_SLICE_X0Y91_COUT = CLBLL_L_X2Y91_SLICE_X0Y91_D_CY;
  assign CLBLL_L_X2Y91_SLICE_X0Y91_A = CLBLL_L_X2Y91_SLICE_X0Y91_AO6;
  assign CLBLL_L_X2Y91_SLICE_X0Y91_B = CLBLL_L_X2Y91_SLICE_X0Y91_BO6;
  assign CLBLL_L_X2Y91_SLICE_X0Y91_C = CLBLL_L_X2Y91_SLICE_X0Y91_CO6;
  assign CLBLL_L_X2Y91_SLICE_X0Y91_D = CLBLL_L_X2Y91_SLICE_X0Y91_DO6;
  assign CLBLL_L_X2Y91_SLICE_X1Y91_COUT = CLBLL_L_X2Y91_SLICE_X1Y91_D_CY;
  assign CLBLL_L_X2Y91_SLICE_X1Y91_A = CLBLL_L_X2Y91_SLICE_X1Y91_AO6;
  assign CLBLL_L_X2Y91_SLICE_X1Y91_B = CLBLL_L_X2Y91_SLICE_X1Y91_BO6;
  assign CLBLL_L_X2Y91_SLICE_X1Y91_C = CLBLL_L_X2Y91_SLICE_X1Y91_CO6;
  assign CLBLL_L_X2Y91_SLICE_X1Y91_D = CLBLL_L_X2Y91_SLICE_X1Y91_DO6;
  assign CLBLL_L_X2Y92_SLICE_X0Y92_COUT = CLBLL_L_X2Y92_SLICE_X0Y92_D_CY;
  assign CLBLL_L_X2Y92_SLICE_X0Y92_A = CLBLL_L_X2Y92_SLICE_X0Y92_AO6;
  assign CLBLL_L_X2Y92_SLICE_X0Y92_B = CLBLL_L_X2Y92_SLICE_X0Y92_BO6;
  assign CLBLL_L_X2Y92_SLICE_X0Y92_C = CLBLL_L_X2Y92_SLICE_X0Y92_CO6;
  assign CLBLL_L_X2Y92_SLICE_X0Y92_D = CLBLL_L_X2Y92_SLICE_X0Y92_DO6;
  assign CLBLL_L_X2Y92_SLICE_X1Y92_COUT = CLBLL_L_X2Y92_SLICE_X1Y92_D_CY;
  assign CLBLL_L_X2Y92_SLICE_X1Y92_A = CLBLL_L_X2Y92_SLICE_X1Y92_AO6;
  assign CLBLL_L_X2Y92_SLICE_X1Y92_B = CLBLL_L_X2Y92_SLICE_X1Y92_BO6;
  assign CLBLL_L_X2Y92_SLICE_X1Y92_C = CLBLL_L_X2Y92_SLICE_X1Y92_CO6;
  assign CLBLL_L_X2Y92_SLICE_X1Y92_D = CLBLL_L_X2Y92_SLICE_X1Y92_DO6;
  assign CLBLL_L_X2Y93_SLICE_X0Y93_COUT = CLBLL_L_X2Y93_SLICE_X0Y93_D_CY;
  assign CLBLL_L_X2Y93_SLICE_X0Y93_A = CLBLL_L_X2Y93_SLICE_X0Y93_AO6;
  assign CLBLL_L_X2Y93_SLICE_X0Y93_B = CLBLL_L_X2Y93_SLICE_X0Y93_BO6;
  assign CLBLL_L_X2Y93_SLICE_X0Y93_C = CLBLL_L_X2Y93_SLICE_X0Y93_CO6;
  assign CLBLL_L_X2Y93_SLICE_X0Y93_D = CLBLL_L_X2Y93_SLICE_X0Y93_DO6;
  assign CLBLL_L_X2Y93_SLICE_X0Y93_AMUX = CLBLL_L_X2Y93_SLICE_X0Y93_F7AMUX_O;
  assign CLBLL_L_X2Y93_SLICE_X0Y93_CMUX = CLBLL_L_X2Y93_SLICE_X0Y93_CO5;
  assign CLBLL_L_X2Y93_SLICE_X0Y93_DMUX = CLBLL_L_X2Y93_SLICE_X0Y93_DO6;
  assign CLBLL_L_X2Y93_SLICE_X1Y93_COUT = CLBLL_L_X2Y93_SLICE_X1Y93_D_CY;
  assign CLBLL_L_X2Y93_SLICE_X1Y93_A = CLBLL_L_X2Y93_SLICE_X1Y93_AO6;
  assign CLBLL_L_X2Y93_SLICE_X1Y93_B = CLBLL_L_X2Y93_SLICE_X1Y93_BO6;
  assign CLBLL_L_X2Y93_SLICE_X1Y93_C = CLBLL_L_X2Y93_SLICE_X1Y93_CO6;
  assign CLBLL_L_X2Y93_SLICE_X1Y93_D = CLBLL_L_X2Y93_SLICE_X1Y93_DO6;
  assign CLBLL_L_X2Y93_SLICE_X1Y93_AMUX = CLBLL_L_X2Y93_SLICE_X1Y93_F7AMUX_O;
  assign CLBLL_L_X2Y93_SLICE_X1Y93_DMUX = CLBLL_L_X2Y93_SLICE_X1Y93_DO6;
  assign CLBLL_L_X2Y94_SLICE_X0Y94_COUT = CLBLL_L_X2Y94_SLICE_X0Y94_D_CY;
  assign CLBLL_L_X2Y94_SLICE_X0Y94_A = CLBLL_L_X2Y94_SLICE_X0Y94_AO6;
  assign CLBLL_L_X2Y94_SLICE_X0Y94_B = CLBLL_L_X2Y94_SLICE_X0Y94_BO6;
  assign CLBLL_L_X2Y94_SLICE_X0Y94_C = CLBLL_L_X2Y94_SLICE_X0Y94_CO6;
  assign CLBLL_L_X2Y94_SLICE_X0Y94_D = CLBLL_L_X2Y94_SLICE_X0Y94_DO6;
  assign CLBLL_L_X2Y94_SLICE_X0Y94_CMUX = CLBLL_L_X2Y94_SLICE_X0Y94_CO6;
  assign CLBLL_L_X2Y94_SLICE_X0Y94_DMUX = CLBLL_L_X2Y94_SLICE_X0Y94_DO6;
  assign CLBLL_L_X2Y94_SLICE_X1Y94_COUT = CLBLL_L_X2Y94_SLICE_X1Y94_D_CY;
  assign CLBLL_L_X2Y94_SLICE_X1Y94_A = CLBLL_L_X2Y94_SLICE_X1Y94_AO6;
  assign CLBLL_L_X2Y94_SLICE_X1Y94_B = CLBLL_L_X2Y94_SLICE_X1Y94_BO6;
  assign CLBLL_L_X2Y94_SLICE_X1Y94_C = CLBLL_L_X2Y94_SLICE_X1Y94_CO6;
  assign CLBLL_L_X2Y94_SLICE_X1Y94_D = CLBLL_L_X2Y94_SLICE_X1Y94_DO6;
  assign CLBLL_L_X2Y94_SLICE_X1Y94_AMUX = CLBLL_L_X2Y94_SLICE_X1Y94_A_XOR;
  assign CLBLL_L_X2Y94_SLICE_X1Y94_BMUX = CLBLL_L_X2Y94_SLICE_X1Y94_B_XOR;
  assign CLBLL_L_X2Y94_SLICE_X1Y94_CMUX = CLBLL_L_X2Y94_SLICE_X1Y94_C_XOR;
  assign CLBLL_L_X2Y94_SLICE_X1Y94_DMUX = CLBLL_L_X2Y94_SLICE_X1Y94_D_XOR;
  assign CLBLL_L_X2Y95_SLICE_X0Y95_COUT = CLBLL_L_X2Y95_SLICE_X0Y95_D_CY;
  assign CLBLL_L_X2Y95_SLICE_X0Y95_A = CLBLL_L_X2Y95_SLICE_X0Y95_AO6;
  assign CLBLL_L_X2Y95_SLICE_X0Y95_B = CLBLL_L_X2Y95_SLICE_X0Y95_BO6;
  assign CLBLL_L_X2Y95_SLICE_X0Y95_C = CLBLL_L_X2Y95_SLICE_X0Y95_CO6;
  assign CLBLL_L_X2Y95_SLICE_X0Y95_D = CLBLL_L_X2Y95_SLICE_X0Y95_DO6;
  assign CLBLL_L_X2Y95_SLICE_X0Y95_DMUX = CLBLL_L_X2Y95_SLICE_X0Y95_D_CY;
  assign CLBLL_L_X2Y95_SLICE_X1Y95_COUT = CLBLL_L_X2Y95_SLICE_X1Y95_D_CY;
  assign CLBLL_L_X2Y95_SLICE_X1Y95_A = CLBLL_L_X2Y95_SLICE_X1Y95_AO6;
  assign CLBLL_L_X2Y95_SLICE_X1Y95_B = CLBLL_L_X2Y95_SLICE_X1Y95_BO6;
  assign CLBLL_L_X2Y95_SLICE_X1Y95_C = CLBLL_L_X2Y95_SLICE_X1Y95_CO6;
  assign CLBLL_L_X2Y95_SLICE_X1Y95_D = CLBLL_L_X2Y95_SLICE_X1Y95_DO6;
  assign CLBLL_L_X2Y95_SLICE_X1Y95_AMUX = CLBLL_L_X2Y95_SLICE_X1Y95_A_XOR;
  assign CLBLL_L_X2Y95_SLICE_X1Y95_BMUX = CLBLL_L_X2Y95_SLICE_X1Y95_B_XOR;
  assign CLBLL_L_X2Y95_SLICE_X1Y95_CMUX = CLBLL_L_X2Y95_SLICE_X1Y95_C_XOR;
  assign CLBLL_L_X2Y95_SLICE_X1Y95_DMUX = CLBLL_L_X2Y95_SLICE_X1Y95_D_XOR;
  assign CLBLL_L_X2Y96_SLICE_X0Y96_COUT = CLBLL_L_X2Y96_SLICE_X0Y96_D_CY;
  assign CLBLL_L_X2Y96_SLICE_X0Y96_A = CLBLL_L_X2Y96_SLICE_X0Y96_AO6;
  assign CLBLL_L_X2Y96_SLICE_X0Y96_B = CLBLL_L_X2Y96_SLICE_X0Y96_BO6;
  assign CLBLL_L_X2Y96_SLICE_X0Y96_C = CLBLL_L_X2Y96_SLICE_X0Y96_CO6;
  assign CLBLL_L_X2Y96_SLICE_X0Y96_D = CLBLL_L_X2Y96_SLICE_X0Y96_DO6;
  assign CLBLL_L_X2Y96_SLICE_X0Y96_BMUX = CLBLL_L_X2Y96_SLICE_X0Y96_BO6;
  assign CLBLL_L_X2Y96_SLICE_X1Y96_COUT = CLBLL_L_X2Y96_SLICE_X1Y96_D_CY;
  assign CLBLL_L_X2Y96_SLICE_X1Y96_A = CLBLL_L_X2Y96_SLICE_X1Y96_AO6;
  assign CLBLL_L_X2Y96_SLICE_X1Y96_B = CLBLL_L_X2Y96_SLICE_X1Y96_BO6;
  assign CLBLL_L_X2Y96_SLICE_X1Y96_C = CLBLL_L_X2Y96_SLICE_X1Y96_CO6;
  assign CLBLL_L_X2Y96_SLICE_X1Y96_D = CLBLL_L_X2Y96_SLICE_X1Y96_DO6;
  assign CLBLL_L_X2Y96_SLICE_X1Y96_AMUX = CLBLL_L_X2Y96_SLICE_X1Y96_AO6;
  assign CLBLL_L_X2Y96_SLICE_X1Y96_DMUX = CLBLL_L_X2Y96_SLICE_X1Y96_DO6;
  assign CLBLL_L_X2Y97_SLICE_X0Y97_COUT = CLBLL_L_X2Y97_SLICE_X0Y97_D_CY;
  assign CLBLL_L_X2Y97_SLICE_X0Y97_A = CLBLL_L_X2Y97_SLICE_X0Y97_AO6;
  assign CLBLL_L_X2Y97_SLICE_X0Y97_B = CLBLL_L_X2Y97_SLICE_X0Y97_BO6;
  assign CLBLL_L_X2Y97_SLICE_X0Y97_C = CLBLL_L_X2Y97_SLICE_X0Y97_CO6;
  assign CLBLL_L_X2Y97_SLICE_X0Y97_D = CLBLL_L_X2Y97_SLICE_X0Y97_DO6;
  assign CLBLL_L_X2Y97_SLICE_X0Y97_AMUX = CLBLL_L_X2Y97_SLICE_X0Y97_AO5;
  assign CLBLL_L_X2Y97_SLICE_X0Y97_DMUX = CLBLL_L_X2Y97_SLICE_X0Y97_DO6;
  assign CLBLL_L_X2Y97_SLICE_X1Y97_COUT = CLBLL_L_X2Y97_SLICE_X1Y97_D_CY;
  assign CLBLL_L_X2Y97_SLICE_X1Y97_A = CLBLL_L_X2Y97_SLICE_X1Y97_AO6;
  assign CLBLL_L_X2Y97_SLICE_X1Y97_B = CLBLL_L_X2Y97_SLICE_X1Y97_BO6;
  assign CLBLL_L_X2Y97_SLICE_X1Y97_C = CLBLL_L_X2Y97_SLICE_X1Y97_CO6;
  assign CLBLL_L_X2Y97_SLICE_X1Y97_D = CLBLL_L_X2Y97_SLICE_X1Y97_DO6;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_COUT = CLBLL_L_X2Y98_SLICE_X0Y98_D_CY;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_A = CLBLL_L_X2Y98_SLICE_X0Y98_AO6;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_B = CLBLL_L_X2Y98_SLICE_X0Y98_BO6;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_C = CLBLL_L_X2Y98_SLICE_X0Y98_CO6;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_D = CLBLL_L_X2Y98_SLICE_X0Y98_DO6;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_COUT = CLBLL_L_X2Y98_SLICE_X1Y98_D_CY;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_A = CLBLL_L_X2Y98_SLICE_X1Y98_AO6;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_B = CLBLL_L_X2Y98_SLICE_X1Y98_BO6;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_C = CLBLL_L_X2Y98_SLICE_X1Y98_CO6;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_D = CLBLL_L_X2Y98_SLICE_X1Y98_DO6;
  assign CLBLL_L_X2Y99_SLICE_X0Y99_COUT = CLBLL_L_X2Y99_SLICE_X0Y99_D_CY;
  assign CLBLL_L_X2Y99_SLICE_X0Y99_A = CLBLL_L_X2Y99_SLICE_X0Y99_AO6;
  assign CLBLL_L_X2Y99_SLICE_X0Y99_B = CLBLL_L_X2Y99_SLICE_X0Y99_BO6;
  assign CLBLL_L_X2Y99_SLICE_X0Y99_C = CLBLL_L_X2Y99_SLICE_X0Y99_CO6;
  assign CLBLL_L_X2Y99_SLICE_X0Y99_D = CLBLL_L_X2Y99_SLICE_X0Y99_DO6;
  assign CLBLL_L_X2Y99_SLICE_X1Y99_COUT = CLBLL_L_X2Y99_SLICE_X1Y99_D_CY;
  assign CLBLL_L_X2Y99_SLICE_X1Y99_A = CLBLL_L_X2Y99_SLICE_X1Y99_AO6;
  assign CLBLL_L_X2Y99_SLICE_X1Y99_B = CLBLL_L_X2Y99_SLICE_X1Y99_BO6;
  assign CLBLL_L_X2Y99_SLICE_X1Y99_C = CLBLL_L_X2Y99_SLICE_X1Y99_CO6;
  assign CLBLL_L_X2Y99_SLICE_X1Y99_D = CLBLL_L_X2Y99_SLICE_X1Y99_DO6;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_COUT = CLBLL_L_X2Y102_SLICE_X0Y102_D_CY;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_A = CLBLL_L_X2Y102_SLICE_X0Y102_AO6;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_B = CLBLL_L_X2Y102_SLICE_X0Y102_BO6;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_C = CLBLL_L_X2Y102_SLICE_X0Y102_CO6;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_D = CLBLL_L_X2Y102_SLICE_X0Y102_DO6;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_COUT = CLBLL_L_X2Y102_SLICE_X1Y102_D_CY;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_A = CLBLL_L_X2Y102_SLICE_X1Y102_AO6;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_B = CLBLL_L_X2Y102_SLICE_X1Y102_BO6;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_C = CLBLL_L_X2Y102_SLICE_X1Y102_CO6;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_D = CLBLL_L_X2Y102_SLICE_X1Y102_DO6;
  assign CLBLL_L_X4Y90_SLICE_X4Y90_COUT = CLBLL_L_X4Y90_SLICE_X4Y90_D_CY;
  assign CLBLL_L_X4Y90_SLICE_X4Y90_A = CLBLL_L_X4Y90_SLICE_X4Y90_AO6;
  assign CLBLL_L_X4Y90_SLICE_X4Y90_B = CLBLL_L_X4Y90_SLICE_X4Y90_BO6;
  assign CLBLL_L_X4Y90_SLICE_X4Y90_C = CLBLL_L_X4Y90_SLICE_X4Y90_CO6;
  assign CLBLL_L_X4Y90_SLICE_X4Y90_D = CLBLL_L_X4Y90_SLICE_X4Y90_DO6;
  assign CLBLL_L_X4Y90_SLICE_X5Y90_COUT = CLBLL_L_X4Y90_SLICE_X5Y90_D_CY;
  assign CLBLL_L_X4Y90_SLICE_X5Y90_A = CLBLL_L_X4Y90_SLICE_X5Y90_AO6;
  assign CLBLL_L_X4Y90_SLICE_X5Y90_B = CLBLL_L_X4Y90_SLICE_X5Y90_BO6;
  assign CLBLL_L_X4Y90_SLICE_X5Y90_C = CLBLL_L_X4Y90_SLICE_X5Y90_CO6;
  assign CLBLL_L_X4Y90_SLICE_X5Y90_D = CLBLL_L_X4Y90_SLICE_X5Y90_DO6;
  assign CLBLL_L_X4Y91_SLICE_X4Y91_COUT = CLBLL_L_X4Y91_SLICE_X4Y91_D_CY;
  assign CLBLL_L_X4Y91_SLICE_X4Y91_A = CLBLL_L_X4Y91_SLICE_X4Y91_AO6;
  assign CLBLL_L_X4Y91_SLICE_X4Y91_B = CLBLL_L_X4Y91_SLICE_X4Y91_BO6;
  assign CLBLL_L_X4Y91_SLICE_X4Y91_C = CLBLL_L_X4Y91_SLICE_X4Y91_CO6;
  assign CLBLL_L_X4Y91_SLICE_X4Y91_D = CLBLL_L_X4Y91_SLICE_X4Y91_DO6;
  assign CLBLL_L_X4Y91_SLICE_X4Y91_AMUX = CLBLL_L_X4Y91_SLICE_X4Y91_AO5;
  assign CLBLL_L_X4Y91_SLICE_X5Y91_COUT = CLBLL_L_X4Y91_SLICE_X5Y91_D_CY;
  assign CLBLL_L_X4Y91_SLICE_X5Y91_A = CLBLL_L_X4Y91_SLICE_X5Y91_AO6;
  assign CLBLL_L_X4Y91_SLICE_X5Y91_B = CLBLL_L_X4Y91_SLICE_X5Y91_BO6;
  assign CLBLL_L_X4Y91_SLICE_X5Y91_C = CLBLL_L_X4Y91_SLICE_X5Y91_CO6;
  assign CLBLL_L_X4Y91_SLICE_X5Y91_D = CLBLL_L_X4Y91_SLICE_X5Y91_DO6;
  assign CLBLL_L_X4Y91_SLICE_X5Y91_AMUX = CLBLL_L_X4Y91_SLICE_X5Y91_F7AMUX_O;
  assign CLBLL_L_X4Y92_SLICE_X4Y92_COUT = CLBLL_L_X4Y92_SLICE_X4Y92_D_CY;
  assign CLBLL_L_X4Y92_SLICE_X4Y92_A = CLBLL_L_X4Y92_SLICE_X4Y92_AO6;
  assign CLBLL_L_X4Y92_SLICE_X4Y92_B = CLBLL_L_X4Y92_SLICE_X4Y92_BO6;
  assign CLBLL_L_X4Y92_SLICE_X4Y92_C = CLBLL_L_X4Y92_SLICE_X4Y92_CO6;
  assign CLBLL_L_X4Y92_SLICE_X4Y92_D = CLBLL_L_X4Y92_SLICE_X4Y92_DO6;
  assign CLBLL_L_X4Y92_SLICE_X4Y92_AMUX = CLBLL_L_X4Y92_SLICE_X4Y92_AO5;
  assign CLBLL_L_X4Y92_SLICE_X4Y92_BMUX = CLBLL_L_X4Y92_SLICE_X4Y92_B5Q;
  assign CLBLL_L_X4Y92_SLICE_X5Y92_COUT = CLBLL_L_X4Y92_SLICE_X5Y92_D_CY;
  assign CLBLL_L_X4Y92_SLICE_X5Y92_A = CLBLL_L_X4Y92_SLICE_X5Y92_AO6;
  assign CLBLL_L_X4Y92_SLICE_X5Y92_B = CLBLL_L_X4Y92_SLICE_X5Y92_BO6;
  assign CLBLL_L_X4Y92_SLICE_X5Y92_C = CLBLL_L_X4Y92_SLICE_X5Y92_CO6;
  assign CLBLL_L_X4Y92_SLICE_X5Y92_D = CLBLL_L_X4Y92_SLICE_X5Y92_DO6;
  assign CLBLL_L_X4Y92_SLICE_X5Y92_AMUX = CLBLL_L_X4Y92_SLICE_X5Y92_F7AMUX_O;
  assign CLBLL_L_X4Y93_SLICE_X4Y93_COUT = CLBLL_L_X4Y93_SLICE_X4Y93_D_CY;
  assign CLBLL_L_X4Y93_SLICE_X4Y93_A = CLBLL_L_X4Y93_SLICE_X4Y93_AO6;
  assign CLBLL_L_X4Y93_SLICE_X4Y93_B = CLBLL_L_X4Y93_SLICE_X4Y93_BO6;
  assign CLBLL_L_X4Y93_SLICE_X4Y93_C = CLBLL_L_X4Y93_SLICE_X4Y93_CO6;
  assign CLBLL_L_X4Y93_SLICE_X4Y93_D = CLBLL_L_X4Y93_SLICE_X4Y93_DO6;
  assign CLBLL_L_X4Y93_SLICE_X4Y93_AMUX = CLBLL_L_X4Y93_SLICE_X4Y93_F7AMUX_O;
  assign CLBLL_L_X4Y93_SLICE_X4Y93_CMUX = CLBLL_L_X4Y93_SLICE_X4Y93_CO5;
  assign CLBLL_L_X4Y93_SLICE_X5Y93_COUT = CLBLL_L_X4Y93_SLICE_X5Y93_D_CY;
  assign CLBLL_L_X4Y93_SLICE_X5Y93_A = CLBLL_L_X4Y93_SLICE_X5Y93_AO6;
  assign CLBLL_L_X4Y93_SLICE_X5Y93_B = CLBLL_L_X4Y93_SLICE_X5Y93_BO6;
  assign CLBLL_L_X4Y93_SLICE_X5Y93_C = CLBLL_L_X4Y93_SLICE_X5Y93_CO6;
  assign CLBLL_L_X4Y93_SLICE_X5Y93_D = CLBLL_L_X4Y93_SLICE_X5Y93_DO6;
  assign CLBLL_L_X4Y93_SLICE_X5Y93_AMUX = CLBLL_L_X4Y93_SLICE_X5Y93_F7AMUX_O;
  assign CLBLL_L_X4Y94_SLICE_X4Y94_COUT = CLBLL_L_X4Y94_SLICE_X4Y94_D_CY;
  assign CLBLL_L_X4Y94_SLICE_X4Y94_A = CLBLL_L_X4Y94_SLICE_X4Y94_AO6;
  assign CLBLL_L_X4Y94_SLICE_X4Y94_B = CLBLL_L_X4Y94_SLICE_X4Y94_BO6;
  assign CLBLL_L_X4Y94_SLICE_X4Y94_C = CLBLL_L_X4Y94_SLICE_X4Y94_CO6;
  assign CLBLL_L_X4Y94_SLICE_X4Y94_D = CLBLL_L_X4Y94_SLICE_X4Y94_DO6;
  assign CLBLL_L_X4Y94_SLICE_X4Y94_CMUX = CLBLL_L_X4Y94_SLICE_X4Y94_CO5;
  assign CLBLL_L_X4Y94_SLICE_X5Y94_COUT = CLBLL_L_X4Y94_SLICE_X5Y94_D_CY;
  assign CLBLL_L_X4Y94_SLICE_X5Y94_A = CLBLL_L_X4Y94_SLICE_X5Y94_AO6;
  assign CLBLL_L_X4Y94_SLICE_X5Y94_B = CLBLL_L_X4Y94_SLICE_X5Y94_BO6;
  assign CLBLL_L_X4Y94_SLICE_X5Y94_C = CLBLL_L_X4Y94_SLICE_X5Y94_CO6;
  assign CLBLL_L_X4Y94_SLICE_X5Y94_D = CLBLL_L_X4Y94_SLICE_X5Y94_DO6;
  assign CLBLL_L_X4Y94_SLICE_X5Y94_AMUX = CLBLL_L_X4Y94_SLICE_X5Y94_F7AMUX_O;
  assign CLBLL_L_X4Y95_SLICE_X4Y95_COUT = CLBLL_L_X4Y95_SLICE_X4Y95_D_CY;
  assign CLBLL_L_X4Y95_SLICE_X4Y95_A = CLBLL_L_X4Y95_SLICE_X4Y95_AO6;
  assign CLBLL_L_X4Y95_SLICE_X4Y95_B = CLBLL_L_X4Y95_SLICE_X4Y95_BO6;
  assign CLBLL_L_X4Y95_SLICE_X4Y95_C = CLBLL_L_X4Y95_SLICE_X4Y95_CO6;
  assign CLBLL_L_X4Y95_SLICE_X4Y95_D = CLBLL_L_X4Y95_SLICE_X4Y95_DO6;
  assign CLBLL_L_X4Y95_SLICE_X5Y95_COUT = CLBLL_L_X4Y95_SLICE_X5Y95_D_CY;
  assign CLBLL_L_X4Y95_SLICE_X5Y95_A = CLBLL_L_X4Y95_SLICE_X5Y95_AO6;
  assign CLBLL_L_X4Y95_SLICE_X5Y95_B = CLBLL_L_X4Y95_SLICE_X5Y95_BO6;
  assign CLBLL_L_X4Y95_SLICE_X5Y95_C = CLBLL_L_X4Y95_SLICE_X5Y95_CO6;
  assign CLBLL_L_X4Y95_SLICE_X5Y95_D = CLBLL_L_X4Y95_SLICE_X5Y95_DO6;
  assign CLBLL_L_X4Y95_SLICE_X5Y95_AMUX = CLBLL_L_X4Y95_SLICE_X5Y95_F7AMUX_O;
  assign CLBLL_L_X4Y96_SLICE_X4Y96_COUT = CLBLL_L_X4Y96_SLICE_X4Y96_D_CY;
  assign CLBLL_L_X4Y96_SLICE_X4Y96_A = CLBLL_L_X4Y96_SLICE_X4Y96_AO6;
  assign CLBLL_L_X4Y96_SLICE_X4Y96_B = CLBLL_L_X4Y96_SLICE_X4Y96_BO6;
  assign CLBLL_L_X4Y96_SLICE_X4Y96_C = CLBLL_L_X4Y96_SLICE_X4Y96_CO6;
  assign CLBLL_L_X4Y96_SLICE_X4Y96_D = CLBLL_L_X4Y96_SLICE_X4Y96_DO6;
  assign CLBLL_L_X4Y96_SLICE_X5Y96_COUT = CLBLL_L_X4Y96_SLICE_X5Y96_D_CY;
  assign CLBLL_L_X4Y96_SLICE_X5Y96_A = CLBLL_L_X4Y96_SLICE_X5Y96_AO6;
  assign CLBLL_L_X4Y96_SLICE_X5Y96_B = CLBLL_L_X4Y96_SLICE_X5Y96_BO6;
  assign CLBLL_L_X4Y96_SLICE_X5Y96_C = CLBLL_L_X4Y96_SLICE_X5Y96_CO6;
  assign CLBLL_L_X4Y96_SLICE_X5Y96_D = CLBLL_L_X4Y96_SLICE_X5Y96_DO6;
  assign CLBLL_L_X4Y97_SLICE_X4Y97_COUT = CLBLL_L_X4Y97_SLICE_X4Y97_D_CY;
  assign CLBLL_L_X4Y97_SLICE_X4Y97_A = CLBLL_L_X4Y97_SLICE_X4Y97_AO6;
  assign CLBLL_L_X4Y97_SLICE_X4Y97_B = CLBLL_L_X4Y97_SLICE_X4Y97_BO6;
  assign CLBLL_L_X4Y97_SLICE_X4Y97_C = CLBLL_L_X4Y97_SLICE_X4Y97_CO6;
  assign CLBLL_L_X4Y97_SLICE_X4Y97_D = CLBLL_L_X4Y97_SLICE_X4Y97_DO6;
  assign CLBLL_L_X4Y97_SLICE_X4Y97_AMUX = CLBLL_L_X4Y97_SLICE_X4Y97_AO5;
  assign CLBLL_L_X4Y97_SLICE_X5Y97_COUT = CLBLL_L_X4Y97_SLICE_X5Y97_D_CY;
  assign CLBLL_L_X4Y97_SLICE_X5Y97_A = CLBLL_L_X4Y97_SLICE_X5Y97_AO6;
  assign CLBLL_L_X4Y97_SLICE_X5Y97_B = CLBLL_L_X4Y97_SLICE_X5Y97_BO6;
  assign CLBLL_L_X4Y97_SLICE_X5Y97_C = CLBLL_L_X4Y97_SLICE_X5Y97_CO6;
  assign CLBLL_L_X4Y97_SLICE_X5Y97_D = CLBLL_L_X4Y97_SLICE_X5Y97_DO6;
  assign CLBLL_L_X4Y97_SLICE_X5Y97_AMUX = CLBLL_L_X4Y97_SLICE_X5Y97_AO5;
  assign CLBLL_L_X4Y98_SLICE_X4Y98_COUT = CLBLL_L_X4Y98_SLICE_X4Y98_D_CY;
  assign CLBLL_L_X4Y98_SLICE_X4Y98_A = CLBLL_L_X4Y98_SLICE_X4Y98_AO6;
  assign CLBLL_L_X4Y98_SLICE_X4Y98_B = CLBLL_L_X4Y98_SLICE_X4Y98_BO6;
  assign CLBLL_L_X4Y98_SLICE_X4Y98_C = CLBLL_L_X4Y98_SLICE_X4Y98_CO6;
  assign CLBLL_L_X4Y98_SLICE_X4Y98_D = CLBLL_L_X4Y98_SLICE_X4Y98_DO6;
  assign CLBLL_L_X4Y98_SLICE_X4Y98_AMUX = CLBLL_L_X4Y98_SLICE_X4Y98_AO6;
  assign CLBLL_L_X4Y98_SLICE_X5Y98_COUT = CLBLL_L_X4Y98_SLICE_X5Y98_D_CY;
  assign CLBLL_L_X4Y98_SLICE_X5Y98_A = CLBLL_L_X4Y98_SLICE_X5Y98_AO6;
  assign CLBLL_L_X4Y98_SLICE_X5Y98_B = CLBLL_L_X4Y98_SLICE_X5Y98_BO6;
  assign CLBLL_L_X4Y98_SLICE_X5Y98_C = CLBLL_L_X4Y98_SLICE_X5Y98_CO6;
  assign CLBLL_L_X4Y98_SLICE_X5Y98_D = CLBLL_L_X4Y98_SLICE_X5Y98_DO6;
  assign CLBLM_L_X8Y89_SLICE_X10Y89_COUT = CLBLM_L_X8Y89_SLICE_X10Y89_D_CY;
  assign CLBLM_L_X8Y89_SLICE_X10Y89_A = CLBLM_L_X8Y89_SLICE_X10Y89_AO6;
  assign CLBLM_L_X8Y89_SLICE_X10Y89_B = CLBLM_L_X8Y89_SLICE_X10Y89_BO6;
  assign CLBLM_L_X8Y89_SLICE_X10Y89_C = CLBLM_L_X8Y89_SLICE_X10Y89_CO6;
  assign CLBLM_L_X8Y89_SLICE_X10Y89_D = CLBLM_L_X8Y89_SLICE_X10Y89_DO6;
  assign CLBLM_L_X8Y89_SLICE_X10Y89_AMUX = CLBLM_L_X8Y89_SLICE_X10Y89_A5Q;
  assign CLBLM_L_X8Y89_SLICE_X11Y89_COUT = CLBLM_L_X8Y89_SLICE_X11Y89_D_CY;
  assign CLBLM_L_X8Y89_SLICE_X11Y89_A = CLBLM_L_X8Y89_SLICE_X11Y89_AO6;
  assign CLBLM_L_X8Y89_SLICE_X11Y89_B = CLBLM_L_X8Y89_SLICE_X11Y89_BO6;
  assign CLBLM_L_X8Y89_SLICE_X11Y89_C = CLBLM_L_X8Y89_SLICE_X11Y89_CO6;
  assign CLBLM_L_X8Y89_SLICE_X11Y89_D = CLBLM_L_X8Y89_SLICE_X11Y89_DO6;
  assign CLBLM_L_X8Y97_SLICE_X10Y97_A = CLBLM_L_X8Y97_SLICE_X10Y97_AO6;
  assign CLBLM_L_X8Y97_SLICE_X10Y97_B = CLBLM_L_X8Y97_SLICE_X10Y97_BO6;
  assign CLBLM_L_X8Y97_SLICE_X10Y97_C = CLBLM_L_X8Y97_SLICE_X10Y97_CO6;
  assign CLBLM_L_X8Y97_SLICE_X10Y97_D = CLBLM_L_X8Y97_SLICE_X10Y97_DO6;
  assign CLBLM_L_X8Y97_SLICE_X11Y97_COUT = CLBLM_L_X8Y97_SLICE_X11Y97_D_CY;
  assign CLBLM_L_X8Y97_SLICE_X11Y97_A = CLBLM_L_X8Y97_SLICE_X11Y97_AO6;
  assign CLBLM_L_X8Y97_SLICE_X11Y97_B = CLBLM_L_X8Y97_SLICE_X11Y97_BO6;
  assign CLBLM_L_X8Y97_SLICE_X11Y97_C = CLBLM_L_X8Y97_SLICE_X11Y97_CO6;
  assign CLBLM_L_X8Y97_SLICE_X11Y97_D = CLBLM_L_X8Y97_SLICE_X11Y97_DO6;
  assign CLBLM_L_X8Y98_SLICE_X10Y98_COUT = CLBLM_L_X8Y98_SLICE_X10Y98_D_CY;
  assign CLBLM_L_X8Y98_SLICE_X10Y98_A = CLBLM_L_X8Y98_SLICE_X10Y98_AO6;
  assign CLBLM_L_X8Y98_SLICE_X10Y98_B = CLBLM_L_X8Y98_SLICE_X10Y98_BO6;
  assign CLBLM_L_X8Y98_SLICE_X10Y98_C = CLBLM_L_X8Y98_SLICE_X10Y98_CO6;
  assign CLBLM_L_X8Y98_SLICE_X10Y98_D = CLBLM_L_X8Y98_SLICE_X10Y98_DO6;
  assign CLBLM_L_X8Y98_SLICE_X10Y98_AMUX = CLBLM_L_X8Y98_SLICE_X10Y98_AO5;
  assign CLBLM_L_X8Y98_SLICE_X11Y98_COUT = CLBLM_L_X8Y98_SLICE_X11Y98_D_CY;
  assign CLBLM_L_X8Y98_SLICE_X11Y98_A = CLBLM_L_X8Y98_SLICE_X11Y98_AO6;
  assign CLBLM_L_X8Y98_SLICE_X11Y98_B = CLBLM_L_X8Y98_SLICE_X11Y98_BO6;
  assign CLBLM_L_X8Y98_SLICE_X11Y98_C = CLBLM_L_X8Y98_SLICE_X11Y98_CO6;
  assign CLBLM_L_X8Y98_SLICE_X11Y98_D = CLBLM_L_X8Y98_SLICE_X11Y98_DO6;
  assign CLBLM_R_X3Y90_SLICE_X2Y90_COUT = CLBLM_R_X3Y90_SLICE_X2Y90_D_CY;
  assign CLBLM_R_X3Y90_SLICE_X2Y90_A = CLBLM_R_X3Y90_SLICE_X2Y90_AO6;
  assign CLBLM_R_X3Y90_SLICE_X2Y90_B = CLBLM_R_X3Y90_SLICE_X2Y90_BO6;
  assign CLBLM_R_X3Y90_SLICE_X2Y90_C = CLBLM_R_X3Y90_SLICE_X2Y90_CO6;
  assign CLBLM_R_X3Y90_SLICE_X2Y90_D = CLBLM_R_X3Y90_SLICE_X2Y90_DO6;
  assign CLBLM_R_X3Y90_SLICE_X3Y90_COUT = CLBLM_R_X3Y90_SLICE_X3Y90_D_CY;
  assign CLBLM_R_X3Y90_SLICE_X3Y90_A = CLBLM_R_X3Y90_SLICE_X3Y90_AO6;
  assign CLBLM_R_X3Y90_SLICE_X3Y90_B = CLBLM_R_X3Y90_SLICE_X3Y90_BO6;
  assign CLBLM_R_X3Y90_SLICE_X3Y90_C = CLBLM_R_X3Y90_SLICE_X3Y90_CO6;
  assign CLBLM_R_X3Y90_SLICE_X3Y90_D = CLBLM_R_X3Y90_SLICE_X3Y90_DO6;
  assign CLBLM_R_X3Y91_SLICE_X2Y91_COUT = CLBLM_R_X3Y91_SLICE_X2Y91_D_CY;
  assign CLBLM_R_X3Y91_SLICE_X2Y91_A = CLBLM_R_X3Y91_SLICE_X2Y91_AO6;
  assign CLBLM_R_X3Y91_SLICE_X2Y91_B = CLBLM_R_X3Y91_SLICE_X2Y91_BO6;
  assign CLBLM_R_X3Y91_SLICE_X2Y91_C = CLBLM_R_X3Y91_SLICE_X2Y91_CO6;
  assign CLBLM_R_X3Y91_SLICE_X2Y91_D = CLBLM_R_X3Y91_SLICE_X2Y91_DO6;
  assign CLBLM_R_X3Y91_SLICE_X2Y91_AMUX = CLBLM_R_X3Y91_SLICE_X2Y91_F7AMUX_O;
  assign CLBLM_R_X3Y91_SLICE_X2Y91_CMUX = CLBLM_R_X3Y91_SLICE_X2Y91_F7BMUX_O;
  assign CLBLM_R_X3Y91_SLICE_X3Y91_COUT = CLBLM_R_X3Y91_SLICE_X3Y91_D_CY;
  assign CLBLM_R_X3Y91_SLICE_X3Y91_A = CLBLM_R_X3Y91_SLICE_X3Y91_AO6;
  assign CLBLM_R_X3Y91_SLICE_X3Y91_B = CLBLM_R_X3Y91_SLICE_X3Y91_BO6;
  assign CLBLM_R_X3Y91_SLICE_X3Y91_C = CLBLM_R_X3Y91_SLICE_X3Y91_CO6;
  assign CLBLM_R_X3Y91_SLICE_X3Y91_D = CLBLM_R_X3Y91_SLICE_X3Y91_DO6;
  assign CLBLM_R_X3Y91_SLICE_X3Y91_AMUX = CLBLM_R_X3Y91_SLICE_X3Y91_F7AMUX_O;
  assign CLBLM_R_X3Y91_SLICE_X3Y91_CMUX = CLBLM_R_X3Y91_SLICE_X3Y91_F7BMUX_O;
  assign CLBLM_R_X3Y92_SLICE_X2Y92_COUT = CLBLM_R_X3Y92_SLICE_X2Y92_D_CY;
  assign CLBLM_R_X3Y92_SLICE_X2Y92_A = CLBLM_R_X3Y92_SLICE_X2Y92_AO6;
  assign CLBLM_R_X3Y92_SLICE_X2Y92_B = CLBLM_R_X3Y92_SLICE_X2Y92_BO6;
  assign CLBLM_R_X3Y92_SLICE_X2Y92_C = CLBLM_R_X3Y92_SLICE_X2Y92_CO6;
  assign CLBLM_R_X3Y92_SLICE_X2Y92_D = CLBLM_R_X3Y92_SLICE_X2Y92_DO6;
  assign CLBLM_R_X3Y92_SLICE_X2Y92_AMUX = CLBLM_R_X3Y92_SLICE_X2Y92_F7AMUX_O;
  assign CLBLM_R_X3Y92_SLICE_X2Y92_CMUX = CLBLM_R_X3Y92_SLICE_X2Y92_F7BMUX_O;
  assign CLBLM_R_X3Y92_SLICE_X3Y92_COUT = CLBLM_R_X3Y92_SLICE_X3Y92_D_CY;
  assign CLBLM_R_X3Y92_SLICE_X3Y92_A = CLBLM_R_X3Y92_SLICE_X3Y92_AO6;
  assign CLBLM_R_X3Y92_SLICE_X3Y92_B = CLBLM_R_X3Y92_SLICE_X3Y92_BO6;
  assign CLBLM_R_X3Y92_SLICE_X3Y92_C = CLBLM_R_X3Y92_SLICE_X3Y92_CO6;
  assign CLBLM_R_X3Y92_SLICE_X3Y92_D = CLBLM_R_X3Y92_SLICE_X3Y92_DO6;
  assign CLBLM_R_X3Y93_SLICE_X2Y93_COUT = CLBLM_R_X3Y93_SLICE_X2Y93_D_CY;
  assign CLBLM_R_X3Y93_SLICE_X2Y93_A = CLBLM_R_X3Y93_SLICE_X2Y93_AO6;
  assign CLBLM_R_X3Y93_SLICE_X2Y93_B = CLBLM_R_X3Y93_SLICE_X2Y93_BO6;
  assign CLBLM_R_X3Y93_SLICE_X2Y93_C = CLBLM_R_X3Y93_SLICE_X2Y93_CO6;
  assign CLBLM_R_X3Y93_SLICE_X2Y93_D = CLBLM_R_X3Y93_SLICE_X2Y93_DO6;
  assign CLBLM_R_X3Y93_SLICE_X2Y93_AMUX = CLBLM_R_X3Y93_SLICE_X2Y93_F7AMUX_O;
  assign CLBLM_R_X3Y93_SLICE_X2Y93_CMUX = CLBLM_R_X3Y93_SLICE_X2Y93_CO5;
  assign CLBLM_R_X3Y93_SLICE_X3Y93_COUT = CLBLM_R_X3Y93_SLICE_X3Y93_D_CY;
  assign CLBLM_R_X3Y93_SLICE_X3Y93_A = CLBLM_R_X3Y93_SLICE_X3Y93_AO6;
  assign CLBLM_R_X3Y93_SLICE_X3Y93_B = CLBLM_R_X3Y93_SLICE_X3Y93_BO6;
  assign CLBLM_R_X3Y93_SLICE_X3Y93_C = CLBLM_R_X3Y93_SLICE_X3Y93_CO6;
  assign CLBLM_R_X3Y93_SLICE_X3Y93_D = CLBLM_R_X3Y93_SLICE_X3Y93_DO6;
  assign CLBLM_R_X3Y93_SLICE_X3Y93_AMUX = CLBLM_R_X3Y93_SLICE_X3Y93_AO6;
  assign CLBLM_R_X3Y94_SLICE_X2Y94_COUT = CLBLM_R_X3Y94_SLICE_X2Y94_D_CY;
  assign CLBLM_R_X3Y94_SLICE_X2Y94_A = CLBLM_R_X3Y94_SLICE_X2Y94_AO6;
  assign CLBLM_R_X3Y94_SLICE_X2Y94_B = CLBLM_R_X3Y94_SLICE_X2Y94_BO6;
  assign CLBLM_R_X3Y94_SLICE_X2Y94_C = CLBLM_R_X3Y94_SLICE_X2Y94_CO6;
  assign CLBLM_R_X3Y94_SLICE_X2Y94_D = CLBLM_R_X3Y94_SLICE_X2Y94_DO6;
  assign CLBLM_R_X3Y94_SLICE_X2Y94_DMUX = CLBLM_R_X3Y94_SLICE_X2Y94_DO5;
  assign CLBLM_R_X3Y94_SLICE_X3Y94_COUT = CLBLM_R_X3Y94_SLICE_X3Y94_D_CY;
  assign CLBLM_R_X3Y94_SLICE_X3Y94_A = CLBLM_R_X3Y94_SLICE_X3Y94_AO6;
  assign CLBLM_R_X3Y94_SLICE_X3Y94_B = CLBLM_R_X3Y94_SLICE_X3Y94_BO6;
  assign CLBLM_R_X3Y94_SLICE_X3Y94_C = CLBLM_R_X3Y94_SLICE_X3Y94_CO6;
  assign CLBLM_R_X3Y94_SLICE_X3Y94_D = CLBLM_R_X3Y94_SLICE_X3Y94_DO6;
  assign CLBLM_R_X3Y94_SLICE_X3Y94_AMUX = CLBLM_R_X3Y94_SLICE_X3Y94_F7AMUX_O;
  assign CLBLM_R_X3Y94_SLICE_X3Y94_CMUX = CLBLM_R_X3Y94_SLICE_X3Y94_F7BMUX_O;
  assign CLBLM_R_X3Y95_SLICE_X2Y95_COUT = CLBLM_R_X3Y95_SLICE_X2Y95_D_CY;
  assign CLBLM_R_X3Y95_SLICE_X2Y95_A = CLBLM_R_X3Y95_SLICE_X2Y95_AO6;
  assign CLBLM_R_X3Y95_SLICE_X2Y95_B = CLBLM_R_X3Y95_SLICE_X2Y95_BO6;
  assign CLBLM_R_X3Y95_SLICE_X2Y95_C = CLBLM_R_X3Y95_SLICE_X2Y95_CO6;
  assign CLBLM_R_X3Y95_SLICE_X2Y95_D = CLBLM_R_X3Y95_SLICE_X2Y95_DO6;
  assign CLBLM_R_X3Y95_SLICE_X3Y95_COUT = CLBLM_R_X3Y95_SLICE_X3Y95_D_CY;
  assign CLBLM_R_X3Y95_SLICE_X3Y95_A = CLBLM_R_X3Y95_SLICE_X3Y95_AO6;
  assign CLBLM_R_X3Y95_SLICE_X3Y95_B = CLBLM_R_X3Y95_SLICE_X3Y95_BO6;
  assign CLBLM_R_X3Y95_SLICE_X3Y95_C = CLBLM_R_X3Y95_SLICE_X3Y95_CO6;
  assign CLBLM_R_X3Y95_SLICE_X3Y95_D = CLBLM_R_X3Y95_SLICE_X3Y95_DO6;
  assign CLBLM_R_X3Y96_SLICE_X2Y96_A = CLBLM_R_X3Y96_SLICE_X2Y96_AO6;
  assign CLBLM_R_X3Y96_SLICE_X2Y96_B = CLBLM_R_X3Y96_SLICE_X2Y96_BO6;
  assign CLBLM_R_X3Y96_SLICE_X2Y96_C = CLBLM_R_X3Y96_SLICE_X2Y96_CO6;
  assign CLBLM_R_X3Y96_SLICE_X2Y96_D = CLBLM_R_X3Y96_SLICE_X2Y96_DO6;
  assign CLBLM_R_X3Y96_SLICE_X3Y96_COUT = CLBLM_R_X3Y96_SLICE_X3Y96_D_CY;
  assign CLBLM_R_X3Y96_SLICE_X3Y96_A = CLBLM_R_X3Y96_SLICE_X3Y96_AO6;
  assign CLBLM_R_X3Y96_SLICE_X3Y96_B = CLBLM_R_X3Y96_SLICE_X3Y96_BO6;
  assign CLBLM_R_X3Y96_SLICE_X3Y96_C = CLBLM_R_X3Y96_SLICE_X3Y96_CO6;
  assign CLBLM_R_X3Y96_SLICE_X3Y96_D = CLBLM_R_X3Y96_SLICE_X3Y96_DO6;
  assign CLBLM_R_X3Y96_SLICE_X3Y96_AMUX = CLBLM_R_X3Y96_SLICE_X3Y96_AO5;
  assign CLBLM_R_X3Y96_SLICE_X3Y96_BMUX = CLBLM_R_X3Y96_SLICE_X3Y96_BO5;
  assign CLBLM_R_X3Y97_SLICE_X2Y97_A = CLBLM_R_X3Y97_SLICE_X2Y97_AO6;
  assign CLBLM_R_X3Y97_SLICE_X2Y97_B = CLBLM_R_X3Y97_SLICE_X2Y97_BO6;
  assign CLBLM_R_X3Y97_SLICE_X2Y97_C = CLBLM_R_X3Y97_SLICE_X2Y97_CO6;
  assign CLBLM_R_X3Y97_SLICE_X2Y97_D = CLBLM_R_X3Y97_SLICE_X2Y97_DO6;
  assign CLBLM_R_X3Y97_SLICE_X3Y97_COUT = CLBLM_R_X3Y97_SLICE_X3Y97_D_CY;
  assign CLBLM_R_X3Y97_SLICE_X3Y97_A = CLBLM_R_X3Y97_SLICE_X3Y97_AO6;
  assign CLBLM_R_X3Y97_SLICE_X3Y97_B = CLBLM_R_X3Y97_SLICE_X3Y97_BO6;
  assign CLBLM_R_X3Y97_SLICE_X3Y97_C = CLBLM_R_X3Y97_SLICE_X3Y97_CO6;
  assign CLBLM_R_X3Y97_SLICE_X3Y97_D = CLBLM_R_X3Y97_SLICE_X3Y97_DO6;
  assign CLBLM_R_X3Y97_SLICE_X3Y97_DMUX = CLBLM_R_X3Y97_SLICE_X3Y97_DO6;
  assign CLBLM_R_X3Y98_SLICE_X2Y98_COUT = CLBLM_R_X3Y98_SLICE_X2Y98_D_CY;
  assign CLBLM_R_X3Y98_SLICE_X2Y98_A = CLBLM_R_X3Y98_SLICE_X2Y98_AO6;
  assign CLBLM_R_X3Y98_SLICE_X2Y98_B = CLBLM_R_X3Y98_SLICE_X2Y98_BO6;
  assign CLBLM_R_X3Y98_SLICE_X2Y98_C = CLBLM_R_X3Y98_SLICE_X2Y98_CO6;
  assign CLBLM_R_X3Y98_SLICE_X2Y98_D = CLBLM_R_X3Y98_SLICE_X2Y98_DO6;
  assign CLBLM_R_X3Y98_SLICE_X2Y98_DMUX = CLBLM_R_X3Y98_SLICE_X2Y98_DO6;
  assign CLBLM_R_X3Y98_SLICE_X3Y98_COUT = CLBLM_R_X3Y98_SLICE_X3Y98_D_CY;
  assign CLBLM_R_X3Y98_SLICE_X3Y98_A = CLBLM_R_X3Y98_SLICE_X3Y98_AO6;
  assign CLBLM_R_X3Y98_SLICE_X3Y98_B = CLBLM_R_X3Y98_SLICE_X3Y98_BO6;
  assign CLBLM_R_X3Y98_SLICE_X3Y98_C = CLBLM_R_X3Y98_SLICE_X3Y98_CO6;
  assign CLBLM_R_X3Y98_SLICE_X3Y98_D = CLBLM_R_X3Y98_SLICE_X3Y98_DO6;
  assign CLBLM_R_X3Y98_SLICE_X3Y98_AMUX = CLBLM_R_X3Y98_SLICE_X3Y98_AO6;
  assign CLBLM_R_X3Y98_SLICE_X3Y98_DMUX = CLBLM_R_X3Y98_SLICE_X3Y98_DO6;
  assign CLBLM_R_X3Y99_SLICE_X2Y99_COUT = CLBLM_R_X3Y99_SLICE_X2Y99_D_CY;
  assign CLBLM_R_X3Y99_SLICE_X2Y99_A = CLBLM_R_X3Y99_SLICE_X2Y99_AO6;
  assign CLBLM_R_X3Y99_SLICE_X2Y99_B = CLBLM_R_X3Y99_SLICE_X2Y99_BO6;
  assign CLBLM_R_X3Y99_SLICE_X2Y99_C = CLBLM_R_X3Y99_SLICE_X2Y99_CO6;
  assign CLBLM_R_X3Y99_SLICE_X2Y99_D = CLBLM_R_X3Y99_SLICE_X2Y99_DO6;
  assign CLBLM_R_X3Y99_SLICE_X2Y99_AMUX = CLBLM_R_X3Y99_SLICE_X2Y99_AO6;
  assign CLBLM_R_X3Y99_SLICE_X3Y99_COUT = CLBLM_R_X3Y99_SLICE_X3Y99_D_CY;
  assign CLBLM_R_X3Y99_SLICE_X3Y99_A = CLBLM_R_X3Y99_SLICE_X3Y99_AO6;
  assign CLBLM_R_X3Y99_SLICE_X3Y99_B = CLBLM_R_X3Y99_SLICE_X3Y99_BO6;
  assign CLBLM_R_X3Y99_SLICE_X3Y99_C = CLBLM_R_X3Y99_SLICE_X3Y99_CO6;
  assign CLBLM_R_X3Y99_SLICE_X3Y99_D = CLBLM_R_X3Y99_SLICE_X3Y99_DO6;
  assign CLBLM_R_X5Y90_SLICE_X6Y90_COUT = CLBLM_R_X5Y90_SLICE_X6Y90_D_CY;
  assign CLBLM_R_X5Y90_SLICE_X6Y90_A = CLBLM_R_X5Y90_SLICE_X6Y90_AO6;
  assign CLBLM_R_X5Y90_SLICE_X6Y90_B = CLBLM_R_X5Y90_SLICE_X6Y90_BO6;
  assign CLBLM_R_X5Y90_SLICE_X6Y90_C = CLBLM_R_X5Y90_SLICE_X6Y90_CO6;
  assign CLBLM_R_X5Y90_SLICE_X6Y90_D = CLBLM_R_X5Y90_SLICE_X6Y90_DO6;
  assign CLBLM_R_X5Y90_SLICE_X6Y90_AMUX = CLBLM_R_X5Y90_SLICE_X6Y90_A5Q;
  assign CLBLM_R_X5Y90_SLICE_X6Y90_BMUX = CLBLM_R_X5Y90_SLICE_X6Y90_B5Q;
  assign CLBLM_R_X5Y90_SLICE_X7Y90_COUT = CLBLM_R_X5Y90_SLICE_X7Y90_D_CY;
  assign CLBLM_R_X5Y90_SLICE_X7Y90_A = CLBLM_R_X5Y90_SLICE_X7Y90_AO6;
  assign CLBLM_R_X5Y90_SLICE_X7Y90_B = CLBLM_R_X5Y90_SLICE_X7Y90_BO6;
  assign CLBLM_R_X5Y90_SLICE_X7Y90_C = CLBLM_R_X5Y90_SLICE_X7Y90_CO6;
  assign CLBLM_R_X5Y90_SLICE_X7Y90_D = CLBLM_R_X5Y90_SLICE_X7Y90_DO6;
  assign CLBLM_R_X5Y90_SLICE_X7Y90_AMUX = CLBLM_R_X5Y90_SLICE_X7Y90_A5Q;
  assign CLBLM_R_X5Y90_SLICE_X7Y90_BMUX = CLBLM_R_X5Y90_SLICE_X7Y90_B5Q;
  assign CLBLM_R_X5Y90_SLICE_X7Y90_CMUX = CLBLM_R_X5Y90_SLICE_X7Y90_C5Q;
  assign CLBLM_R_X5Y91_SLICE_X6Y91_COUT = CLBLM_R_X5Y91_SLICE_X6Y91_D_CY;
  assign CLBLM_R_X5Y91_SLICE_X6Y91_A = CLBLM_R_X5Y91_SLICE_X6Y91_AO6;
  assign CLBLM_R_X5Y91_SLICE_X6Y91_B = CLBLM_R_X5Y91_SLICE_X6Y91_BO6;
  assign CLBLM_R_X5Y91_SLICE_X6Y91_C = CLBLM_R_X5Y91_SLICE_X6Y91_CO6;
  assign CLBLM_R_X5Y91_SLICE_X6Y91_D = CLBLM_R_X5Y91_SLICE_X6Y91_DO6;
  assign CLBLM_R_X5Y91_SLICE_X7Y91_COUT = CLBLM_R_X5Y91_SLICE_X7Y91_D_CY;
  assign CLBLM_R_X5Y91_SLICE_X7Y91_A = CLBLM_R_X5Y91_SLICE_X7Y91_AO6;
  assign CLBLM_R_X5Y91_SLICE_X7Y91_B = CLBLM_R_X5Y91_SLICE_X7Y91_BO6;
  assign CLBLM_R_X5Y91_SLICE_X7Y91_C = CLBLM_R_X5Y91_SLICE_X7Y91_CO6;
  assign CLBLM_R_X5Y91_SLICE_X7Y91_D = CLBLM_R_X5Y91_SLICE_X7Y91_DO6;
  assign CLBLM_R_X5Y92_SLICE_X6Y92_COUT = CLBLM_R_X5Y92_SLICE_X6Y92_D_CY;
  assign CLBLM_R_X5Y92_SLICE_X6Y92_A = CLBLM_R_X5Y92_SLICE_X6Y92_AO6;
  assign CLBLM_R_X5Y92_SLICE_X6Y92_B = CLBLM_R_X5Y92_SLICE_X6Y92_BO6;
  assign CLBLM_R_X5Y92_SLICE_X6Y92_C = CLBLM_R_X5Y92_SLICE_X6Y92_CO6;
  assign CLBLM_R_X5Y92_SLICE_X6Y92_D = CLBLM_R_X5Y92_SLICE_X6Y92_DO6;
  assign CLBLM_R_X5Y92_SLICE_X7Y92_COUT = CLBLM_R_X5Y92_SLICE_X7Y92_D_CY;
  assign CLBLM_R_X5Y92_SLICE_X7Y92_A = CLBLM_R_X5Y92_SLICE_X7Y92_AO6;
  assign CLBLM_R_X5Y92_SLICE_X7Y92_B = CLBLM_R_X5Y92_SLICE_X7Y92_BO6;
  assign CLBLM_R_X5Y92_SLICE_X7Y92_C = CLBLM_R_X5Y92_SLICE_X7Y92_CO6;
  assign CLBLM_R_X5Y92_SLICE_X7Y92_D = CLBLM_R_X5Y92_SLICE_X7Y92_DO6;
  assign CLBLM_R_X5Y93_SLICE_X6Y93_COUT = CLBLM_R_X5Y93_SLICE_X6Y93_D_CY;
  assign CLBLM_R_X5Y93_SLICE_X6Y93_A = CLBLM_R_X5Y93_SLICE_X6Y93_AO6;
  assign CLBLM_R_X5Y93_SLICE_X6Y93_B = CLBLM_R_X5Y93_SLICE_X6Y93_BO6;
  assign CLBLM_R_X5Y93_SLICE_X6Y93_C = CLBLM_R_X5Y93_SLICE_X6Y93_CO6;
  assign CLBLM_R_X5Y93_SLICE_X6Y93_D = CLBLM_R_X5Y93_SLICE_X6Y93_DO6;
  assign CLBLM_R_X5Y93_SLICE_X6Y93_AMUX = CLBLM_R_X5Y93_SLICE_X6Y93_F7AMUX_O;
  assign CLBLM_R_X5Y93_SLICE_X7Y93_COUT = CLBLM_R_X5Y93_SLICE_X7Y93_D_CY;
  assign CLBLM_R_X5Y93_SLICE_X7Y93_A = CLBLM_R_X5Y93_SLICE_X7Y93_AO6;
  assign CLBLM_R_X5Y93_SLICE_X7Y93_B = CLBLM_R_X5Y93_SLICE_X7Y93_BO6;
  assign CLBLM_R_X5Y93_SLICE_X7Y93_C = CLBLM_R_X5Y93_SLICE_X7Y93_CO6;
  assign CLBLM_R_X5Y93_SLICE_X7Y93_D = CLBLM_R_X5Y93_SLICE_X7Y93_DO6;
  assign CLBLM_R_X5Y94_SLICE_X6Y94_COUT = CLBLM_R_X5Y94_SLICE_X6Y94_D_CY;
  assign CLBLM_R_X5Y94_SLICE_X6Y94_A = CLBLM_R_X5Y94_SLICE_X6Y94_AO6;
  assign CLBLM_R_X5Y94_SLICE_X6Y94_B = CLBLM_R_X5Y94_SLICE_X6Y94_BO6;
  assign CLBLM_R_X5Y94_SLICE_X6Y94_C = CLBLM_R_X5Y94_SLICE_X6Y94_CO6;
  assign CLBLM_R_X5Y94_SLICE_X6Y94_D = CLBLM_R_X5Y94_SLICE_X6Y94_DO6;
  assign CLBLM_R_X5Y94_SLICE_X6Y94_AMUX = CLBLM_R_X5Y94_SLICE_X6Y94_AO6;
  assign CLBLM_R_X5Y94_SLICE_X7Y94_COUT = CLBLM_R_X5Y94_SLICE_X7Y94_D_CY;
  assign CLBLM_R_X5Y94_SLICE_X7Y94_A = CLBLM_R_X5Y94_SLICE_X7Y94_AO6;
  assign CLBLM_R_X5Y94_SLICE_X7Y94_B = CLBLM_R_X5Y94_SLICE_X7Y94_BO6;
  assign CLBLM_R_X5Y94_SLICE_X7Y94_C = CLBLM_R_X5Y94_SLICE_X7Y94_CO6;
  assign CLBLM_R_X5Y94_SLICE_X7Y94_D = CLBLM_R_X5Y94_SLICE_X7Y94_DO6;
  assign CLBLM_R_X5Y94_SLICE_X7Y94_AMUX = CLBLM_R_X5Y94_SLICE_X7Y94_AO5;
  assign CLBLM_R_X5Y95_SLICE_X6Y95_COUT = CLBLM_R_X5Y95_SLICE_X6Y95_D_CY;
  assign CLBLM_R_X5Y95_SLICE_X6Y95_A = CLBLM_R_X5Y95_SLICE_X6Y95_AO6;
  assign CLBLM_R_X5Y95_SLICE_X6Y95_B = CLBLM_R_X5Y95_SLICE_X6Y95_BO6;
  assign CLBLM_R_X5Y95_SLICE_X6Y95_C = CLBLM_R_X5Y95_SLICE_X6Y95_CO6;
  assign CLBLM_R_X5Y95_SLICE_X6Y95_D = CLBLM_R_X5Y95_SLICE_X6Y95_DO6;
  assign CLBLM_R_X5Y95_SLICE_X6Y95_BMUX = CLBLM_R_X5Y95_SLICE_X6Y95_BO5;
  assign CLBLM_R_X5Y95_SLICE_X7Y95_COUT = CLBLM_R_X5Y95_SLICE_X7Y95_D_CY;
  assign CLBLM_R_X5Y95_SLICE_X7Y95_A = CLBLM_R_X5Y95_SLICE_X7Y95_AO6;
  assign CLBLM_R_X5Y95_SLICE_X7Y95_B = CLBLM_R_X5Y95_SLICE_X7Y95_BO6;
  assign CLBLM_R_X5Y95_SLICE_X7Y95_C = CLBLM_R_X5Y95_SLICE_X7Y95_CO6;
  assign CLBLM_R_X5Y95_SLICE_X7Y95_D = CLBLM_R_X5Y95_SLICE_X7Y95_DO6;
  assign CLBLM_R_X5Y96_SLICE_X6Y96_COUT = CLBLM_R_X5Y96_SLICE_X6Y96_D_CY;
  assign CLBLM_R_X5Y96_SLICE_X6Y96_A = CLBLM_R_X5Y96_SLICE_X6Y96_AO6;
  assign CLBLM_R_X5Y96_SLICE_X6Y96_B = CLBLM_R_X5Y96_SLICE_X6Y96_BO6;
  assign CLBLM_R_X5Y96_SLICE_X6Y96_C = CLBLM_R_X5Y96_SLICE_X6Y96_CO6;
  assign CLBLM_R_X5Y96_SLICE_X6Y96_D = CLBLM_R_X5Y96_SLICE_X6Y96_DO6;
  assign CLBLM_R_X5Y96_SLICE_X7Y96_COUT = CLBLM_R_X5Y96_SLICE_X7Y96_D_CY;
  assign CLBLM_R_X5Y96_SLICE_X7Y96_A = CLBLM_R_X5Y96_SLICE_X7Y96_AO6;
  assign CLBLM_R_X5Y96_SLICE_X7Y96_B = CLBLM_R_X5Y96_SLICE_X7Y96_BO6;
  assign CLBLM_R_X5Y96_SLICE_X7Y96_C = CLBLM_R_X5Y96_SLICE_X7Y96_CO6;
  assign CLBLM_R_X5Y96_SLICE_X7Y96_D = CLBLM_R_X5Y96_SLICE_X7Y96_DO6;
  assign CLBLM_R_X5Y96_SLICE_X7Y96_CMUX = CLBLM_R_X5Y96_SLICE_X7Y96_CO5;
  assign CLBLM_R_X5Y97_SLICE_X6Y97_A = CLBLM_R_X5Y97_SLICE_X6Y97_AO6;
  assign CLBLM_R_X5Y97_SLICE_X6Y97_B = CLBLM_R_X5Y97_SLICE_X6Y97_BO6;
  assign CLBLM_R_X5Y97_SLICE_X6Y97_C = CLBLM_R_X5Y97_SLICE_X6Y97_CO6;
  assign CLBLM_R_X5Y97_SLICE_X6Y97_D = CLBLM_R_X5Y97_SLICE_X6Y97_DO6;
  assign CLBLM_R_X5Y97_SLICE_X6Y97_AMUX = CLBLM_R_X5Y97_SLICE_X6Y97_AO6;
  assign CLBLM_R_X5Y97_SLICE_X6Y97_BMUX = CLBLM_R_X5Y97_SLICE_X6Y97_BO6;
  assign CLBLM_R_X5Y97_SLICE_X7Y97_COUT = CLBLM_R_X5Y97_SLICE_X7Y97_D_CY;
  assign CLBLM_R_X5Y97_SLICE_X7Y97_A = CLBLM_R_X5Y97_SLICE_X7Y97_AO6;
  assign CLBLM_R_X5Y97_SLICE_X7Y97_B = CLBLM_R_X5Y97_SLICE_X7Y97_BO6;
  assign CLBLM_R_X5Y97_SLICE_X7Y97_C = CLBLM_R_X5Y97_SLICE_X7Y97_CO6;
  assign CLBLM_R_X5Y97_SLICE_X7Y97_D = CLBLM_R_X5Y97_SLICE_X7Y97_DO6;
  assign CLBLM_R_X5Y97_SLICE_X7Y97_AMUX = CLBLM_R_X5Y97_SLICE_X7Y97_AO5;
  assign CLBLM_R_X5Y98_SLICE_X6Y98_A = CLBLM_R_X5Y98_SLICE_X6Y98_AO6;
  assign CLBLM_R_X5Y98_SLICE_X6Y98_B = CLBLM_R_X5Y98_SLICE_X6Y98_BO6;
  assign CLBLM_R_X5Y98_SLICE_X6Y98_C = CLBLM_R_X5Y98_SLICE_X6Y98_CO6;
  assign CLBLM_R_X5Y98_SLICE_X6Y98_D = CLBLM_R_X5Y98_SLICE_X6Y98_DO6;
  assign CLBLM_R_X5Y98_SLICE_X6Y98_CMUX = CLBLM_R_X5Y98_SLICE_X6Y98_CO6;
  assign CLBLM_R_X5Y98_SLICE_X6Y98_DMUX = CLBLM_R_X5Y98_SLICE_X6Y98_DO6;
  assign CLBLM_R_X5Y98_SLICE_X7Y98_COUT = CLBLM_R_X5Y98_SLICE_X7Y98_D_CY;
  assign CLBLM_R_X5Y98_SLICE_X7Y98_A = CLBLM_R_X5Y98_SLICE_X7Y98_AO6;
  assign CLBLM_R_X5Y98_SLICE_X7Y98_B = CLBLM_R_X5Y98_SLICE_X7Y98_BO6;
  assign CLBLM_R_X5Y98_SLICE_X7Y98_C = CLBLM_R_X5Y98_SLICE_X7Y98_CO6;
  assign CLBLM_R_X5Y98_SLICE_X7Y98_D = CLBLM_R_X5Y98_SLICE_X7Y98_DO6;
  assign CLBLM_R_X5Y98_SLICE_X7Y98_AMUX = CLBLM_R_X5Y98_SLICE_X7Y98_AO5;
  assign CLBLM_R_X5Y99_SLICE_X6Y99_COUT = CLBLM_R_X5Y99_SLICE_X6Y99_D_CY;
  assign CLBLM_R_X5Y99_SLICE_X6Y99_A = CLBLM_R_X5Y99_SLICE_X6Y99_AO6;
  assign CLBLM_R_X5Y99_SLICE_X6Y99_B = CLBLM_R_X5Y99_SLICE_X6Y99_BO6;
  assign CLBLM_R_X5Y99_SLICE_X6Y99_C = CLBLM_R_X5Y99_SLICE_X6Y99_CO6;
  assign CLBLM_R_X5Y99_SLICE_X6Y99_D = CLBLM_R_X5Y99_SLICE_X6Y99_DO6;
  assign CLBLM_R_X5Y99_SLICE_X7Y99_COUT = CLBLM_R_X5Y99_SLICE_X7Y99_D_CY;
  assign CLBLM_R_X5Y99_SLICE_X7Y99_A = CLBLM_R_X5Y99_SLICE_X7Y99_AO6;
  assign CLBLM_R_X5Y99_SLICE_X7Y99_B = CLBLM_R_X5Y99_SLICE_X7Y99_BO6;
  assign CLBLM_R_X5Y99_SLICE_X7Y99_C = CLBLM_R_X5Y99_SLICE_X7Y99_CO6;
  assign CLBLM_R_X5Y99_SLICE_X7Y99_D = CLBLM_R_X5Y99_SLICE_X7Y99_DO6;
  assign CLBLM_R_X5Y99_SLICE_X7Y99_BMUX = CLBLM_R_X5Y99_SLICE_X7Y99_BO5;
  assign CLBLM_R_X7Y87_SLICE_X8Y87_COUT = CLBLM_R_X7Y87_SLICE_X8Y87_D_CY;
  assign CLBLM_R_X7Y87_SLICE_X8Y87_A = CLBLM_R_X7Y87_SLICE_X8Y87_AO6;
  assign CLBLM_R_X7Y87_SLICE_X8Y87_B = CLBLM_R_X7Y87_SLICE_X8Y87_BO6;
  assign CLBLM_R_X7Y87_SLICE_X8Y87_C = CLBLM_R_X7Y87_SLICE_X8Y87_CO6;
  assign CLBLM_R_X7Y87_SLICE_X8Y87_D = CLBLM_R_X7Y87_SLICE_X8Y87_DO6;
  assign CLBLM_R_X7Y87_SLICE_X9Y87_COUT = CLBLM_R_X7Y87_SLICE_X9Y87_D_CY;
  assign CLBLM_R_X7Y87_SLICE_X9Y87_A = CLBLM_R_X7Y87_SLICE_X9Y87_AO6;
  assign CLBLM_R_X7Y87_SLICE_X9Y87_B = CLBLM_R_X7Y87_SLICE_X9Y87_BO6;
  assign CLBLM_R_X7Y87_SLICE_X9Y87_C = CLBLM_R_X7Y87_SLICE_X9Y87_CO6;
  assign CLBLM_R_X7Y87_SLICE_X9Y87_D = CLBLM_R_X7Y87_SLICE_X9Y87_DO6;
  assign CLBLM_R_X7Y88_SLICE_X8Y88_COUT = CLBLM_R_X7Y88_SLICE_X8Y88_D_CY;
  assign CLBLM_R_X7Y88_SLICE_X8Y88_A = CLBLM_R_X7Y88_SLICE_X8Y88_AO6;
  assign CLBLM_R_X7Y88_SLICE_X8Y88_B = CLBLM_R_X7Y88_SLICE_X8Y88_BO6;
  assign CLBLM_R_X7Y88_SLICE_X8Y88_C = CLBLM_R_X7Y88_SLICE_X8Y88_CO6;
  assign CLBLM_R_X7Y88_SLICE_X8Y88_D = CLBLM_R_X7Y88_SLICE_X8Y88_DO6;
  assign CLBLM_R_X7Y88_SLICE_X9Y88_COUT = CLBLM_R_X7Y88_SLICE_X9Y88_D_CY;
  assign CLBLM_R_X7Y88_SLICE_X9Y88_A = CLBLM_R_X7Y88_SLICE_X9Y88_AO6;
  assign CLBLM_R_X7Y88_SLICE_X9Y88_B = CLBLM_R_X7Y88_SLICE_X9Y88_BO6;
  assign CLBLM_R_X7Y88_SLICE_X9Y88_C = CLBLM_R_X7Y88_SLICE_X9Y88_CO6;
  assign CLBLM_R_X7Y88_SLICE_X9Y88_D = CLBLM_R_X7Y88_SLICE_X9Y88_DO6;
  assign CLBLM_R_X7Y89_SLICE_X8Y89_COUT = CLBLM_R_X7Y89_SLICE_X8Y89_D_CY;
  assign CLBLM_R_X7Y89_SLICE_X8Y89_A = CLBLM_R_X7Y89_SLICE_X8Y89_AO6;
  assign CLBLM_R_X7Y89_SLICE_X8Y89_B = CLBLM_R_X7Y89_SLICE_X8Y89_BO6;
  assign CLBLM_R_X7Y89_SLICE_X8Y89_C = CLBLM_R_X7Y89_SLICE_X8Y89_CO6;
  assign CLBLM_R_X7Y89_SLICE_X8Y89_D = CLBLM_R_X7Y89_SLICE_X8Y89_DO6;
  assign CLBLM_R_X7Y89_SLICE_X8Y89_BMUX = CLBLM_R_X7Y89_SLICE_X8Y89_B5Q;
  assign CLBLM_R_X7Y89_SLICE_X9Y89_COUT = CLBLM_R_X7Y89_SLICE_X9Y89_D_CY;
  assign CLBLM_R_X7Y89_SLICE_X9Y89_A = CLBLM_R_X7Y89_SLICE_X9Y89_AO6;
  assign CLBLM_R_X7Y89_SLICE_X9Y89_B = CLBLM_R_X7Y89_SLICE_X9Y89_BO6;
  assign CLBLM_R_X7Y89_SLICE_X9Y89_C = CLBLM_R_X7Y89_SLICE_X9Y89_CO6;
  assign CLBLM_R_X7Y89_SLICE_X9Y89_D = CLBLM_R_X7Y89_SLICE_X9Y89_DO6;
  assign CLBLM_R_X7Y89_SLICE_X9Y89_AMUX = CLBLM_R_X7Y89_SLICE_X9Y89_AO5;
  assign CLBLM_R_X7Y90_SLICE_X8Y90_COUT = CLBLM_R_X7Y90_SLICE_X8Y90_D_CY;
  assign CLBLM_R_X7Y90_SLICE_X8Y90_A = CLBLM_R_X7Y90_SLICE_X8Y90_AO6;
  assign CLBLM_R_X7Y90_SLICE_X8Y90_B = CLBLM_R_X7Y90_SLICE_X8Y90_BO6;
  assign CLBLM_R_X7Y90_SLICE_X8Y90_C = CLBLM_R_X7Y90_SLICE_X8Y90_CO6;
  assign CLBLM_R_X7Y90_SLICE_X8Y90_D = CLBLM_R_X7Y90_SLICE_X8Y90_DO6;
  assign CLBLM_R_X7Y90_SLICE_X9Y90_COUT = CLBLM_R_X7Y90_SLICE_X9Y90_D_CY;
  assign CLBLM_R_X7Y90_SLICE_X9Y90_A = CLBLM_R_X7Y90_SLICE_X9Y90_AO6;
  assign CLBLM_R_X7Y90_SLICE_X9Y90_B = CLBLM_R_X7Y90_SLICE_X9Y90_BO6;
  assign CLBLM_R_X7Y90_SLICE_X9Y90_C = CLBLM_R_X7Y90_SLICE_X9Y90_CO6;
  assign CLBLM_R_X7Y90_SLICE_X9Y90_D = CLBLM_R_X7Y90_SLICE_X9Y90_DO6;
  assign CLBLM_R_X7Y90_SLICE_X9Y90_AMUX = CLBLM_R_X7Y90_SLICE_X9Y90_A5Q;
  assign CLBLM_R_X7Y91_SLICE_X8Y91_COUT = CLBLM_R_X7Y91_SLICE_X8Y91_D_CY;
  assign CLBLM_R_X7Y91_SLICE_X8Y91_A = CLBLM_R_X7Y91_SLICE_X8Y91_AO6;
  assign CLBLM_R_X7Y91_SLICE_X8Y91_B = CLBLM_R_X7Y91_SLICE_X8Y91_BO6;
  assign CLBLM_R_X7Y91_SLICE_X8Y91_C = CLBLM_R_X7Y91_SLICE_X8Y91_CO6;
  assign CLBLM_R_X7Y91_SLICE_X8Y91_D = CLBLM_R_X7Y91_SLICE_X8Y91_DO6;
  assign CLBLM_R_X7Y91_SLICE_X9Y91_COUT = CLBLM_R_X7Y91_SLICE_X9Y91_D_CY;
  assign CLBLM_R_X7Y91_SLICE_X9Y91_A = CLBLM_R_X7Y91_SLICE_X9Y91_AO6;
  assign CLBLM_R_X7Y91_SLICE_X9Y91_B = CLBLM_R_X7Y91_SLICE_X9Y91_BO6;
  assign CLBLM_R_X7Y91_SLICE_X9Y91_C = CLBLM_R_X7Y91_SLICE_X9Y91_CO6;
  assign CLBLM_R_X7Y91_SLICE_X9Y91_D = CLBLM_R_X7Y91_SLICE_X9Y91_DO6;
  assign CLBLM_R_X7Y93_SLICE_X8Y93_COUT = CLBLM_R_X7Y93_SLICE_X8Y93_D_CY;
  assign CLBLM_R_X7Y93_SLICE_X8Y93_A = CLBLM_R_X7Y93_SLICE_X8Y93_AO6;
  assign CLBLM_R_X7Y93_SLICE_X8Y93_B = CLBLM_R_X7Y93_SLICE_X8Y93_BO6;
  assign CLBLM_R_X7Y93_SLICE_X8Y93_C = CLBLM_R_X7Y93_SLICE_X8Y93_CO6;
  assign CLBLM_R_X7Y93_SLICE_X8Y93_D = CLBLM_R_X7Y93_SLICE_X8Y93_DO6;
  assign CLBLM_R_X7Y93_SLICE_X9Y93_COUT = CLBLM_R_X7Y93_SLICE_X9Y93_D_CY;
  assign CLBLM_R_X7Y93_SLICE_X9Y93_A = CLBLM_R_X7Y93_SLICE_X9Y93_AO6;
  assign CLBLM_R_X7Y93_SLICE_X9Y93_B = CLBLM_R_X7Y93_SLICE_X9Y93_BO6;
  assign CLBLM_R_X7Y93_SLICE_X9Y93_C = CLBLM_R_X7Y93_SLICE_X9Y93_CO6;
  assign CLBLM_R_X7Y93_SLICE_X9Y93_D = CLBLM_R_X7Y93_SLICE_X9Y93_DO6;
  assign CLBLM_R_X7Y94_SLICE_X8Y94_COUT = CLBLM_R_X7Y94_SLICE_X8Y94_D_CY;
  assign CLBLM_R_X7Y94_SLICE_X8Y94_A = CLBLM_R_X7Y94_SLICE_X8Y94_AO6;
  assign CLBLM_R_X7Y94_SLICE_X8Y94_B = CLBLM_R_X7Y94_SLICE_X8Y94_BO6;
  assign CLBLM_R_X7Y94_SLICE_X8Y94_C = CLBLM_R_X7Y94_SLICE_X8Y94_CO6;
  assign CLBLM_R_X7Y94_SLICE_X8Y94_D = CLBLM_R_X7Y94_SLICE_X8Y94_DO6;
  assign CLBLM_R_X7Y94_SLICE_X9Y94_COUT = CLBLM_R_X7Y94_SLICE_X9Y94_D_CY;
  assign CLBLM_R_X7Y94_SLICE_X9Y94_A = CLBLM_R_X7Y94_SLICE_X9Y94_AO6;
  assign CLBLM_R_X7Y94_SLICE_X9Y94_B = CLBLM_R_X7Y94_SLICE_X9Y94_BO6;
  assign CLBLM_R_X7Y94_SLICE_X9Y94_C = CLBLM_R_X7Y94_SLICE_X9Y94_CO6;
  assign CLBLM_R_X7Y94_SLICE_X9Y94_D = CLBLM_R_X7Y94_SLICE_X9Y94_DO6;
  assign CLBLM_R_X7Y96_SLICE_X8Y96_COUT = CLBLM_R_X7Y96_SLICE_X8Y96_D_CY;
  assign CLBLM_R_X7Y96_SLICE_X8Y96_A = CLBLM_R_X7Y96_SLICE_X8Y96_AO6;
  assign CLBLM_R_X7Y96_SLICE_X8Y96_B = CLBLM_R_X7Y96_SLICE_X8Y96_BO6;
  assign CLBLM_R_X7Y96_SLICE_X8Y96_C = CLBLM_R_X7Y96_SLICE_X8Y96_CO6;
  assign CLBLM_R_X7Y96_SLICE_X8Y96_D = CLBLM_R_X7Y96_SLICE_X8Y96_DO6;
  assign CLBLM_R_X7Y96_SLICE_X8Y96_BMUX = CLBLM_R_X7Y96_SLICE_X8Y96_BO5;
  assign CLBLM_R_X7Y96_SLICE_X8Y96_CMUX = CLBLM_R_X7Y96_SLICE_X8Y96_CO6;
  assign CLBLM_R_X7Y96_SLICE_X9Y96_COUT = CLBLM_R_X7Y96_SLICE_X9Y96_D_CY;
  assign CLBLM_R_X7Y96_SLICE_X9Y96_A = CLBLM_R_X7Y96_SLICE_X9Y96_AO6;
  assign CLBLM_R_X7Y96_SLICE_X9Y96_B = CLBLM_R_X7Y96_SLICE_X9Y96_BO6;
  assign CLBLM_R_X7Y96_SLICE_X9Y96_C = CLBLM_R_X7Y96_SLICE_X9Y96_CO6;
  assign CLBLM_R_X7Y96_SLICE_X9Y96_D = CLBLM_R_X7Y96_SLICE_X9Y96_DO6;
  assign CLBLM_R_X7Y97_SLICE_X8Y97_COUT = CLBLM_R_X7Y97_SLICE_X8Y97_D_CY;
  assign CLBLM_R_X7Y97_SLICE_X8Y97_A = CLBLM_R_X7Y97_SLICE_X8Y97_AO6;
  assign CLBLM_R_X7Y97_SLICE_X8Y97_B = CLBLM_R_X7Y97_SLICE_X8Y97_BO6;
  assign CLBLM_R_X7Y97_SLICE_X8Y97_C = CLBLM_R_X7Y97_SLICE_X8Y97_CO6;
  assign CLBLM_R_X7Y97_SLICE_X8Y97_D = CLBLM_R_X7Y97_SLICE_X8Y97_DO6;
  assign CLBLM_R_X7Y97_SLICE_X8Y97_BMUX = CLBLM_R_X7Y97_SLICE_X8Y97_BO5;
  assign CLBLM_R_X7Y97_SLICE_X8Y97_DMUX = CLBLM_R_X7Y97_SLICE_X8Y97_DO6;
  assign CLBLM_R_X7Y97_SLICE_X9Y97_COUT = CLBLM_R_X7Y97_SLICE_X9Y97_D_CY;
  assign CLBLM_R_X7Y97_SLICE_X9Y97_A = CLBLM_R_X7Y97_SLICE_X9Y97_AO6;
  assign CLBLM_R_X7Y97_SLICE_X9Y97_B = CLBLM_R_X7Y97_SLICE_X9Y97_BO6;
  assign CLBLM_R_X7Y97_SLICE_X9Y97_C = CLBLM_R_X7Y97_SLICE_X9Y97_CO6;
  assign CLBLM_R_X7Y97_SLICE_X9Y97_D = CLBLM_R_X7Y97_SLICE_X9Y97_DO6;
  assign CLBLM_R_X7Y97_SLICE_X9Y97_AMUX = CLBLM_R_X7Y97_SLICE_X9Y97_A5Q;
  assign CLBLM_R_X7Y97_SLICE_X9Y97_BMUX = CLBLM_R_X7Y97_SLICE_X9Y97_B5Q;
  assign CLBLM_R_X7Y97_SLICE_X9Y97_CMUX = CLBLM_R_X7Y97_SLICE_X9Y97_CO6;
  assign CLBLM_R_X7Y98_SLICE_X8Y98_COUT = CLBLM_R_X7Y98_SLICE_X8Y98_D_CY;
  assign CLBLM_R_X7Y98_SLICE_X8Y98_A = CLBLM_R_X7Y98_SLICE_X8Y98_AO6;
  assign CLBLM_R_X7Y98_SLICE_X8Y98_B = CLBLM_R_X7Y98_SLICE_X8Y98_BO6;
  assign CLBLM_R_X7Y98_SLICE_X8Y98_C = CLBLM_R_X7Y98_SLICE_X8Y98_CO6;
  assign CLBLM_R_X7Y98_SLICE_X8Y98_D = CLBLM_R_X7Y98_SLICE_X8Y98_DO6;
  assign CLBLM_R_X7Y98_SLICE_X8Y98_AMUX = CLBLM_R_X7Y98_SLICE_X8Y98_F7AMUX_O;
  assign CLBLM_R_X7Y98_SLICE_X9Y98_COUT = CLBLM_R_X7Y98_SLICE_X9Y98_D_CY;
  assign CLBLM_R_X7Y98_SLICE_X9Y98_A = CLBLM_R_X7Y98_SLICE_X9Y98_AO6;
  assign CLBLM_R_X7Y98_SLICE_X9Y98_B = CLBLM_R_X7Y98_SLICE_X9Y98_BO6;
  assign CLBLM_R_X7Y98_SLICE_X9Y98_C = CLBLM_R_X7Y98_SLICE_X9Y98_CO6;
  assign CLBLM_R_X7Y98_SLICE_X9Y98_D = CLBLM_R_X7Y98_SLICE_X9Y98_DO6;
  assign CLBLM_R_X7Y99_SLICE_X8Y99_COUT = CLBLM_R_X7Y99_SLICE_X8Y99_D_CY;
  assign CLBLM_R_X7Y99_SLICE_X8Y99_A = CLBLM_R_X7Y99_SLICE_X8Y99_AO6;
  assign CLBLM_R_X7Y99_SLICE_X8Y99_B = CLBLM_R_X7Y99_SLICE_X8Y99_BO6;
  assign CLBLM_R_X7Y99_SLICE_X8Y99_C = CLBLM_R_X7Y99_SLICE_X8Y99_CO6;
  assign CLBLM_R_X7Y99_SLICE_X8Y99_D = CLBLM_R_X7Y99_SLICE_X8Y99_DO6;
  assign CLBLM_R_X7Y99_SLICE_X9Y99_COUT = CLBLM_R_X7Y99_SLICE_X9Y99_D_CY;
  assign CLBLM_R_X7Y99_SLICE_X9Y99_A = CLBLM_R_X7Y99_SLICE_X9Y99_AO6;
  assign CLBLM_R_X7Y99_SLICE_X9Y99_B = CLBLM_R_X7Y99_SLICE_X9Y99_BO6;
  assign CLBLM_R_X7Y99_SLICE_X9Y99_C = CLBLM_R_X7Y99_SLICE_X9Y99_CO6;
  assign CLBLM_R_X7Y99_SLICE_X9Y99_D = CLBLM_R_X7Y99_SLICE_X9Y99_DO6;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_OQ = CLBLL_L_X4Y90_SLICE_X5Y90_AQ;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_TQ = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_OQ = CLBLM_R_X7Y91_SLICE_X8Y91_CO6;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_OQ = CLBLL_L_X2Y102_SLICE_X0Y102_AQ;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_OQ = CLBLM_R_X7Y91_SLICE_X8Y91_DO6;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_TQ = 1'b1;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_O = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_O = LIOB33_X0Y105_IOB_X0Y105_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_O = LIOB33_X0Y109_IOB_X0Y109_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y128_O = LIOB33_X0Y127_IOB_X0Y128_I;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ = CLBLM_R_X7Y91_SLICE_X8Y91_BO6;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O = LIOB33_X0Y107_IOB_X0Y107_I;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ENARDENL = CLBLM_R_X5Y93_SLICE_X7Y93_CQ;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ENARDENU = CLBLM_R_X5Y93_SLICE_X7Y93_CQ;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ENBWRENL = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ENBWRENU = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_REGCEAREGCEL = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_REGCEAREGCEU = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_REGCEBL = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_REGCEBU = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_REGCLKARDRCLKL = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_REGCLKARDRCLKU = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_REGCLKBL = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_REGCLKBU = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_RSTRAMARSTRAMLRST = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_RSTRAMARSTRAMU = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_RSTRAMBL = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_RSTRAMBU = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_RSTREGARSTREGL = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_RSTREGARSTREGU = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_RSTREGBL = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_RSTREGBU = 1'b1;
  assign CLBLM_R_X7Y87_SLICE_X9Y87_A1 = 1'b1;
  assign CLBLM_R_X7Y87_SLICE_X9Y87_A2 = 1'b1;
  assign CLBLM_R_X7Y87_SLICE_X9Y87_A3 = 1'b1;
  assign CLBLM_R_X7Y87_SLICE_X9Y87_A4 = 1'b1;
  assign CLBLM_R_X7Y87_SLICE_X9Y87_A5 = 1'b1;
  assign CLBLM_R_X7Y87_SLICE_X9Y87_A6 = 1'b1;
  assign CLBLM_R_X7Y87_SLICE_X9Y87_B1 = 1'b1;
  assign CLBLM_R_X7Y87_SLICE_X9Y87_B2 = 1'b1;
  assign CLBLM_R_X7Y87_SLICE_X9Y87_B3 = 1'b1;
  assign CLBLM_R_X7Y87_SLICE_X9Y87_B4 = 1'b1;
  assign CLBLM_R_X7Y87_SLICE_X9Y87_B5 = 1'b1;
  assign CLBLM_R_X7Y87_SLICE_X9Y87_B6 = 1'b1;
  assign CLBLM_R_X7Y87_SLICE_X9Y87_C1 = 1'b1;
  assign CLBLM_R_X7Y87_SLICE_X9Y87_C2 = 1'b1;
  assign CLBLM_R_X7Y87_SLICE_X9Y87_C3 = 1'b1;
  assign CLBLM_R_X7Y87_SLICE_X9Y87_C4 = 1'b1;
  assign CLBLM_R_X7Y87_SLICE_X9Y87_C5 = 1'b1;
  assign CLBLM_R_X7Y87_SLICE_X9Y87_C6 = 1'b1;
  assign CLBLM_R_X7Y87_SLICE_X9Y87_D1 = 1'b1;
  assign CLBLM_R_X7Y87_SLICE_X9Y87_D2 = 1'b1;
  assign CLBLM_R_X7Y87_SLICE_X9Y87_D3 = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_WEAL0 = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_WEAL1 = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_WEAL2 = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_WEAL3 = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_WEAU0 = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_WEAU1 = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_WEAU2 = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_WEAU3 = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_WEBWEL0 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_WEBWEL1 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_WEBWEL2 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_WEBWEL3 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_WEBWEL4 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_WEBWEL5 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_WEBWEL6 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_WEBWEL7 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_WEBWEU0 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_WEBWEU1 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_WEBWEU2 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_WEBWEU3 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_WEBWEU4 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_WEBWEU5 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_WEBWEU6 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_WEBWEU7 = 1'b0;
  assign CLBLM_R_X3Y93_SLICE_X3Y93_B6 = CLBLM_R_X5Y94_SLICE_X7Y94_DO6;
  assign CLBLM_R_X3Y93_SLICE_X3Y93_BX = CLBLM_R_X3Y94_SLICE_X2Y94_DO5;
  assign CLBLM_R_X3Y93_SLICE_X3Y93_C1 = CLBLL_L_X2Y93_SLICE_X0Y93_CO6;
  assign CLBLM_R_X3Y93_SLICE_X3Y93_C2 = 1'b1;
  assign CLBLM_R_X3Y93_SLICE_X3Y93_C3 = CLBLL_L_X4Y94_SLICE_X5Y94_DO6;
  assign CLBLM_R_X3Y93_SLICE_X3Y93_C4 = CLBLM_R_X5Y94_SLICE_X7Y94_DO6;
  assign CLBLM_R_X3Y93_SLICE_X3Y93_C5 = 1'b1;
  assign CLBLM_R_X3Y93_SLICE_X3Y93_C6 = CLBLM_R_X5Y94_SLICE_X6Y94_BO6;
  assign CLBLM_R_X3Y93_SLICE_X3Y93_CE = CLBLM_R_X3Y93_SLICE_X3Y93_BO6;
  assign CLBLM_R_X3Y93_SLICE_X3Y93_CX = CLBLL_L_X4Y93_SLICE_X4Y93_CO6;
  assign CLBLM_R_X3Y93_SLICE_X3Y93_D1 = 1'b1;
  assign CLBLM_R_X3Y93_SLICE_X3Y93_D2 = 1'b1;
  assign CLBLM_R_X3Y93_SLICE_X3Y93_D3 = 1'b1;
  assign CLBLM_R_X3Y93_SLICE_X3Y93_D4 = 1'b1;
  assign CLBLM_R_X3Y93_SLICE_X3Y93_D5 = 1'b1;
  assign CLBLM_R_X3Y93_SLICE_X3Y93_D6 = 1'b1;
  assign CLBLM_R_X7Y87_SLICE_X8Y87_C1 = 1'b1;
  assign CLBLM_R_X7Y87_SLICE_X8Y87_C2 = 1'b1;
  assign CLBLM_R_X3Y93_SLICE_X3Y93_DX = CLBLL_L_X4Y94_SLICE_X4Y94_CO6;
  assign CLBLM_R_X7Y87_SLICE_X8Y87_C4 = 1'b1;
  assign CLBLM_R_X7Y87_SLICE_X8Y87_C5 = 1'b1;
  assign CLBLM_R_X7Y87_SLICE_X8Y87_C6 = 1'b1;
  assign CLBLM_R_X7Y87_SLICE_X8Y87_CLK = CLBLM_R_X7Y88_SLICE_X8Y88_AQ;
  assign CLBLM_R_X3Y93_SLICE_X2Y93_A1 = CLBLL_L_X2Y93_SLICE_X0Y93_BQ;
  assign CLBLM_R_X3Y93_SLICE_X2Y93_A2 = CLBLM_R_X3Y93_SLICE_X2Y93_BQ;
  assign CLBLM_R_X3Y93_SLICE_X2Y93_A3 = CLBLM_R_X3Y92_SLICE_X2Y92_BQ;
  assign CLBLM_R_X3Y93_SLICE_X2Y93_A4 = CLBLL_L_X4Y91_SLICE_X4Y91_AO6;
  assign CLBLM_R_X3Y93_SLICE_X2Y93_A5 = CLBLL_L_X2Y93_SLICE_X1Y93_BQ;
  assign CLBLM_R_X3Y93_SLICE_X2Y93_A6 = CLBLM_R_X3Y96_SLICE_X3Y96_AO6;
  assign CLBLM_R_X7Y87_SLICE_X8Y87_D1 = 1'b1;
  assign CLBLM_R_X7Y87_SLICE_X8Y87_D2 = 1'b1;
  assign CLBLM_R_X3Y93_SLICE_X2Y93_AX = CLBLL_L_X4Y95_SLICE_X5Y95_DO6;
  assign CLBLM_R_X7Y87_SLICE_X8Y87_D3 = 1'b1;
  assign CLBLM_R_X3Y93_SLICE_X2Y93_B1 = CLBLL_L_X2Y91_SLICE_X1Y91_AQ;
  assign CLBLM_R_X3Y93_SLICE_X2Y93_B2 = CLBLL_L_X4Y91_SLICE_X4Y91_AO6;
  assign CLBLM_R_X3Y93_SLICE_X2Y93_B3 = CLBLL_L_X2Y92_SLICE_X1Y92_AQ;
  assign CLBLM_R_X3Y93_SLICE_X2Y93_B4 = CLBLM_R_X3Y96_SLICE_X3Y96_AO6;
  assign CLBLM_R_X3Y93_SLICE_X2Y93_B5 = CLBLL_L_X2Y94_SLICE_X1Y94_BQ;
  assign CLBLM_R_X3Y93_SLICE_X2Y93_B6 = CLBLM_R_X3Y94_SLICE_X2Y94_AQ;
  assign CLBLM_R_X7Y87_SLICE_X8Y87_SR = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y93_SLICE_X2Y93_BX = CLBLM_R_X3Y94_SLICE_X2Y94_DO6;
  assign CLBLM_R_X3Y93_SLICE_X2Y93_C1 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X3Y93_SLICE_X2Y93_C2 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X3Y93_SLICE_X2Y93_C3 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X3Y93_SLICE_X2Y93_C4 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X3Y93_SLICE_X2Y93_C5 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLM_R_X3Y93_SLICE_X2Y93_C6 = 1'b1;
  assign CLBLM_R_X3Y93_SLICE_X2Y93_CE = CLBLM_R_X3Y93_SLICE_X3Y93_BO6;
  assign CLBLM_R_X3Y93_SLICE_X2Y93_CX = CLBLL_L_X4Y94_SLICE_X4Y94_CO5;
  assign CLBLM_R_X3Y93_SLICE_X2Y93_D1 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO15;
  assign CLBLM_R_X3Y93_SLICE_X2Y93_D2 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO10;
  assign CLBLM_R_X3Y93_SLICE_X2Y93_D3 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO12;
  assign CLBLM_R_X3Y93_SLICE_X2Y93_D4 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO13;
  assign CLBLM_R_X3Y93_SLICE_X2Y93_D5 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO14;
  assign CLBLM_R_X3Y93_SLICE_X2Y93_D6 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO11;
  assign LIOI3_X0Y127_ILOGIC_X0Y128_D = LIOB33_X0Y127_IOB_X0Y128_I;
  assign CLBLM_R_X7Y88_SLICE_X9Y88_A1 = 1'b1;
  assign CLBLM_R_X7Y88_SLICE_X9Y88_A2 = 1'b1;
  assign CLBLM_R_X7Y88_SLICE_X9Y88_A3 = 1'b1;
  assign CLBLM_R_X7Y88_SLICE_X9Y88_A4 = 1'b1;
  assign CLBLM_R_X7Y88_SLICE_X9Y88_A5 = 1'b1;
  assign CLBLM_R_X7Y88_SLICE_X9Y88_A6 = 1'b1;
  assign CLBLM_R_X7Y88_SLICE_X9Y88_B1 = 1'b1;
  assign CLBLM_R_X7Y88_SLICE_X9Y88_B2 = 1'b1;
  assign CLBLM_R_X7Y88_SLICE_X9Y88_B3 = 1'b1;
  assign CLBLM_R_X7Y88_SLICE_X9Y88_B4 = 1'b1;
  assign CLBLM_R_X7Y88_SLICE_X9Y88_B5 = 1'b1;
  assign CLBLM_R_X7Y88_SLICE_X9Y88_B6 = 1'b1;
  assign CLBLM_R_X7Y88_SLICE_X9Y88_C1 = 1'b1;
  assign CLBLM_R_X7Y88_SLICE_X9Y88_C2 = 1'b1;
  assign CLBLM_R_X7Y88_SLICE_X9Y88_C3 = 1'b1;
  assign CLBLM_R_X7Y88_SLICE_X9Y88_C4 = 1'b1;
  assign CLBLM_R_X7Y88_SLICE_X9Y88_C5 = 1'b1;
  assign CLBLM_R_X7Y88_SLICE_X9Y88_C6 = 1'b1;
  assign CLBLM_R_X7Y93_SLICE_X8Y93_D3 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO15;
  assign CLBLM_R_X7Y88_SLICE_X9Y88_D1 = 1'b1;
  assign CLBLM_R_X7Y88_SLICE_X9Y88_D2 = 1'b1;
  assign CLBLM_R_X7Y88_SLICE_X9Y88_D3 = 1'b1;
  assign CLBLM_R_X3Y94_SLICE_X3Y94_A1 = CLBLM_R_X5Y93_SLICE_X6Y93_F7AMUX_O;
  assign CLBLM_R_X3Y94_SLICE_X3Y94_A2 = CLBLM_R_X3Y94_SLICE_X3Y94_BQ;
  assign CLBLM_R_X3Y94_SLICE_X3Y94_A3 = CLBLL_L_X4Y91_SLICE_X5Y91_F7AMUX_O;
  assign CLBLM_R_X3Y94_SLICE_X3Y94_A4 = CLBLM_R_X3Y93_SLICE_X3Y93_BQ;
  assign CLBLM_R_X3Y94_SLICE_X3Y94_A5 = CLBLM_R_X3Y92_SLICE_X3Y92_AQ;
  assign CLBLM_R_X3Y94_SLICE_X3Y94_A6 = CLBLL_L_X2Y93_SLICE_X0Y93_CQ;
  assign CLBLM_R_X7Y88_SLICE_X9Y88_D4 = 1'b1;
  assign CLBLM_R_X7Y88_SLICE_X9Y88_D5 = 1'b1;
  assign CLBLM_R_X3Y94_SLICE_X3Y94_AX = CLBLL_L_X2Y93_SLICE_X0Y93_F7AMUX_O;
  assign CLBLM_R_X7Y88_SLICE_X9Y88_D6 = 1'b1;
  assign CLBLM_R_X3Y94_SLICE_X3Y94_B1 = CLBLM_R_X5Y93_SLICE_X6Y93_F7AMUX_O;
  assign CLBLM_R_X3Y94_SLICE_X3Y94_B2 = CLBLL_L_X2Y94_SLICE_X1Y94_CQ;
  assign CLBLM_R_X3Y94_SLICE_X3Y94_B3 = CLBLL_L_X4Y91_SLICE_X5Y91_F7AMUX_O;
  assign CLBLM_R_X3Y94_SLICE_X3Y94_B4 = CLBLM_R_X3Y94_SLICE_X2Y94_BQ;
  assign CLBLM_R_X3Y94_SLICE_X3Y94_B5 = CLBLL_L_X4Y93_SLICE_X4Y93_BQ;
  assign CLBLM_R_X3Y94_SLICE_X3Y94_B6 = CLBLL_L_X4Y92_SLICE_X4Y92_BQ;
  assign CLBLM_R_X7Y88_SLICE_X8Y88_A1 = 1'b1;
  assign CLBLM_R_X7Y88_SLICE_X8Y88_A2 = 1'b1;
  assign CLBLM_R_X3Y94_SLICE_X3Y94_BX = CLBLM_R_X3Y94_SLICE_X2Y94_DO5;
  assign CLBLM_R_X7Y88_SLICE_X8Y88_A3 = CLBLM_R_X7Y88_SLICE_X8Y88_AQ;
  assign CLBLM_R_X3Y94_SLICE_X3Y94_C1 = CLBLM_R_X3Y96_SLICE_X3Y96_AO6;
  assign CLBLM_R_X3Y94_SLICE_X3Y94_C2 = CLBLL_L_X2Y93_SLICE_X0Y93_CQ;
  assign CLBLM_R_X3Y94_SLICE_X3Y94_C3 = CLBLM_R_X3Y94_SLICE_X3Y94_BQ;
  assign CLBLM_R_X3Y94_SLICE_X3Y94_C4 = CLBLL_L_X4Y91_SLICE_X4Y91_AO6;
  assign CLBLM_R_X3Y94_SLICE_X3Y94_C5 = CLBLM_R_X3Y92_SLICE_X3Y92_AQ;
  assign CLBLM_R_X3Y94_SLICE_X3Y94_C6 = CLBLM_R_X3Y93_SLICE_X3Y93_BQ;
  assign CLBLM_R_X3Y94_SLICE_X3Y94_CE = CLBLM_R_X3Y93_SLICE_X3Y93_CO6;
  assign CLBLM_R_X7Y88_SLICE_X8Y88_B1 = CLBLM_R_X7Y90_SLICE_X8Y90_DO6;
  assign CLBLM_R_X7Y88_SLICE_X8Y88_B2 = CLBLM_R_X7Y87_SLICE_X8Y87_BQ;
  assign CLBLM_R_X7Y88_SLICE_X8Y88_B3 = CLBLM_R_X7Y87_SLICE_X8Y87_AQ;
  assign CLBLM_R_X7Y88_SLICE_X8Y88_B4 = 1'b1;
  assign CLBLM_R_X3Y94_SLICE_X3Y94_CX = CLBLL_L_X4Y95_SLICE_X5Y95_DO6;
  assign CLBLM_R_X7Y88_SLICE_X8Y88_B5 = CLBLM_R_X7Y91_SLICE_X9Y91_AQ;
  assign CLBLM_R_X3Y94_SLICE_X3Y94_D1 = CLBLL_L_X4Y93_SLICE_X4Y93_BQ;
  assign CLBLM_R_X3Y94_SLICE_X3Y94_D2 = CLBLL_L_X4Y92_SLICE_X4Y92_BQ;
  assign CLBLM_R_X3Y94_SLICE_X3Y94_D3 = CLBLM_R_X3Y96_SLICE_X3Y96_AO6;
  assign CLBLM_R_X3Y94_SLICE_X3Y94_D4 = CLBLL_L_X2Y94_SLICE_X1Y94_CQ;
  assign CLBLM_R_X3Y94_SLICE_X3Y94_D5 = CLBLL_L_X4Y91_SLICE_X4Y91_AO6;
  assign CLBLM_R_X3Y94_SLICE_X3Y94_D6 = CLBLM_R_X3Y94_SLICE_X2Y94_BQ;
  assign CLBLM_R_X7Y88_SLICE_X8Y88_C1 = 1'b1;
  assign CLBLM_R_X7Y88_SLICE_X8Y88_C2 = 1'b1;
  assign CLBLM_R_X7Y88_SLICE_X8Y88_C4 = 1'b1;
  assign CLBLM_R_X7Y88_SLICE_X8Y88_C5 = 1'b1;
  assign CLBLM_R_X7Y88_SLICE_X8Y88_C6 = 1'b1;
  assign CLBLM_R_X3Y94_SLICE_X2Y94_A1 = CLBLM_R_X3Y98_SLICE_X2Y98_BO6;
  assign CLBLM_R_X3Y94_SLICE_X2Y94_A2 = CLBLM_R_X5Y94_SLICE_X6Y94_BO6;
  assign CLBLM_R_X3Y94_SLICE_X2Y94_A3 = CLBLM_R_X3Y93_SLICE_X2Y93_CO6;
  assign CLBLM_R_X3Y94_SLICE_X2Y94_A4 = CLBLM_R_X5Y94_SLICE_X7Y94_DO6;
  assign CLBLM_R_X3Y94_SLICE_X2Y94_A5 = CLBLL_L_X2Y97_SLICE_X1Y97_AO6;
  assign CLBLM_R_X3Y94_SLICE_X2Y94_A6 = CLBLL_L_X4Y94_SLICE_X5Y94_DO6;
  assign CLBLM_R_X7Y88_SLICE_X8Y88_D1 = 1'b1;
  assign CLBLM_R_X7Y88_SLICE_X8Y88_D2 = 1'b1;
  assign CLBLM_R_X7Y88_SLICE_X8Y88_D3 = 1'b1;
  assign CLBLM_R_X3Y94_SLICE_X2Y94_B1 = CLBLM_R_X3Y99_SLICE_X2Y99_DO6;
  assign CLBLM_R_X3Y94_SLICE_X2Y94_B2 = CLBLL_L_X4Y94_SLICE_X5Y94_DO6;
  assign CLBLM_R_X3Y94_SLICE_X2Y94_B3 = CLBLM_R_X3Y93_SLICE_X2Y93_CO6;
  assign CLBLM_R_X3Y94_SLICE_X2Y94_B4 = CLBLM_R_X5Y94_SLICE_X7Y94_DO6;
  assign CLBLM_R_X3Y94_SLICE_X2Y94_B5 = CLBLM_R_X5Y94_SLICE_X6Y94_BO6;
  assign CLBLM_R_X3Y94_SLICE_X2Y94_B6 = CLBLL_L_X2Y97_SLICE_X0Y97_CO6;
  assign CLBLM_R_X7Y88_SLICE_X8Y88_SR = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y94_SLICE_X2Y94_C1 = CLBLM_R_X5Y94_SLICE_X6Y94_BO6;
  assign CLBLM_R_X3Y94_SLICE_X2Y94_C2 = CLBLL_L_X4Y94_SLICE_X5Y94_DO6;
  assign CLBLM_R_X3Y94_SLICE_X2Y94_C3 = CLBLL_L_X2Y96_SLICE_X1Y96_DO6;
  assign CLBLM_R_X3Y94_SLICE_X2Y94_C4 = CLBLM_R_X3Y93_SLICE_X2Y93_CO6;
  assign CLBLM_R_X3Y94_SLICE_X2Y94_C5 = CLBLM_R_X3Y96_SLICE_X3Y96_DO6;
  assign CLBLM_R_X3Y94_SLICE_X2Y94_C6 = CLBLM_R_X5Y94_SLICE_X7Y94_DO6;
  assign CLBLM_R_X3Y94_SLICE_X2Y94_D1 = CLBLL_L_X2Y97_SLICE_X1Y97_AO6;
  assign CLBLM_R_X3Y94_SLICE_X2Y94_D2 = CLBLL_L_X2Y97_SLICE_X0Y97_CO6;
  assign CLBLM_R_X3Y94_SLICE_X2Y94_D3 = CLBLM_R_X3Y99_SLICE_X2Y99_DO6;
  assign CLBLM_R_X3Y94_SLICE_X2Y94_D4 = CLBLM_R_X3Y93_SLICE_X2Y93_CO6;
  assign CLBLM_R_X3Y94_SLICE_X2Y94_D5 = CLBLM_R_X3Y98_SLICE_X2Y98_BO6;
  assign CLBLM_R_X3Y94_SLICE_X2Y94_D6 = 1'b1;
  assign CLBLM_R_X3Y94_SLICE_X2Y94_SR = CLBLM_R_X5Y92_SLICE_X7Y92_AO6;
  assign CLBLM_R_X7Y93_SLICE_X8Y93_D4 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO13;
  assign CLBLM_R_X7Y99_SLICE_X9Y99_B1 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X7Y99_SLICE_X9Y99_B5 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLL_L_X4Y98_SLICE_X5Y98_B5 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLL_L_X4Y98_SLICE_X5Y98_C2 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO15;
  assign CLBLL_L_X4Y98_SLICE_X5Y98_C3 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO4;
  assign CLBLM_R_X7Y93_SLICE_X8Y93_D5 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO12;
  assign CLBLM_R_X7Y89_SLICE_X9Y89_A1 = CLBLM_L_X8Y89_SLICE_X10Y89_CQ;
  assign CLBLM_R_X7Y89_SLICE_X9Y89_A2 = CLBLM_L_X8Y89_SLICE_X10Y89_A5Q;
  assign CLBLM_R_X7Y89_SLICE_X9Y89_A3 = CLBLM_L_X8Y89_SLICE_X10Y89_AQ;
  assign CLBLM_R_X7Y89_SLICE_X9Y89_A4 = CLBLM_R_X7Y89_SLICE_X9Y89_AQ;
  assign CLBLM_R_X7Y89_SLICE_X9Y89_A5 = CLBLM_L_X8Y89_SLICE_X10Y89_BQ;
  assign CLBLM_R_X7Y89_SLICE_X9Y89_A6 = 1'b1;
  assign CLBLM_R_X7Y89_SLICE_X9Y89_B1 = CLBLM_L_X8Y89_SLICE_X10Y89_CQ;
  assign CLBLM_R_X7Y89_SLICE_X9Y89_B2 = CLBLM_L_X8Y89_SLICE_X10Y89_A5Q;
  assign CLBLM_R_X7Y89_SLICE_X9Y89_B3 = CLBLM_L_X8Y89_SLICE_X10Y89_AQ;
  assign CLBLM_R_X7Y89_SLICE_X9Y89_B4 = CLBLM_R_X7Y89_SLICE_X9Y89_AQ;
  assign CLBLM_R_X7Y89_SLICE_X9Y89_B5 = CLBLM_L_X8Y89_SLICE_X10Y89_BQ;
  assign CLBLM_R_X7Y89_SLICE_X9Y89_B6 = CLBLM_R_X7Y89_SLICE_X9Y89_BQ;
  assign CLBLM_R_X7Y89_SLICE_X9Y89_C1 = CLBLM_L_X8Y89_SLICE_X10Y89_BQ;
  assign CLBLM_R_X7Y89_SLICE_X9Y89_C2 = CLBLM_L_X8Y89_SLICE_X10Y89_A5Q;
  assign CLBLM_R_X7Y89_SLICE_X9Y89_C3 = CLBLM_L_X8Y89_SLICE_X10Y89_CQ;
  assign CLBLM_R_X7Y89_SLICE_X9Y89_C4 = CLBLM_R_X7Y89_SLICE_X9Y89_BQ;
  assign CLBLM_R_X7Y89_SLICE_X9Y89_C5 = CLBLM_L_X8Y89_SLICE_X10Y89_AQ;
  assign CLBLM_R_X7Y89_SLICE_X9Y89_C6 = CLBLM_R_X7Y89_SLICE_X9Y89_AQ;
  assign CLBLM_R_X7Y89_SLICE_X9Y89_CE = CLBLM_R_X7Y88_SLICE_X8Y88_BO6;
  assign CLBLM_R_X7Y89_SLICE_X9Y89_CLK = CLBLM_R_X7Y88_SLICE_X8Y88_AQ;
  assign CLBLM_R_X7Y89_SLICE_X9Y89_D1 = CLBLM_L_X8Y89_SLICE_X10Y89_BQ;
  assign CLBLM_R_X7Y89_SLICE_X9Y89_D2 = CLBLM_R_X7Y89_SLICE_X9Y89_AQ;
  assign CLBLM_R_X7Y89_SLICE_X9Y89_D3 = CLBLM_R_X7Y89_SLICE_X8Y89_B5Q;
  assign CLBLM_R_X3Y95_SLICE_X3Y95_A1 = CLBLL_L_X4Y91_SLICE_X4Y91_AO5;
  assign CLBLM_R_X3Y95_SLICE_X3Y95_A2 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X3Y95_SLICE_X3Y95_A3 = CLBLM_R_X3Y91_SLICE_X2Y91_F7BMUX_O;
  assign CLBLM_R_X3Y95_SLICE_X3Y95_A4 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X3Y95_SLICE_X3Y95_A5 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X3Y95_SLICE_X3Y95_A6 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO4;
  assign CLBLM_R_X7Y89_SLICE_X9Y89_D4 = CLBLM_L_X8Y89_SLICE_X10Y89_CQ;
  assign CLBLM_R_X7Y89_SLICE_X9Y89_D5 = CLBLM_L_X8Y89_SLICE_X10Y89_AQ;
  assign CLBLM_R_X7Y89_SLICE_X9Y89_D6 = CLBLM_L_X8Y89_SLICE_X10Y89_A5Q;
  assign CLBLM_R_X3Y95_SLICE_X3Y95_B1 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO7;
  assign CLBLM_R_X3Y95_SLICE_X3Y95_B2 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X3Y95_SLICE_X3Y95_B3 = CLBLM_R_X3Y92_SLICE_X2Y92_F7BMUX_O;
  assign CLBLM_R_X3Y95_SLICE_X3Y95_B4 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X3Y95_SLICE_X3Y95_B5 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X3Y95_SLICE_X3Y95_B6 = CLBLL_L_X4Y91_SLICE_X4Y91_AO5;
  assign CLBLM_R_X7Y89_SLICE_X8Y89_A1 = CLBLM_R_X7Y89_SLICE_X9Y89_BQ;
  assign CLBLM_R_X7Y89_SLICE_X8Y89_A2 = CLBLM_R_X7Y89_SLICE_X9Y89_AQ;
  assign CLBLM_R_X7Y89_SLICE_X8Y89_A3 = CLBLM_R_X7Y89_SLICE_X8Y89_AQ;
  assign CLBLM_R_X3Y95_SLICE_X3Y95_C1 = CLBLM_R_X3Y95_SLICE_X3Y95_AO6;
  assign CLBLM_R_X3Y95_SLICE_X3Y95_C2 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X3Y95_SLICE_X3Y95_C3 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X3Y95_SLICE_X3Y95_C4 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X3Y95_SLICE_X3Y95_C5 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X3Y95_SLICE_X3Y95_C6 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLM_R_X7Y89_SLICE_X8Y89_B1 = CLBLM_R_X7Y89_SLICE_X8Y89_B5Q;
  assign CLBLM_R_X7Y89_SLICE_X8Y89_B2 = CLBLM_R_X7Y89_SLICE_X8Y89_BQ;
  assign CLBLM_R_X7Y89_SLICE_X8Y89_B3 = CLBLM_R_X7Y89_SLICE_X8Y89_AQ;
  assign CLBLM_R_X7Y89_SLICE_X8Y89_B4 = CLBLM_R_X7Y89_SLICE_X9Y89_CO6;
  assign CLBLM_R_X7Y89_SLICE_X8Y89_B5 = 1'b1;
  assign CLBLM_R_X7Y89_SLICE_X8Y89_B6 = 1'b1;
  assign CLBLM_R_X3Y95_SLICE_X3Y95_D1 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X3Y95_SLICE_X3Y95_D2 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO2;
  assign CLBLM_R_X3Y95_SLICE_X3Y95_D3 = CLBLM_R_X3Y94_SLICE_X3Y94_F7BMUX_O;
  assign CLBLM_R_X3Y95_SLICE_X3Y95_D4 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X3Y95_SLICE_X3Y95_D5 = CLBLL_L_X4Y91_SLICE_X4Y91_AO5;
  assign CLBLM_R_X3Y95_SLICE_X3Y95_D6 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X7Y89_SLICE_X8Y89_C1 = CLBLM_R_X7Y89_SLICE_X8Y89_BQ;
  assign CLBLM_R_X7Y89_SLICE_X8Y89_C2 = CLBLM_R_X7Y89_SLICE_X8Y89_AQ;
  assign CLBLM_R_X7Y89_SLICE_X8Y89_C4 = 1'b1;
  assign CLBLM_R_X7Y89_SLICE_X8Y89_C5 = CLBLM_R_X7Y89_SLICE_X8Y89_B5Q;
  assign CLBLM_R_X7Y89_SLICE_X8Y89_C6 = CLBLM_R_X7Y89_SLICE_X9Y89_BQ;
  assign CLBLM_R_X7Y89_SLICE_X8Y89_CE = CLBLM_R_X7Y88_SLICE_X8Y88_BO6;
  assign CLBLM_R_X3Y95_SLICE_X2Y95_A1 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X3Y95_SLICE_X2Y95_A2 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLM_R_X3Y95_SLICE_X2Y95_A3 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X3Y95_SLICE_X2Y95_A4 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X3Y95_SLICE_X2Y95_A5 = CLBLL_L_X4Y91_SLICE_X4Y91_BO6;
  assign CLBLM_R_X3Y95_SLICE_X2Y95_A6 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X7Y89_SLICE_X8Y89_D1 = 1'b1;
  assign CLBLM_R_X7Y89_SLICE_X8Y89_D2 = 1'b1;
  assign CLBLM_R_X7Y89_SLICE_X8Y89_D3 = 1'b1;
  assign CLBLM_R_X3Y95_SLICE_X2Y95_B1 = CLBLM_R_X3Y93_SLICE_X2Y93_CO5;
  assign CLBLM_R_X3Y95_SLICE_X2Y95_B2 = CLBLL_L_X2Y94_SLICE_X1Y94_D_XOR;
  assign CLBLM_R_X3Y95_SLICE_X2Y95_B3 = CLBLL_L_X4Y95_SLICE_X4Y95_BO6;
  assign CLBLM_R_X3Y95_SLICE_X2Y95_B4 = CLBLL_L_X4Y93_SLICE_X4Y93_F7AMUX_O;
  assign CLBLM_R_X3Y95_SLICE_X2Y95_B5 = CLBLL_L_X2Y93_SLICE_X0Y93_CO5;
  assign CLBLM_R_X3Y95_SLICE_X2Y95_B6 = CLBLL_L_X2Y97_SLICE_X0Y97_AO6;
  assign CLBLM_R_X7Y89_SLICE_X8Y89_SR = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y94_SLICE_X9Y94_A5 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X7Y94_SLICE_X9Y94_A6 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLM_R_X3Y95_SLICE_X2Y95_C1 = CLBLL_L_X2Y93_SLICE_X0Y93_CO5;
  assign CLBLM_R_X3Y95_SLICE_X2Y95_C2 = CLBLM_R_X3Y93_SLICE_X2Y93_CO5;
  assign CLBLM_R_X3Y95_SLICE_X2Y95_C3 = CLBLM_R_X3Y95_SLICE_X3Y95_AO6;
  assign CLBLM_R_X3Y95_SLICE_X2Y95_C4 = CLBLL_L_X2Y97_SLICE_X0Y97_AO6;
  assign CLBLM_R_X3Y95_SLICE_X2Y95_C5 = CLBLL_L_X2Y95_SLICE_X1Y95_A_XOR;
  assign CLBLM_R_X3Y95_SLICE_X2Y95_C6 = CLBLM_R_X3Y91_SLICE_X2Y91_F7AMUX_O;
  assign CLBLM_R_X7Y99_SLICE_X8Y99_B1 = CLBLM_R_X7Y99_SLICE_X8Y99_DO6;
  assign CLBLM_R_X7Y99_SLICE_X8Y99_B2 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X7Y99_SLICE_X8Y99_B3 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO0;
  assign CLBLM_R_X7Y99_SLICE_X8Y99_B4 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X3Y95_SLICE_X2Y95_D1 = CLBLL_L_X4Y91_SLICE_X4Y91_BO6;
  assign CLBLM_R_X3Y95_SLICE_X2Y95_D2 = CLBLM_R_X3Y93_SLICE_X2Y93_CO5;
  assign CLBLM_R_X3Y95_SLICE_X2Y95_D3 = CLBLL_L_X2Y93_SLICE_X0Y93_CO5;
  assign CLBLM_R_X3Y95_SLICE_X2Y95_D4 = CLBLL_L_X2Y95_SLICE_X1Y95_B_XOR;
  assign CLBLM_R_X3Y95_SLICE_X2Y95_D5 = CLBLL_L_X2Y97_SLICE_X0Y97_AO6;
  assign CLBLM_R_X3Y95_SLICE_X2Y95_D6 = CLBLM_R_X3Y91_SLICE_X3Y91_F7AMUX_O;
  assign CLBLM_R_X7Y99_SLICE_X8Y99_B6 = CLBLM_R_X5Y95_SLICE_X6Y95_AQ;
  assign CLBLM_R_X7Y94_SLICE_X9Y94_B4 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X7Y94_SLICE_X9Y94_B5 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X7Y94_SLICE_X9Y94_B6 = CLBLM_R_X7Y94_SLICE_X9Y94_CO6;
  assign CLBLM_R_X7Y99_SLICE_X8Y99_C4 = CLBLL_L_X4Y97_SLICE_X4Y97_BQ;
  assign CLBLM_R_X7Y94_SLICE_X9Y94_A3 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X7Y99_SLICE_X8Y99_C5 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X7Y99_SLICE_X8Y99_C6 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X7Y99_SLICE_X8Y99_CE = CLBLM_R_X7Y99_SLICE_X9Y99_DO6;
  assign CLBLM_R_X7Y94_SLICE_X9Y94_C5 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO14;
  assign CLBLM_R_X7Y94_SLICE_X9Y94_A4 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X7Y94_SLICE_X9Y94_CE = CLBLM_R_X7Y94_SLICE_X8Y94_CO6;
  assign CLBLM_R_X5Y96_SLICE_X7Y96_A5 = CLBLM_R_X5Y96_SLICE_X7Y96_CO5;
  assign CLBLM_R_X5Y96_SLICE_X7Y96_A6 = CLBLM_R_X7Y98_SLICE_X8Y98_F7AMUX_O;
  assign CLBLM_R_X7Y94_SLICE_X9Y94_D6 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO11;
  assign CLBLM_R_X7Y94_SLICE_X9Y94_SR = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y90_SLICE_X9Y90_C1 = CLBLM_R_X7Y91_SLICE_X9Y91_AQ;
  assign CLBLM_R_X3Y96_SLICE_X3Y96_C1 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRL3 = CLBLM_R_X5Y90_SLICE_X7Y90_BQ;
  assign CLBLM_R_X3Y96_SLICE_X3Y96_C2 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLM_R_X3Y96_SLICE_X3Y96_C3 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X3Y96_SLICE_X3Y96_C4 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X3Y96_SLICE_X3Y96_C5 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRL4 = CLBLM_R_X5Y90_SLICE_X7Y90_CQ;
  assign CLBLM_R_X3Y96_SLICE_X3Y96_D1 = CLBLM_R_X3Y98_SLICE_X3Y98_AO6;
  assign CLBLM_R_X3Y96_SLICE_X3Y96_D2 = CLBLM_R_X3Y96_SLICE_X2Y96_CO6;
  assign CLBLM_R_X3Y96_SLICE_X3Y96_D3 = CLBLL_L_X4Y97_SLICE_X4Y97_AO6;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRL5 = CLBLM_R_X5Y90_SLICE_X7Y90_DQ;
  assign CLBLM_R_X3Y96_SLICE_X3Y96_D4 = CLBLM_R_X3Y96_SLICE_X3Y96_CO6;
  assign CLBLM_R_X3Y96_SLICE_X3Y96_D5 = CLBLL_L_X4Y97_SLICE_X4Y97_CO6;
  assign CLBLM_R_X3Y96_SLICE_X3Y96_D6 = CLBLL_L_X4Y98_SLICE_X4Y98_AO6;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRL6 = CLBLM_R_X5Y90_SLICE_X7Y90_A5Q;
  assign CLBLM_R_X7Y90_SLICE_X8Y90_C5 = CLBLM_R_X7Y90_SLICE_X9Y90_AQ;
  assign CLBLM_R_X7Y90_SLICE_X8Y90_C6 = CLBLM_R_X7Y90_SLICE_X9Y90_BQ;
  assign CLBLM_R_X7Y90_SLICE_X8Y90_CLK = CLBLM_R_X7Y88_SLICE_X8Y88_AQ;
  assign CLBLM_R_X3Y96_SLICE_X2Y96_A1 = CLBLM_R_X3Y97_SLICE_X3Y97_CO6;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRL7 = CLBLM_R_X5Y90_SLICE_X7Y90_B5Q;
  assign CLBLM_R_X3Y96_SLICE_X2Y96_A2 = CLBLL_L_X4Y98_SLICE_X4Y98_DO6;
  assign CLBLM_R_X3Y96_SLICE_X2Y96_A3 = CLBLM_R_X3Y97_SLICE_X3Y97_DO6;
  assign CLBLM_R_X3Y96_SLICE_X2Y96_A4 = CLBLM_R_X3Y98_SLICE_X3Y98_DO6;
  assign CLBLM_R_X3Y96_SLICE_X2Y96_A5 = CLBLL_L_X4Y98_SLICE_X5Y98_DO6;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRL8 = CLBLM_R_X5Y90_SLICE_X7Y90_C5Q;
  assign CLBLM_R_X3Y96_SLICE_X2Y96_A6 = 1'b1;
  assign CLBLM_R_X7Y90_SLICE_X8Y90_D1 = CLBLM_R_X7Y91_SLICE_X9Y91_CQ;
  assign CLBLM_R_X3Y96_SLICE_X2Y96_AX = CLBLL_L_X2Y96_SLICE_X1Y96_BO6;
  assign CLBLM_R_X7Y90_SLICE_X8Y90_D2 = CLBLM_R_X7Y90_SLICE_X9Y90_A5Q;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRL9 = CLBLM_R_X5Y90_SLICE_X6Y90_AQ;
  assign CLBLM_R_X3Y96_SLICE_X2Y96_B1 = CLBLM_R_X3Y97_SLICE_X3Y97_CO6;
  assign CLBLM_R_X3Y96_SLICE_X2Y96_B2 = CLBLL_L_X4Y98_SLICE_X4Y98_DO6;
  assign CLBLM_R_X3Y96_SLICE_X2Y96_B3 = CLBLM_R_X3Y97_SLICE_X3Y97_DO6;
  assign CLBLM_R_X3Y96_SLICE_X2Y96_B4 = CLBLM_R_X3Y98_SLICE_X3Y98_DO6;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRL10 = CLBLM_R_X5Y90_SLICE_X6Y90_BQ;
  assign CLBLM_R_X3Y96_SLICE_X2Y96_B5 = CLBLL_L_X4Y98_SLICE_X5Y98_DO6;
  assign CLBLM_R_X3Y96_SLICE_X2Y96_B6 = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRL11 = CLBLM_R_X5Y90_SLICE_X6Y90_CQ;
  assign CLBLM_R_X3Y96_SLICE_X2Y96_BX = CLBLL_L_X2Y97_SLICE_X1Y97_CO6;
  assign CLBLM_R_X3Y96_SLICE_X2Y96_C1 = CLBLM_R_X3Y97_SLICE_X3Y97_CO6;
  assign CLBLM_R_X3Y96_SLICE_X2Y96_C2 = CLBLL_L_X4Y98_SLICE_X4Y98_DO6;
  assign CLBLM_R_X3Y96_SLICE_X2Y96_C3 = CLBLM_R_X3Y97_SLICE_X3Y97_DO6;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRL12 = CLBLM_R_X5Y90_SLICE_X6Y90_DQ;
  assign CLBLM_R_X3Y96_SLICE_X2Y96_C4 = CLBLM_R_X3Y98_SLICE_X3Y98_DO6;
  assign CLBLM_R_X3Y96_SLICE_X2Y96_C5 = CLBLL_L_X4Y98_SLICE_X5Y98_DO6;
  assign CLBLM_R_X3Y96_SLICE_X2Y96_C6 = 1'b1;
  assign CLBLM_R_X3Y96_SLICE_X2Y96_CE = CLBLM_R_X5Y94_SLICE_X6Y94_CO6;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRL13 = CLBLM_R_X5Y90_SLICE_X6Y90_A5Q;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRU0 = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRU1 = 1'b1;
  assign CLBLM_R_X3Y96_SLICE_X2Y96_DX = CLBLL_L_X2Y96_SLICE_X1Y96_AO6;
  assign CLBLM_R_X7Y94_SLICE_X8Y94_C4 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRU2 = CLBLM_R_X5Y90_SLICE_X7Y90_AQ;
  assign CLBLM_R_X7Y94_SLICE_X8Y94_C5 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X7Y94_SLICE_X8Y94_C6 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRU3 = CLBLM_R_X5Y90_SLICE_X7Y90_BQ;
  assign CLBLM_R_X7Y94_SLICE_X8Y94_CE = CLBLM_R_X7Y94_SLICE_X8Y94_CO6;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRU4 = CLBLM_R_X5Y90_SLICE_X7Y90_CQ;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRU5 = CLBLM_R_X5Y90_SLICE_X7Y90_DQ;
  assign CLBLM_R_X5Y96_SLICE_X7Y96_SR = LIOB33_X0Y107_IOB_X0Y107_I;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRU6 = CLBLM_R_X5Y90_SLICE_X7Y90_A5Q;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRU7 = CLBLM_R_X5Y90_SLICE_X7Y90_B5Q;
  assign CLBLM_L_X8Y97_SLICE_X11Y97_A1 = CLBLL_L_X4Y97_SLICE_X4Y97_BQ;
  assign CLBLM_L_X8Y97_SLICE_X11Y97_A2 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO7;
  assign CLBLM_L_X8Y97_SLICE_X11Y97_A3 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRU8 = CLBLM_R_X5Y90_SLICE_X7Y90_C5Q;
  assign CLBLM_L_X8Y97_SLICE_X11Y97_A4 = CLBLM_L_X8Y97_SLICE_X11Y97_BO6;
  assign CLBLM_L_X8Y97_SLICE_X11Y97_A5 = CLBLM_L_X8Y97_SLICE_X10Y97_DO6;
  assign CLBLM_L_X8Y97_SLICE_X11Y97_A6 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRU9 = CLBLM_R_X5Y90_SLICE_X6Y90_AQ;
  assign CLBLM_L_X8Y97_SLICE_X11Y97_AX = CLBLM_R_X7Y99_SLICE_X9Y99_DO6;
  assign CLBLM_L_X8Y97_SLICE_X11Y97_B1 = 1'b1;
  assign CLBLM_L_X8Y97_SLICE_X11Y97_B2 = CLBLM_R_X5Y97_SLICE_X6Y97_CO6;
  assign CLBLM_L_X8Y97_SLICE_X11Y97_B3 = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRU10 = CLBLM_R_X5Y90_SLICE_X6Y90_BQ;
  assign CLBLM_L_X8Y97_SLICE_X11Y97_B4 = 1'b1;
  assign CLBLM_L_X8Y97_SLICE_X11Y97_B5 = 1'b1;
  assign CLBLM_L_X8Y97_SLICE_X11Y97_B6 = CLBLM_R_X5Y97_SLICE_X7Y97_DO6;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRU11 = CLBLM_R_X5Y90_SLICE_X6Y90_CQ;
  assign CLBLM_L_X8Y97_SLICE_X11Y97_C1 = 1'b1;
  assign CLBLM_L_X8Y97_SLICE_X11Y97_C2 = 1'b1;
  assign CLBLM_L_X8Y97_SLICE_X11Y97_C3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y97_SLICE_X11Y97_C4 = 1'b1;
  assign CLBLM_L_X8Y97_SLICE_X11Y97_C5 = CLBLM_L_X8Y97_SLICE_X11Y97_AQ;
  assign CLBLM_L_X8Y97_SLICE_X11Y97_C6 = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRU12 = CLBLM_R_X5Y90_SLICE_X6Y90_DQ;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRU13 = CLBLM_R_X5Y90_SLICE_X6Y90_A5Q;
  assign CLBLM_R_X7Y94_SLICE_X8Y94_D1 = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRU14 = CLBLM_R_X5Y90_SLICE_X6Y90_B5Q;
  assign CLBLM_L_X8Y97_SLICE_X11Y97_D1 = 1'b1;
  assign CLBLM_L_X8Y97_SLICE_X11Y97_D2 = 1'b1;
  assign CLBLM_L_X8Y97_SLICE_X11Y97_D3 = 1'b1;
  assign CLBLM_L_X8Y97_SLICE_X11Y97_D4 = 1'b1;
  assign CLBLM_L_X8Y97_SLICE_X11Y97_D5 = 1'b1;
  assign CLBLM_L_X8Y97_SLICE_X11Y97_D6 = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRL0 = 1'b1;
  assign CLBLM_R_X7Y94_SLICE_X8Y94_D2 = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRL1 = 1'b1;
  assign CLBLM_R_X7Y94_SLICE_X8Y94_D3 = 1'b1;
  assign CLBLM_R_X7Y94_SLICE_X8Y94_D4 = 1'b1;
  assign CLBLM_L_X8Y97_SLICE_X10Y97_A1 = CLBLM_R_X7Y97_SLICE_X9Y97_AQ;
  assign CLBLM_L_X8Y97_SLICE_X10Y97_A2 = CLBLM_R_X7Y97_SLICE_X9Y97_A5Q;
  assign CLBLM_L_X8Y97_SLICE_X10Y97_A3 = CLBLM_R_X7Y97_SLICE_X9Y97_BQ;
  assign CLBLM_L_X8Y97_SLICE_X10Y97_A4 = CLBLM_R_X7Y97_SLICE_X9Y97_B5Q;
  assign CLBLM_L_X8Y97_SLICE_X10Y97_A5 = 1'b0;
  assign CLBLM_L_X8Y97_SLICE_X10Y97_A6 = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRL2 = CLBLM_R_X7Y90_SLICE_X9Y90_A5Q;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRL3 = CLBLM_R_X7Y90_SLICE_X9Y90_BQ;
  assign CLBLM_R_X7Y94_SLICE_X8Y94_D5 = 1'b1;
  assign CLBLM_L_X8Y97_SLICE_X10Y97_AX = CLBLM_R_X7Y98_SLICE_X9Y98_AQ;
  assign CLBLM_L_X8Y97_SLICE_X10Y97_B1 = CLBLM_R_X7Y97_SLICE_X9Y97_AQ;
  assign CLBLM_L_X8Y97_SLICE_X10Y97_B2 = CLBLM_R_X7Y97_SLICE_X9Y97_A5Q;
  assign CLBLM_L_X8Y97_SLICE_X10Y97_B3 = CLBLM_R_X7Y97_SLICE_X9Y97_BQ;
  assign CLBLM_L_X8Y97_SLICE_X10Y97_B4 = CLBLM_R_X7Y97_SLICE_X9Y97_B5Q;
  assign CLBLM_L_X8Y97_SLICE_X10Y97_B5 = 1'b0;
  assign CLBLM_L_X8Y97_SLICE_X10Y97_B6 = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRL5 = CLBLM_R_X7Y91_SLICE_X9Y91_AQ;
  assign CLBLM_R_X5Y96_SLICE_X6Y96_B1 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_L_X8Y97_SLICE_X10Y97_BX = CLBLM_R_X7Y99_SLICE_X9Y99_AQ;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRL6 = CLBLM_R_X7Y87_SLICE_X8Y87_BQ;
  assign CLBLM_L_X8Y97_SLICE_X10Y97_C1 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO6;
  assign CLBLM_L_X8Y97_SLICE_X10Y97_C2 = CLBLM_R_X5Y97_SLICE_X7Y97_DO6;
  assign CLBLM_L_X8Y97_SLICE_X10Y97_C3 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_L_X8Y97_SLICE_X10Y97_C4 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_L_X8Y97_SLICE_X10Y97_C5 = CLBLL_L_X4Y97_SLICE_X4Y97_BQ;
  assign CLBLM_L_X8Y97_SLICE_X10Y97_C6 = CLBLM_R_X5Y97_SLICE_X6Y97_CO6;
  assign CLBLM_L_X8Y97_SLICE_X10Y97_CE = CLBLL_L_X4Y97_SLICE_X5Y97_DO6;
  assign CLBLM_R_X5Y96_SLICE_X6Y96_B2 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X5Y96_SLICE_X6Y96_B3 = CLBLL_L_X4Y97_SLICE_X4Y97_BQ;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRL8 = CLBLM_R_X7Y87_SLICE_X8Y87_AQ;
  assign CLBLM_R_X7Y89_SLICE_X9Y89_SR = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y97_SLICE_X10Y97_D1 = CLBLM_R_X7Y97_SLICE_X9Y97_AQ;
  assign CLBLM_L_X8Y97_SLICE_X10Y97_D2 = CLBLM_R_X7Y97_SLICE_X9Y97_A5Q;
  assign CLBLM_L_X8Y97_SLICE_X10Y97_D3 = CLBLM_R_X7Y97_SLICE_X9Y97_BQ;
  assign CLBLM_L_X8Y97_SLICE_X10Y97_D4 = CLBLM_R_X7Y97_SLICE_X9Y97_B5Q;
  assign CLBLM_L_X8Y97_SLICE_X10Y97_D5 = 1'b0;
  assign CLBLM_L_X8Y97_SLICE_X10Y97_DI = 1'b1;
  assign CLBLM_L_X8Y97_SLICE_X10Y97_DX = CLBLM_R_X7Y96_SLICE_X9Y96_AQ;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRL12 = CLBLM_R_X7Y89_SLICE_X8Y89_AQ;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRL13 = CLBLM_R_X7Y89_SLICE_X8Y89_BQ;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRL15 = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRU0 = 1'b1;
  assign CLBLM_R_X7Y89_SLICE_X8Y89_A4 = CLBLM_L_X8Y89_SLICE_X10Y89_A5Q;
  assign CLBLM_R_X5Y96_SLICE_X6Y96_C1 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRU1 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X1Y91_D6 = 1'b1;
  assign CLBLM_R_X7Y89_SLICE_X8Y89_A5 = CLBLM_L_X8Y89_SLICE_X10Y89_AQ;
  assign CLBLM_R_X5Y96_SLICE_X6Y96_C2 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRU2 = CLBLM_R_X7Y90_SLICE_X9Y90_A5Q;
  assign CLBLM_R_X7Y89_SLICE_X8Y89_A6 = CLBLM_L_X8Y89_SLICE_X10Y89_BO6;
  assign CLBLM_R_X5Y96_SLICE_X6Y96_C3 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO5;
  assign CLBLM_R_X5Y96_SLICE_X6Y96_C4 = CLBLM_R_X5Y95_SLICE_X6Y95_AQ;
  assign CLBLM_R_X5Y96_SLICE_X6Y96_C5 = CLBLL_L_X4Y97_SLICE_X4Y97_BQ;
  assign CLBLM_R_X5Y91_SLICE_X7Y91_C2 = 1'b1;
  assign CLBLM_R_X7Y91_SLICE_X9Y91_A1 = CLBLM_R_X7Y90_SLICE_X8Y90_CO6;
  assign CLBLM_R_X5Y96_SLICE_X6Y96_C6 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X7Y91_SLICE_X9Y91_A2 = CLBLM_R_X7Y87_SLICE_X8Y87_AQ;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRU6 = CLBLM_R_X7Y87_SLICE_X8Y87_BQ;
  assign CLBLM_R_X7Y91_SLICE_X9Y91_A3 = CLBLM_R_X7Y91_SLICE_X9Y91_AQ;
  assign CLBLM_R_X7Y91_SLICE_X9Y91_A4 = CLBLM_R_X7Y90_SLICE_X9Y90_CQ;
  assign CLBLM_R_X5Y96_SLICE_X6Y96_CE = CLBLM_R_X7Y99_SLICE_X9Y99_DO6;
  assign CLBLM_R_X7Y91_SLICE_X9Y91_A5 = CLBLM_R_X7Y91_SLICE_X8Y91_AQ;
  assign CLBLM_R_X7Y91_SLICE_X9Y91_A6 = CLBLM_R_X7Y87_SLICE_X8Y87_BQ;
  assign CLBLM_R_X7Y91_SLICE_X9Y91_B1 = CLBLM_R_X7Y87_SLICE_X8Y87_AQ;
  assign CLBLM_R_X7Y91_SLICE_X9Y91_B2 = CLBLM_R_X7Y91_SLICE_X9Y91_BQ;
  assign CLBLM_R_X7Y91_SLICE_X9Y91_B3 = CLBLM_R_X7Y91_SLICE_X9Y91_AQ;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRU8 = CLBLM_R_X7Y87_SLICE_X8Y87_AQ;
  assign CLBLM_R_X5Y91_SLICE_X7Y91_C5 = 1'b1;
  assign CLBLM_R_X7Y91_SLICE_X9Y91_B4 = CLBLM_R_X7Y87_SLICE_X8Y87_BQ;
  assign CLBLM_R_X7Y91_SLICE_X9Y91_B5 = CLBLM_R_X7Y90_SLICE_X9Y90_CQ;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRU9 = CLBLM_L_X8Y89_SLICE_X10Y89_A5Q;
  assign CLBLM_R_X7Y91_SLICE_X9Y91_B6 = CLBLM_R_X7Y91_SLICE_X8Y91_AQ;
  assign CLBLM_R_X7Y91_SLICE_X9Y91_C1 = 1'b1;
  assign CLBLM_R_X7Y91_SLICE_X9Y91_C2 = CLBLM_R_X7Y91_SLICE_X9Y91_CQ;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRU10 = CLBLM_R_X7Y89_SLICE_X9Y89_AQ;
  assign CLBLM_R_X7Y91_SLICE_X9Y91_C3 = CLBLM_R_X7Y91_SLICE_X9Y91_BQ;
  assign CLBLM_R_X7Y91_SLICE_X9Y91_C4 = 1'b1;
  assign CLBLM_R_X7Y91_SLICE_X9Y91_C5 = CLBLM_R_X7Y91_SLICE_X9Y91_DO6;
  assign CLBLM_R_X7Y91_SLICE_X9Y91_C6 = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRU11 = CLBLM_R_X7Y89_SLICE_X9Y89_BQ;
  assign CLBLM_R_X7Y91_SLICE_X9Y91_CLK = CLBLM_R_X7Y88_SLICE_X8Y88_AQ;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRU12 = CLBLM_R_X7Y89_SLICE_X8Y89_AQ;
  assign CLBLM_R_X7Y91_SLICE_X9Y91_D1 = CLBLM_R_X7Y90_SLICE_X9Y90_CQ;
  assign CLBLM_R_X7Y91_SLICE_X9Y91_D2 = CLBLM_R_X7Y87_SLICE_X8Y87_AQ;
  assign CLBLM_R_X7Y91_SLICE_X9Y91_D3 = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRU13 = CLBLM_R_X7Y89_SLICE_X8Y89_BQ;
  assign CLBLM_R_X3Y97_SLICE_X3Y97_A1 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO13;
  assign CLBLM_R_X3Y97_SLICE_X3Y97_A2 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO15;
  assign CLBLM_R_X3Y97_SLICE_X3Y97_A3 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO12;
  assign CLBLM_R_X3Y97_SLICE_X3Y97_A4 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO11;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRU14 = CLBLM_R_X7Y89_SLICE_X8Y89_B5Q;
  assign CLBLM_R_X3Y97_SLICE_X3Y97_A5 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO14;
  assign CLBLM_R_X3Y97_SLICE_X3Y97_A6 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO0;
  assign CLBLM_R_X7Y91_SLICE_X9Y91_D4 = CLBLM_R_X7Y91_SLICE_X8Y91_AQ;
  assign CLBLM_R_X3Y97_SLICE_X3Y97_B1 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO13;
  assign CLBLM_R_X3Y97_SLICE_X3Y97_B2 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO15;
  assign CLBLM_R_X3Y97_SLICE_X3Y97_B3 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO12;
  assign CLBLM_R_X3Y97_SLICE_X3Y97_B4 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO11;
  assign CLBLM_R_X3Y97_SLICE_X3Y97_B5 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO14;
  assign CLBLM_R_X3Y97_SLICE_X3Y97_B6 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO2;
  assign CLBLM_R_X7Y91_SLICE_X8Y91_A1 = CLBLM_R_X7Y90_SLICE_X8Y90_CO6;
  assign CLBLM_R_X7Y91_SLICE_X8Y91_A2 = CLBLM_R_X7Y90_SLICE_X9Y90_CQ;
  assign CLBLM_R_X3Y97_SLICE_X3Y97_C1 = CLBLM_R_X3Y97_SLICE_X3Y97_AO6;
  assign CLBLM_R_X3Y97_SLICE_X3Y97_C2 = CLBLL_L_X4Y97_SLICE_X5Y97_AO6;
  assign CLBLM_R_X3Y97_SLICE_X3Y97_C3 = CLBLM_R_X3Y96_SLICE_X3Y96_AO5;
  assign CLBLM_R_X3Y97_SLICE_X3Y97_C4 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO0;
  assign CLBLM_R_X3Y97_SLICE_X3Y97_C5 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X3Y97_SLICE_X3Y97_C6 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLM_R_X7Y91_SLICE_X8Y91_B1 = 1'b1;
  assign CLBLM_R_X7Y91_SLICE_X8Y91_B2 = CLBLM_R_X7Y87_SLICE_X8Y87_BQ;
  assign CLBLM_R_X7Y91_SLICE_X8Y91_B3 = CLBLM_R_X7Y91_SLICE_X8Y91_AQ;
  assign CLBLM_R_X3Y93_SLICE_X3Y93_A1 = CLBLM_R_X3Y95_SLICE_X3Y95_DO6;
  assign CLBLM_R_X7Y91_SLICE_X8Y91_B4 = CLBLM_R_X7Y89_SLICE_X8Y89_CO6;
  assign CLBLM_R_X7Y91_SLICE_X8Y91_B5 = BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO0;
  assign CLBLM_R_X7Y91_SLICE_X8Y91_B6 = CLBLM_R_X7Y87_SLICE_X8Y87_AQ;
  assign CLBLM_R_X3Y93_SLICE_X3Y93_A2 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLM_R_X3Y97_SLICE_X3Y97_D1 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLM_R_X3Y97_SLICE_X3Y97_D2 = CLBLL_L_X4Y97_SLICE_X5Y97_AO6;
  assign CLBLM_R_X3Y97_SLICE_X3Y97_D3 = CLBLM_R_X3Y96_SLICE_X3Y96_AO5;
  assign CLBLM_R_X3Y97_SLICE_X3Y97_D4 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X3Y93_SLICE_X3Y93_A3 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X3Y97_SLICE_X3Y97_D5 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO2;
  assign CLBLM_R_X3Y97_SLICE_X3Y97_D6 = CLBLM_R_X3Y97_SLICE_X3Y97_BO6;
  assign CLBLM_R_X7Y89_SLICE_X8Y89_C3 = 1'b1;
  assign CLBLM_R_X3Y93_SLICE_X3Y93_A4 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X7Y91_SLICE_X8Y91_C5 = 1'b1;
  assign CLBLM_R_X7Y91_SLICE_X8Y91_C6 = CLBLM_R_X7Y89_SLICE_X8Y89_CO6;
  assign CLBLM_R_X7Y91_SLICE_X8Y91_CLK = CLBLM_R_X7Y88_SLICE_X8Y88_AQ;
  assign CLBLM_R_X3Y97_SLICE_X2Y97_A1 = CLBLM_R_X3Y97_SLICE_X3Y97_CO6;
  assign CLBLM_R_X3Y93_SLICE_X3Y93_A5 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X3Y97_SLICE_X2Y97_A2 = CLBLL_L_X4Y98_SLICE_X4Y98_DO6;
  assign CLBLM_R_X3Y97_SLICE_X2Y97_A3 = CLBLM_R_X3Y97_SLICE_X3Y97_DO6;
  assign CLBLM_R_X3Y97_SLICE_X2Y97_A4 = CLBLM_R_X3Y98_SLICE_X3Y98_DO6;
  assign CLBLM_R_X3Y97_SLICE_X2Y97_A5 = CLBLL_L_X4Y98_SLICE_X5Y98_DO6;
  assign CLBLM_R_X3Y93_SLICE_X3Y93_A6 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X3Y97_SLICE_X2Y97_A6 = 1'b1;
  assign CLBLM_R_X3Y97_SLICE_X2Y97_AX = CLBLL_L_X2Y97_SLICE_X1Y97_AO6;
  assign CLBLM_R_X3Y98_SLICE_X2Y98_B1 = CLBLM_R_X3Y98_SLICE_X2Y98_DO6;
  assign CLBLM_R_X3Y97_SLICE_X2Y97_B1 = CLBLM_R_X3Y97_SLICE_X3Y97_CO6;
  assign CLBLM_R_X3Y97_SLICE_X2Y97_B2 = CLBLL_L_X4Y98_SLICE_X4Y98_DO6;
  assign CLBLM_R_X3Y97_SLICE_X2Y97_B3 = CLBLM_R_X3Y97_SLICE_X3Y97_DO6;
  assign CLBLM_R_X3Y97_SLICE_X2Y97_B4 = CLBLM_R_X3Y98_SLICE_X3Y98_DO6;
  assign CLBLM_R_X3Y97_SLICE_X2Y97_B5 = CLBLL_L_X4Y98_SLICE_X5Y98_DO6;
  assign CLBLM_R_X3Y97_SLICE_X2Y97_B6 = 1'b1;
  assign CLBLM_R_X7Y91_SLICE_X8Y91_SR = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y97_SLICE_X2Y97_BX = CLBLL_L_X2Y97_SLICE_X0Y97_CO6;
  assign CLBLM_R_X3Y93_SLICE_X3Y93_AX = CLBLL_L_X4Y93_SLICE_X4Y93_CO5;
  assign CLBLM_R_X3Y97_SLICE_X2Y97_C1 = CLBLM_R_X3Y97_SLICE_X3Y97_CO6;
  assign CLBLM_R_X3Y97_SLICE_X2Y97_C2 = CLBLL_L_X4Y98_SLICE_X4Y98_DO6;
  assign CLBLM_R_X3Y97_SLICE_X2Y97_C3 = CLBLM_R_X3Y97_SLICE_X3Y97_DO6;
  assign CLBLM_R_X3Y97_SLICE_X2Y97_C4 = CLBLM_R_X3Y98_SLICE_X3Y98_DO6;
  assign CLBLM_R_X3Y97_SLICE_X2Y97_C5 = CLBLL_L_X4Y98_SLICE_X5Y98_DO6;
  assign CLBLM_R_X3Y97_SLICE_X2Y97_C6 = 1'b1;
  assign CLBLM_R_X3Y97_SLICE_X2Y97_CE = CLBLM_R_X5Y94_SLICE_X6Y94_CO6;
  assign CLBLM_R_X3Y98_SLICE_X2Y98_B3 = CLBLM_R_X3Y97_SLICE_X2Y97_AO6;
  assign CLBLM_R_X3Y93_SLICE_X3Y93_B1 = 1'b1;
  assign CLBLM_R_X7Y89_SLICE_X8Y89_CLK = CLBLM_R_X7Y88_SLICE_X8Y88_AQ;
  assign CLBLM_R_X3Y93_SLICE_X3Y93_B2 = CLBLL_L_X2Y93_SLICE_X0Y93_CO6;
  assign CLBLM_R_X3Y97_SLICE_X2Y97_CX = CLBLL_L_X2Y97_SLICE_X1Y97_BO6;
  assign CLBLM_R_X3Y97_SLICE_X2Y97_D1 = CLBLM_R_X3Y97_SLICE_X3Y97_CO6;
  assign CLBLM_R_X3Y97_SLICE_X2Y97_D2 = CLBLL_L_X4Y98_SLICE_X4Y98_DO6;
  assign CLBLM_R_X3Y97_SLICE_X2Y97_D3 = CLBLM_R_X3Y97_SLICE_X3Y97_DO6;
  assign CLBLM_R_X3Y93_SLICE_X3Y93_B3 = 1'b1;
  assign CLBLM_R_X3Y97_SLICE_X2Y97_D4 = CLBLM_R_X3Y98_SLICE_X3Y98_DO6;
  assign CLBLM_R_X3Y97_SLICE_X2Y97_D5 = CLBLL_L_X4Y98_SLICE_X5Y98_DO6;
  assign CLBLM_R_X3Y97_SLICE_X2Y97_D6 = 1'b1;
  assign CLBLM_R_X3Y97_SLICE_X2Y97_DI = 1'b1;
  assign CLBLM_R_X3Y93_SLICE_X3Y93_B4 = CLBLL_L_X4Y94_SLICE_X5Y94_DO6;
  assign CLBLM_R_X3Y97_SLICE_X2Y97_DX = CLBLL_L_X2Y97_SLICE_X0Y97_BO6;
  assign CLBLM_R_X3Y93_SLICE_X3Y93_B5 = CLBLM_R_X5Y94_SLICE_X6Y94_BO6;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIADI10 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIADI14 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIADI16 = 1'b0;
  assign CLBLM_R_X3Y98_SLICE_X2Y98_C2 = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIADI18 = 1'b0;
  assign CLBLM_R_X3Y98_SLICE_X2Y98_C3 = CLBLL_L_X2Y99_SLICE_X1Y99_AQ;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIADI20 = 1'b0;
  assign CLBLM_R_X7Y89_SLICE_X8Y89_D4 = 1'b1;
  assign CLBLM_R_X3Y98_SLICE_X2Y98_C4 = CLBLM_R_X3Y97_SLICE_X2Y97_CO6;
  assign CLBLM_L_X8Y98_SLICE_X11Y98_A1 = 1'b1;
  assign CLBLM_L_X8Y98_SLICE_X11Y98_A2 = 1'b1;
  assign CLBLM_L_X8Y98_SLICE_X11Y98_A3 = 1'b1;
  assign CLBLM_L_X8Y98_SLICE_X11Y98_A4 = 1'b1;
  assign CLBLM_L_X8Y98_SLICE_X11Y98_A5 = 1'b1;
  assign CLBLM_L_X8Y98_SLICE_X11Y98_A6 = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIADI22 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIADI24 = 1'b0;
  assign CLBLM_R_X7Y89_SLICE_X8Y89_D5 = 1'b1;
  assign CLBLM_L_X8Y98_SLICE_X11Y98_B1 = 1'b1;
  assign CLBLM_L_X8Y98_SLICE_X11Y98_B2 = 1'b1;
  assign CLBLM_L_X8Y98_SLICE_X11Y98_B3 = 1'b1;
  assign CLBLM_L_X8Y98_SLICE_X11Y98_B4 = 1'b1;
  assign CLBLM_L_X8Y98_SLICE_X11Y98_B5 = 1'b1;
  assign CLBLM_L_X8Y98_SLICE_X11Y98_B6 = 1'b1;
  assign CLBLM_L_X8Y98_SLICE_X11Y98_C1 = 1'b1;
  assign CLBLM_L_X8Y98_SLICE_X11Y98_C2 = 1'b1;
  assign CLBLM_L_X8Y98_SLICE_X11Y98_C3 = 1'b1;
  assign CLBLM_L_X8Y98_SLICE_X11Y98_C4 = 1'b1;
  assign CLBLM_L_X8Y98_SLICE_X11Y98_C5 = 1'b1;
  assign CLBLM_L_X8Y98_SLICE_X11Y98_C6 = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIADI1 = CLBLM_R_X5Y93_SLICE_X7Y93_AQ;
  assign CLBLM_L_X8Y98_SLICE_X11Y98_D1 = 1'b1;
  assign CLBLM_L_X8Y98_SLICE_X11Y98_D2 = 1'b1;
  assign CLBLM_L_X8Y98_SLICE_X11Y98_D3 = 1'b1;
  assign CLBLM_L_X8Y98_SLICE_X11Y98_D4 = 1'b1;
  assign CLBLM_L_X8Y98_SLICE_X11Y98_D5 = 1'b1;
  assign CLBLM_L_X8Y98_SLICE_X11Y98_D6 = 1'b1;
  assign CLBLM_L_X8Y98_SLICE_X10Y98_A1 = CLBLM_R_X5Y97_SLICE_X7Y97_DO6;
  assign CLBLM_L_X8Y98_SLICE_X10Y98_A2 = CLBLM_R_X5Y97_SLICE_X6Y97_CO6;
  assign CLBLM_L_X8Y98_SLICE_X10Y98_A3 = CLBLM_L_X8Y97_SLICE_X10Y97_AO6;
  assign CLBLM_L_X8Y98_SLICE_X10Y98_A4 = CLBLM_L_X8Y97_SLICE_X10Y97_DO6;
  assign CLBLM_L_X8Y98_SLICE_X10Y98_A5 = 1'b1;
  assign CLBLM_L_X8Y98_SLICE_X10Y98_A6 = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIADI11 = 1'b0;
  assign CLBLM_L_X8Y98_SLICE_X10Y98_B1 = CLBLM_R_X5Y97_SLICE_X6Y97_CO6;
  assign CLBLM_L_X8Y98_SLICE_X10Y98_B2 = CLBLM_R_X5Y98_SLICE_X6Y98_AO6;
  assign CLBLM_L_X8Y98_SLICE_X10Y98_B3 = CLBLM_L_X8Y97_SLICE_X10Y97_AO6;
  assign CLBLM_L_X8Y98_SLICE_X10Y98_B4 = CLBLM_L_X8Y97_SLICE_X10Y97_DO6;
  assign CLBLM_L_X8Y98_SLICE_X10Y98_B5 = CLBLM_L_X8Y97_SLICE_X10Y97_BO6;
  assign CLBLM_L_X8Y98_SLICE_X10Y98_B6 = CLBLM_R_X5Y97_SLICE_X7Y97_DO6;
  assign CLBLM_R_X7Y97_SLICE_X8Y97_B3 = CLBLM_R_X7Y99_SLICE_X9Y99_AQ;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_D1 = CLBLL_L_X4Y90_SLICE_X5Y90_AQ;
  assign CLBLM_L_X8Y98_SLICE_X10Y98_C1 = CLBLM_L_X8Y97_SLICE_X10Y97_AO6;
  assign CLBLM_L_X8Y98_SLICE_X10Y98_C2 = CLBLL_L_X4Y97_SLICE_X4Y97_BQ;
  assign CLBLM_L_X8Y98_SLICE_X10Y98_C3 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_L_X8Y98_SLICE_X10Y98_C4 = CLBLM_L_X8Y98_SLICE_X10Y98_AO5;
  assign CLBLM_L_X8Y98_SLICE_X10Y98_C5 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO8;
  assign CLBLM_L_X8Y98_SLICE_X10Y98_C6 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIADI21 = 1'b0;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_T1 = 1'b1;
  assign CLBLM_L_X8Y98_SLICE_X10Y98_D1 = CLBLM_L_X8Y98_SLICE_X10Y98_AO6;
  assign CLBLM_L_X8Y98_SLICE_X10Y98_D2 = CLBLM_L_X8Y97_SLICE_X10Y97_BO6;
  assign CLBLM_L_X8Y98_SLICE_X10Y98_D3 = CLBLL_L_X4Y97_SLICE_X4Y97_BQ;
  assign CLBLM_L_X8Y98_SLICE_X10Y98_D4 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_L_X8Y98_SLICE_X10Y98_D5 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_L_X8Y98_SLICE_X10Y98_D6 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO9;
  assign CLBLM_R_X7Y97_SLICE_X8Y97_B4 = CLBLM_R_X7Y98_SLICE_X9Y98_AQ;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_D1 = CLBLM_R_X7Y91_SLICE_X8Y91_CO6;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_T1 = 1'b1;
  assign LIOB33_X0Y101_IOB_X0Y102_O = CLBLL_L_X4Y90_SLICE_X5Y90_AQ;
  assign LIOB33_X0Y101_IOB_X0Y101_O = CLBLM_R_X7Y91_SLICE_X8Y91_CO6;
  assign CLBLL_L_X2Y90_SLICE_X0Y90_A1 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X0Y90_A2 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X0Y90_A3 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X0Y90_A4 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X0Y90_A5 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X0Y90_A6 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X0Y90_B1 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X0Y90_B2 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X0Y90_B3 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X0Y90_B4 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X0Y90_B5 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X0Y90_B6 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X0Y90_C1 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X0Y90_C2 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X0Y90_C3 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X0Y90_C4 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X0Y90_C5 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X0Y90_C6 = 1'b1;
  assign CLBLM_R_X3Y98_SLICE_X3Y98_A1 = CLBLM_R_X3Y96_SLICE_X3Y96_AO5;
  assign CLBLM_R_X3Y98_SLICE_X3Y98_A2 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO7;
  assign CLBLM_R_X3Y98_SLICE_X3Y98_A3 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLM_R_X3Y98_SLICE_X3Y98_A4 = CLBLM_R_X3Y98_SLICE_X3Y98_BO6;
  assign CLBLM_R_X3Y98_SLICE_X3Y98_A5 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X3Y98_SLICE_X3Y98_A6 = CLBLL_L_X4Y97_SLICE_X5Y97_AO6;
  assign CLBLL_L_X2Y90_SLICE_X0Y90_D1 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X0Y90_D2 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X0Y90_D3 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X0Y90_D4 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X0Y90_D5 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X0Y90_D6 = 1'b1;
  assign CLBLM_R_X3Y98_SLICE_X3Y98_B1 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO12;
  assign CLBLM_R_X3Y98_SLICE_X3Y98_B2 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO7;
  assign CLBLM_R_X3Y98_SLICE_X3Y98_B3 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO11;
  assign CLBLM_R_X3Y98_SLICE_X3Y98_B4 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO15;
  assign CLBLM_R_X3Y98_SLICE_X3Y98_B5 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO13;
  assign CLBLM_R_X3Y98_SLICE_X3Y98_B6 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO14;
  assign CLBLM_R_X3Y98_SLICE_X3Y98_C1 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO13;
  assign CLBLM_R_X3Y98_SLICE_X3Y98_C2 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO14;
  assign CLBLM_R_X3Y98_SLICE_X3Y98_C3 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO3;
  assign CLBLM_R_X3Y98_SLICE_X3Y98_C4 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO11;
  assign CLBLM_R_X3Y98_SLICE_X3Y98_C5 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO12;
  assign CLBLM_R_X3Y98_SLICE_X3Y98_C6 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO15;
  assign CLBLM_R_X3Y98_SLICE_X3Y98_D1 = CLBLL_L_X4Y97_SLICE_X5Y97_AO6;
  assign CLBLM_R_X3Y98_SLICE_X3Y98_D2 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLM_R_X3Y98_SLICE_X3Y98_D3 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO3;
  assign CLBLM_R_X3Y98_SLICE_X3Y98_D4 = CLBLM_R_X3Y98_SLICE_X3Y98_CO6;
  assign CLBLM_R_X3Y98_SLICE_X3Y98_D5 = CLBLM_R_X3Y96_SLICE_X3Y96_AO5;
  assign CLBLM_R_X3Y98_SLICE_X3Y98_D6 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLL_L_X2Y90_SLICE_X1Y90_A1 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X1Y90_A2 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X1Y90_A3 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X1Y90_A4 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X1Y90_A5 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X1Y90_A6 = 1'b1;
  assign CLBLM_R_X3Y98_SLICE_X2Y98_A1 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO3;
  assign CLBLM_R_X3Y98_SLICE_X2Y98_A2 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLL_L_X2Y90_SLICE_X1Y90_AX = CLBLL_L_X4Y92_SLICE_X4Y92_AO6;
  assign CLBLM_R_X3Y98_SLICE_X2Y98_A3 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLL_L_X2Y90_SLICE_X1Y90_B1 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X1Y90_B2 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X1Y90_B3 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X1Y90_B4 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X1Y90_B5 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X1Y90_B6 = 1'b1;
  assign CLBLM_R_X3Y98_SLICE_X2Y98_A4 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X3Y98_SLICE_X2Y98_A5 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X3Y98_SLICE_X2Y98_A6 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLL_L_X2Y90_SLICE_X1Y90_C1 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X1Y90_C2 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X1Y90_C3 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X1Y90_C4 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X1Y90_C5 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X1Y90_C6 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X1Y90_CE = CLBLL_L_X2Y92_SLICE_X1Y92_AO6;
  assign CLBLM_R_X3Y98_SLICE_X2Y98_B2 = CLBLL_L_X4Y98_SLICE_X5Y98_BO6;
  assign CLBLM_R_X3Y98_SLICE_X2Y98_B4 = CLBLL_L_X2Y98_SLICE_X0Y98_AQ;
  assign CLBLM_R_X3Y98_SLICE_X2Y98_B5 = CLBLL_L_X4Y97_SLICE_X4Y97_AO6;
  assign CLBLM_R_X3Y98_SLICE_X2Y98_B6 = 1'b1;
  assign CLBLM_R_X3Y98_SLICE_X2Y98_C1 = CLBLM_R_X3Y98_SLICE_X2Y98_AO6;
  assign CLBLL_L_X2Y90_SLICE_X1Y90_D1 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X1Y90_D2 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X1Y90_D3 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X1Y90_D4 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X1Y90_D5 = 1'b1;
  assign CLBLL_L_X2Y90_SLICE_X1Y90_D6 = 1'b1;
  assign CLBLM_R_X3Y98_SLICE_X2Y98_C5 = CLBLL_L_X4Y97_SLICE_X4Y97_AO6;
  assign CLBLM_R_X3Y98_SLICE_X2Y98_C6 = CLBLM_R_X3Y98_SLICE_X2Y98_DO6;
  assign CLBLM_R_X3Y98_SLICE_X2Y98_D1 = 1'b1;
  assign CLBLM_R_X3Y98_SLICE_X2Y98_D3 = CLBLL_L_X4Y97_SLICE_X4Y97_CO6;
  assign CLBLM_R_X3Y98_SLICE_X2Y98_D4 = 1'b1;
  assign CLBLM_R_X3Y98_SLICE_X2Y98_D5 = 1'b1;
  assign CLBLM_R_X3Y98_SLICE_X2Y98_D6 = CLBLL_L_X4Y98_SLICE_X4Y98_AO6;
  assign CLBLM_R_X3Y98_SLICE_X2Y98_D2 = CLBLM_R_X3Y98_SLICE_X3Y98_AO6;
  assign CLBLM_R_X7Y96_SLICE_X8Y96_B2 = 1'b1;
  assign LIOB33_X0Y103_IOB_X0Y104_O = CLBLL_L_X2Y102_SLICE_X0Y102_AQ;
  assign LIOB33_X0Y103_IOB_X0Y103_O = CLBLM_R_X7Y91_SLICE_X8Y91_DO6;
  assign CLBLL_L_X2Y91_SLICE_X0Y91_A1 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X0Y91_A2 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X0Y91_A3 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X0Y91_A4 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X0Y91_A5 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X0Y91_A6 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X0Y91_AX = CLBLL_L_X4Y92_SLICE_X4Y92_AO6;
  assign CLBLL_L_X2Y91_SLICE_X0Y91_B1 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X0Y91_B2 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X0Y91_B3 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X0Y91_B4 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X0Y91_B5 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X0Y91_B6 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X0Y91_C1 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X0Y91_C2 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X0Y91_C3 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X0Y91_C4 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X0Y91_C5 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X0Y91_C6 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X0Y91_CE = CLBLL_L_X2Y93_SLICE_X0Y93_DO6;
  assign CLBLL_L_X2Y91_SLICE_X0Y91_D1 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X0Y91_D2 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X0Y91_D3 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X0Y91_D4 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X0Y91_D5 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X0Y91_D6 = 1'b1;
  assign CLBLM_R_X3Y99_SLICE_X3Y99_B2 = 1'b1;
  assign CLBLM_R_X3Y99_SLICE_X3Y99_B3 = 1'b1;
  assign CLBLM_R_X3Y99_SLICE_X3Y99_B4 = 1'b1;
  assign CLBLM_R_X3Y99_SLICE_X3Y99_B5 = 1'b1;
  assign CLBLM_R_X3Y99_SLICE_X3Y99_B6 = 1'b1;
  assign CLBLM_R_X3Y99_SLICE_X3Y99_C1 = 1'b1;
  assign CLBLM_R_X3Y99_SLICE_X3Y99_C2 = 1'b1;
  assign CLBLM_R_X3Y99_SLICE_X3Y99_C3 = 1'b1;
  assign CLBLM_R_X3Y99_SLICE_X3Y99_C4 = 1'b1;
  assign CLBLM_R_X3Y99_SLICE_X3Y99_C5 = 1'b1;
  assign CLBLM_R_X3Y99_SLICE_X3Y99_C6 = 1'b1;
  assign CLBLM_R_X7Y93_SLICE_X8Y93_C1 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO11;
  assign CLBLM_R_X3Y99_SLICE_X3Y99_D1 = 1'b1;
  assign CLBLM_R_X3Y99_SLICE_X3Y99_D2 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X1Y91_A1 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X1Y91_A2 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X1Y91_A3 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X1Y91_A4 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X1Y91_A5 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X1Y91_A6 = 1'b1;
  assign CLBLM_R_X3Y99_SLICE_X3Y99_D3 = 1'b1;
  assign CLBLM_R_X3Y99_SLICE_X3Y99_D4 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X1Y91_AX = CLBLM_R_X3Y94_SLICE_X2Y94_DO6;
  assign CLBLM_R_X3Y99_SLICE_X3Y99_D5 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X1Y91_B1 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X1Y91_B2 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X1Y91_B3 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X1Y91_B4 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X1Y91_B5 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X1Y91_B6 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X1Y91_BX = CLBLL_L_X4Y92_SLICE_X4Y92_AO6;
  assign CLBLM_R_X3Y99_SLICE_X2Y99_A1 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLL_L_X2Y91_SLICE_X1Y91_C1 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X1Y91_C2 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X1Y91_C3 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X1Y91_C4 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X1Y91_C5 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X1Y91_C6 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X1Y91_CE = CLBLL_L_X2Y93_SLICE_X1Y93_CO6;
  assign CLBLM_R_X3Y99_SLICE_X2Y99_AX = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X2Y91_SLICE_X1Y91_CX = CLBLL_L_X4Y94_SLICE_X4Y94_CO5;
  assign CLBLL_L_X2Y91_SLICE_X1Y91_D1 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X1Y91_D2 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X1Y91_D3 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X1Y91_D4 = 1'b1;
  assign CLBLL_L_X2Y91_SLICE_X1Y91_D5 = 1'b1;
  assign CLBLM_R_X3Y99_SLICE_X2Y99_D1 = CLBLL_L_X4Y97_SLICE_X4Y97_AO6;
  assign CLBLM_R_X3Y99_SLICE_X2Y99_D2 = CLBLM_R_X3Y99_SLICE_X2Y99_AQ;
  assign CLBLM_R_X3Y99_SLICE_X2Y99_D3 = CLBLM_R_X3Y97_SLICE_X2Y97_BO6;
  assign CLBLM_R_X3Y99_SLICE_X2Y99_D4 = CLBLM_R_X3Y98_SLICE_X2Y98_DO6;
  assign CLBLM_R_X3Y99_SLICE_X2Y99_D5 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRL0 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRL1 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRL2 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRL3 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRL4 = CLBLM_R_X7Y99_SLICE_X8Y99_AQ;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRL5 = CLBLM_R_X5Y99_SLICE_X7Y99_AQ;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRL6 = CLBLM_R_X5Y99_SLICE_X6Y99_AQ;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRL7 = CLBLM_R_X5Y96_SLICE_X7Y96_AQ;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRL8 = CLBLM_R_X5Y96_SLICE_X7Y96_BQ;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRL9 = CLBLM_R_X5Y96_SLICE_X6Y96_AQ;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRL10 = CLBLM_R_X7Y96_SLICE_X8Y96_AQ;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRL11 = CLBLM_R_X7Y96_SLICE_X9Y96_AQ;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRL12 = CLBLM_R_X7Y98_SLICE_X9Y98_AQ;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRL13 = CLBLM_R_X7Y99_SLICE_X9Y99_AQ;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRL14 = CLBLM_R_X7Y97_SLICE_X8Y97_AQ;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRL15 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRU0 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRU1 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRU2 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRU3 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRU4 = CLBLM_R_X7Y99_SLICE_X8Y99_AQ;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRU5 = CLBLM_R_X5Y99_SLICE_X7Y99_AQ;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRU6 = CLBLM_R_X5Y99_SLICE_X6Y99_AQ;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRU7 = CLBLM_R_X5Y96_SLICE_X7Y96_AQ;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRU8 = CLBLM_R_X5Y96_SLICE_X7Y96_BQ;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRU9 = CLBLM_R_X5Y96_SLICE_X6Y96_AQ;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRU10 = CLBLM_R_X7Y96_SLICE_X8Y96_AQ;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRU11 = CLBLM_R_X7Y96_SLICE_X9Y96_AQ;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRU12 = CLBLM_R_X7Y98_SLICE_X9Y98_AQ;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRU13 = CLBLM_R_X7Y99_SLICE_X9Y99_AQ;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRARDADDRU14 = CLBLM_R_X7Y97_SLICE_X8Y97_AQ;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRL0 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRL1 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRL2 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRL3 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRL4 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRL5 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRL6 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRL7 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRL8 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRL9 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRL10 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRL11 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRL12 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRL13 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRL14 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRL15 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRU0 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRU1 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRU2 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRU3 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRU4 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRU5 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRU6 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRU7 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRU8 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRU9 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRU10 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRU11 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRU12 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRU13 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ADDRBWRADDRU14 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_CLKBWRCLKL = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_CLKBWRCLKU = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIADI0 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIADI2 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIADI4 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIADI6 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIADI8 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIADI10 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIADI12 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIADI14 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIADI16 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIADI18 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIADI20 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIADI22 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIADI24 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIADI26 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIADI28 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIADI30 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIADI1 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIADI3 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIADI5 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIADI7 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIADI9 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIADI11 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIADI13 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIADI15 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIADI17 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIADI19 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIADI21 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIADI23 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIADI25 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIADI27 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIADI29 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIADI31 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI0 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI2 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI4 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI6 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI8 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI10 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI12 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI14 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI16 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI18 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI20 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI22 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI24 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI26 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI28 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI30 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI1 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI3 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI5 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI7 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI9 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI11 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI13 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI15 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI17 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI19 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI21 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI23 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI25 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI27 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI29 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIBDI31 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIPADIP0 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIPADIP2 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIPADIP1 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIPADIP3 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIPBDIP0 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIPBDIP2 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIPBDIP1 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_DIPBDIP3 = 1'b1;
  assign CLBLL_L_X2Y92_SLICE_X0Y92_A1 = 1'b1;
  assign CLBLL_L_X2Y92_SLICE_X0Y92_A2 = 1'b1;
  assign CLBLL_L_X2Y92_SLICE_X0Y92_A3 = 1'b1;
  assign CLBLL_L_X2Y92_SLICE_X0Y92_A4 = 1'b1;
  assign CLBLL_L_X2Y92_SLICE_X0Y92_A5 = 1'b1;
  assign CLBLL_L_X2Y92_SLICE_X0Y92_A6 = 1'b1;
  assign CLBLM_R_X7Y94_SLICE_X9Y94_A1 = CLBLM_R_X7Y94_SLICE_X9Y94_DO6;
  assign CLBLM_R_X7Y94_SLICE_X9Y94_A2 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLL_L_X2Y92_SLICE_X0Y92_AX = CLBLL_L_X4Y94_SLICE_X4Y94_CO5;
  assign CLBLL_L_X2Y92_SLICE_X0Y92_B1 = 1'b1;
  assign CLBLL_L_X2Y92_SLICE_X0Y92_B2 = 1'b1;
  assign CLBLL_L_X2Y92_SLICE_X0Y92_B3 = 1'b1;
  assign CLBLL_L_X2Y92_SLICE_X0Y92_B4 = 1'b1;
  assign CLBLL_L_X2Y92_SLICE_X0Y92_B5 = 1'b1;
  assign CLBLL_L_X2Y92_SLICE_X0Y92_B6 = 1'b1;
  assign CLBLM_R_X7Y94_SLICE_X9Y94_B1 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLM_R_X7Y94_SLICE_X9Y94_B2 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X7Y94_SLICE_X9Y94_B3 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLL_L_X2Y92_SLICE_X0Y92_C1 = 1'b1;
  assign CLBLL_L_X2Y92_SLICE_X0Y92_C2 = 1'b1;
  assign CLBLL_L_X2Y92_SLICE_X0Y92_C3 = 1'b1;
  assign CLBLL_L_X2Y92_SLICE_X0Y92_C4 = 1'b1;
  assign CLBLL_L_X2Y92_SLICE_X0Y92_C5 = 1'b1;
  assign CLBLL_L_X2Y92_SLICE_X0Y92_C6 = 1'b1;
  assign CLBLL_L_X2Y92_SLICE_X0Y92_CE = CLBLL_L_X2Y93_SLICE_X0Y93_DO6;
  assign CLBLM_R_X7Y94_SLICE_X9Y94_C1 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X7Y94_SLICE_X9Y94_C2 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO11;
  assign CLBLM_R_X7Y94_SLICE_X9Y94_C3 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO15;
  assign CLBLM_R_X7Y94_SLICE_X9Y94_C4 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO13;
  assign CLBLM_R_X7Y94_SLICE_X9Y94_C6 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO12;
  assign CLBLL_L_X2Y92_SLICE_X0Y92_D1 = 1'b1;
  assign CLBLL_L_X2Y92_SLICE_X0Y92_D2 = 1'b1;
  assign CLBLL_L_X2Y92_SLICE_X0Y92_D3 = 1'b1;
  assign CLBLL_L_X2Y92_SLICE_X0Y92_D4 = 1'b1;
  assign CLBLL_L_X2Y92_SLICE_X0Y92_D5 = 1'b1;
  assign CLBLL_L_X2Y92_SLICE_X0Y92_D6 = 1'b1;
  assign CLBLM_R_X7Y94_SLICE_X9Y94_D1 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X7Y94_SLICE_X9Y94_D2 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO12;
  assign CLBLM_R_X7Y94_SLICE_X9Y94_D3 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO15;
  assign CLBLM_R_X7Y94_SLICE_X9Y94_D4 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO13;
  assign CLBLM_R_X7Y94_SLICE_X9Y94_D5 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO14;
  assign CLBLM_R_X7Y94_SLICE_X8Y94_A1 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ENARDENL = CLBLM_L_X8Y97_SLICE_X11Y97_CO6;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ENARDENU = CLBLM_L_X8Y97_SLICE_X11Y97_CO6;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ENBWRENL = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_ENBWRENU = 1'b1;
  assign CLBLM_R_X7Y94_SLICE_X8Y94_A2 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLM_R_X7Y94_SLICE_X8Y94_A3 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X7Y94_SLICE_X8Y94_A4 = CLBLM_R_X7Y94_SLICE_X8Y94_BO6;
  assign CLBLM_R_X7Y94_SLICE_X8Y94_A5 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X7Y94_SLICE_X8Y94_A6 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X7Y94_SLICE_X8Y94_B1 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO15;
  assign CLBLM_R_X7Y94_SLICE_X8Y94_B2 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO14;
  assign CLBLM_R_X7Y94_SLICE_X8Y94_B3 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X7Y94_SLICE_X8Y94_B4 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO11;
  assign CLBLM_R_X7Y94_SLICE_X8Y94_B5 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO12;
  assign CLBLM_R_X7Y94_SLICE_X8Y94_B6 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO13;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_D1 = CLBLM_R_X7Y91_SLICE_X8Y91_DO6;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_REGCEAREGCEL = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_REGCEAREGCEU = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_REGCEBL = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_REGCEBU = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_REGCLKARDRCLKL = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_REGCLKARDRCLKU = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_REGCLKBL = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_REGCLKBU = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_RSTRAMARSTRAMLRST = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_RSTRAMARSTRAMU = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_RSTRAMBL = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_RSTRAMBU = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_RSTREGARSTREGL = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_RSTREGARSTREGU = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_RSTREGBL = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_RSTREGBU = 1'b1;
  assign CLBLL_L_X2Y92_SLICE_X1Y92_AX = CLBLM_R_X3Y94_SLICE_X2Y94_DO6;
  assign CLBLL_L_X2Y92_SLICE_X1Y92_B1 = 1'b1;
  assign CLBLL_L_X2Y92_SLICE_X1Y92_B2 = 1'b1;
  assign CLBLL_L_X2Y92_SLICE_X1Y92_B3 = 1'b1;
  assign CLBLL_L_X2Y92_SLICE_X1Y92_B4 = 1'b1;
  assign CLBLL_L_X2Y92_SLICE_X1Y92_B6 = 1'b1;
  assign CLBLL_L_X2Y92_SLICE_X1Y92_BX = CLBLL_L_X4Y92_SLICE_X4Y92_AO6;
  assign CLBLL_L_X2Y92_SLICE_X1Y92_C1 = 1'b1;
  assign CLBLL_L_X2Y92_SLICE_X1Y92_C2 = 1'b1;
  assign CLBLL_L_X2Y92_SLICE_X1Y92_C3 = 1'b1;
  assign CLBLL_L_X2Y92_SLICE_X1Y92_C4 = 1'b1;
  assign CLBLL_L_X2Y92_SLICE_X1Y92_C5 = 1'b1;
  assign CLBLL_L_X2Y92_SLICE_X1Y92_C6 = 1'b1;
  assign CLBLL_L_X2Y92_SLICE_X1Y92_CE = CLBLL_L_X4Y92_SLICE_X4Y92_BO6;
  assign CLBLM_R_X7Y94_SLICE_X8Y94_SR = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X2Y92_SLICE_X1Y92_CX = CLBLL_L_X4Y94_SLICE_X4Y94_CO5;
  assign CLBLL_L_X2Y92_SLICE_X1Y92_D1 = 1'b1;
  assign CLBLL_L_X2Y92_SLICE_X1Y92_D2 = 1'b1;
  assign CLBLL_L_X2Y92_SLICE_X1Y92_D3 = 1'b1;
  assign CLBLL_L_X2Y92_SLICE_X1Y92_D4 = 1'b1;
  assign CLBLL_L_X2Y92_SLICE_X1Y92_D5 = 1'b1;
  assign CLBLL_L_X2Y92_SLICE_X1Y92_D6 = 1'b1;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_WEAL0 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_WEAL1 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_WEAL2 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_WEAL3 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_WEAU0 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_WEAU1 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_WEAU2 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_WEAU3 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_WEBWEL0 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_WEBWEL1 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_WEBWEL2 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_WEBWEL3 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_WEBWEL4 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_WEBWEL5 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_WEBWEL6 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_WEBWEL7 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_WEBWEU0 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_WEBWEU1 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_WEBWEU2 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_WEBWEU3 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_WEBWEU4 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_WEBWEU5 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_WEBWEU6 = 1'b0;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_WEBWEU7 = 1'b0;
  assign CLBLM_R_X7Y93_SLICE_X8Y93_B1 = 1'b1;
  assign CLBLL_L_X2Y93_SLICE_X0Y93_A1 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLL_L_X2Y93_SLICE_X0Y93_A2 = 1'b1;
  assign CLBLL_L_X2Y93_SLICE_X0Y93_A3 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLL_L_X2Y93_SLICE_X0Y93_A4 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO10;
  assign CLBLL_L_X2Y93_SLICE_X0Y93_A5 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLL_L_X2Y93_SLICE_X0Y93_A6 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X7Y94_SLICE_X8Y94_C1 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLL_L_X2Y93_SLICE_X0Y93_AX = CLBLL_L_X4Y91_SLICE_X5Y91_CO6;
  assign CLBLL_L_X2Y93_SLICE_X0Y93_B1 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLL_L_X2Y93_SLICE_X0Y93_B2 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLL_L_X2Y93_SLICE_X0Y93_B3 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLL_L_X2Y93_SLICE_X0Y93_B4 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLL_L_X2Y93_SLICE_X0Y93_B5 = CLBLM_R_X3Y93_SLICE_X2Y93_DO6;
  assign CLBLL_L_X2Y93_SLICE_X0Y93_B6 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO10;
  assign CLBLL_L_X2Y93_SLICE_X0Y93_BX = CLBLM_R_X3Y94_SLICE_X2Y94_DO6;
  assign CLBLL_L_X2Y93_SLICE_X0Y93_C1 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLL_L_X2Y93_SLICE_X0Y93_C2 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLL_L_X2Y93_SLICE_X0Y93_C3 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLL_L_X2Y93_SLICE_X0Y93_C4 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLL_L_X2Y93_SLICE_X0Y93_C5 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLL_L_X2Y93_SLICE_X0Y93_C6 = 1'b1;
  assign CLBLL_L_X2Y93_SLICE_X0Y93_CE = CLBLL_L_X2Y93_SLICE_X0Y93_DO6;
  assign CLBLM_R_X7Y93_SLICE_X8Y93_B2 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X7Y94_SLICE_X8Y94_C2 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLL_L_X2Y93_SLICE_X0Y93_CX = CLBLM_R_X3Y94_SLICE_X2Y94_DO5;
  assign CLBLL_L_X2Y93_SLICE_X0Y93_D1 = 1'b1;
  assign CLBLL_L_X2Y93_SLICE_X0Y93_D2 = CLBLM_R_X5Y94_SLICE_X7Y94_DO6;
  assign CLBLL_L_X2Y93_SLICE_X0Y93_D3 = CLBLL_L_X4Y94_SLICE_X5Y94_DO6;
  assign CLBLL_L_X2Y93_SLICE_X0Y93_D4 = CLBLL_L_X2Y93_SLICE_X0Y93_CO6;
  assign CLBLL_L_X2Y93_SLICE_X0Y93_D5 = CLBLM_R_X5Y94_SLICE_X6Y94_BO6;
  assign CLBLL_L_X2Y93_SLICE_X0Y93_D6 = 1'b1;
  assign CLBLM_R_X7Y93_SLICE_X8Y93_B3 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X7Y90_SLICE_X9Y90_A1 = CLBLM_R_X7Y91_SLICE_X9Y91_DO6;
  assign CLBLM_R_X7Y90_SLICE_X9Y90_A2 = CLBLM_R_X7Y91_SLICE_X9Y91_BQ;
  assign CLBLM_R_X7Y90_SLICE_X9Y90_A3 = CLBLM_R_X7Y90_SLICE_X9Y90_AQ;
  assign CLBLM_R_X7Y94_SLICE_X8Y94_C3 = 1'b1;
  assign CLBLM_R_X7Y90_SLICE_X9Y90_A4 = CLBLM_R_X7Y91_SLICE_X9Y91_CQ;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1 = CLBLM_R_X7Y91_SLICE_X8Y91_BO6;
  assign CLBLM_R_X7Y90_SLICE_X9Y90_A5 = CLBLM_R_X7Y90_SLICE_X9Y90_A5Q;
  assign CLBLL_L_X2Y93_SLICE_X1Y93_A1 = CLBLM_R_X5Y93_SLICE_X6Y93_F7AMUX_O;
  assign CLBLL_L_X2Y93_SLICE_X1Y93_A2 = CLBLL_L_X2Y93_SLICE_X1Y93_BQ;
  assign CLBLL_L_X2Y93_SLICE_X1Y93_A3 = CLBLL_L_X4Y91_SLICE_X5Y91_F7AMUX_O;
  assign CLBLL_L_X2Y93_SLICE_X1Y93_A4 = CLBLL_L_X2Y93_SLICE_X0Y93_BQ;
  assign CLBLL_L_X2Y93_SLICE_X1Y93_A5 = CLBLM_R_X3Y92_SLICE_X2Y92_BQ;
  assign CLBLL_L_X2Y93_SLICE_X1Y93_A6 = CLBLM_R_X3Y93_SLICE_X2Y93_BQ;
  assign CLBLM_R_X7Y90_SLICE_X9Y90_A6 = 1'b1;
  assign CLBLM_R_X7Y93_SLICE_X8Y93_B4 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLL_L_X2Y93_SLICE_X1Y93_AX = CLBLL_L_X2Y93_SLICE_X0Y93_F7AMUX_O;
  assign CLBLL_L_X2Y93_SLICE_X1Y93_B1 = CLBLL_L_X2Y94_SLICE_X1Y94_BQ;
  assign CLBLL_L_X2Y93_SLICE_X1Y93_B2 = CLBLL_L_X4Y91_SLICE_X5Y91_F7AMUX_O;
  assign CLBLL_L_X2Y92_SLICE_X1Y92_A1 = CLBLM_R_X5Y94_SLICE_X7Y94_DO6;
  assign CLBLL_L_X2Y93_SLICE_X1Y93_B3 = CLBLL_L_X2Y91_SLICE_X1Y91_AQ;
  assign CLBLL_L_X2Y93_SLICE_X1Y93_B4 = CLBLL_L_X2Y92_SLICE_X1Y92_AQ;
  assign CLBLL_L_X2Y93_SLICE_X1Y93_B5 = CLBLM_R_X3Y94_SLICE_X2Y94_AQ;
  assign CLBLL_L_X2Y93_SLICE_X1Y93_B6 = CLBLM_R_X5Y93_SLICE_X6Y93_F7AMUX_O;
  assign CLBLL_L_X2Y92_SLICE_X1Y92_A2 = 1'b1;
  assign CLBLL_L_X2Y93_SLICE_X1Y93_BX = CLBLM_R_X3Y94_SLICE_X2Y94_DO6;
  assign CLBLL_L_X2Y93_SLICE_X1Y93_C1 = 1'b1;
  assign CLBLL_L_X2Y93_SLICE_X1Y93_C2 = CLBLL_L_X2Y93_SLICE_X0Y93_CO6;
  assign CLBLL_L_X2Y93_SLICE_X1Y93_C3 = CLBLM_R_X5Y94_SLICE_X6Y94_BO6;
  assign CLBLL_L_X2Y92_SLICE_X1Y92_A3 = 1'b1;
  assign CLBLL_L_X2Y93_SLICE_X1Y93_C4 = CLBLM_R_X5Y94_SLICE_X7Y94_DO6;
  assign CLBLL_L_X2Y93_SLICE_X1Y93_C5 = CLBLL_L_X4Y94_SLICE_X5Y94_DO6;
  assign CLBLL_L_X2Y93_SLICE_X1Y93_C6 = 1'b1;
  assign CLBLL_L_X2Y93_SLICE_X1Y93_CE = CLBLL_L_X2Y93_SLICE_X1Y93_DO6;
  assign CLBLL_L_X2Y92_SLICE_X1Y92_A4 = CLBLM_R_X5Y94_SLICE_X6Y94_BO6;
  assign CLBLM_R_X7Y90_SLICE_X9Y90_B1 = CLBLM_R_X7Y91_SLICE_X9Y91_DO6;
  assign CLBLM_R_X7Y93_SLICE_X8Y93_B5 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLM_R_X7Y90_SLICE_X9Y90_B2 = CLBLM_R_X7Y90_SLICE_X9Y90_BQ;
  assign CLBLL_L_X2Y92_SLICE_X1Y92_A5 = CLBLL_L_X4Y94_SLICE_X5Y94_DO6;
  assign CLBLL_L_X2Y93_SLICE_X1Y93_D1 = 1'b1;
  assign CLBLL_L_X2Y93_SLICE_X1Y93_D2 = CLBLL_L_X2Y93_SLICE_X0Y93_CO6;
  assign CLBLL_L_X2Y93_SLICE_X1Y93_D3 = CLBLM_R_X5Y94_SLICE_X6Y94_BO6;
  assign CLBLL_L_X2Y92_SLICE_X1Y92_A6 = CLBLL_L_X2Y93_SLICE_X0Y93_CO6;
  assign CLBLL_L_X2Y93_SLICE_X1Y93_D4 = CLBLM_R_X5Y94_SLICE_X7Y94_DO6;
  assign CLBLL_L_X2Y93_SLICE_X1Y93_D5 = CLBLL_L_X4Y94_SLICE_X5Y94_DO6;
  assign CLBLL_L_X2Y93_SLICE_X1Y93_D6 = 1'b1;
  assign CLBLM_R_X7Y90_SLICE_X9Y90_B3 = CLBLM_R_X7Y90_SLICE_X9Y90_AQ;
  assign CLBLM_R_X7Y90_SLICE_X9Y90_B4 = CLBLM_R_X7Y91_SLICE_X9Y91_BQ;
  assign CLBLM_R_X7Y90_SLICE_X9Y90_B5 = CLBLM_R_X7Y90_SLICE_X9Y90_A5Q;
  assign CLBLM_R_X7Y90_SLICE_X9Y90_B6 = CLBLM_R_X7Y91_SLICE_X9Y91_CQ;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1 = 1'b1;
  assign CLBLM_R_X3Y99_SLICE_X3Y99_A1 = 1'b1;
  assign CLBLM_R_X3Y99_SLICE_X3Y99_A2 = 1'b1;
  assign CLBLM_R_X3Y99_SLICE_X3Y99_A3 = 1'b1;
  assign CLBLM_R_X3Y99_SLICE_X3Y99_A4 = 1'b1;
  assign CLBLM_R_X3Y99_SLICE_X3Y99_A5 = 1'b1;
  assign CLBLL_L_X2Y92_SLICE_X1Y92_B5 = 1'b1;
  assign CLBLM_R_X3Y99_SLICE_X3Y99_A6 = 1'b1;
  assign CLBLM_R_X5Y97_SLICE_X7Y97_D6 = CLBLM_R_X5Y98_SLICE_X6Y98_DO6;
  assign CLBLM_R_X7Y90_SLICE_X9Y90_C2 = CLBLM_R_X7Y90_SLICE_X9Y90_CQ;
  assign CLBLM_R_X7Y90_SLICE_X9Y90_C3 = CLBLM_R_X7Y91_SLICE_X8Y91_AQ;
  assign CLBLM_R_X7Y90_SLICE_X9Y90_C4 = CLBLM_R_X7Y87_SLICE_X8Y87_AQ;
  assign CLBLM_R_X7Y90_SLICE_X9Y90_C5 = CLBLM_R_X7Y90_SLICE_X9Y90_DO6;
  assign CLBLM_R_X7Y90_SLICE_X9Y90_C6 = CLBLM_R_X7Y87_SLICE_X8Y87_BQ;
  assign CLBLM_R_X3Y99_SLICE_X3Y99_B1 = 1'b1;
  assign CLBLM_R_X7Y90_SLICE_X9Y90_CLK = CLBLM_R_X7Y88_SLICE_X8Y88_AQ;
  assign CLBLM_R_X5Y97_SLICE_X6Y97_A4 = CLBLM_R_X7Y97_SLICE_X9Y97_B5Q;
  assign CLBLM_R_X5Y97_SLICE_X6Y97_A5 = 1'b0;
  assign CLBLM_R_X5Y97_SLICE_X6Y97_A6 = 1'b1;
  assign CLBLM_R_X7Y90_SLICE_X9Y90_D1 = CLBLM_R_X7Y90_SLICE_X9Y90_BQ;
  assign CLBLM_R_X7Y90_SLICE_X9Y90_D2 = CLBLM_R_X7Y91_SLICE_X9Y91_CQ;
  assign CLBLM_R_X7Y90_SLICE_X9Y90_D3 = 1'b1;
  assign CLBLM_R_X7Y90_SLICE_X9Y90_D4 = CLBLM_R_X7Y90_SLICE_X9Y90_A5Q;
  assign CLBLM_R_X7Y90_SLICE_X9Y90_D5 = CLBLM_R_X7Y90_SLICE_X9Y90_AQ;
  assign CLBLM_R_X7Y90_SLICE_X9Y90_D6 = CLBLM_R_X7Y91_SLICE_X9Y91_BQ;
  assign CLBLM_R_X7Y90_SLICE_X9Y90_SR = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y97_SLICE_X6Y97_B6 = 1'b1;
  assign CLBLM_R_X7Y90_SLICE_X8Y90_A1 = CLBLM_R_X7Y87_SLICE_X8Y87_BQ;
  assign CLBLM_R_X7Y90_SLICE_X8Y90_A2 = CLBLM_R_X7Y91_SLICE_X9Y91_AQ;
  assign CLBLM_R_X5Y97_SLICE_X6Y97_BX = CLBLM_R_X5Y96_SLICE_X6Y96_AQ;
  assign CLBLM_R_X7Y90_SLICE_X8Y90_A3 = CLBLM_R_X7Y87_SLICE_X8Y87_AQ;
  assign CLBLM_R_X7Y90_SLICE_X8Y90_A4 = CLBLM_R_X7Y90_SLICE_X9Y90_BQ;
  assign CLBLM_R_X7Y90_SLICE_X8Y90_A5 = CLBLM_R_X7Y90_SLICE_X9Y90_CQ;
  assign CLBLL_L_X2Y94_SLICE_X0Y94_A1 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLL_L_X2Y94_SLICE_X0Y94_A2 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLL_L_X2Y94_SLICE_X0Y94_A3 = CLBLL_L_X4Y95_SLICE_X4Y95_BO6;
  assign CLBLL_L_X2Y94_SLICE_X0Y94_A4 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLL_L_X2Y94_SLICE_X0Y94_A5 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLL_L_X2Y94_SLICE_X0Y94_A6 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X7Y90_SLICE_X8Y90_A6 = CLBLM_R_X7Y91_SLICE_X8Y91_AQ;
  assign CLBLL_L_X2Y94_SLICE_X0Y94_B1 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLL_L_X2Y94_SLICE_X0Y94_B2 = CLBLL_L_X4Y95_SLICE_X4Y95_CO6;
  assign CLBLL_L_X2Y94_SLICE_X0Y94_B3 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLL_L_X2Y94_SLICE_X0Y94_B4 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLL_L_X2Y94_SLICE_X0Y94_B5 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLL_L_X2Y94_SLICE_X0Y94_B6 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLM_R_X7Y96_SLICE_X9Y96_A1 = CLBLM_R_X7Y96_SLICE_X9Y96_DO6;
  assign CLBLM_R_X7Y96_SLICE_X9Y96_A2 = CLBLM_R_X7Y96_SLICE_X8Y96_BO5;
  assign CLBLM_R_X7Y96_SLICE_X9Y96_A3 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLL_L_X2Y94_SLICE_X0Y94_C1 = CLBLL_L_X2Y93_SLICE_X0Y93_CO5;
  assign CLBLL_L_X2Y94_SLICE_X0Y94_C2 = CLBLM_R_X3Y93_SLICE_X2Y93_CO5;
  assign CLBLL_L_X2Y94_SLICE_X0Y94_C3 = CLBLL_L_X2Y94_SLICE_X1Y94_B_XOR;
  assign CLBLL_L_X2Y94_SLICE_X0Y94_C4 = CLBLL_L_X2Y93_SLICE_X1Y93_F7AMUX_O;
  assign CLBLL_L_X2Y94_SLICE_X0Y94_C5 = CLBLL_L_X2Y97_SLICE_X0Y97_AO6;
  assign CLBLL_L_X2Y94_SLICE_X0Y94_C6 = CLBLL_L_X4Y95_SLICE_X4Y95_CO6;
  assign CLBLM_R_X3Y99_SLICE_X3Y99_D6 = 1'b1;
  assign CLBLM_R_X7Y96_SLICE_X9Y96_B1 = CLBLM_L_X8Y97_SLICE_X10Y97_CO6;
  assign CLBLM_R_X7Y96_SLICE_X9Y96_C1 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X7Y96_SLICE_X9Y96_C2 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO7;
  assign CLBLM_R_X7Y96_SLICE_X9Y96_C3 = CLBLM_L_X8Y97_SLICE_X11Y97_AO6;
  assign CLBLM_R_X7Y90_SLICE_X8Y90_B1 = CLBLM_R_X7Y89_SLICE_X9Y89_DO6;
  assign CLBLL_L_X2Y94_SLICE_X0Y94_D1 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLL_L_X2Y94_SLICE_X0Y94_D2 = 1'b1;
  assign CLBLL_L_X2Y94_SLICE_X0Y94_D3 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLL_L_X2Y94_SLICE_X0Y94_D4 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLL_L_X2Y94_SLICE_X0Y94_D5 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLL_L_X2Y94_SLICE_X0Y94_D6 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X7Y90_SLICE_X8Y90_B2 = CLBLM_R_X7Y89_SLICE_X9Y89_BQ;
  assign CLBLM_R_X7Y90_SLICE_X8Y90_B3 = CLBLM_R_X7Y89_SLICE_X8Y89_AQ;
  assign CLBLM_R_X7Y96_SLICE_X9Y96_CE = CLBLM_R_X7Y99_SLICE_X9Y99_DO6;
  assign CLBLM_R_X7Y96_SLICE_X9Y96_D1 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X7Y90_SLICE_X8Y90_B4 = CLBLM_R_X7Y89_SLICE_X8Y89_B5Q;
  assign CLBLM_R_X7Y96_SLICE_X9Y96_D2 = CLBLM_R_X5Y95_SLICE_X6Y95_AQ;
  assign CLBLM_R_X7Y96_SLICE_X9Y96_D3 = CLBLL_L_X4Y97_SLICE_X4Y97_BQ;
  assign CLBLM_R_X7Y96_SLICE_X9Y96_D4 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X7Y96_SLICE_X9Y96_D5 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X7Y90_SLICE_X8Y90_B5 = CLBLM_R_X7Y89_SLICE_X8Y89_BQ;
  assign CLBLM_R_X7Y96_SLICE_X9Y96_D6 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO7;
  assign CLBLM_R_X7Y96_SLICE_X9Y96_SR = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y96_SLICE_X8Y96_A1 = CLBLM_R_X7Y96_SLICE_X8Y96_DO6;
  assign CLBLM_R_X7Y90_SLICE_X8Y90_B6 = CLBLM_R_X7Y89_SLICE_X9Y89_AO5;
  assign CLBLM_R_X7Y96_SLICE_X8Y96_A2 = CLBLM_R_X7Y96_SLICE_X9Y96_BO6;
  assign CLBLM_R_X7Y96_SLICE_X8Y96_A3 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLM_R_X7Y96_SLICE_X8Y96_A4 = CLBLM_R_X7Y96_SLICE_X8Y96_BO6;
  assign CLBLM_R_X7Y96_SLICE_X8Y96_A5 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X7Y96_SLICE_X8Y96_A6 = CLBLM_R_X7Y98_SLICE_X8Y98_F7AMUX_O;
  assign CLBLM_R_X3Y99_SLICE_X2Y99_A2 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X7Y96_SLICE_X8Y96_B1 = CLBLM_R_X7Y96_SLICE_X9Y96_AQ;
  assign CLBLL_L_X2Y94_SLICE_X1Y94_A1 = 1'b1;
  assign CLBLL_L_X2Y94_SLICE_X1Y94_A2 = CLBLL_L_X2Y94_SLICE_X0Y94_DO6;
  assign CLBLL_L_X2Y94_SLICE_X1Y94_A3 = 1'b1;
  assign CLBLL_L_X2Y94_SLICE_X1Y94_A4 = 1'b1;
  assign CLBLL_L_X2Y94_SLICE_X1Y94_A5 = CLBLL_L_X2Y96_SLICE_X0Y96_AO6;
  assign CLBLL_L_X2Y94_SLICE_X1Y94_A6 = 1'b1;
  assign CLBLM_R_X3Y99_SLICE_X2Y99_A3 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X3Y99_SLICE_X2Y99_A4 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLL_L_X2Y94_SLICE_X1Y94_AX = CLBLL_L_X4Y93_SLICE_X4Y93_DO6;
  assign CLBLL_L_X2Y94_SLICE_X1Y94_B1 = CLBLM_R_X3Y94_SLICE_X2Y94_DO6;
  assign CLBLL_L_X2Y94_SLICE_X1Y94_B2 = CLBLL_L_X2Y97_SLICE_X0Y97_AO6;
  assign CLBLL_L_X2Y94_SLICE_X1Y94_B3 = CLBLM_R_X3Y93_SLICE_X2Y93_CO5;
  assign CLBLL_L_X2Y94_SLICE_X1Y94_B4 = CLBLL_L_X4Y95_SLICE_X4Y95_CO6;
  assign CLBLL_L_X2Y94_SLICE_X1Y94_B5 = CLBLL_L_X2Y93_SLICE_X1Y93_F7AMUX_O;
  assign CLBLL_L_X2Y94_SLICE_X1Y94_B6 = 1'b1;
  assign CLBLM_R_X3Y99_SLICE_X2Y99_A5 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X3Y99_SLICE_X2Y99_A6 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO0;
  assign CLBLL_L_X2Y94_SLICE_X1Y94_BX = CLBLL_L_X2Y94_SLICE_X0Y94_BO6;
  assign CLBLM_R_X7Y90_SLICE_X8Y90_C1 = CLBLM_R_X7Y91_SLICE_X9Y91_CQ;
  assign CLBLL_L_X2Y94_SLICE_X1Y94_C1 = CLBLM_R_X3Y94_SLICE_X2Y94_DO5;
  assign CLBLL_L_X2Y94_SLICE_X1Y94_C2 = CLBLM_R_X3Y94_SLICE_X3Y94_F7AMUX_O;
  assign CLBLL_L_X2Y94_SLICE_X1Y94_C3 = CLBLM_R_X3Y95_SLICE_X3Y95_DO6;
  assign CLBLL_L_X2Y94_SLICE_X1Y94_C4 = CLBLL_L_X2Y97_SLICE_X0Y97_AO6;
  assign CLBLL_L_X2Y94_SLICE_X1Y94_C5 = CLBLM_R_X3Y93_SLICE_X2Y93_CO5;
  assign CLBLL_L_X2Y94_SLICE_X1Y94_C6 = 1'b1;
  assign CLBLL_L_X2Y94_SLICE_X1Y94_CE = CLBLL_L_X2Y92_SLICE_X1Y92_AO6;
  assign CLBLM_R_X7Y90_SLICE_X8Y90_C2 = CLBLM_R_X7Y90_SLICE_X9Y90_A5Q;
  assign CLBLM_R_X7Y90_SLICE_X8Y90_C3 = CLBLM_R_X7Y91_SLICE_X9Y91_BQ;
  assign CLBLM_R_X7Y96_SLICE_X8Y96_D1 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO6;
  assign CLBLM_R_X7Y96_SLICE_X8Y96_D2 = CLBLM_R_X5Y95_SLICE_X6Y95_AQ;
  assign CLBLL_L_X2Y94_SLICE_X1Y94_CX = CLBLM_R_X3Y93_SLICE_X3Y93_AO6;
  assign CLBLM_R_X7Y90_SLICE_X8Y90_C4 = CLBLM_R_X7Y90_SLICE_X9Y90_CQ;
  assign CLBLL_L_X2Y94_SLICE_X1Y94_D1 = CLBLL_L_X4Y94_SLICE_X4Y94_CO5;
  assign CLBLL_L_X2Y94_SLICE_X1Y94_D2 = CLBLL_L_X2Y97_SLICE_X0Y97_AO6;
  assign CLBLL_L_X2Y94_SLICE_X1Y94_D3 = CLBLL_L_X4Y95_SLICE_X4Y95_BO6;
  assign CLBLL_L_X2Y94_SLICE_X1Y94_D4 = CLBLL_L_X4Y93_SLICE_X4Y93_F7AMUX_O;
  assign CLBLL_L_X2Y94_SLICE_X1Y94_D5 = CLBLM_R_X3Y93_SLICE_X2Y93_CO5;
  assign CLBLL_L_X2Y94_SLICE_X1Y94_D6 = 1'b1;
  assign CLBLM_R_X7Y96_SLICE_X8Y96_SR = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X2Y94_SLICE_X1Y94_DX = CLBLL_L_X2Y94_SLICE_X0Y94_AO6;
  assign CLBLM_R_X3Y99_SLICE_X2Y99_B1 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLM_R_X3Y99_SLICE_X2Y99_B2 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X3Y99_SLICE_X2Y99_B3 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X3Y99_SLICE_X2Y99_B4 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X3Y99_SLICE_X2Y99_B5 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO2;
  assign CLBLM_R_X3Y99_SLICE_X2Y99_B6 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X3Y99_SLICE_X2Y99_C1 = CLBLL_L_X4Y97_SLICE_X4Y97_AO6;
  assign CLBLM_R_X3Y99_SLICE_X2Y99_C2 = 1'b1;
  assign CLBLM_R_X7Y90_SLICE_X8Y90_D3 = CLBLM_R_X7Y91_SLICE_X9Y91_BQ;
  assign CLBLM_R_X3Y99_SLICE_X2Y99_C3 = CLBLM_R_X3Y97_SLICE_X2Y97_DO6;
  assign CLBLM_R_X7Y90_SLICE_X8Y90_D4 = CLBLM_R_X7Y90_SLICE_X9Y90_CQ;
  assign CLBLM_R_X3Y99_SLICE_X2Y99_C4 = CLBLM_R_X3Y99_SLICE_X2Y99_AO6;
  assign CLBLM_R_X7Y90_SLICE_X8Y90_D5 = CLBLM_R_X7Y90_SLICE_X9Y90_AQ;
  assign CLBLM_R_X3Y99_SLICE_X2Y99_C5 = CLBLL_L_X2Y99_SLICE_X0Y99_AQ;
  assign CLBLM_R_X7Y90_SLICE_X8Y90_D6 = CLBLM_R_X7Y90_SLICE_X9Y90_BQ;
  assign CLBLM_R_X3Y99_SLICE_X2Y99_C6 = CLBLM_R_X3Y98_SLICE_X2Y98_DO6;
  assign CLBLM_R_X3Y99_SLICE_X2Y99_CE = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y90_SLICE_X8Y90_SR = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y94_SLICE_X8Y94_D6 = 1'b1;
  assign CLBLM_R_X3Y99_SLICE_X2Y99_D6 = CLBLM_R_X3Y99_SLICE_X2Y99_BO6;
  assign CLBLM_R_X3Y99_SLICE_X2Y99_SR = CLBLL_L_X2Y98_SLICE_X1Y98_BO6;
  assign CLBLL_L_X2Y95_SLICE_X0Y95_A1 = CLBLL_L_X4Y95_SLICE_X4Y95_DO6;
  assign CLBLL_L_X2Y95_SLICE_X0Y95_A2 = CLBLL_L_X2Y93_SLICE_X1Y93_F7AMUX_O;
  assign CLBLL_L_X2Y95_SLICE_X0Y95_A3 = 1'b1;
  assign CLBLL_L_X2Y95_SLICE_X0Y95_A4 = CLBLL_L_X4Y95_SLICE_X4Y95_CO6;
  assign CLBLL_L_X2Y95_SLICE_X0Y95_A5 = CLBLL_L_X4Y93_SLICE_X4Y93_DO6;
  assign CLBLL_L_X2Y95_SLICE_X0Y95_A6 = 1'b1;
  assign CLBLM_R_X5Y95_SLICE_X6Y95_A5 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLL_L_X2Y95_SLICE_X0Y95_B1 = CLBLM_R_X3Y95_SLICE_X3Y95_DO6;
  assign CLBLL_L_X2Y95_SLICE_X0Y95_B2 = CLBLM_R_X3Y94_SLICE_X3Y94_F7AMUX_O;
  assign CLBLL_L_X2Y95_SLICE_X0Y95_B3 = 1'b1;
  assign CLBLL_L_X2Y95_SLICE_X0Y95_B4 = CLBLL_L_X4Y93_SLICE_X4Y93_F7AMUX_O;
  assign CLBLL_L_X2Y95_SLICE_X0Y95_B5 = CLBLL_L_X4Y95_SLICE_X4Y95_BO6;
  assign CLBLL_L_X2Y95_SLICE_X0Y95_B6 = 1'b1;
  assign CLBLM_R_X7Y97_SLICE_X9Y97_A1 = CLBLM_R_X7Y97_SLICE_X9Y97_DO6;
  assign CLBLM_R_X7Y97_SLICE_X9Y97_A2 = CLBLM_R_X7Y97_SLICE_X9Y97_BQ;
  assign CLBLM_R_X7Y97_SLICE_X9Y97_A3 = CLBLM_R_X7Y97_SLICE_X9Y97_AQ;
  assign CLBLM_R_X7Y97_SLICE_X9Y97_A4 = CLBLM_R_X7Y97_SLICE_X9Y97_B5Q;
  assign CLBLL_L_X2Y95_SLICE_X0Y95_C1 = CLBLL_L_X4Y91_SLICE_X4Y91_BO6;
  assign CLBLL_L_X2Y95_SLICE_X0Y95_C2 = CLBLM_R_X3Y91_SLICE_X2Y91_F7AMUX_O;
  assign CLBLL_L_X2Y95_SLICE_X0Y95_C3 = CLBLM_R_X3Y91_SLICE_X3Y91_F7AMUX_O;
  assign CLBLL_L_X2Y95_SLICE_X0Y95_C4 = CLBLM_R_X3Y95_SLICE_X3Y95_AO6;
  assign CLBLL_L_X2Y95_SLICE_X0Y95_C5 = 1'b1;
  assign CLBLL_L_X2Y95_SLICE_X0Y95_C6 = 1'b1;
  assign CLBLM_R_X5Y95_SLICE_X6Y95_A6 = CLBLL_L_X2Y95_SLICE_X0Y95_D_CY;
  assign CLBLM_R_X7Y97_SLICE_X9Y97_A5 = CLBLM_R_X7Y97_SLICE_X9Y97_A5Q;
  assign CLBLM_R_X7Y97_SLICE_X9Y97_A6 = 1'b1;
  assign CLBLM_R_X7Y97_SLICE_X9Y97_B1 = CLBLM_R_X7Y97_SLICE_X9Y97_DO6;
  assign CLBLM_R_X7Y97_SLICE_X9Y97_B2 = CLBLM_R_X7Y97_SLICE_X9Y97_BQ;
  assign CLBLM_R_X7Y97_SLICE_X9Y97_B3 = CLBLM_R_X7Y97_SLICE_X9Y97_AQ;
  assign CLBLM_R_X7Y97_SLICE_X9Y97_B4 = CLBLM_R_X7Y97_SLICE_X9Y97_B5Q;
  assign CLBLM_R_X7Y97_SLICE_X9Y97_B5 = CLBLM_R_X7Y97_SLICE_X9Y97_A5Q;
  assign CLBLL_L_X2Y95_SLICE_X0Y95_D1 = 1'b1;
  assign CLBLL_L_X2Y95_SLICE_X0Y95_D2 = CLBLM_R_X3Y95_SLICE_X3Y95_BO6;
  assign CLBLL_L_X2Y95_SLICE_X0Y95_D3 = CLBLL_L_X4Y95_SLICE_X5Y95_CO6;
  assign CLBLL_L_X2Y95_SLICE_X0Y95_D4 = CLBLL_L_X4Y94_SLICE_X5Y94_F7AMUX_O;
  assign CLBLL_L_X2Y95_SLICE_X0Y95_D5 = CLBLM_R_X3Y92_SLICE_X2Y92_F7AMUX_O;
  assign CLBLL_L_X2Y95_SLICE_X0Y95_D6 = 1'b1;
  assign CLBLM_R_X7Y97_SLICE_X9Y97_C1 = CLBLM_R_X5Y95_SLICE_X6Y95_BO5;
  assign CLBLM_R_X7Y97_SLICE_X9Y97_C2 = CLBLL_L_X4Y97_SLICE_X5Y97_DO6;
  assign CLBLM_R_X7Y97_SLICE_X9Y97_C3 = CLBLM_R_X7Y97_SLICE_X9Y97_BQ;
  assign CLBLM_R_X7Y97_SLICE_X9Y97_C4 = CLBLM_R_X7Y97_SLICE_X9Y97_A5Q;
  assign CLBLM_R_X7Y97_SLICE_X9Y97_C5 = CLBLM_R_X7Y97_SLICE_X9Y97_B5Q;
  assign CLBLM_R_X7Y97_SLICE_X9Y97_C6 = CLBLM_R_X7Y97_SLICE_X9Y97_AQ;
  assign CLBLM_R_X7Y97_SLICE_X9Y97_CE = CLBLM_R_X7Y97_SLICE_X9Y97_CO6;
  assign CLBLM_R_X7Y97_SLICE_X9Y97_D1 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLM_R_X7Y97_SLICE_X9Y97_D2 = CLBLM_R_X5Y95_SLICE_X6Y95_CO6;
  assign CLBLM_R_X7Y97_SLICE_X9Y97_D3 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X7Y97_SLICE_X9Y97_D4 = CLBLL_L_X4Y97_SLICE_X5Y97_DO6;
  assign CLBLM_R_X7Y97_SLICE_X9Y97_D5 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X7Y97_SLICE_X9Y97_D6 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_D = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y97_SLICE_X9Y97_SR = LIOB33_X0Y107_IOB_X0Y107_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_D = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X7Y97_SLICE_X8Y97_A1 = CLBLM_R_X7Y98_SLICE_X8Y98_CO6;
  assign CLBLM_R_X7Y97_SLICE_X8Y97_A2 = CLBLM_R_X7Y98_SLICE_X8Y98_F7AMUX_O;
  assign CLBLM_R_X7Y97_SLICE_X8Y97_A3 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLM_R_X7Y97_SLICE_X8Y97_A4 = CLBLM_R_X7Y97_SLICE_X8Y97_DO6;
  assign CLBLM_R_X7Y97_SLICE_X8Y97_A5 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X7Y97_SLICE_X8Y97_A6 = CLBLM_R_X7Y97_SLICE_X8Y97_CO6;
  assign CLBLL_L_X2Y95_SLICE_X1Y95_A1 = 1'b1;
  assign CLBLL_L_X2Y95_SLICE_X1Y95_A2 = CLBLM_R_X3Y93_SLICE_X2Y93_CO5;
  assign CLBLL_L_X2Y95_SLICE_X1Y95_A3 = CLBLM_R_X3Y95_SLICE_X3Y95_AO6;
  assign CLBLL_L_X2Y95_SLICE_X1Y95_A4 = CLBLM_R_X3Y91_SLICE_X2Y91_F7AMUX_O;
  assign CLBLL_L_X2Y95_SLICE_X1Y95_A5 = CLBLL_L_X2Y97_SLICE_X0Y97_AO6;
  assign CLBLL_L_X2Y95_SLICE_X1Y95_A6 = 1'b1;
  assign CLBLM_R_X7Y97_SLICE_X8Y97_B1 = CLBLM_R_X7Y96_SLICE_X9Y96_AQ;
  assign CLBLL_L_X2Y95_SLICE_X1Y95_AX = CLBLM_R_X3Y95_SLICE_X3Y95_CO6;
  assign CLBLM_R_X7Y97_SLICE_X8Y97_B2 = CLBLM_R_X7Y96_SLICE_X8Y96_CO6;
  assign CLBLL_L_X2Y95_SLICE_X1Y95_B1 = CLBLM_R_X3Y91_SLICE_X3Y91_F7AMUX_O;
  assign CLBLL_L_X2Y95_SLICE_X1Y95_B2 = CLBLM_R_X3Y93_SLICE_X2Y93_CO5;
  assign CLBLL_L_X2Y95_SLICE_X1Y95_B3 = CLBLL_L_X4Y91_SLICE_X4Y91_BO6;
  assign CLBLL_L_X2Y95_SLICE_X1Y95_B4 = 1'b1;
  assign CLBLL_L_X2Y95_SLICE_X1Y95_B5 = CLBLL_L_X2Y97_SLICE_X0Y97_AO6;
  assign CLBLL_L_X2Y95_SLICE_X1Y95_B6 = 1'b1;
  assign CLBLM_R_X7Y93_SLICE_X8Y93_D2 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X7Y97_SLICE_X8Y97_B5 = CLBLM_R_X7Y96_SLICE_X8Y96_AQ;
  assign CLBLL_L_X2Y95_SLICE_X1Y95_BX = CLBLM_R_X3Y95_SLICE_X2Y95_AO6;
  assign CLBLL_L_X2Y95_SLICE_X1Y95_C1 = CLBLL_L_X2Y97_SLICE_X0Y97_AO6;
  assign CLBLL_L_X2Y95_SLICE_X1Y95_C2 = CLBLL_L_X4Y94_SLICE_X5Y94_F7AMUX_O;
  assign CLBLL_L_X2Y95_SLICE_X1Y95_C3 = CLBLM_R_X3Y93_SLICE_X2Y93_CO5;
  assign CLBLL_L_X2Y95_SLICE_X1Y95_C4 = CLBLL_L_X4Y95_SLICE_X5Y95_CO6;
  assign CLBLL_L_X2Y95_SLICE_X1Y95_C5 = 1'b1;
  assign CLBLL_L_X2Y95_SLICE_X1Y95_C6 = 1'b1;
  assign CLBLM_R_X7Y97_SLICE_X8Y97_C3 = CLBLM_R_X7Y98_SLICE_X8Y98_DO6;
  assign CLBLL_L_X2Y95_SLICE_X1Y95_CIN = CLBLL_L_X2Y94_SLICE_X1Y94_D_CY;
  assign CLBLM_R_X7Y97_SLICE_X8Y97_C5 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X7Y97_SLICE_X8Y97_C6 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X7Y97_SLICE_X8Y97_CE = CLBLM_R_X7Y99_SLICE_X9Y99_DO6;
  assign CLBLM_R_X7Y97_SLICE_X8Y97_D2 = CLBLM_R_X7Y97_SLICE_X8Y97_AQ;
  assign CLBLL_L_X2Y95_SLICE_X1Y95_CX = CLBLL_L_X4Y95_SLICE_X4Y95_AO6;
  assign CLBLM_R_X7Y97_SLICE_X8Y97_D3 = CLBLM_R_X7Y96_SLICE_X8Y96_AQ;
  assign CLBLL_L_X2Y95_SLICE_X1Y95_D1 = 1'b1;
  assign CLBLL_L_X2Y95_SLICE_X1Y95_D2 = CLBLM_R_X3Y95_SLICE_X3Y95_BO6;
  assign CLBLL_L_X2Y95_SLICE_X1Y95_D3 = CLBLM_R_X3Y93_SLICE_X2Y93_CO5;
  assign CLBLL_L_X2Y95_SLICE_X1Y95_D4 = CLBLL_L_X2Y97_SLICE_X0Y97_AO6;
  assign CLBLL_L_X2Y95_SLICE_X1Y95_D5 = 1'b1;
  assign CLBLL_L_X2Y95_SLICE_X1Y95_D6 = CLBLM_R_X3Y92_SLICE_X2Y92_F7AMUX_O;
  assign CLBLM_R_X7Y93_SLICE_X8Y93_D6 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO14;
  assign CLBLM_R_X5Y95_SLICE_X6Y95_B3 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X5Y95_SLICE_X6Y95_B4 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X5Y95_SLICE_X6Y95_B5 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X5Y95_SLICE_X6Y95_B6 = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_D1 = CLBLL_L_X2Y102_SLICE_X0Y102_AQ;
  assign CLBLM_R_X7Y93_SLICE_X8Y93_SR = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X2Y96_SLICE_X0Y96_A1 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLL_L_X2Y96_SLICE_X0Y96_A2 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLL_L_X2Y96_SLICE_X0Y96_A3 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLL_L_X2Y96_SLICE_X0Y96_A4 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLL_L_X2Y96_SLICE_X0Y96_A5 = CLBLL_L_X4Y95_SLICE_X4Y95_DO6;
  assign CLBLL_L_X2Y96_SLICE_X0Y96_A6 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLL_L_X2Y96_SLICE_X0Y96_B1 = CLBLL_L_X2Y93_SLICE_X0Y93_CO5;
  assign CLBLL_L_X2Y96_SLICE_X0Y96_B2 = CLBLM_R_X3Y92_SLICE_X2Y92_F7AMUX_O;
  assign CLBLL_L_X2Y96_SLICE_X0Y96_B3 = CLBLM_R_X3Y95_SLICE_X3Y95_BO6;
  assign CLBLL_L_X2Y96_SLICE_X0Y96_B4 = CLBLL_L_X2Y97_SLICE_X0Y97_AO6;
  assign CLBLL_L_X2Y96_SLICE_X0Y96_B5 = CLBLL_L_X2Y95_SLICE_X1Y95_D_XOR;
  assign CLBLL_L_X2Y96_SLICE_X0Y96_B6 = CLBLM_R_X3Y93_SLICE_X2Y93_CO5;
  assign CLBLL_L_X2Y96_SLICE_X0Y96_C1 = CLBLL_L_X4Y95_SLICE_X4Y95_DO6;
  assign CLBLL_L_X2Y96_SLICE_X0Y96_C2 = CLBLL_L_X2Y93_SLICE_X0Y93_CO5;
  assign CLBLL_L_X2Y96_SLICE_X0Y96_C3 = CLBLL_L_X4Y93_SLICE_X4Y93_DO6;
  assign CLBLL_L_X2Y96_SLICE_X0Y96_C4 = CLBLM_R_X3Y93_SLICE_X2Y93_CO5;
  assign CLBLL_L_X2Y96_SLICE_X0Y96_C5 = CLBLL_L_X2Y97_SLICE_X0Y97_AO6;
  assign CLBLL_L_X2Y96_SLICE_X0Y96_C6 = CLBLL_L_X2Y94_SLICE_X1Y94_A_XOR;
  assign CLBLM_R_X7Y98_SLICE_X9Y98_A1 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLM_R_X7Y98_SLICE_X9Y98_A2 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X7Y98_SLICE_X9Y98_A3 = CLBLM_R_X7Y98_SLICE_X8Y98_F7AMUX_O;
  assign CLBLM_R_X7Y98_SLICE_X9Y98_A4 = CLBLM_R_X7Y98_SLICE_X9Y98_BO6;
  assign CLBLM_R_X7Y98_SLICE_X9Y98_A5 = CLBLM_R_X7Y97_SLICE_X8Y97_BO6;
  assign CLBLM_R_X7Y98_SLICE_X9Y98_A6 = CLBLM_R_X7Y98_SLICE_X9Y98_CO6;
  assign CLBLM_R_X7Y98_SLICE_X9Y98_B1 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLL_L_X2Y96_SLICE_X0Y96_D1 = CLBLL_L_X2Y97_SLICE_X0Y97_AO6;
  assign CLBLL_L_X2Y96_SLICE_X0Y96_D2 = CLBLM_R_X3Y95_SLICE_X3Y95_DO6;
  assign CLBLL_L_X2Y96_SLICE_X0Y96_D3 = CLBLL_L_X2Y93_SLICE_X0Y93_CO5;
  assign CLBLL_L_X2Y96_SLICE_X0Y96_D4 = CLBLM_R_X3Y93_SLICE_X2Y93_CO5;
  assign CLBLL_L_X2Y96_SLICE_X0Y96_D5 = CLBLL_L_X2Y94_SLICE_X1Y94_C_XOR;
  assign CLBLL_L_X2Y96_SLICE_X0Y96_D6 = CLBLM_R_X3Y94_SLICE_X3Y94_F7AMUX_O;
  assign CLBLM_R_X7Y98_SLICE_X9Y98_B3 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X7Y98_SLICE_X9Y98_B4 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X7Y98_SLICE_X9Y98_B6 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO8;
  assign CLBLM_R_X7Y98_SLICE_X9Y98_C1 = CLBLL_L_X4Y97_SLICE_X4Y97_BQ;
  assign CLBLM_R_X7Y98_SLICE_X9Y98_C2 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X7Y98_SLICE_X9Y98_C3 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X7Y98_SLICE_X9Y98_C4 = CLBLM_R_X5Y95_SLICE_X6Y95_AQ;
  assign CLBLM_R_X7Y98_SLICE_X9Y98_C5 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO8;
  assign CLBLM_R_X7Y98_SLICE_X9Y98_C6 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X7Y98_SLICE_X9Y98_CE = CLBLM_R_X7Y99_SLICE_X9Y99_DO6;
  assign CLBLM_R_X7Y98_SLICE_X9Y98_D1 = 1'b1;
  assign CLBLM_R_X7Y98_SLICE_X9Y98_D2 = 1'b1;
  assign CLBLM_R_X7Y98_SLICE_X9Y98_D3 = 1'b1;
  assign CLBLM_R_X7Y98_SLICE_X9Y98_D4 = 1'b1;
  assign CLBLM_R_X7Y98_SLICE_X9Y98_D5 = 1'b1;
  assign CLBLM_R_X7Y98_SLICE_X9Y98_D6 = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_T1 = 1'b1;
  assign CLBLM_R_X7Y98_SLICE_X9Y98_SR = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y98_SLICE_X8Y98_A1 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X7Y98_SLICE_X8Y98_A2 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLL_L_X2Y96_SLICE_X1Y96_A1 = CLBLM_R_X3Y96_SLICE_X3Y96_BO5;
  assign CLBLL_L_X2Y96_SLICE_X1Y96_A2 = CLBLM_R_X3Y95_SLICE_X2Y95_CO6;
  assign CLBLL_L_X2Y96_SLICE_X1Y96_A3 = CLBLM_R_X3Y95_SLICE_X2Y95_DO6;
  assign CLBLL_L_X2Y96_SLICE_X1Y96_A4 = CLBLM_R_X3Y95_SLICE_X2Y95_BO6;
  assign CLBLL_L_X2Y96_SLICE_X1Y96_A5 = CLBLL_L_X2Y97_SLICE_X0Y97_AO5;
  assign CLBLL_L_X2Y96_SLICE_X1Y96_A6 = CLBLM_R_X3Y96_SLICE_X3Y96_BO6;
  assign CLBLM_R_X7Y98_SLICE_X8Y98_A3 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X7Y98_SLICE_X8Y98_A4 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X7Y98_SLICE_X8Y98_A5 = CLBLL_L_X4Y97_SLICE_X4Y97_BQ;
  assign CLBLL_L_X2Y96_SLICE_X1Y96_B1 = CLBLM_R_X3Y96_SLICE_X3Y96_BO5;
  assign CLBLL_L_X2Y96_SLICE_X1Y96_B2 = CLBLM_R_X3Y95_SLICE_X2Y95_CO6;
  assign CLBLL_L_X2Y96_SLICE_X1Y96_B3 = CLBLM_R_X3Y95_SLICE_X2Y95_DO6;
  assign CLBLL_L_X2Y96_SLICE_X1Y96_B4 = CLBLL_L_X2Y97_SLICE_X0Y97_AO5;
  assign CLBLL_L_X2Y96_SLICE_X1Y96_B5 = CLBLM_R_X3Y96_SLICE_X3Y96_BO6;
  assign CLBLL_L_X2Y96_SLICE_X1Y96_B6 = CLBLL_L_X2Y96_SLICE_X1Y96_CO6;
  assign CLBLM_R_X7Y98_SLICE_X8Y98_AX = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLM_R_X7Y98_SLICE_X8Y98_B1 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X7Y98_SLICE_X8Y98_B2 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLL_L_X2Y96_SLICE_X1Y96_C1 = CLBLL_L_X2Y95_SLICE_X1Y95_C_XOR;
  assign CLBLL_L_X2Y96_SLICE_X1Y96_C2 = CLBLL_L_X4Y95_SLICE_X5Y95_CO6;
  assign CLBLL_L_X2Y96_SLICE_X1Y96_C3 = CLBLL_L_X2Y97_SLICE_X0Y97_AO6;
  assign CLBLL_L_X2Y96_SLICE_X1Y96_C4 = CLBLL_L_X4Y94_SLICE_X5Y94_F7AMUX_O;
  assign CLBLL_L_X2Y96_SLICE_X1Y96_C5 = CLBLL_L_X2Y93_SLICE_X0Y93_CO5;
  assign CLBLL_L_X2Y96_SLICE_X1Y96_C6 = CLBLM_R_X3Y93_SLICE_X2Y93_CO5;
  assign CLBLM_R_X7Y98_SLICE_X8Y98_C1 = CLBLL_L_X4Y97_SLICE_X4Y97_BQ;
  assign CLBLM_R_X7Y98_SLICE_X8Y98_C2 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO10;
  assign CLBLM_R_X7Y98_SLICE_X8Y98_C3 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X7Y98_SLICE_X8Y98_C4 = CLBLM_R_X5Y95_SLICE_X6Y95_AQ;
  assign CLBLM_R_X7Y98_SLICE_X8Y98_C5 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X7Y98_SLICE_X8Y98_C6 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLL_L_X2Y96_SLICE_X1Y96_D1 = CLBLM_R_X3Y96_SLICE_X3Y96_BO5;
  assign CLBLL_L_X2Y96_SLICE_X1Y96_D2 = CLBLM_R_X3Y96_SLICE_X3Y96_BO6;
  assign CLBLL_L_X2Y96_SLICE_X1Y96_D3 = CLBLL_L_X2Y96_SLICE_X0Y96_BO6;
  assign CLBLL_L_X2Y96_SLICE_X1Y96_D4 = CLBLL_L_X2Y96_SLICE_X1Y96_CO6;
  assign CLBLL_L_X2Y96_SLICE_X1Y96_D5 = CLBLL_L_X2Y96_SLICE_X0Y96_CO6;
  assign CLBLL_L_X2Y96_SLICE_X1Y96_D6 = CLBLL_L_X2Y97_SLICE_X0Y97_AO5;
  assign CLBLM_R_X7Y98_SLICE_X8Y98_D1 = CLBLL_L_X4Y97_SLICE_X4Y97_BQ;
  assign CLBLM_R_X7Y98_SLICE_X8Y98_D2 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO10;
  assign CLBLM_R_X7Y98_SLICE_X8Y98_D3 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X7Y98_SLICE_X8Y98_D4 = CLBLM_L_X8Y98_SLICE_X10Y98_BO6;
  assign CLBLM_R_X7Y98_SLICE_X8Y98_D5 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X7Y98_SLICE_X8Y98_D6 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_T1 = 1'b1;
  assign CLBLM_R_X5Y90_SLICE_X7Y90_C4 = 1'b1;
  assign CLBLL_L_X2Y97_SLICE_X0Y97_A1 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLL_L_X2Y97_SLICE_X0Y97_A2 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLL_L_X2Y97_SLICE_X0Y97_A3 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLL_L_X2Y97_SLICE_X0Y97_A4 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLL_L_X2Y97_SLICE_X0Y97_A5 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLL_L_X2Y97_SLICE_X0Y97_A6 = 1'b1;
  assign CLBLL_L_X2Y97_SLICE_X0Y97_B1 = CLBLL_L_X2Y96_SLICE_X0Y96_CO6;
  assign CLBLL_L_X2Y97_SLICE_X0Y97_B2 = CLBLM_R_X3Y96_SLICE_X3Y96_BO6;
  assign CLBLL_L_X2Y97_SLICE_X0Y97_B3 = CLBLL_L_X2Y94_SLICE_X0Y94_CO6;
  assign CLBLL_L_X2Y97_SLICE_X0Y97_B4 = CLBLL_L_X2Y96_SLICE_X0Y96_BO6;
  assign CLBLL_L_X2Y97_SLICE_X0Y97_B5 = CLBLM_R_X3Y96_SLICE_X3Y96_BO5;
  assign CLBLL_L_X2Y97_SLICE_X0Y97_B6 = CLBLL_L_X2Y97_SLICE_X0Y97_AO5;
  assign CLBLM_R_X5Y90_SLICE_X7Y90_C5 = 1'b1;
  assign CLBLL_L_X2Y97_SLICE_X0Y97_C1 = CLBLL_L_X2Y97_SLICE_X0Y97_AO5;
  assign CLBLL_L_X2Y97_SLICE_X0Y97_C2 = CLBLL_L_X2Y94_SLICE_X0Y94_CO6;
  assign CLBLL_L_X2Y97_SLICE_X0Y97_C3 = CLBLM_R_X3Y96_SLICE_X3Y96_BO5;
  assign CLBLL_L_X2Y97_SLICE_X0Y97_C4 = CLBLL_L_X2Y96_SLICE_X0Y96_DO6;
  assign CLBLL_L_X2Y97_SLICE_X0Y97_C5 = CLBLM_R_X3Y96_SLICE_X3Y96_BO6;
  assign CLBLL_L_X2Y97_SLICE_X0Y97_C6 = CLBLM_R_X3Y95_SLICE_X2Y95_BO6;
  assign CLBLM_R_X7Y99_SLICE_X9Y99_A1 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLM_R_X7Y99_SLICE_X9Y99_A2 = CLBLM_R_X7Y97_SLICE_X8Y97_BO5;
  assign CLBLM_R_X7Y99_SLICE_X9Y99_A3 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X7Y99_SLICE_X9Y99_A4 = CLBLM_R_X7Y99_SLICE_X9Y99_BO6;
  assign CLBLM_R_X7Y99_SLICE_X9Y99_A5 = CLBLM_R_X7Y98_SLICE_X8Y98_F7AMUX_O;
  assign CLBLM_R_X7Y99_SLICE_X9Y99_A6 = CLBLM_R_X7Y99_SLICE_X9Y99_CO6;
  assign CLBLL_L_X2Y97_SLICE_X0Y97_D1 = CLBLL_L_X2Y94_SLICE_X0Y94_CO6;
  assign CLBLL_L_X2Y97_SLICE_X0Y97_D2 = CLBLL_L_X2Y96_SLICE_X0Y96_CO6;
  assign CLBLL_L_X2Y97_SLICE_X0Y97_D3 = 1'b1;
  assign CLBLL_L_X2Y97_SLICE_X0Y97_D5 = 1'b1;
  assign CLBLL_L_X2Y97_SLICE_X0Y97_D6 = CLBLM_R_X3Y95_SLICE_X2Y95_BO6;
  assign CLBLL_L_X2Y97_SLICE_X0Y97_D4 = CLBLL_L_X2Y96_SLICE_X0Y96_DO6;
  assign CLBLM_R_X5Y90_SLICE_X7Y90_C6 = CLBLL_L_X2Y97_SLICE_X0Y97_CO6;
  assign CLBLM_R_X7Y99_SLICE_X9Y99_B2 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO9;
  assign CLBLM_R_X7Y99_SLICE_X9Y99_B3 = CLBLM_L_X8Y98_SLICE_X10Y98_DO6;
  assign CLBLM_R_X7Y99_SLICE_X9Y99_B4 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X7Y99_SLICE_X9Y99_B6 = CLBLM_R_X5Y95_SLICE_X6Y95_AQ;
  assign CLBLM_R_X7Y99_SLICE_X9Y99_C1 = CLBLL_L_X4Y97_SLICE_X4Y97_BQ;
  assign CLBLM_R_X7Y99_SLICE_X9Y99_C2 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO9;
  assign CLBLM_R_X7Y99_SLICE_X9Y99_C3 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X7Y99_SLICE_X9Y99_C4 = CLBLM_R_X5Y95_SLICE_X6Y95_AQ;
  assign CLBLM_R_X7Y99_SLICE_X9Y99_C5 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X7Y99_SLICE_X9Y99_C6 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X7Y99_SLICE_X9Y99_CE = CLBLM_R_X7Y99_SLICE_X9Y99_DO6;
  assign CLBLM_R_X7Y99_SLICE_X9Y99_D1 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X7Y99_SLICE_X9Y99_D2 = 1'b1;
  assign CLBLM_R_X7Y99_SLICE_X9Y99_D3 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLM_R_X7Y99_SLICE_X9Y99_D4 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X7Y99_SLICE_X9Y99_D5 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X7Y99_SLICE_X9Y99_D6 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X7Y99_SLICE_X9Y99_SR = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X2Y97_SLICE_X1Y97_A1 = CLBLL_L_X2Y96_SLICE_X0Y96_CO6;
  assign CLBLL_L_X2Y97_SLICE_X1Y97_A2 = CLBLL_L_X2Y96_SLICE_X0Y96_DO6;
  assign CLBLL_L_X2Y97_SLICE_X1Y97_A3 = CLBLL_L_X2Y97_SLICE_X0Y97_AO5;
  assign CLBLL_L_X2Y97_SLICE_X1Y97_A4 = CLBLM_R_X3Y96_SLICE_X3Y96_BO6;
  assign CLBLL_L_X2Y97_SLICE_X1Y97_A5 = CLBLL_L_X2Y94_SLICE_X0Y94_CO6;
  assign CLBLL_L_X2Y97_SLICE_X1Y97_A6 = CLBLM_R_X3Y96_SLICE_X3Y96_BO5;
  assign CLBLM_R_X7Y99_SLICE_X8Y99_A1 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLM_R_X7Y99_SLICE_X8Y99_A2 = CLBLM_R_X7Y98_SLICE_X8Y98_F7AMUX_O;
  assign CLBLL_L_X2Y97_SLICE_X1Y97_B1 = CLBLM_R_X3Y96_SLICE_X3Y96_BO5;
  assign CLBLL_L_X2Y97_SLICE_X1Y97_B2 = CLBLL_L_X2Y96_SLICE_X0Y96_DO6;
  assign CLBLL_L_X2Y97_SLICE_X1Y97_B3 = CLBLL_L_X2Y97_SLICE_X0Y97_AO5;
  assign CLBLL_L_X2Y97_SLICE_X1Y97_B4 = CLBLM_R_X3Y95_SLICE_X2Y95_CO6;
  assign CLBLL_L_X2Y97_SLICE_X1Y97_B5 = CLBLM_R_X3Y96_SLICE_X3Y96_BO6;
  assign CLBLL_L_X2Y97_SLICE_X1Y97_B6 = CLBLM_R_X3Y95_SLICE_X2Y95_BO6;
  assign CLBLM_R_X7Y99_SLICE_X8Y99_A6 = CLBLM_R_X7Y99_SLICE_X8Y99_CO6;
  assign CLBLL_L_X2Y97_SLICE_X1Y97_C1 = CLBLM_R_X3Y96_SLICE_X3Y96_BO6;
  assign CLBLL_L_X2Y97_SLICE_X1Y97_C2 = CLBLL_L_X2Y96_SLICE_X1Y96_CO6;
  assign CLBLL_L_X2Y97_SLICE_X1Y97_C3 = CLBLL_L_X2Y96_SLICE_X0Y96_BO6;
  assign CLBLL_L_X2Y97_SLICE_X1Y97_C4 = CLBLM_R_X3Y96_SLICE_X3Y96_BO5;
  assign CLBLL_L_X2Y97_SLICE_X1Y97_C5 = CLBLM_R_X3Y95_SLICE_X2Y95_DO6;
  assign CLBLL_L_X2Y97_SLICE_X1Y97_C6 = CLBLL_L_X2Y97_SLICE_X0Y97_AO5;
  assign CLBLM_R_X7Y99_SLICE_X8Y99_B5 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X7Y99_SLICE_X8Y99_C1 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO0;
  assign CLBLM_R_X7Y99_SLICE_X8Y99_C2 = CLBLM_R_X5Y95_SLICE_X6Y95_AQ;
  assign CLBLM_R_X7Y99_SLICE_X8Y99_C3 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLL_L_X2Y97_SLICE_X1Y97_D1 = 1'b1;
  assign CLBLL_L_X2Y97_SLICE_X1Y97_D2 = CLBLM_R_X3Y95_SLICE_X2Y95_CO6;
  assign CLBLL_L_X2Y97_SLICE_X1Y97_D3 = CLBLL_L_X2Y96_SLICE_X0Y96_BO6;
  assign CLBLL_L_X2Y97_SLICE_X1Y97_D4 = CLBLL_L_X2Y96_SLICE_X1Y96_CO6;
  assign CLBLL_L_X2Y97_SLICE_X1Y97_D5 = CLBLM_R_X3Y95_SLICE_X2Y95_DO6;
  assign CLBLL_L_X2Y97_SLICE_X1Y97_D6 = 1'b1;
  assign CLBLM_R_X7Y99_SLICE_X8Y99_D1 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO0;
  assign CLBLM_R_X7Y99_SLICE_X8Y99_D2 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X7Y99_SLICE_X8Y99_D3 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X7Y99_SLICE_X8Y99_D4 = CLBLL_L_X4Y97_SLICE_X4Y97_BQ;
  assign CLBLM_R_X7Y99_SLICE_X8Y99_D5 = CLBLM_R_X5Y98_SLICE_X6Y98_DO6;
  assign CLBLM_R_X5Y91_SLICE_X7Y91_D5 = 1'b1;
  assign CLBLM_R_X7Y99_SLICE_X8Y99_D6 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X7Y99_SLICE_X8Y99_SR = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y96_SLICE_X9Y96_A4 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X7Y96_SLICE_X9Y96_A5 = CLBLM_R_X7Y98_SLICE_X8Y98_F7AMUX_O;
  assign CLBLM_R_X5Y91_SLICE_X7Y91_D6 = 1'b1;
  assign CLBLM_R_X7Y96_SLICE_X9Y96_A6 = CLBLM_R_X7Y96_SLICE_X9Y96_CO6;
  assign CLBLM_R_X7Y99_SLICE_X8Y99_A3 = CLBLM_R_X7Y99_SLICE_X8Y99_AQ;
  assign CLBLM_R_X7Y96_SLICE_X9Y96_B2 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_D = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y96_SLICE_X9Y96_B3 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X7Y96_SLICE_X9Y96_B4 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X7Y96_SLICE_X9Y96_B5 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO6;
  assign CLBLM_R_X7Y96_SLICE_X9Y96_B6 = CLBLM_R_X5Y95_SLICE_X6Y95_AQ;
  assign CLBLM_R_X3Y92_SLICE_X3Y92_A1 = 1'b1;
  assign CLBLM_R_X3Y92_SLICE_X3Y92_A2 = 1'b1;
  assign CLBLM_R_X7Y96_SLICE_X9Y96_C4 = CLBLM_R_X5Y95_SLICE_X6Y95_AQ;
  assign CLBLM_R_X7Y96_SLICE_X9Y96_C5 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X7Y96_SLICE_X9Y96_C6 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X5Y90_SLICE_X7Y90_D1 = 1'b1;
  assign CLBLM_R_X7Y99_SLICE_X8Y99_A4 = CLBLM_R_X7Y99_SLICE_X8Y99_BO6;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_A1 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_A2 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_A3 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_A4 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_A5 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_A6 = 1'b1;
  assign CLBLM_R_X5Y90_SLICE_X7Y90_D2 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_AX = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_B1 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_B2 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_B3 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_B4 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_B5 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_B6 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_C1 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_C2 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_C3 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_C4 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_C5 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_C6 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_CE = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_D1 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_D2 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_D3 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_D4 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_D5 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_D6 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_SR = CLBLL_L_X2Y98_SLICE_X1Y98_BO6;
  assign CLBLM_R_X5Y90_SLICE_X7Y90_A1 = CLBLM_R_X3Y98_SLICE_X3Y98_AO6;
  assign CLBLM_R_X5Y90_SLICE_X7Y90_A2 = CLBLL_L_X4Y98_SLICE_X4Y98_AO6;
  assign CLBLM_R_X5Y90_SLICE_X7Y90_A3 = CLBLM_R_X5Y94_SLICE_X6Y94_CO6;
  assign CLBLM_R_X5Y90_SLICE_X7Y90_A4 = CLBLL_L_X2Y97_SLICE_X0Y97_BO6;
  assign CLBLM_R_X5Y90_SLICE_X7Y90_A5 = CLBLL_L_X4Y97_SLICE_X4Y97_CO6;
  assign CLBLM_R_X5Y90_SLICE_X7Y90_A6 = 1'b1;
  assign CLBLM_R_X5Y90_SLICE_X7Y90_AX = CLBLL_L_X2Y96_SLICE_X1Y96_AO6;
  assign CLBLM_R_X5Y90_SLICE_X7Y90_B1 = 1'b1;
  assign CLBLM_R_X5Y90_SLICE_X7Y90_B2 = 1'b1;
  assign CLBLM_R_X5Y90_SLICE_X7Y90_B3 = 1'b1;
  assign CLBLM_R_X5Y90_SLICE_X7Y90_B4 = 1'b1;
  assign CLBLM_R_X5Y90_SLICE_X7Y90_B5 = 1'b1;
  assign CLBLM_R_X5Y90_SLICE_X7Y90_B6 = CLBLL_L_X2Y97_SLICE_X1Y97_AO6;
  assign CLBLM_R_X5Y90_SLICE_X7Y90_BX = CLBLL_L_X2Y96_SLICE_X1Y96_BO6;
  assign CLBLL_L_X4Y90_SLICE_X4Y90_C3 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_A1 = CLBLM_R_X3Y98_SLICE_X3Y98_AO6;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_A2 = CLBLL_L_X2Y97_SLICE_X0Y97_BO6;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_A3 = CLBLL_L_X2Y98_SLICE_X1Y98_AQ;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_A4 = CLBLL_L_X4Y97_SLICE_X4Y97_CO6;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_A5 = CLBLM_R_X5Y94_SLICE_X6Y94_CO6;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_A6 = CLBLL_L_X4Y98_SLICE_X4Y98_AO6;
  assign CLBLL_L_X4Y90_SLICE_X4Y90_C4 = 1'b1;
  assign CLBLM_R_X5Y90_SLICE_X7Y90_C1 = 1'b1;
  assign CLBLM_R_X5Y90_SLICE_X7Y90_C2 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_B1 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_B2 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_B3 = CLBLL_L_X2Y98_SLICE_X1Y98_AQ;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_B4 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_B5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_B6 = 1'b1;
  assign CLBLL_L_X4Y90_SLICE_X4Y90_C5 = 1'b1;
  assign CLBLM_R_X5Y90_SLICE_X7Y90_CX = CLBLL_L_X2Y97_SLICE_X1Y97_CO6;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_C1 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_C2 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_C3 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_C4 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_C5 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_C6 = 1'b1;
  assign CLBLM_R_X5Y90_SLICE_X7Y90_D3 = 1'b1;
  assign CLBLM_R_X5Y90_SLICE_X7Y90_D4 = 1'b1;
  assign CLBLM_R_X5Y90_SLICE_X6Y90_A1 = CLBLM_R_X3Y98_SLICE_X3Y98_AO6;
  assign CLBLM_R_X5Y90_SLICE_X6Y90_A2 = CLBLL_L_X2Y97_SLICE_X0Y97_BO6;
  assign CLBLM_R_X5Y90_SLICE_X6Y90_A3 = CLBLL_L_X4Y97_SLICE_X4Y97_CO6;
  assign CLBLM_R_X5Y90_SLICE_X6Y90_A4 = CLBLL_L_X4Y98_SLICE_X4Y98_AO6;
  assign CLBLM_R_X5Y90_SLICE_X6Y90_A5 = CLBLM_R_X5Y94_SLICE_X6Y94_CO6;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_D1 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_D2 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_D3 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_D4 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_D5 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_D6 = 1'b1;
  assign CLBLM_R_X5Y90_SLICE_X6Y90_A6 = 1'b1;
  assign CLBLM_R_X5Y90_SLICE_X6Y90_AX = CLBLL_L_X2Y96_SLICE_X1Y96_AO6;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_SR = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y90_SLICE_X6Y90_B1 = 1'b1;
  assign CLBLM_R_X5Y90_SLICE_X6Y90_B2 = 1'b1;
  assign CLBLM_R_X5Y90_SLICE_X6Y90_B3 = 1'b1;
  assign CLBLM_R_X5Y90_SLICE_X6Y90_B4 = 1'b1;
  assign CLBLM_R_X5Y90_SLICE_X6Y90_B5 = 1'b1;
  assign CLBLM_R_X5Y90_SLICE_X6Y90_B6 = CLBLL_L_X2Y97_SLICE_X1Y97_AO6;
  assign CLBLM_R_X5Y90_SLICE_X6Y90_BX = CLBLL_L_X2Y96_SLICE_X1Y96_BO6;
  assign CLBLM_R_X5Y90_SLICE_X6Y90_C1 = 1'b1;
  assign CLBLM_R_X5Y90_SLICE_X6Y90_C2 = 1'b1;
  assign CLBLM_R_X5Y90_SLICE_X6Y90_C3 = 1'b1;
  assign CLBLM_R_X5Y90_SLICE_X6Y90_C4 = 1'b1;
  assign CLBLM_R_X5Y90_SLICE_X6Y90_C5 = 1'b1;
  assign CLBLM_R_X5Y90_SLICE_X6Y90_C6 = 1'b1;
  assign CLBLM_R_X5Y90_SLICE_X6Y90_CE = CLBLM_R_X5Y90_SLICE_X6Y90_AO6;
  assign CLBLM_R_X7Y96_SLICE_X8Y96_B3 = CLBLM_R_X7Y96_SLICE_X8Y96_AQ;
  assign CLBLM_R_X7Y96_SLICE_X8Y96_B4 = 1'b1;
  assign CLBLM_R_X7Y96_SLICE_X8Y96_B5 = CLBLM_R_X7Y96_SLICE_X8Y96_CO6;
  assign CLBLM_R_X5Y90_SLICE_X6Y90_CX = CLBLL_L_X2Y97_SLICE_X0Y97_CO6;
  assign CLBLM_R_X5Y90_SLICE_X6Y90_D1 = 1'b1;
  assign CLBLM_R_X5Y90_SLICE_X6Y90_D2 = 1'b1;
  assign CLBLM_R_X5Y90_SLICE_X6Y90_D3 = 1'b1;
  assign CLBLM_R_X5Y90_SLICE_X6Y90_D4 = 1'b1;
  assign CLBLM_R_X5Y90_SLICE_X6Y90_D5 = 1'b1;
  assign CLBLM_R_X5Y90_SLICE_X6Y90_D6 = 1'b1;
  assign CLBLM_R_X7Y96_SLICE_X8Y96_B6 = 1'b1;
  assign CLBLM_R_X5Y90_SLICE_X6Y90_DX = CLBLL_L_X2Y97_SLICE_X1Y97_BO6;
  assign CLBLM_R_X5Y90_SLICE_X6Y90_SR = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0 = LIOB33_X0Y127_IOB_X0Y128_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1 = 1'b1;
  assign CLBLM_R_X7Y96_SLICE_X8Y96_C1 = CLBLM_R_X5Y96_SLICE_X6Y96_AQ;
  assign CLBLM_R_X7Y96_SLICE_X8Y96_C2 = CLBLM_R_X5Y99_SLICE_X7Y99_AQ;
  assign CLBLM_R_X5Y98_SLICE_X7Y98_D3 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X7Y96_SLICE_X8Y96_C3 = CLBLM_R_X5Y96_SLICE_X7Y96_AQ;
  assign CLBLM_R_X7Y87_SLICE_X8Y87_B6 = CLBLM_R_X7Y90_SLICE_X8Y90_CO6;
  assign CLBLM_R_X5Y90_SLICE_X7Y90_DX = CLBLL_L_X2Y97_SLICE_X1Y97_BO6;
  assign CLBLM_R_X5Y98_SLICE_X7Y98_D4 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X7Y96_SLICE_X8Y96_C4 = CLBLM_R_X7Y99_SLICE_X8Y99_AQ;
  assign CLBLM_R_X5Y98_SLICE_X7Y98_D5 = CLBLM_R_X5Y95_SLICE_X6Y95_AQ;
  assign CLBLM_R_X7Y96_SLICE_X8Y96_C5 = CLBLM_R_X5Y99_SLICE_X6Y99_AQ;
  assign CLBLM_R_X5Y98_SLICE_X7Y98_D6 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X7Y96_SLICE_X8Y96_C6 = CLBLM_R_X5Y96_SLICE_X7Y96_BQ;
  assign CLBLM_R_X7Y96_SLICE_X8Y96_CE = CLBLM_R_X7Y99_SLICE_X9Y99_DO6;
  assign CLBLM_R_X5Y90_SLICE_X7Y90_SR = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y98_SLICE_X6Y98_A4 = CLBLM_R_X7Y97_SLICE_X9Y97_B5Q;
  assign CLBLM_R_X5Y98_SLICE_X6Y98_A5 = 1'b0;
  assign CLBLM_R_X5Y98_SLICE_X6Y98_A6 = 1'b1;
  assign CLBLM_R_X7Y96_SLICE_X8Y96_D3 = CLBLL_L_X4Y97_SLICE_X4Y97_BQ;
  assign CLBLM_R_X7Y96_SLICE_X8Y96_D4 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X7Y96_SLICE_X8Y96_D5 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X7Y96_SLICE_X8Y96_D6 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X5Y98_SLICE_X6Y98_AX = CLBLM_R_X7Y97_SLICE_X8Y97_AQ;
  assign CLBLM_R_X7Y91_SLICE_X9Y91_D5 = CLBLM_R_X7Y91_SLICE_X9Y91_AQ;
  assign CLBLM_R_X7Y91_SLICE_X9Y91_D6 = CLBLM_R_X7Y87_SLICE_X8Y87_BQ;
  assign CLBLM_R_X7Y91_SLICE_X9Y91_SR = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X2Y99_SLICE_X0Y99_A1 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X0Y99_A2 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X0Y99_A3 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X0Y99_A4 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X0Y99_A5 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X0Y99_A6 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X0Y99_AX = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X2Y99_SLICE_X0Y99_B1 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X0Y99_B2 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X0Y99_B3 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X0Y99_B4 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X0Y99_B5 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X0Y99_B6 = 1'b1;
  assign CLBLM_R_X7Y89_SLICE_X8Y89_D6 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X0Y99_C1 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X0Y99_C2 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X0Y99_C3 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X0Y99_C4 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X0Y99_C5 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X0Y99_C6 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X0Y99_CE = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y91_SLICE_X8Y91_A3 = CLBLM_R_X7Y91_SLICE_X8Y91_AQ;
  assign CLBLM_R_X7Y91_SLICE_X8Y91_A4 = CLBLM_R_X7Y87_SLICE_X8Y87_BQ;
  assign CLBLM_R_X7Y91_SLICE_X8Y91_A5 = CLBLM_R_X7Y91_SLICE_X9Y91_AQ;
  assign CLBLL_L_X2Y99_SLICE_X0Y99_D1 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X0Y99_D2 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X0Y99_D3 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X0Y99_D4 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X0Y99_D5 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X0Y99_D6 = 1'b1;
  assign CLBLM_R_X7Y91_SLICE_X8Y91_A6 = CLBLM_R_X7Y87_SLICE_X8Y87_AQ;
  assign CLBLL_L_X2Y99_SLICE_X0Y99_SR = CLBLL_L_X2Y98_SLICE_X1Y98_BO6;
  assign CLBLM_R_X5Y91_SLICE_X7Y91_A1 = 1'b1;
  assign CLBLM_R_X5Y91_SLICE_X7Y91_A2 = 1'b1;
  assign CLBLM_R_X5Y91_SLICE_X7Y91_A3 = 1'b1;
  assign CLBLM_R_X5Y91_SLICE_X7Y91_A4 = 1'b1;
  assign CLBLM_R_X5Y91_SLICE_X7Y91_A5 = 1'b1;
  assign CLBLM_R_X5Y91_SLICE_X7Y91_A6 = 1'b1;
  assign CLBLM_R_X5Y91_SLICE_X7Y91_B1 = 1'b1;
  assign CLBLM_R_X5Y91_SLICE_X7Y91_B2 = 1'b1;
  assign CLBLM_R_X5Y91_SLICE_X7Y91_B3 = 1'b1;
  assign CLBLM_R_X5Y91_SLICE_X7Y91_B4 = 1'b1;
  assign CLBLM_R_X5Y91_SLICE_X7Y91_B5 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X1Y99_A1 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X1Y99_A2 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X1Y99_A3 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X1Y99_A4 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X1Y99_A5 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X1Y99_A6 = 1'b1;
  assign CLBLM_R_X5Y91_SLICE_X7Y91_B6 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X1Y99_AX = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y91_SLICE_X7Y91_C1 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X1Y99_B1 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X1Y99_B2 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X1Y99_B3 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X1Y99_B4 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X1Y99_B5 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X1Y99_B6 = 1'b1;
  assign CLBLM_R_X5Y91_SLICE_X7Y91_C3 = 1'b1;
  assign CLBLM_R_X5Y91_SLICE_X7Y91_C4 = 1'b1;
  assign CLBLM_R_X5Y91_SLICE_X7Y91_C6 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X1Y99_C1 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X1Y99_C2 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X1Y99_C3 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X1Y99_C4 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X1Y99_C5 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X1Y99_C6 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X1Y99_CE = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y91_SLICE_X7Y91_D1 = 1'b1;
  assign CLBLM_R_X5Y91_SLICE_X7Y91_D2 = 1'b1;
  assign CLBLM_R_X5Y91_SLICE_X7Y91_D3 = 1'b1;
  assign CLBLM_R_X5Y91_SLICE_X7Y91_D4 = 1'b1;
  assign CLBLM_R_X5Y91_SLICE_X6Y91_A1 = CLBLM_R_X5Y94_SLICE_X6Y94_CO6;
  assign CLBLL_L_X2Y99_SLICE_X1Y99_D1 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X1Y99_D2 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X1Y99_D3 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X1Y99_D4 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X1Y99_D5 = 1'b1;
  assign CLBLL_L_X2Y99_SLICE_X1Y99_D6 = 1'b1;
  assign CLBLM_R_X5Y91_SLICE_X6Y91_A2 = CLBLL_L_X4Y98_SLICE_X4Y98_AO6;
  assign CLBLM_R_X5Y91_SLICE_X6Y91_A3 = CLBLM_R_X5Y91_SLICE_X6Y91_AQ;
  assign CLBLL_L_X2Y99_SLICE_X1Y99_SR = CLBLL_L_X2Y98_SLICE_X1Y98_BO6;
  assign CLBLM_R_X5Y91_SLICE_X6Y91_A4 = CLBLL_L_X2Y97_SLICE_X0Y97_CO6;
  assign CLBLM_R_X5Y91_SLICE_X6Y91_A5 = CLBLL_L_X4Y97_SLICE_X4Y97_CO6;
  assign CLBLM_R_X5Y91_SLICE_X6Y91_A6 = CLBLM_R_X3Y98_SLICE_X3Y98_AO6;
  assign CLBLM_R_X5Y91_SLICE_X6Y91_B1 = 1'b1;
  assign CLBLM_R_X5Y91_SLICE_X6Y91_B2 = 1'b1;
  assign CLBLM_R_X5Y91_SLICE_X6Y91_B3 = 1'b1;
  assign CLBLM_R_X5Y91_SLICE_X6Y91_B4 = 1'b1;
  assign CLBLM_R_X5Y91_SLICE_X6Y91_B5 = 1'b1;
  assign CLBLM_R_X5Y91_SLICE_X6Y91_B6 = 1'b1;
  assign CLBLM_R_X5Y91_SLICE_X6Y91_C1 = 1'b1;
  assign CLBLM_R_X5Y91_SLICE_X6Y91_C2 = 1'b1;
  assign CLBLM_R_X5Y91_SLICE_X6Y91_C3 = 1'b1;
  assign CLBLM_R_X5Y91_SLICE_X6Y91_C4 = 1'b1;
  assign CLBLM_R_X5Y91_SLICE_X6Y91_C5 = 1'b1;
  assign CLBLM_R_X5Y91_SLICE_X6Y91_C6 = 1'b1;
  assign CLBLM_R_X7Y91_SLICE_X8Y91_C1 = CLBLM_R_X7Y87_SLICE_X8Y87_BQ;
  assign CLBLM_R_X7Y91_SLICE_X8Y91_C2 = CLBLM_R_X7Y91_SLICE_X8Y91_AQ;
  assign CLBLM_R_X7Y91_SLICE_X8Y91_C3 = BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO1;
  assign CLBLM_R_X7Y91_SLICE_X8Y91_C4 = CLBLM_R_X7Y87_SLICE_X8Y87_AQ;
  assign CLBLM_R_X5Y91_SLICE_X6Y91_D1 = 1'b1;
  assign CLBLM_R_X5Y91_SLICE_X6Y91_D2 = 1'b1;
  assign CLBLM_R_X5Y91_SLICE_X6Y91_D3 = 1'b1;
  assign CLBLM_R_X5Y91_SLICE_X6Y91_D4 = 1'b1;
  assign CLBLM_R_X5Y91_SLICE_X6Y91_D5 = 1'b1;
  assign CLBLM_R_X5Y91_SLICE_X6Y91_D6 = 1'b1;
  assign CLBLM_R_X5Y91_SLICE_X6Y91_SR = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y92_SLICE_X3Y92_C5 = 1'b1;
  assign CLBLM_R_X7Y91_SLICE_X8Y91_D1 = CLBLM_R_X7Y87_SLICE_X8Y87_BQ;
  assign CLBLM_R_X7Y91_SLICE_X8Y91_D2 = CLBLM_R_X7Y91_SLICE_X8Y91_AQ;
  assign CLBLM_R_X7Y91_SLICE_X8Y91_D3 = BRAM_L_X6Y90_RAMB36_X0Y18_DOBDO2;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0 = 1'b1;
  assign CLBLM_R_X7Y91_SLICE_X8Y91_D4 = CLBLM_R_X7Y89_SLICE_X8Y89_CO6;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1 = 1'b1;
  assign CLBLM_R_X7Y91_SLICE_X8Y91_D5 = 1'b1;
  assign CLBLM_R_X7Y88_SLICE_X8Y88_D4 = 1'b1;
  assign CLBLM_R_X7Y91_SLICE_X8Y91_D6 = CLBLM_R_X7Y87_SLICE_X8Y87_AQ;
  assign CLBLM_R_X7Y88_SLICE_X8Y88_D5 = 1'b1;
  assign CLBLM_R_X7Y88_SLICE_X8Y88_D6 = 1'b1;
  assign CLBLM_R_X7Y93_SLICE_X9Y93_A2 = 1'b1;
  assign CLBLM_R_X5Y92_SLICE_X7Y92_A1 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLM_R_X5Y92_SLICE_X7Y92_A2 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X5Y92_SLICE_X7Y92_A3 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X5Y92_SLICE_X7Y92_A4 = 1'b1;
  assign CLBLM_R_X5Y92_SLICE_X7Y92_A5 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X5Y92_SLICE_X7Y92_A6 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X5Y92_SLICE_X7Y92_B1 = 1'b1;
  assign CLBLM_R_X5Y92_SLICE_X7Y92_B2 = 1'b1;
  assign CLBLM_R_X5Y92_SLICE_X7Y92_B3 = 1'b1;
  assign CLBLM_R_X5Y92_SLICE_X7Y92_B4 = 1'b1;
  assign CLBLM_R_X5Y92_SLICE_X7Y92_B5 = 1'b1;
  assign CLBLM_R_X5Y92_SLICE_X7Y92_B6 = 1'b1;
  assign CLBLM_R_X5Y92_SLICE_X7Y92_C1 = 1'b1;
  assign CLBLM_R_X5Y92_SLICE_X7Y92_C2 = 1'b1;
  assign CLBLM_R_X5Y92_SLICE_X7Y92_C3 = 1'b1;
  assign CLBLM_R_X5Y92_SLICE_X7Y92_C4 = 1'b1;
  assign CLBLM_R_X5Y92_SLICE_X7Y92_C5 = 1'b1;
  assign CLBLM_R_X5Y92_SLICE_X7Y92_C6 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X3Y90_A3 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X3Y90_A4 = 1'b1;
  assign CLBLM_R_X5Y92_SLICE_X7Y92_D1 = 1'b1;
  assign CLBLM_R_X5Y92_SLICE_X7Y92_D2 = 1'b1;
  assign CLBLM_R_X5Y92_SLICE_X7Y92_D3 = 1'b1;
  assign CLBLM_R_X5Y92_SLICE_X7Y92_D4 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X3Y90_A5 = 1'b1;
  assign CLBLM_R_X5Y92_SLICE_X7Y92_D5 = 1'b1;
  assign CLBLM_R_X5Y92_SLICE_X7Y92_D6 = 1'b1;
  assign CLBLM_R_X5Y92_SLICE_X6Y92_A1 = CLBLM_R_X5Y94_SLICE_X7Y94_DO6;
  assign CLBLM_R_X5Y92_SLICE_X6Y92_A2 = CLBLL_L_X4Y94_SLICE_X5Y94_DO6;
  assign CLBLM_R_X5Y92_SLICE_X6Y92_A3 = CLBLL_L_X2Y96_SLICE_X1Y96_AO6;
  assign CLBLM_R_X5Y92_SLICE_X6Y92_A4 = CLBLM_R_X5Y94_SLICE_X6Y94_BO6;
  assign CLBLM_R_X5Y92_SLICE_X6Y92_A5 = CLBLM_R_X3Y93_SLICE_X2Y93_CO6;
  assign CLBLM_R_X5Y92_SLICE_X6Y92_A6 = CLBLL_L_X4Y96_SLICE_X4Y96_AO6;
  assign CLBLM_R_X5Y92_SLICE_X6Y92_B1 = CLBLM_R_X5Y94_SLICE_X7Y94_DO6;
  assign CLBLM_R_X5Y92_SLICE_X6Y92_B2 = CLBLL_L_X2Y96_SLICE_X1Y96_BO6;
  assign CLBLM_R_X5Y92_SLICE_X6Y92_B3 = CLBLL_L_X4Y96_SLICE_X5Y96_AO6;
  assign CLBLM_R_X5Y92_SLICE_X6Y92_B4 = CLBLL_L_X4Y94_SLICE_X5Y94_DO6;
  assign CLBLM_R_X5Y92_SLICE_X6Y92_B5 = CLBLM_R_X3Y93_SLICE_X2Y93_CO6;
  assign CLBLM_R_X5Y92_SLICE_X6Y92_B6 = CLBLM_R_X5Y94_SLICE_X6Y94_BO6;
  assign CLBLM_R_X5Y92_SLICE_X6Y92_C1 = CLBLM_R_X3Y93_SLICE_X2Y93_CO6;
  assign CLBLM_R_X5Y92_SLICE_X6Y92_C2 = CLBLM_R_X5Y94_SLICE_X7Y94_DO6;
  assign CLBLM_R_X5Y92_SLICE_X6Y92_C3 = CLBLM_R_X3Y99_SLICE_X2Y99_CO6;
  assign CLBLM_R_X5Y92_SLICE_X6Y92_C4 = CLBLL_L_X4Y94_SLICE_X5Y94_DO6;
  assign CLBLM_R_X5Y92_SLICE_X6Y92_C5 = CLBLL_L_X2Y97_SLICE_X0Y97_BO6;
  assign CLBLM_R_X5Y92_SLICE_X6Y92_C6 = CLBLM_R_X5Y94_SLICE_X6Y94_BO6;
  assign CLBLM_R_X5Y92_SLICE_X6Y92_D1 = 1'b1;
  assign CLBLM_R_X5Y92_SLICE_X6Y92_D2 = 1'b1;
  assign CLBLM_R_X5Y92_SLICE_X6Y92_D3 = 1'b1;
  assign CLBLM_R_X5Y92_SLICE_X6Y92_D4 = 1'b1;
  assign CLBLM_R_X5Y92_SLICE_X6Y92_D5 = 1'b1;
  assign CLBLM_R_X5Y92_SLICE_X6Y92_D6 = 1'b1;
  assign CLBLM_R_X5Y92_SLICE_X6Y92_SR = CLBLM_R_X5Y92_SLICE_X7Y92_AO6;
  assign CLBLM_R_X5Y90_SLICE_X7Y90_D5 = 1'b1;
  assign CLBLM_R_X7Y99_SLICE_X8Y99_A5 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X5Y90_SLICE_X7Y90_D6 = 1'b1;
  assign CLBLM_R_X7Y88_SLICE_X8Y88_C3 = 1'b1;
  assign CLBLM_R_X5Y93_SLICE_X7Y93_A1 = CLBLM_R_X5Y93_SLICE_X7Y93_AQ;
  assign CLBLM_R_X5Y93_SLICE_X7Y93_A2 = CLBLL_L_X2Y97_SLICE_X1Y97_AO6;
  assign CLBLM_R_X5Y93_SLICE_X7Y93_A3 = CLBLM_R_X5Y94_SLICE_X6Y94_CO6;
  assign CLBLM_R_X5Y93_SLICE_X7Y93_A4 = CLBLL_L_X4Y97_SLICE_X4Y97_CO6;
  assign CLBLM_R_X5Y93_SLICE_X7Y93_A5 = CLBLL_L_X4Y98_SLICE_X4Y98_AO6;
  assign CLBLM_R_X5Y93_SLICE_X7Y93_A6 = CLBLM_R_X3Y98_SLICE_X3Y98_AO6;
  assign CLBLM_R_X5Y93_SLICE_X7Y93_B1 = CLBLL_L_X2Y97_SLICE_X0Y97_BO6;
  assign CLBLM_R_X5Y93_SLICE_X7Y93_B2 = CLBLM_R_X5Y93_SLICE_X7Y93_BQ;
  assign CLBLM_R_X5Y93_SLICE_X7Y93_B3 = CLBLM_R_X5Y94_SLICE_X6Y94_CO6;
  assign CLBLM_R_X5Y93_SLICE_X7Y93_B4 = CLBLL_L_X4Y98_SLICE_X4Y98_AO6;
  assign CLBLM_R_X5Y93_SLICE_X7Y93_B5 = CLBLL_L_X4Y97_SLICE_X4Y97_CO6;
  assign CLBLM_R_X5Y93_SLICE_X7Y93_B6 = CLBLM_R_X3Y98_SLICE_X3Y98_AO6;
  assign CLBLM_R_X5Y93_SLICE_X7Y93_C1 = CLBLL_L_X4Y97_SLICE_X4Y97_CO6;
  assign CLBLM_R_X5Y93_SLICE_X7Y93_C2 = CLBLM_R_X5Y94_SLICE_X6Y94_CO6;
  assign CLBLM_R_X5Y93_SLICE_X7Y93_C3 = CLBLL_L_X4Y98_SLICE_X4Y98_AO6;
  assign CLBLM_R_X5Y93_SLICE_X7Y93_C4 = CLBLM_R_X3Y98_SLICE_X3Y98_AO6;
  assign CLBLM_R_X5Y93_SLICE_X7Y93_C5 = CLBLM_R_X5Y93_SLICE_X7Y93_CQ;
  assign CLBLM_R_X5Y93_SLICE_X7Y93_C6 = CLBLL_L_X2Y97_SLICE_X0Y97_BO6;
  assign CLBLM_R_X5Y93_SLICE_X7Y93_D1 = 1'b1;
  assign CLBLM_R_X5Y93_SLICE_X7Y93_D2 = 1'b1;
  assign CLBLM_R_X5Y93_SLICE_X7Y93_D3 = 1'b1;
  assign CLBLM_R_X5Y93_SLICE_X7Y93_D4 = 1'b1;
  assign CLBLM_R_X5Y93_SLICE_X7Y93_D5 = 1'b1;
  assign CLBLM_R_X5Y93_SLICE_X7Y93_D6 = 1'b1;
  assign CLBLM_R_X5Y93_SLICE_X7Y93_SR = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y93_SLICE_X6Y93_A1 = 1'b1;
  assign CLBLM_R_X5Y93_SLICE_X6Y93_A2 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X5Y93_SLICE_X6Y93_A3 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X5Y93_SLICE_X6Y93_A4 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO9;
  assign CLBLM_R_X5Y93_SLICE_X6Y93_A5 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X5Y93_SLICE_X6Y93_A6 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X5Y93_SLICE_X6Y93_AX = CLBLL_L_X4Y91_SLICE_X5Y91_CO6;
  assign CLBLM_R_X5Y93_SLICE_X6Y93_B1 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X5Y93_SLICE_X6Y93_B2 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X5Y93_SLICE_X6Y93_B3 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X5Y93_SLICE_X6Y93_B4 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO9;
  assign CLBLM_R_X5Y93_SLICE_X6Y93_B5 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X5Y93_SLICE_X6Y93_B6 = CLBLM_R_X5Y93_SLICE_X6Y93_CO6;
  assign CLBLM_R_X5Y93_SLICE_X6Y93_BX = CLBLL_L_X4Y93_SLICE_X4Y93_CO6;
  assign CLBLM_R_X5Y93_SLICE_X6Y93_C1 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO12;
  assign CLBLM_R_X5Y93_SLICE_X6Y93_C2 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO13;
  assign CLBLM_R_X5Y93_SLICE_X6Y93_C3 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO15;
  assign CLBLM_R_X5Y93_SLICE_X6Y93_C4 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO9;
  assign CLBLM_R_X5Y93_SLICE_X6Y93_C5 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO14;
  assign CLBLM_R_X5Y93_SLICE_X6Y93_C6 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO11;
  assign CLBLM_R_X5Y93_SLICE_X6Y93_CE = CLBLL_L_X2Y93_SLICE_X0Y93_DO6;
  assign CLBLM_R_X5Y93_SLICE_X6Y93_D1 = 1'b1;
  assign CLBLM_R_X5Y93_SLICE_X6Y93_D2 = 1'b1;
  assign CLBLM_R_X5Y93_SLICE_X6Y93_D3 = 1'b1;
  assign CLBLM_R_X5Y93_SLICE_X6Y93_D4 = 1'b1;
  assign CLBLM_R_X5Y93_SLICE_X6Y93_D5 = 1'b1;
  assign CLBLM_R_X5Y93_SLICE_X6Y93_D6 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_A1 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_A2 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_A3 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_A4 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_A5 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_A6 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_AX = CLBLM_R_X7Y90_SLICE_X8Y90_BQ;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_B1 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_B2 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_B3 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_B4 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_B5 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_B6 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_C1 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_C2 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_C3 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_C4 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_C5 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_C6 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_D1 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_D2 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_D3 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_D4 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_D5 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_D6 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_SR = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y90_SLICE_X4Y90_A1 = 1'b1;
  assign CLBLL_L_X4Y90_SLICE_X4Y90_A2 = 1'b1;
  assign CLBLL_L_X4Y90_SLICE_X4Y90_A3 = 1'b1;
  assign CLBLL_L_X4Y90_SLICE_X4Y90_A4 = 1'b1;
  assign CLBLL_L_X4Y90_SLICE_X4Y90_A5 = 1'b1;
  assign CLBLL_L_X4Y90_SLICE_X4Y90_A6 = 1'b1;
  assign CLBLL_L_X4Y90_SLICE_X4Y90_B1 = 1'b1;
  assign CLBLL_L_X4Y90_SLICE_X4Y90_B2 = 1'b1;
  assign CLBLL_L_X4Y90_SLICE_X4Y90_B3 = 1'b1;
  assign CLBLL_L_X4Y90_SLICE_X4Y90_B4 = 1'b1;
  assign CLBLL_L_X4Y90_SLICE_X4Y90_B5 = 1'b1;
  assign CLBLL_L_X4Y90_SLICE_X4Y90_B6 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_A1 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_A2 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_A3 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_A4 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_A5 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_A6 = 1'b1;
  assign CLBLL_L_X4Y90_SLICE_X4Y90_C1 = 1'b1;
  assign CLBLL_L_X4Y90_SLICE_X4Y90_C2 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_B1 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_B2 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_B3 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_B4 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_B5 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_B6 = 1'b1;
  assign CLBLL_L_X4Y90_SLICE_X4Y90_C6 = 1'b1;
  assign CLBLL_L_X4Y90_SLICE_X4Y90_D1 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_C1 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_C2 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_C3 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_C4 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_C5 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_C6 = 1'b1;
  assign CLBLL_L_X4Y90_SLICE_X4Y90_D2 = 1'b1;
  assign CLBLL_L_X4Y90_SLICE_X4Y90_D3 = 1'b1;
  assign CLBLL_L_X4Y90_SLICE_X4Y90_D4 = 1'b1;
  assign CLBLL_L_X4Y90_SLICE_X4Y90_D5 = 1'b1;
  assign CLBLL_L_X4Y90_SLICE_X4Y90_D6 = 1'b1;
  assign CLBLM_R_X5Y94_SLICE_X7Y94_C4 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO8;
  assign CLBLM_R_X5Y94_SLICE_X7Y94_C6 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO11;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_D1 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_D2 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_D3 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_D4 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_D5 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_D6 = 1'b1;
  assign CLBLM_R_X5Y94_SLICE_X7Y94_D4 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLM_R_X5Y94_SLICE_X7Y94_D5 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X5Y94_SLICE_X7Y94_D6 = CLBLM_R_X5Y94_SLICE_X7Y94_BO6;
  assign CLBLM_R_X5Y94_SLICE_X7Y94_D3 = CLBLM_R_X5Y94_SLICE_X7Y94_AO5;
  assign CLBLM_R_X5Y94_SLICE_X6Y94_A1 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X5Y94_SLICE_X6Y94_A2 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X5Y94_SLICE_X6Y94_A3 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO9;
  assign CLBLM_R_X5Y94_SLICE_X6Y94_A4 = CLBLM_R_X5Y95_SLICE_X6Y95_DO6;
  assign CLBLL_L_X4Y90_SLICE_X5Y90_A1 = 1'b1;
  assign CLBLL_L_X4Y90_SLICE_X5Y90_A2 = 1'b1;
  assign CLBLL_L_X4Y90_SLICE_X5Y90_A3 = 1'b1;
  assign CLBLL_L_X4Y90_SLICE_X5Y90_A4 = 1'b1;
  assign CLBLL_L_X4Y90_SLICE_X5Y90_A5 = 1'b1;
  assign CLBLL_L_X4Y90_SLICE_X5Y90_A6 = 1'b1;
  assign CLBLM_R_X5Y94_SLICE_X6Y94_A5 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X5Y94_SLICE_X6Y94_A6 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLL_L_X4Y90_SLICE_X5Y90_AX = CLBLM_R_X7Y90_SLICE_X8Y90_AQ;
  assign CLBLM_R_X5Y94_SLICE_X6Y94_AX = CLBLL_L_X4Y93_SLICE_X4Y93_CO5;
  assign CLBLL_L_X4Y90_SLICE_X5Y90_B1 = 1'b1;
  assign CLBLL_L_X4Y90_SLICE_X5Y90_B2 = 1'b1;
  assign CLBLL_L_X4Y90_SLICE_X5Y90_B3 = 1'b1;
  assign CLBLL_L_X4Y90_SLICE_X5Y90_B4 = 1'b1;
  assign CLBLL_L_X4Y90_SLICE_X5Y90_B5 = 1'b1;
  assign CLBLL_L_X4Y90_SLICE_X5Y90_B6 = 1'b1;
  assign CLBLM_R_X5Y94_SLICE_X6Y94_B1 = CLBLM_R_X5Y94_SLICE_X7Y94_AO5;
  assign CLBLM_R_X5Y94_SLICE_X6Y94_B2 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X5Y94_SLICE_X6Y94_B4 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLL_L_X4Y90_SLICE_X5Y90_C1 = 1'b1;
  assign CLBLL_L_X4Y90_SLICE_X5Y90_C2 = 1'b1;
  assign CLBLL_L_X4Y90_SLICE_X5Y90_C3 = 1'b1;
  assign CLBLL_L_X4Y90_SLICE_X5Y90_C4 = 1'b1;
  assign CLBLL_L_X4Y90_SLICE_X5Y90_C5 = 1'b1;
  assign CLBLL_L_X4Y90_SLICE_X5Y90_C6 = 1'b1;
  assign CLBLM_R_X5Y94_SLICE_X6Y94_C1 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X5Y94_SLICE_X6Y94_C2 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X5Y94_SLICE_X6Y94_C3 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLM_R_X5Y94_SLICE_X6Y94_C4 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X5Y94_SLICE_X6Y94_C5 = 1'b1;
  assign CLBLM_R_X5Y94_SLICE_X6Y94_C6 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLL_L_X4Y90_SLICE_X5Y90_D1 = 1'b1;
  assign CLBLL_L_X4Y90_SLICE_X5Y90_D2 = 1'b1;
  assign CLBLL_L_X4Y90_SLICE_X5Y90_D3 = 1'b1;
  assign CLBLL_L_X4Y90_SLICE_X5Y90_D4 = 1'b1;
  assign CLBLL_L_X4Y90_SLICE_X5Y90_D5 = 1'b1;
  assign CLBLL_L_X4Y90_SLICE_X5Y90_D6 = 1'b1;
  assign CLBLM_R_X5Y94_SLICE_X6Y94_D1 = 1'b1;
  assign CLBLL_L_X4Y90_SLICE_X5Y90_SR = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y94_SLICE_X6Y94_D3 = 1'b1;
  assign CLBLM_R_X5Y94_SLICE_X6Y94_D4 = 1'b1;
  assign CLBLM_R_X5Y94_SLICE_X6Y94_D5 = 1'b1;
  assign CLBLM_R_X5Y94_SLICE_X6Y94_D6 = 1'b1;
  assign CLBLM_R_X7Y97_SLICE_X9Y97_B6 = 1'b1;
  assign CLBLL_L_X4Y96_SLICE_X5Y96_B3 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLL_L_X4Y96_SLICE_X5Y96_B4 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO5;
  assign CLBLL_L_X4Y96_SLICE_X5Y96_B5 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLL_L_X4Y96_SLICE_X5Y96_B6 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X7Y98_SLICE_X8Y98_A6 = CLBLM_R_X5Y95_SLICE_X6Y95_AQ;
  assign CLBLL_L_X4Y96_SLICE_X5Y96_C2 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLL_L_X4Y96_SLICE_X5Y96_C3 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLL_L_X4Y91_SLICE_X4Y91_A1 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLL_L_X4Y91_SLICE_X4Y91_A2 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO5;
  assign CLBLL_L_X4Y91_SLICE_X4Y91_A3 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLL_L_X4Y91_SLICE_X4Y91_A4 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLL_L_X4Y91_SLICE_X4Y91_A5 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLL_L_X4Y91_SLICE_X4Y91_A6 = 1'b1;
  assign CLBLL_L_X4Y91_SLICE_X4Y91_AX = CLBLL_L_X4Y93_SLICE_X4Y93_CO5;
  assign CLBLL_L_X4Y91_SLICE_X4Y91_B1 = CLBLM_R_X3Y91_SLICE_X3Y91_F7BMUX_O;
  assign CLBLL_L_X4Y91_SLICE_X4Y91_B2 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLL_L_X4Y91_SLICE_X4Y91_B3 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLL_L_X4Y91_SLICE_X4Y91_B4 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLL_L_X4Y91_SLICE_X4Y91_B5 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO5;
  assign CLBLL_L_X4Y91_SLICE_X4Y91_B6 = CLBLL_L_X4Y91_SLICE_X4Y91_AO5;
  assign CLBLL_L_X4Y91_SLICE_X4Y91_BX = CLBLL_L_X4Y92_SLICE_X4Y92_AO5;
  assign CLBLL_L_X4Y91_SLICE_X4Y91_C1 = 1'b1;
  assign CLBLL_L_X4Y91_SLICE_X4Y91_C2 = 1'b1;
  assign CLBLL_L_X4Y91_SLICE_X4Y91_C3 = 1'b1;
  assign CLBLL_L_X4Y91_SLICE_X4Y91_C4 = 1'b1;
  assign CLBLL_L_X4Y91_SLICE_X4Y91_C5 = 1'b1;
  assign CLBLL_L_X4Y91_SLICE_X4Y91_C6 = 1'b1;
  assign CLBLL_L_X4Y91_SLICE_X4Y91_CE = CLBLL_L_X2Y93_SLICE_X1Y93_CO6;
  assign CLBLM_R_X5Y95_SLICE_X7Y95_A1 = 1'b1;
  assign CLBLM_R_X5Y95_SLICE_X7Y95_A2 = 1'b1;
  assign CLBLM_R_X5Y95_SLICE_X7Y95_A3 = 1'b1;
  assign CLBLM_R_X5Y95_SLICE_X7Y95_A4 = 1'b1;
  assign CLBLM_R_X5Y95_SLICE_X7Y95_A5 = 1'b1;
  assign CLBLM_R_X5Y95_SLICE_X7Y95_A6 = 1'b1;
  assign CLBLL_L_X4Y91_SLICE_X4Y91_D1 = 1'b1;
  assign CLBLL_L_X4Y91_SLICE_X4Y91_D2 = 1'b1;
  assign CLBLL_L_X4Y91_SLICE_X4Y91_D3 = 1'b1;
  assign CLBLL_L_X4Y91_SLICE_X4Y91_D4 = 1'b1;
  assign CLBLL_L_X4Y91_SLICE_X4Y91_D5 = 1'b1;
  assign CLBLL_L_X4Y91_SLICE_X4Y91_D6 = 1'b1;
  assign CLBLM_R_X5Y95_SLICE_X7Y95_B1 = 1'b1;
  assign CLBLM_R_X5Y95_SLICE_X7Y95_B2 = 1'b1;
  assign CLBLM_R_X5Y95_SLICE_X7Y95_B3 = 1'b1;
  assign CLBLM_R_X5Y95_SLICE_X7Y95_B4 = 1'b1;
  assign CLBLM_R_X5Y95_SLICE_X7Y95_B5 = 1'b1;
  assign CLBLM_R_X5Y95_SLICE_X7Y95_B6 = 1'b1;
  assign CLBLM_R_X5Y95_SLICE_X7Y95_C1 = 1'b1;
  assign CLBLM_R_X5Y95_SLICE_X7Y95_C2 = 1'b1;
  assign CLBLM_R_X5Y95_SLICE_X7Y95_C3 = 1'b1;
  assign CLBLM_R_X5Y95_SLICE_X7Y95_C4 = 1'b1;
  assign CLBLM_R_X5Y95_SLICE_X7Y95_C5 = 1'b1;
  assign CLBLM_R_X5Y95_SLICE_X7Y95_C6 = 1'b1;
  assign CLBLM_R_X5Y95_SLICE_X7Y95_D1 = 1'b1;
  assign CLBLM_R_X5Y95_SLICE_X7Y95_D2 = 1'b1;
  assign CLBLM_R_X5Y95_SLICE_X7Y95_D3 = 1'b1;
  assign CLBLL_L_X4Y96_SLICE_X5Y96_D3 = 1'b1;
  assign CLBLM_R_X5Y95_SLICE_X7Y95_D4 = 1'b1;
  assign CLBLM_R_X5Y95_SLICE_X7Y95_D5 = 1'b1;
  assign CLBLM_R_X5Y95_SLICE_X7Y95_D6 = 1'b1;
  assign CLBLL_L_X4Y96_SLICE_X5Y96_D4 = 1'b1;
  assign CLBLL_L_X4Y91_SLICE_X5Y91_A1 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLL_L_X4Y91_SLICE_X5Y91_A2 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLL_L_X4Y91_SLICE_X5Y91_A3 = 1'b1;
  assign CLBLL_L_X4Y91_SLICE_X5Y91_A4 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLL_L_X4Y91_SLICE_X5Y91_A5 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLL_L_X4Y91_SLICE_X5Y91_A6 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO8;
  assign CLBLM_R_X5Y95_SLICE_X6Y95_A1 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X5Y95_SLICE_X6Y95_A2 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLL_L_X4Y91_SLICE_X5Y91_AX = CLBLL_L_X4Y91_SLICE_X5Y91_CO6;
  assign CLBLM_R_X5Y95_SLICE_X6Y95_A3 = CLBLM_R_X5Y95_SLICE_X6Y95_AQ;
  assign CLBLL_L_X4Y91_SLICE_X5Y91_B1 = CLBLL_L_X4Y94_SLICE_X5Y94_CO6;
  assign CLBLL_L_X4Y91_SLICE_X5Y91_B2 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLL_L_X4Y91_SLICE_X5Y91_B3 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLL_L_X4Y91_SLICE_X5Y91_B4 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLL_L_X4Y91_SLICE_X5Y91_B5 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLL_L_X4Y91_SLICE_X5Y91_B6 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO8;
  assign CLBLM_R_X5Y95_SLICE_X6Y95_B1 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLL_L_X4Y91_SLICE_X5Y91_BX = CLBLL_L_X4Y92_SLICE_X4Y92_AO5;
  assign CLBLM_R_X5Y95_SLICE_X6Y95_B2 = CLBLM_R_X5Y95_SLICE_X6Y95_CO6;
  assign CLBLL_L_X4Y91_SLICE_X5Y91_C1 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLL_L_X4Y91_SLICE_X5Y91_C2 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLL_L_X4Y91_SLICE_X5Y91_C3 = 1'b1;
  assign CLBLL_L_X4Y91_SLICE_X5Y91_C4 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLL_L_X4Y91_SLICE_X5Y91_C5 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLL_L_X4Y91_SLICE_X5Y91_C6 = 1'b1;
  assign CLBLL_L_X4Y91_SLICE_X5Y91_CE = CLBLL_L_X2Y93_SLICE_X0Y93_DO6;
  assign CLBLM_R_X5Y95_SLICE_X6Y95_C1 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X5Y95_SLICE_X6Y95_C2 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO13;
  assign CLBLM_R_X5Y95_SLICE_X6Y95_C3 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO15;
  assign CLBLM_R_X5Y95_SLICE_X6Y95_C4 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO14;
  assign CLBLM_R_X5Y95_SLICE_X6Y95_C5 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO12;
  assign CLBLL_L_X4Y91_SLICE_X5Y91_D1 = 1'b1;
  assign CLBLL_L_X4Y91_SLICE_X5Y91_D2 = 1'b1;
  assign CLBLL_L_X4Y91_SLICE_X5Y91_D3 = 1'b1;
  assign CLBLL_L_X4Y91_SLICE_X5Y91_D4 = 1'b1;
  assign CLBLL_L_X4Y91_SLICE_X5Y91_D5 = 1'b1;
  assign CLBLL_L_X4Y91_SLICE_X5Y91_D6 = 1'b1;
  assign CLBLM_R_X5Y95_SLICE_X6Y95_D1 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO13;
  assign CLBLM_R_X5Y95_SLICE_X6Y95_D2 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO14;
  assign CLBLM_R_X5Y95_SLICE_X6Y95_D3 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO15;
  assign CLBLM_R_X5Y95_SLICE_X6Y95_D4 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO9;
  assign CLBLM_R_X5Y95_SLICE_X6Y95_D5 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO12;
  assign CLBLM_R_X5Y95_SLICE_X6Y95_D6 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO11;
  assign CLBLM_R_X5Y95_SLICE_X6Y95_SR = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y97_SLICE_X8Y97_B6 = 1'b1;
  assign CLBLM_R_X7Y97_SLICE_X8Y97_C1 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X7Y97_SLICE_X8Y97_C2 = CLBLM_R_X5Y95_SLICE_X6Y95_AQ;
  assign CLBLM_R_X7Y97_SLICE_X8Y97_C4 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO10;
  assign CLBLM_R_X5Y99_SLICE_X7Y99_D5 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X5Y99_SLICE_X7Y99_D6 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X5Y99_SLICE_X7Y99_SR = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y97_SLICE_X8Y97_D1 = CLBLM_R_X7Y99_SLICE_X9Y99_AQ;
  assign CLBLM_R_X7Y93_SLICE_X9Y93_A3 = 1'b1;
  assign CLBLM_R_X5Y94_SLICE_X7Y94_A1 = 1'b1;
  assign CLBLM_R_X5Y94_SLICE_X7Y94_A2 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X7Y97_SLICE_X8Y97_D4 = CLBLM_R_X7Y96_SLICE_X8Y96_CO6;
  assign CLBLM_R_X5Y94_SLICE_X7Y94_A3 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X7Y97_SLICE_X8Y97_D5 = CLBLM_R_X7Y96_SLICE_X9Y96_AQ;
  assign CLBLM_R_X5Y94_SLICE_X7Y94_A4 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X7Y97_SLICE_X8Y97_D6 = CLBLM_R_X7Y98_SLICE_X9Y98_AQ;
  assign CLBLM_R_X5Y94_SLICE_X7Y94_A5 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X5Y94_SLICE_X7Y94_A6 = 1'b1;
  assign CLBLM_R_X7Y97_SLICE_X8Y97_SR = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y94_SLICE_X7Y94_B1 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO8;
  assign CLBLM_R_X5Y94_SLICE_X7Y94_B2 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X5Y94_SLICE_X7Y94_B3 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X5Y94_SLICE_X7Y94_B4 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLL_L_X4Y92_SLICE_X4Y92_A1 = CLBLM_R_X3Y93_SLICE_X2Y93_CO6;
  assign CLBLL_L_X4Y92_SLICE_X4Y92_A2 = CLBLL_L_X2Y96_SLICE_X1Y96_AO6;
  assign CLBLL_L_X4Y92_SLICE_X4Y92_A3 = CLBLL_L_X4Y96_SLICE_X4Y96_AO6;
  assign CLBLL_L_X4Y92_SLICE_X4Y92_A4 = CLBLL_L_X4Y96_SLICE_X5Y96_AO6;
  assign CLBLL_L_X4Y92_SLICE_X4Y92_A5 = CLBLL_L_X2Y96_SLICE_X1Y96_BO6;
  assign CLBLL_L_X4Y92_SLICE_X4Y92_A6 = 1'b1;
  assign CLBLM_R_X5Y94_SLICE_X7Y94_B5 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X5Y94_SLICE_X7Y94_B6 = CLBLM_R_X5Y94_SLICE_X7Y94_CO6;
  assign CLBLL_L_X4Y92_SLICE_X4Y92_AX = CLBLL_L_X4Y93_SLICE_X4Y93_CO5;
  assign CLBLL_L_X4Y92_SLICE_X4Y92_B1 = CLBLM_R_X5Y94_SLICE_X7Y94_DO6;
  assign CLBLL_L_X4Y92_SLICE_X4Y92_B2 = CLBLL_L_X2Y93_SLICE_X0Y93_CO6;
  assign CLBLL_L_X4Y92_SLICE_X4Y92_B3 = CLBLL_L_X4Y94_SLICE_X5Y94_DO6;
  assign CLBLL_L_X4Y92_SLICE_X4Y92_B4 = CLBLM_R_X3Y94_SLICE_X2Y94_DO5;
  assign CLBLL_L_X4Y92_SLICE_X4Y92_B5 = CLBLM_R_X5Y94_SLICE_X6Y94_BO6;
  assign CLBLL_L_X4Y92_SLICE_X4Y92_B6 = 1'b1;
  assign CLBLL_L_X4Y92_SLICE_X4Y92_BX = CLBLL_L_X4Y94_SLICE_X4Y94_CO6;
  assign CLBLL_L_X4Y92_SLICE_X4Y92_C1 = 1'b1;
  assign CLBLL_L_X4Y92_SLICE_X4Y92_C2 = 1'b1;
  assign CLBLL_L_X4Y92_SLICE_X4Y92_C3 = 1'b1;
  assign CLBLL_L_X4Y92_SLICE_X4Y92_C4 = 1'b1;
  assign CLBLL_L_X4Y92_SLICE_X4Y92_C5 = 1'b1;
  assign CLBLL_L_X4Y92_SLICE_X4Y92_C6 = 1'b1;
  assign CLBLL_L_X4Y92_SLICE_X4Y92_CE = CLBLL_L_X4Y92_SLICE_X4Y92_BO6;
  assign CLBLM_R_X5Y96_SLICE_X7Y96_A1 = CLBLM_R_X5Y96_SLICE_X7Y96_DO6;
  assign CLBLM_R_X5Y94_SLICE_X7Y94_C1 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO12;
  assign CLBLM_R_X5Y96_SLICE_X7Y96_A2 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X5Y96_SLICE_X7Y96_A3 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLL_L_X4Y92_SLICE_X4Y92_CX = CLBLL_L_X4Y93_SLICE_X4Y93_CO6;
  assign CLBLM_R_X5Y96_SLICE_X7Y96_A4 = CLBLM_R_X5Y97_SLICE_X7Y97_BO6;
  assign CLBLL_L_X4Y92_SLICE_X4Y92_D1 = 1'b1;
  assign CLBLL_L_X4Y92_SLICE_X4Y92_D2 = 1'b1;
  assign CLBLL_L_X4Y92_SLICE_X4Y92_D3 = 1'b1;
  assign CLBLL_L_X4Y92_SLICE_X4Y92_D4 = 1'b1;
  assign CLBLL_L_X4Y92_SLICE_X4Y92_D5 = 1'b1;
  assign CLBLL_L_X4Y92_SLICE_X4Y92_D6 = 1'b1;
  assign CLBLM_R_X5Y94_SLICE_X7Y94_C2 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO14;
  assign CLBLM_R_X5Y94_SLICE_X7Y94_C3 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO13;
  assign CLBLL_L_X4Y92_SLICE_X4Y92_DX = CLBLL_L_X4Y92_SLICE_X4Y92_AO5;
  assign CLBLM_R_X5Y96_SLICE_X7Y96_B1 = CLBLM_R_X7Y98_SLICE_X8Y98_F7AMUX_O;
  assign CLBLM_R_X5Y96_SLICE_X7Y96_B2 = CLBLM_R_X5Y96_SLICE_X6Y96_BO6;
  assign CLBLM_R_X5Y96_SLICE_X7Y96_B3 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLM_R_X5Y96_SLICE_X7Y96_B4 = CLBLM_R_X5Y98_SLICE_X7Y98_DO6;
  assign CLBLM_R_X5Y96_SLICE_X7Y96_B5 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X5Y94_SLICE_X7Y94_C5 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO15;
  assign CLBLM_R_X5Y96_SLICE_X7Y96_B6 = CLBLM_R_X5Y96_SLICE_X7Y96_CO6;
  assign CLBLM_R_X5Y96_SLICE_X7Y96_C1 = CLBLM_R_X7Y99_SLICE_X8Y99_AQ;
  assign CLBLM_R_X5Y96_SLICE_X7Y96_C2 = CLBLM_R_X5Y99_SLICE_X6Y99_AQ;
  assign CLBLM_R_X5Y96_SLICE_X7Y96_C3 = CLBLM_R_X5Y99_SLICE_X7Y99_AQ;
  assign CLBLM_R_X5Y96_SLICE_X7Y96_C4 = CLBLM_R_X5Y96_SLICE_X7Y96_BQ;
  assign CLBLM_R_X5Y96_SLICE_X7Y96_C5 = CLBLM_R_X5Y96_SLICE_X7Y96_AQ;
  assign CLBLM_R_X5Y96_SLICE_X7Y96_C6 = 1'b1;
  assign CLBLM_R_X5Y96_SLICE_X7Y96_CE = CLBLM_R_X7Y99_SLICE_X9Y99_DO6;
  assign CLBLM_R_X5Y96_SLICE_X7Y96_D1 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X5Y96_SLICE_X7Y96_D2 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO3;
  assign CLBLM_R_X5Y96_SLICE_X7Y96_D3 = CLBLL_L_X4Y97_SLICE_X4Y97_BQ;
  assign CLBLM_R_X5Y96_SLICE_X7Y96_D4 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X5Y96_SLICE_X7Y96_D5 = CLBLM_R_X5Y95_SLICE_X6Y95_AQ;
  assign CLBLM_R_X5Y96_SLICE_X7Y96_D6 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLL_L_X4Y92_SLICE_X5Y92_A1 = CLBLM_R_X3Y93_SLICE_X3Y93_AQ;
  assign CLBLL_L_X4Y92_SLICE_X5Y92_A2 = CLBLL_L_X4Y92_SLICE_X5Y92_BQ;
  assign CLBLL_L_X4Y92_SLICE_X5Y92_A3 = CLBLL_L_X4Y94_SLICE_X5Y94_BQ;
  assign CLBLL_L_X4Y92_SLICE_X5Y92_A4 = CLBLM_R_X3Y96_SLICE_X3Y96_AO6;
  assign CLBLL_L_X4Y92_SLICE_X5Y92_A5 = CLBLL_L_X4Y91_SLICE_X4Y91_AO6;
  assign CLBLL_L_X4Y92_SLICE_X5Y92_A6 = CLBLL_L_X4Y93_SLICE_X5Y93_BQ;
  assign CLBLM_R_X5Y96_SLICE_X6Y96_A1 = CLBLM_R_X5Y96_SLICE_X6Y96_DO6;
  assign CLBLM_R_X5Y96_SLICE_X6Y96_A2 = CLBLM_R_X7Y98_SLICE_X8Y98_F7AMUX_O;
  assign CLBLL_L_X4Y92_SLICE_X5Y92_AX = CLBLL_L_X4Y95_SLICE_X5Y95_DO6;
  assign CLBLM_R_X5Y96_SLICE_X6Y96_A3 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLL_L_X4Y92_SLICE_X5Y92_B1 = CLBLM_R_X5Y92_SLICE_X6Y92_CQ;
  assign CLBLL_L_X4Y92_SLICE_X5Y92_B2 = CLBLM_R_X5Y94_SLICE_X6Y94_AQ;
  assign CLBLL_L_X4Y92_SLICE_X5Y92_B3 = CLBLL_L_X4Y91_SLICE_X4Y91_AQ;
  assign CLBLL_L_X4Y92_SLICE_X5Y92_B4 = CLBLM_R_X3Y96_SLICE_X3Y96_AO6;
  assign CLBLL_L_X4Y92_SLICE_X5Y92_B5 = CLBLL_L_X4Y92_SLICE_X4Y92_AQ;
  assign CLBLL_L_X4Y92_SLICE_X5Y92_B6 = CLBLL_L_X4Y91_SLICE_X4Y91_AO6;
  assign CLBLM_R_X5Y96_SLICE_X6Y96_A4 = CLBLL_L_X4Y97_SLICE_X5Y97_BO6;
  assign CLBLM_R_X5Y96_SLICE_X6Y96_A5 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLL_L_X4Y92_SLICE_X5Y92_BX = CLBLL_L_X4Y93_SLICE_X4Y93_CO5;
  assign CLBLM_R_X5Y96_SLICE_X6Y96_A6 = CLBLM_R_X5Y96_SLICE_X6Y96_CO6;
  assign CLBLL_L_X4Y92_SLICE_X5Y92_C1 = CLBLL_L_X4Y91_SLICE_X5Y91_CO6;
  assign CLBLL_L_X4Y92_SLICE_X5Y92_C2 = CLBLM_R_X5Y94_SLICE_X7Y94_AO5;
  assign CLBLL_L_X4Y92_SLICE_X5Y92_C3 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO8;
  assign CLBLL_L_X4Y92_SLICE_X5Y92_C4 = CLBLL_L_X4Y93_SLICE_X5Y93_BQ;
  assign CLBLL_L_X4Y92_SLICE_X5Y92_C5 = CLBLL_L_X4Y91_SLICE_X5Y91_BO6;
  assign CLBLL_L_X4Y92_SLICE_X5Y92_C6 = CLBLL_L_X4Y92_SLICE_X5Y92_BQ;
  assign CLBLL_L_X4Y92_SLICE_X5Y92_CE = CLBLL_L_X2Y93_SLICE_X0Y93_DO6;
  assign CLBLM_R_X5Y96_SLICE_X6Y96_B4 = CLBLM_R_X5Y95_SLICE_X6Y95_AQ;
  assign CLBLM_R_X5Y96_SLICE_X6Y96_B5 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X5Y96_SLICE_X6Y96_B6 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO4;
  assign CLBLL_L_X4Y92_SLICE_X5Y92_CX = CLBLL_L_X4Y94_SLICE_X4Y94_CO6;
  assign CLBLM_R_X3Y96_SLICE_X3Y96_A1 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO6;
  assign CLBLL_L_X4Y92_SLICE_X5Y92_D1 = CLBLL_L_X4Y92_SLICE_X4Y92_AQ;
  assign CLBLL_L_X4Y92_SLICE_X5Y92_D2 = CLBLM_R_X5Y94_SLICE_X7Y94_AO5;
  assign CLBLL_L_X4Y92_SLICE_X5Y92_D3 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO8;
  assign CLBLL_L_X4Y92_SLICE_X5Y92_D4 = CLBLM_R_X5Y92_SLICE_X6Y92_CQ;
  assign CLBLL_L_X4Y92_SLICE_X5Y92_D5 = CLBLL_L_X4Y91_SLICE_X5Y91_BO6;
  assign CLBLL_L_X4Y92_SLICE_X5Y92_D6 = CLBLL_L_X4Y91_SLICE_X5Y91_CO6;
  assign CLBLM_R_X3Y96_SLICE_X3Y96_A2 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLM_R_X5Y94_SLICE_X7Y94_D1 = CLBLM_R_X5Y94_SLICE_X7Y94_AO6;
  assign CLBLM_R_X3Y96_SLICE_X3Y96_A3 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X5Y94_SLICE_X7Y94_D2 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO8;
  assign CLBLM_R_X5Y96_SLICE_X6Y96_D1 = CLBLM_R_X5Y96_SLICE_X7Y96_AQ;
  assign CLBLM_R_X3Y96_SLICE_X3Y96_A4 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X5Y96_SLICE_X6Y96_D2 = CLBLM_R_X5Y96_SLICE_X7Y96_BQ;
  assign CLBLM_R_X5Y96_SLICE_X6Y96_D3 = CLBLM_R_X7Y99_SLICE_X8Y99_AQ;
  assign CLBLM_R_X5Y96_SLICE_X6Y96_D4 = CLBLM_R_X5Y96_SLICE_X6Y96_AQ;
  assign CLBLM_R_X5Y96_SLICE_X6Y96_D5 = CLBLM_R_X5Y99_SLICE_X7Y99_AQ;
  assign CLBLM_R_X3Y96_SLICE_X3Y96_A5 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X5Y96_SLICE_X6Y96_D6 = CLBLM_R_X5Y99_SLICE_X6Y99_AQ;
  assign CLBLM_R_X5Y96_SLICE_X6Y96_SR = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y96_SLICE_X3Y96_A6 = 1'b1;
  assign CLBLM_R_X3Y96_SLICE_X3Y96_B1 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X3Y96_SLICE_X3Y96_B2 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLM_R_X3Y96_SLICE_X3Y96_B3 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X3Y96_SLICE_X3Y96_B4 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X3Y96_SLICE_X3Y96_B5 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X3Y96_SLICE_X3Y96_B6 = 1'b1;
  assign CLBLM_R_X7Y87_SLICE_X9Y87_D4 = 1'b1;
  assign CLBLM_R_X7Y87_SLICE_X9Y87_D5 = 1'b1;
  assign CLBLM_R_X7Y87_SLICE_X9Y87_D6 = 1'b1;
  assign CLBLM_R_X3Y96_SLICE_X3Y96_C6 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO7;
  assign CLBLM_R_X5Y94_SLICE_X6Y94_B3 = CLBLM_R_X5Y94_SLICE_X7Y94_AO6;
  assign CLBLM_R_X5Y94_SLICE_X6Y94_B5 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO9;
  assign CLBLM_R_X5Y94_SLICE_X6Y94_B6 = CLBLM_R_X5Y94_SLICE_X6Y94_AO6;
  assign CLBLM_R_X7Y87_SLICE_X8Y87_A1 = CLBLM_R_X7Y90_SLICE_X9Y90_CQ;
  assign CLBLM_R_X7Y87_SLICE_X8Y87_A2 = CLBLM_R_X7Y87_SLICE_X8Y87_BQ;
  assign CLBLM_R_X5Y94_SLICE_X6Y94_BX = CLBLL_L_X4Y94_SLICE_X4Y94_CO6;
  assign CLBLM_R_X7Y87_SLICE_X8Y87_A3 = CLBLM_R_X7Y87_SLICE_X8Y87_AQ;
  assign CLBLM_R_X7Y87_SLICE_X8Y87_A4 = CLBLM_R_X7Y91_SLICE_X8Y91_AQ;
  assign CLBLM_R_X7Y87_SLICE_X8Y87_A5 = CLBLM_R_X7Y91_SLICE_X9Y91_AQ;
  assign CLBLM_R_X7Y87_SLICE_X8Y87_A6 = CLBLM_R_X7Y90_SLICE_X8Y90_CO6;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRL14 = CLBLM_R_X5Y90_SLICE_X6Y90_B5Q;
  assign CLBLL_L_X4Y93_SLICE_X4Y93_A1 = CLBLM_R_X5Y93_SLICE_X6Y93_F7AMUX_O;
  assign CLBLL_L_X4Y93_SLICE_X4Y93_A2 = CLBLM_R_X5Y93_SLICE_X6Y93_BQ;
  assign CLBLL_L_X4Y93_SLICE_X4Y93_A3 = CLBLL_L_X4Y91_SLICE_X5Y91_F7AMUX_O;
  assign CLBLL_L_X4Y93_SLICE_X4Y93_A4 = CLBLM_R_X3Y93_SLICE_X3Y93_CQ;
  assign CLBLL_L_X4Y93_SLICE_X4Y93_A5 = CLBLL_L_X4Y93_SLICE_X5Y93_CQ;
  assign CLBLL_L_X4Y93_SLICE_X4Y93_A6 = CLBLL_L_X4Y94_SLICE_X5Y94_CQ;
  assign CLBLM_R_X5Y94_SLICE_X6Y94_CE = CLBLL_L_X2Y92_SLICE_X1Y92_AO6;
  assign CLBLL_L_X4Y93_SLICE_X4Y93_AX = CLBLL_L_X2Y93_SLICE_X0Y93_F7AMUX_O;
  assign CLBLM_R_X7Y87_SLICE_X8Y87_B1 = 1'b1;
  assign CLBLL_L_X4Y93_SLICE_X4Y93_B1 = CLBLM_R_X5Y93_SLICE_X6Y93_F7AMUX_O;
  assign CLBLL_L_X4Y93_SLICE_X4Y93_B2 = CLBLL_L_X4Y95_SLICE_X4Y95_AQ;
  assign CLBLL_L_X4Y93_SLICE_X4Y93_B3 = CLBLL_L_X4Y92_SLICE_X4Y92_CQ;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRL15 = 1'b1;
  assign CLBLL_L_X4Y93_SLICE_X4Y93_B4 = CLBLL_L_X4Y93_SLICE_X4Y93_CQ;
  assign CLBLL_L_X4Y93_SLICE_X4Y93_B6 = CLBLL_L_X4Y91_SLICE_X5Y91_F7AMUX_O;
  assign CLBLL_L_X4Y93_SLICE_X4Y93_B5 = CLBLL_L_X4Y94_SLICE_X4Y94_AQ;
  assign CLBLM_R_X7Y87_SLICE_X8Y87_B2 = CLBLM_R_X7Y87_SLICE_X8Y87_BQ;
  assign CLBLL_L_X4Y93_SLICE_X4Y93_BX = CLBLM_R_X3Y94_SLICE_X2Y94_DO5;
  assign CLBLM_R_X7Y87_SLICE_X8Y87_B3 = CLBLM_R_X7Y87_SLICE_X8Y87_AQ;
  assign CLBLL_L_X4Y93_SLICE_X4Y93_C1 = CLBLL_L_X2Y97_SLICE_X0Y97_BO6;
  assign CLBLL_L_X4Y93_SLICE_X4Y93_C2 = CLBLM_R_X3Y98_SLICE_X2Y98_CO6;
  assign CLBLL_L_X4Y93_SLICE_X4Y93_C3 = CLBLL_L_X2Y97_SLICE_X1Y97_BO6;
  assign CLBLL_L_X4Y93_SLICE_X4Y93_C4 = CLBLM_R_X3Y93_SLICE_X2Y93_CO6;
  assign CLBLL_L_X4Y93_SLICE_X4Y93_C5 = CLBLM_R_X3Y99_SLICE_X2Y99_CO6;
  assign CLBLL_L_X4Y93_SLICE_X4Y93_C6 = 1'b1;
  assign CLBLL_L_X4Y93_SLICE_X4Y93_CE = CLBLL_L_X2Y93_SLICE_X1Y93_CO6;
  assign CLBLM_R_X7Y87_SLICE_X8Y87_B4 = CLBLM_R_X7Y91_SLICE_X8Y91_AQ;
  assign CLBLM_R_X7Y87_SLICE_X8Y87_B5 = CLBLM_R_X7Y91_SLICE_X9Y91_AQ;
  assign CLBLM_R_X5Y97_SLICE_X7Y97_A1 = CLBLM_R_X5Y98_SLICE_X6Y98_BO6;
  assign CLBLL_L_X4Y93_SLICE_X4Y93_D1 = CLBLM_R_X5Y93_SLICE_X6Y93_F7AMUX_O;
  assign CLBLL_L_X4Y93_SLICE_X4Y93_D2 = CLBLL_L_X4Y93_SLICE_X5Y93_CO6;
  assign CLBLL_L_X4Y93_SLICE_X4Y93_D3 = CLBLL_L_X4Y93_SLICE_X5Y93_DO6;
  assign CLBLL_L_X4Y93_SLICE_X4Y93_D4 = CLBLL_L_X4Y92_SLICE_X5Y92_CO6;
  assign CLBLL_L_X4Y93_SLICE_X4Y93_D5 = CLBLL_L_X2Y93_SLICE_X0Y93_F7AMUX_O;
  assign CLBLL_L_X4Y93_SLICE_X4Y93_D6 = CLBLL_L_X4Y92_SLICE_X5Y92_DO6;
  assign CLBLM_R_X5Y97_SLICE_X7Y97_A2 = CLBLM_R_X5Y98_SLICE_X6Y98_CO6;
  assign CLBLM_R_X5Y97_SLICE_X7Y97_A3 = CLBLM_R_X5Y97_SLICE_X6Y97_AO6;
  assign CLBLL_L_X4Y93_SLICE_X4Y93_DX = CLBLL_L_X4Y94_SLICE_X4Y94_CO6;
  assign CLBLM_R_X5Y97_SLICE_X7Y97_A4 = CLBLM_R_X5Y98_SLICE_X6Y98_DO6;
  assign CLBLM_R_X5Y97_SLICE_X7Y97_A5 = CLBLM_R_X5Y97_SLICE_X6Y97_DO6;
  assign CLBLM_R_X5Y97_SLICE_X7Y97_A6 = 1'b1;
  assign CLBLM_R_X5Y97_SLICE_X7Y97_B1 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X5Y97_SLICE_X7Y97_B2 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X5Y97_SLICE_X7Y97_B3 = CLBLM_R_X5Y95_SLICE_X6Y95_AQ;
  assign CLBLM_R_X5Y97_SLICE_X7Y97_B4 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X5Y97_SLICE_X7Y97_B5 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO3;
  assign CLBLM_R_X5Y97_SLICE_X7Y97_B6 = CLBLM_R_X5Y98_SLICE_X7Y98_CO6;
  assign CLBLM_R_X5Y97_SLICE_X7Y97_C1 = CLBLM_R_X5Y97_SLICE_X7Y97_AO6;
  assign CLBLM_R_X5Y97_SLICE_X7Y97_C2 = CLBLM_R_X5Y97_SLICE_X6Y97_AO6;
  assign CLBLM_R_X5Y94_SLICE_X6Y94_D2 = 1'b1;
  assign CLBLM_R_X5Y97_SLICE_X7Y97_C3 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X5Y97_SLICE_X7Y97_C4 = CLBLL_L_X4Y97_SLICE_X4Y97_BQ;
  assign CLBLM_R_X5Y97_SLICE_X7Y97_C5 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X5Y97_SLICE_X7Y97_C6 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO4;
  assign CLBLM_R_X5Y97_SLICE_X7Y97_D1 = CLBLM_R_X5Y97_SLICE_X6Y97_DO6;
  assign CLBLM_R_X5Y97_SLICE_X7Y97_D2 = CLBLM_R_X5Y97_SLICE_X6Y97_AO6;
  assign CLBLL_L_X4Y93_SLICE_X5Y93_A1 = CLBLM_R_X3Y96_SLICE_X3Y96_AO6;
  assign CLBLL_L_X4Y93_SLICE_X5Y93_A2 = CLBLM_R_X3Y93_SLICE_X3Y93_CQ;
  assign CLBLL_L_X4Y93_SLICE_X5Y93_A3 = CLBLL_L_X4Y93_SLICE_X5Y93_CQ;
  assign CLBLL_L_X4Y93_SLICE_X5Y93_A4 = CLBLM_R_X5Y93_SLICE_X6Y93_BQ;
  assign CLBLL_L_X4Y93_SLICE_X5Y93_A5 = CLBLL_L_X4Y91_SLICE_X4Y91_AO6;
  assign CLBLL_L_X4Y93_SLICE_X5Y93_A6 = CLBLL_L_X4Y94_SLICE_X5Y94_CQ;
  assign CLBLM_R_X5Y97_SLICE_X7Y97_D3 = CLBLM_R_X5Y97_SLICE_X6Y97_BO6;
  assign CLBLM_R_X5Y97_SLICE_X7Y97_D4 = CLBLM_R_X5Y98_SLICE_X6Y98_CO6;
  assign CLBLL_L_X4Y93_SLICE_X5Y93_AX = CLBLL_L_X4Y95_SLICE_X5Y95_DO6;
  assign CLBLM_R_X5Y97_SLICE_X7Y97_D5 = CLBLM_R_X5Y98_SLICE_X6Y98_BO6;
  assign CLBLL_L_X4Y93_SLICE_X5Y93_B1 = CLBLM_R_X3Y96_SLICE_X3Y96_AO6;
  assign CLBLL_L_X4Y93_SLICE_X5Y93_B2 = CLBLL_L_X4Y93_SLICE_X4Y93_CQ;
  assign CLBLL_L_X4Y93_SLICE_X5Y93_B3 = CLBLL_L_X4Y94_SLICE_X4Y94_AQ;
  assign CLBLL_L_X4Y93_SLICE_X5Y93_B4 = CLBLL_L_X4Y92_SLICE_X4Y92_CQ;
  assign CLBLL_L_X4Y93_SLICE_X5Y93_B5 = CLBLL_L_X4Y95_SLICE_X4Y95_AQ;
  assign CLBLL_L_X4Y93_SLICE_X5Y93_B6 = CLBLL_L_X4Y91_SLICE_X4Y91_AO6;
  assign CLBLM_R_X5Y97_SLICE_X6Y97_A1 = CLBLM_R_X7Y97_SLICE_X9Y97_AQ;
  assign CLBLM_R_X5Y97_SLICE_X6Y97_A2 = CLBLM_R_X7Y97_SLICE_X9Y97_A5Q;
  assign CLBLL_L_X4Y93_SLICE_X5Y93_BX = CLBLL_L_X4Y93_SLICE_X4Y93_CO5;
  assign CLBLM_R_X5Y97_SLICE_X6Y97_A3 = CLBLM_R_X7Y97_SLICE_X9Y97_BQ;
  assign CLBLL_L_X4Y93_SLICE_X5Y93_C1 = CLBLL_L_X4Y91_SLICE_X5Y91_BO6;
  assign CLBLL_L_X4Y93_SLICE_X5Y93_C2 = CLBLL_L_X4Y91_SLICE_X5Y91_CO6;
  assign CLBLL_L_X4Y93_SLICE_X5Y93_C3 = CLBLM_R_X3Y93_SLICE_X3Y93_AQ;
  assign CLBLL_L_X4Y93_SLICE_X5Y93_C4 = CLBLM_R_X5Y94_SLICE_X7Y94_AO5;
  assign CLBLL_L_X4Y93_SLICE_X5Y93_C5 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO8;
  assign CLBLL_L_X4Y93_SLICE_X5Y93_C6 = CLBLL_L_X4Y94_SLICE_X5Y94_BQ;
  assign CLBLL_L_X4Y93_SLICE_X5Y93_CE = CLBLL_L_X2Y93_SLICE_X1Y93_DO6;
  assign CLBLM_R_X5Y97_SLICE_X6Y97_AX = CLBLM_R_X5Y96_SLICE_X7Y96_BQ;
  assign CLBLM_R_X5Y97_SLICE_X6Y97_B1 = CLBLM_R_X7Y97_SLICE_X9Y97_AQ;
  assign CLBLM_R_X5Y97_SLICE_X6Y97_B2 = CLBLM_R_X7Y97_SLICE_X9Y97_A5Q;
  assign CLBLM_R_X5Y97_SLICE_X6Y97_B3 = CLBLM_R_X7Y97_SLICE_X9Y97_BQ;
  assign CLBLM_R_X5Y97_SLICE_X6Y97_B4 = CLBLM_R_X7Y97_SLICE_X9Y97_B5Q;
  assign CLBLL_L_X4Y93_SLICE_X5Y93_CX = CLBLL_L_X4Y93_SLICE_X4Y93_CO6;
  assign CLBLM_R_X5Y97_SLICE_X6Y97_B5 = 1'b0;
  assign CLBLL_L_X4Y93_SLICE_X5Y93_D1 = CLBLL_L_X4Y91_SLICE_X4Y91_AQ;
  assign CLBLL_L_X4Y93_SLICE_X5Y93_D2 = CLBLL_L_X4Y91_SLICE_X5Y91_CO6;
  assign CLBLL_L_X4Y93_SLICE_X5Y93_D3 = CLBLM_R_X5Y94_SLICE_X6Y94_AQ;
  assign CLBLL_L_X4Y93_SLICE_X5Y93_D4 = CLBLM_R_X5Y94_SLICE_X7Y94_AO5;
  assign CLBLL_L_X4Y93_SLICE_X5Y93_D5 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO8;
  assign CLBLL_L_X4Y93_SLICE_X5Y93_D6 = CLBLL_L_X4Y91_SLICE_X5Y91_BO6;
  assign CLBLM_R_X5Y97_SLICE_X6Y97_C1 = CLBLM_R_X7Y97_SLICE_X9Y97_AQ;
  assign CLBLM_R_X5Y97_SLICE_X6Y97_C2 = CLBLM_R_X7Y97_SLICE_X9Y97_A5Q;
  assign CLBLL_L_X4Y93_SLICE_X5Y93_DX = CLBLL_L_X4Y94_SLICE_X4Y94_CO6;
  assign CLBLM_R_X5Y97_SLICE_X6Y97_C3 = CLBLM_R_X7Y97_SLICE_X9Y97_BQ;
  assign CLBLM_R_X5Y97_SLICE_X6Y97_C4 = CLBLM_R_X7Y97_SLICE_X9Y97_B5Q;
  assign CLBLM_R_X5Y97_SLICE_X6Y97_C5 = 1'b0;
  assign CLBLM_R_X5Y97_SLICE_X6Y97_C6 = 1'b1;
  assign CLBLM_R_X5Y97_SLICE_X6Y97_CE = CLBLL_L_X4Y97_SLICE_X5Y97_DO6;
  assign CLBLM_R_X5Y97_SLICE_X6Y97_CX = CLBLM_R_X7Y96_SLICE_X8Y96_AQ;
  assign CLBLM_R_X5Y97_SLICE_X6Y97_D1 = CLBLM_R_X7Y97_SLICE_X9Y97_AQ;
  assign CLBLM_R_X5Y97_SLICE_X6Y97_D2 = CLBLM_R_X7Y97_SLICE_X9Y97_A5Q;
  assign CLBLM_R_X5Y97_SLICE_X6Y97_D3 = CLBLM_R_X7Y97_SLICE_X9Y97_BQ;
  assign CLBLM_R_X5Y97_SLICE_X6Y97_D4 = CLBLM_R_X7Y97_SLICE_X9Y97_B5Q;
  assign CLBLM_R_X5Y97_SLICE_X6Y97_D5 = 1'b0;
  assign CLBLM_R_X5Y97_SLICE_X6Y97_D6 = 1'b1;
  assign CLBLM_R_X5Y97_SLICE_X6Y97_DI = CLBLM_R_X5Y98_SLICE_X6Y98_CO6;
  assign CLBLM_R_X5Y97_SLICE_X6Y97_DX = CLBLM_R_X5Y96_SLICE_X7Y96_AQ;
  assign CLBLM_R_X7Y87_SLICE_X8Y87_D4 = 1'b1;
  assign CLBLM_R_X7Y87_SLICE_X8Y87_D5 = 1'b1;
  assign CLBLM_R_X7Y87_SLICE_X8Y87_D6 = 1'b1;
  assign CLBLM_R_X3Y96_SLICE_X2Y96_CX = CLBLL_L_X2Y96_SLICE_X1Y96_DO6;
  assign CLBLM_R_X3Y96_SLICE_X2Y96_D1 = CLBLM_R_X3Y97_SLICE_X3Y97_CO6;
  assign CLBLM_R_X3Y96_SLICE_X2Y96_D2 = CLBLL_L_X4Y98_SLICE_X4Y98_DO6;
  assign CLBLM_R_X3Y96_SLICE_X2Y96_D3 = CLBLM_R_X3Y97_SLICE_X3Y97_DO6;
  assign CLBLM_R_X3Y96_SLICE_X2Y96_D4 = CLBLM_R_X3Y98_SLICE_X3Y98_DO6;
  assign CLBLM_R_X3Y96_SLICE_X2Y96_D5 = CLBLL_L_X4Y98_SLICE_X5Y98_DO6;
  assign CLBLM_R_X3Y96_SLICE_X2Y96_D6 = 1'b1;
  assign CLBLM_R_X3Y96_SLICE_X2Y96_DI = CLBLL_L_X4Y98_SLICE_X4Y98_DO6;
  assign CLBLL_L_X4Y94_SLICE_X4Y94_A1 = CLBLM_R_X5Y94_SLICE_X7Y94_DO6;
  assign CLBLL_L_X4Y94_SLICE_X4Y94_A2 = CLBLL_L_X2Y97_SLICE_X1Y97_BO6;
  assign CLBLL_L_X4Y94_SLICE_X4Y94_A3 = CLBLL_L_X4Y94_SLICE_X5Y94_DO6;
  assign CLBLL_L_X4Y94_SLICE_X4Y94_A4 = CLBLM_R_X3Y98_SLICE_X2Y98_CO6;
  assign CLBLL_L_X4Y94_SLICE_X4Y94_A5 = CLBLM_R_X3Y93_SLICE_X2Y93_CO6;
  assign CLBLL_L_X4Y94_SLICE_X4Y94_A6 = CLBLM_R_X5Y94_SLICE_X6Y94_BO6;
  assign CLBLL_L_X4Y94_SLICE_X4Y94_B1 = CLBLM_R_X5Y94_SLICE_X7Y94_DO6;
  assign CLBLL_L_X4Y94_SLICE_X4Y94_B2 = CLBLL_L_X4Y94_SLICE_X5Y94_DO6;
  assign CLBLL_L_X4Y94_SLICE_X4Y94_B3 = CLBLM_R_X3Y93_SLICE_X2Y93_CO6;
  assign CLBLL_L_X4Y94_SLICE_X4Y94_B4 = CLBLL_L_X2Y97_SLICE_X1Y97_CO6;
  assign CLBLL_L_X4Y94_SLICE_X4Y94_B5 = CLBLL_L_X4Y96_SLICE_X4Y96_CO6;
  assign CLBLL_L_X4Y94_SLICE_X4Y94_B6 = CLBLM_R_X5Y94_SLICE_X6Y94_BO6;
  assign CLBLL_L_X4Y94_SLICE_X4Y94_C1 = CLBLM_R_X3Y93_SLICE_X2Y93_CO6;
  assign CLBLL_L_X4Y94_SLICE_X4Y94_C2 = CLBLL_L_X2Y97_SLICE_X1Y97_CO6;
  assign CLBLL_L_X4Y94_SLICE_X4Y94_C3 = CLBLL_L_X2Y96_SLICE_X1Y96_DO6;
  assign CLBLL_L_X4Y94_SLICE_X4Y94_C4 = CLBLL_L_X4Y96_SLICE_X4Y96_CO6;
  assign CLBLL_L_X4Y94_SLICE_X4Y94_C5 = CLBLM_R_X3Y96_SLICE_X3Y96_DO6;
  assign CLBLL_L_X4Y94_SLICE_X4Y94_C6 = 1'b1;
  assign CLBLL_L_X4Y94_SLICE_X4Y94_D1 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLL_L_X4Y94_SLICE_X4Y94_D2 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO10;
  assign CLBLL_L_X4Y94_SLICE_X4Y94_D3 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLL_L_X4Y94_SLICE_X4Y94_D4 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLL_L_X4Y94_SLICE_X4Y94_D5 = CLBLL_L_X4Y96_SLICE_X4Y96_DO6;
  assign CLBLL_L_X4Y94_SLICE_X4Y94_D6 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X5Y98_SLICE_X7Y98_A1 = 1'b1;
  assign CLBLM_R_X5Y98_SLICE_X7Y98_A2 = CLBLM_R_X5Y98_SLICE_X6Y98_BO6;
  assign CLBLL_L_X4Y94_SLICE_X4Y94_SR = CLBLM_R_X5Y92_SLICE_X7Y92_AO6;
  assign CLBLM_R_X5Y98_SLICE_X7Y98_A3 = CLBLM_R_X5Y98_SLICE_X6Y98_CO6;
  assign CLBLM_R_X5Y98_SLICE_X7Y98_A4 = CLBLM_R_X5Y98_SLICE_X6Y98_DO6;
  assign CLBLM_R_X5Y98_SLICE_X7Y98_A5 = 1'b1;
  assign CLBLM_R_X5Y98_SLICE_X7Y98_A6 = 1'b1;
  assign CLBLM_R_X5Y98_SLICE_X7Y98_B1 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X5Y98_SLICE_X7Y98_B2 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X5Y98_SLICE_X7Y98_B3 = CLBLM_R_X5Y98_SLICE_X6Y98_CO6;
  assign CLBLM_R_X5Y98_SLICE_X7Y98_B4 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO2;
  assign CLBLM_R_X5Y98_SLICE_X7Y98_B5 = CLBLM_R_X5Y98_SLICE_X7Y98_AO6;
  assign CLBLM_R_X5Y98_SLICE_X7Y98_B6 = CLBLL_L_X4Y97_SLICE_X4Y97_BQ;
  assign CLBLM_R_X5Y98_SLICE_X7Y98_C1 = CLBLL_L_X4Y97_SLICE_X4Y97_BQ;
  assign CLBLM_R_X5Y98_SLICE_X7Y98_C2 = CLBLM_R_X5Y97_SLICE_X6Y97_DO6;
  assign CLBLM_R_X5Y98_SLICE_X7Y98_C3 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO3;
  assign CLBLM_R_X5Y98_SLICE_X7Y98_C4 = CLBLM_R_X5Y98_SLICE_X7Y98_AO5;
  assign CLBLM_R_X5Y98_SLICE_X7Y98_C5 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X5Y98_SLICE_X7Y98_C6 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLL_L_X4Y94_SLICE_X5Y94_A1 = CLBLL_L_X4Y93_SLICE_X5Y93_DQ;
  assign CLBLL_L_X4Y94_SLICE_X5Y94_A2 = CLBLL_L_X4Y94_SLICE_X5Y94_DQ;
  assign CLBLL_L_X4Y94_SLICE_X5Y94_A3 = CLBLM_R_X5Y93_SLICE_X6Y93_F7AMUX_O;
  assign CLBLL_L_X4Y94_SLICE_X5Y94_A4 = CLBLM_R_X3Y93_SLICE_X3Y93_DQ;
  assign CLBLL_L_X4Y94_SLICE_X5Y94_A5 = CLBLL_L_X4Y91_SLICE_X5Y91_F7AMUX_O;
  assign CLBLL_L_X4Y94_SLICE_X5Y94_A6 = CLBLL_L_X4Y92_SLICE_X5Y92_CQ;
  assign CLBLM_R_X5Y98_SLICE_X7Y98_D1 = CLBLM_R_X5Y97_SLICE_X7Y97_CO6;
  assign CLBLL_L_X4Y94_SLICE_X5Y94_AX = CLBLL_L_X2Y93_SLICE_X0Y93_F7AMUX_O;
  assign CLBLM_R_X5Y98_SLICE_X7Y98_D2 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO4;
  assign CLBLL_L_X4Y94_SLICE_X5Y94_B1 = CLBLL_L_X4Y92_SLICE_X4Y92_B5Q;
  assign CLBLL_L_X4Y94_SLICE_X5Y94_B2 = CLBLL_L_X4Y93_SLICE_X4Y93_DQ;
  assign CLBLL_L_X4Y94_SLICE_X5Y94_B3 = CLBLM_R_X5Y93_SLICE_X6Y93_F7AMUX_O;
  assign CLBLL_L_X4Y94_SLICE_X5Y94_B4 = CLBLL_L_X4Y94_SLICE_X4Y94_BQ;
  assign CLBLL_L_X4Y94_SLICE_X5Y94_B5 = CLBLL_L_X4Y91_SLICE_X5Y91_F7AMUX_O;
  assign CLBLL_L_X4Y94_SLICE_X5Y94_B6 = CLBLM_R_X5Y94_SLICE_X6Y94_BQ;
  assign CLBLM_R_X5Y98_SLICE_X6Y98_A1 = CLBLM_R_X7Y97_SLICE_X9Y97_AQ;
  assign CLBLM_R_X5Y98_SLICE_X6Y98_A2 = CLBLM_R_X7Y97_SLICE_X9Y97_A5Q;
  assign CLBLL_L_X4Y94_SLICE_X5Y94_BX = CLBLL_L_X4Y93_SLICE_X4Y93_CO5;
  assign CLBLM_R_X5Y98_SLICE_X6Y98_A3 = CLBLM_R_X7Y97_SLICE_X9Y97_BQ;
  assign CLBLL_L_X4Y94_SLICE_X5Y94_C1 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO14;
  assign CLBLL_L_X4Y94_SLICE_X5Y94_C2 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO11;
  assign CLBLL_L_X4Y94_SLICE_X5Y94_C3 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO15;
  assign CLBLL_L_X4Y94_SLICE_X5Y94_C4 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO13;
  assign CLBLL_L_X4Y94_SLICE_X5Y94_C5 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO12;
  assign CLBLL_L_X4Y94_SLICE_X5Y94_C6 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO8;
  assign CLBLL_L_X4Y94_SLICE_X5Y94_CE = CLBLM_R_X3Y93_SLICE_X3Y93_CO6;
  assign CLBLM_R_X5Y98_SLICE_X6Y98_B1 = CLBLM_R_X7Y97_SLICE_X9Y97_AQ;
  assign CLBLM_R_X5Y98_SLICE_X6Y98_B2 = CLBLM_R_X7Y97_SLICE_X9Y97_A5Q;
  assign CLBLM_R_X5Y98_SLICE_X6Y98_B3 = CLBLM_R_X7Y97_SLICE_X9Y97_BQ;
  assign CLBLM_R_X5Y98_SLICE_X6Y98_B4 = CLBLM_R_X7Y97_SLICE_X9Y97_B5Q;
  assign CLBLM_R_X5Y98_SLICE_X6Y98_B5 = 1'b0;
  assign CLBLL_L_X4Y94_SLICE_X5Y94_CX = CLBLL_L_X4Y93_SLICE_X4Y93_CO6;
  assign CLBLM_R_X5Y98_SLICE_X6Y98_B6 = 1'b1;
  assign CLBLL_L_X4Y94_SLICE_X5Y94_D1 = CLBLM_R_X5Y94_SLICE_X7Y94_AO6;
  assign CLBLL_L_X4Y94_SLICE_X5Y94_D2 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLL_L_X4Y94_SLICE_X5Y94_D3 = CLBLL_L_X4Y94_SLICE_X4Y94_DO6;
  assign CLBLL_L_X4Y94_SLICE_X5Y94_D4 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO10;
  assign CLBLL_L_X4Y94_SLICE_X5Y94_D5 = CLBLM_R_X5Y94_SLICE_X7Y94_AO5;
  assign CLBLL_L_X4Y94_SLICE_X5Y94_D6 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLM_R_X5Y98_SLICE_X6Y98_BX = CLBLM_R_X5Y99_SLICE_X7Y99_AQ;
  assign CLBLM_R_X5Y98_SLICE_X6Y98_C1 = CLBLM_R_X7Y97_SLICE_X9Y97_AQ;
  assign CLBLL_L_X4Y94_SLICE_X5Y94_DX = CLBLL_L_X4Y94_SLICE_X4Y94_CO6;
  assign CLBLM_R_X5Y98_SLICE_X6Y98_C2 = CLBLM_R_X7Y97_SLICE_X9Y97_A5Q;
  assign CLBLM_R_X5Y98_SLICE_X6Y98_C3 = CLBLM_R_X7Y97_SLICE_X9Y97_BQ;
  assign CLBLM_R_X5Y98_SLICE_X6Y98_C4 = CLBLM_R_X7Y97_SLICE_X9Y97_B5Q;
  assign CLBLM_R_X5Y98_SLICE_X6Y98_C5 = 1'b0;
  assign CLBLM_R_X5Y98_SLICE_X6Y98_C6 = 1'b1;
  assign CLBLM_R_X5Y98_SLICE_X6Y98_CE = CLBLL_L_X4Y97_SLICE_X5Y97_DO6;
  assign CLBLM_R_X5Y98_SLICE_X6Y98_CX = CLBLM_R_X5Y99_SLICE_X6Y99_AQ;
  assign CLBLM_R_X5Y98_SLICE_X6Y98_D1 = CLBLM_R_X7Y97_SLICE_X9Y97_AQ;
  assign CLBLM_R_X5Y98_SLICE_X6Y98_D2 = CLBLM_R_X7Y97_SLICE_X9Y97_A5Q;
  assign CLBLM_R_X5Y98_SLICE_X6Y98_D3 = CLBLM_R_X7Y97_SLICE_X9Y97_BQ;
  assign CLBLM_R_X5Y98_SLICE_X6Y98_D4 = CLBLM_R_X7Y97_SLICE_X9Y97_B5Q;
  assign CLBLM_R_X5Y98_SLICE_X6Y98_D5 = 1'b0;
  assign CLBLM_R_X5Y98_SLICE_X6Y98_D6 = 1'b1;
  assign CLBLM_R_X5Y98_SLICE_X6Y98_DI = CLBLL_L_X4Y97_SLICE_X5Y97_DO6;
  assign CLBLM_R_X5Y98_SLICE_X6Y98_DX = CLBLM_R_X7Y99_SLICE_X8Y99_AQ;
  assign CLBLM_L_X8Y89_SLICE_X11Y89_A1 = 1'b1;
  assign CLBLM_L_X8Y89_SLICE_X11Y89_A2 = 1'b1;
  assign CLBLM_L_X8Y89_SLICE_X11Y89_A3 = 1'b1;
  assign CLBLM_L_X8Y89_SLICE_X11Y89_A4 = 1'b1;
  assign CLBLM_L_X8Y89_SLICE_X11Y89_A5 = 1'b1;
  assign CLBLM_L_X8Y89_SLICE_X11Y89_A6 = 1'b1;
  assign CLBLM_L_X8Y89_SLICE_X11Y89_B1 = 1'b1;
  assign CLBLM_L_X8Y89_SLICE_X11Y89_B2 = 1'b1;
  assign CLBLM_L_X8Y89_SLICE_X11Y89_B3 = 1'b1;
  assign CLBLM_L_X8Y89_SLICE_X11Y89_B4 = 1'b1;
  assign CLBLM_L_X8Y89_SLICE_X11Y89_B5 = 1'b1;
  assign CLBLM_L_X8Y89_SLICE_X11Y89_B6 = 1'b1;
  assign CLBLM_L_X8Y89_SLICE_X11Y89_C1 = 1'b1;
  assign CLBLM_L_X8Y89_SLICE_X11Y89_C2 = 1'b1;
  assign CLBLM_L_X8Y89_SLICE_X11Y89_C3 = 1'b1;
  assign CLBLM_L_X8Y89_SLICE_X11Y89_C4 = 1'b1;
  assign CLBLM_L_X8Y89_SLICE_X11Y89_C5 = 1'b1;
  assign CLBLM_L_X8Y89_SLICE_X11Y89_C6 = 1'b1;
  assign CLBLM_L_X8Y89_SLICE_X11Y89_D1 = 1'b1;
  assign CLBLM_L_X8Y89_SLICE_X11Y89_D2 = 1'b1;
  assign CLBLM_L_X8Y89_SLICE_X11Y89_D3 = 1'b1;
  assign CLBLM_L_X8Y89_SLICE_X11Y89_D4 = 1'b1;
  assign CLBLM_L_X8Y89_SLICE_X11Y89_D5 = 1'b1;
  assign CLBLM_L_X8Y89_SLICE_X11Y89_D6 = 1'b1;
  assign CLBLM_L_X8Y89_SLICE_X10Y89_A1 = CLBLM_L_X8Y89_SLICE_X10Y89_CQ;
  assign CLBLM_L_X8Y89_SLICE_X10Y89_A2 = CLBLM_L_X8Y89_SLICE_X10Y89_BQ;
  assign CLBLM_L_X8Y89_SLICE_X10Y89_A3 = CLBLM_L_X8Y89_SLICE_X10Y89_AQ;
  assign CLBLM_L_X8Y89_SLICE_X10Y89_A4 = 1'b1;
  assign CLBLM_L_X8Y89_SLICE_X10Y89_A5 = CLBLM_L_X8Y89_SLICE_X10Y89_A5Q;
  assign CLBLM_L_X8Y89_SLICE_X10Y89_A6 = 1'b1;
  assign CLBLM_L_X8Y89_SLICE_X10Y89_B1 = CLBLM_L_X8Y89_SLICE_X10Y89_CQ;
  assign CLBLM_L_X8Y89_SLICE_X10Y89_B2 = CLBLM_L_X8Y89_SLICE_X10Y89_BQ;
  assign CLBLM_L_X8Y89_SLICE_X10Y89_B3 = 1'b1;
  assign CLBLM_L_X8Y89_SLICE_X10Y89_B4 = 1'b1;
  assign CLBLM_L_X8Y89_SLICE_X10Y89_B5 = 1'b1;
  assign CLBLM_L_X8Y89_SLICE_X10Y89_B6 = 1'b1;
  assign CLBLM_L_X8Y89_SLICE_X10Y89_C1 = 1'b1;
  assign CLBLM_L_X8Y89_SLICE_X10Y89_C2 = CLBLM_L_X8Y89_SLICE_X10Y89_CQ;
  assign CLBLM_L_X8Y89_SLICE_X10Y89_C3 = 1'b1;
  assign CLBLM_L_X8Y89_SLICE_X10Y89_C4 = 1'b1;
  assign CLBLM_L_X8Y89_SLICE_X10Y89_C5 = 1'b1;
  assign CLBLM_L_X8Y89_SLICE_X10Y89_C6 = 1'b1;
  assign CLBLM_L_X8Y89_SLICE_X10Y89_CE = CLBLM_R_X7Y88_SLICE_X8Y88_BO6;
  assign CLBLM_L_X8Y89_SLICE_X10Y89_CLK = CLBLM_R_X7Y88_SLICE_X8Y88_AQ;
  assign LIOB33_SING_X0Y100_IOB_X0Y100_O = CLBLM_R_X7Y91_SLICE_X8Y91_BO6;
  assign CLBLM_L_X8Y89_SLICE_X10Y89_D1 = 1'b1;
  assign CLBLM_L_X8Y89_SLICE_X10Y89_D2 = 1'b1;
  assign CLBLM_L_X8Y89_SLICE_X10Y89_D3 = 1'b1;
  assign CLBLM_L_X8Y89_SLICE_X10Y89_D4 = 1'b1;
  assign CLBLM_L_X8Y89_SLICE_X10Y89_D5 = 1'b1;
  assign CLBLM_L_X8Y89_SLICE_X10Y89_D6 = 1'b1;
  assign CLBLM_L_X8Y89_SLICE_X10Y89_SR = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y95_SLICE_X4Y95_A1 = CLBLL_L_X4Y95_SLICE_X5Y95_CO6;
  assign CLBLL_L_X4Y95_SLICE_X4Y95_A2 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLL_L_X4Y95_SLICE_X4Y95_A3 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLL_L_X4Y95_SLICE_X4Y95_A4 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLL_L_X4Y95_SLICE_X4Y95_A5 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLL_L_X4Y95_SLICE_X4Y95_A6 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLL_L_X4Y95_SLICE_X4Y95_AX = CLBLL_L_X4Y93_SLICE_X4Y93_CO6;
  assign CLBLL_L_X4Y95_SLICE_X4Y95_B1 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLL_L_X4Y95_SLICE_X4Y95_B2 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLL_L_X4Y95_SLICE_X4Y95_B3 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLL_L_X4Y95_SLICE_X4Y95_B4 = CLBLL_L_X4Y91_SLICE_X4Y91_AO5;
  assign CLBLL_L_X4Y95_SLICE_X4Y95_B5 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO3;
  assign CLBLL_L_X4Y95_SLICE_X4Y95_B6 = CLBLL_L_X4Y93_SLICE_X5Y93_F7AMUX_O;
  assign CLBLL_L_X4Y95_SLICE_X4Y95_C1 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLL_L_X4Y95_SLICE_X4Y95_C2 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLL_L_X4Y95_SLICE_X4Y95_C3 = CLBLM_R_X3Y93_SLICE_X2Y93_F7AMUX_O;
  assign CLBLL_L_X4Y95_SLICE_X4Y95_C4 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLL_L_X4Y95_SLICE_X4Y95_C5 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO1;
  assign CLBLL_L_X4Y95_SLICE_X4Y95_C6 = CLBLL_L_X4Y91_SLICE_X4Y91_AO5;
  assign CLBLL_L_X4Y95_SLICE_X4Y95_CE = CLBLL_L_X2Y92_SLICE_X1Y92_AO6;
  assign CLBLL_L_X4Y95_SLICE_X4Y95_D1 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLL_L_X4Y95_SLICE_X4Y95_D2 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLL_L_X4Y95_SLICE_X4Y95_D3 = CLBLL_L_X4Y92_SLICE_X5Y92_F7AMUX_O;
  assign CLBLL_L_X4Y95_SLICE_X4Y95_D4 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO0;
  assign CLBLL_L_X4Y95_SLICE_X4Y95_D5 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLL_L_X4Y95_SLICE_X4Y95_D6 = CLBLL_L_X4Y91_SLICE_X4Y91_AO5;
  assign CLBLM_R_X5Y99_SLICE_X7Y99_A1 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLM_R_X5Y99_SLICE_X7Y99_A2 = CLBLM_R_X5Y99_SLICE_X6Y99_BO6;
  assign CLBLM_R_X5Y99_SLICE_X7Y99_A3 = CLBLM_R_X7Y98_SLICE_X8Y98_F7AMUX_O;
  assign CLBLM_R_X5Y99_SLICE_X7Y99_A4 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X5Y99_SLICE_X7Y99_A5 = CLBLM_R_X5Y99_SLICE_X7Y99_BO5;
  assign CLBLM_R_X5Y99_SLICE_X7Y99_A6 = CLBLM_R_X5Y99_SLICE_X7Y99_CO6;
  assign CLBLM_R_X5Y99_SLICE_X7Y99_B1 = 1'b1;
  assign CLBLM_R_X5Y99_SLICE_X7Y99_B2 = 1'b1;
  assign CLBLM_R_X5Y99_SLICE_X7Y99_B3 = CLBLM_R_X5Y99_SLICE_X7Y99_AQ;
  assign CLBLM_R_X5Y99_SLICE_X7Y99_B4 = CLBLM_R_X7Y99_SLICE_X8Y99_AQ;
  assign CLBLM_R_X5Y99_SLICE_X7Y99_B5 = CLBLM_R_X5Y99_SLICE_X6Y99_AQ;
  assign CLBLM_R_X5Y99_SLICE_X7Y99_B6 = 1'b1;
  assign CLBLM_R_X5Y99_SLICE_X7Y99_C1 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X5Y99_SLICE_X7Y99_C2 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO1;
  assign CLBLM_R_X5Y99_SLICE_X7Y99_C3 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X5Y99_SLICE_X7Y99_C4 = CLBLM_R_X5Y95_SLICE_X6Y95_AQ;
  assign CLBLM_R_X5Y99_SLICE_X7Y99_C5 = CLBLM_R_X5Y99_SLICE_X7Y99_DO6;
  assign CLBLM_R_X5Y99_SLICE_X7Y99_C6 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X5Y99_SLICE_X7Y99_CE = CLBLM_R_X7Y99_SLICE_X9Y99_DO6;
  assign CLBLL_L_X4Y95_SLICE_X5Y95_A1 = CLBLL_L_X4Y93_SLICE_X5Y93_DQ;
  assign CLBLL_L_X4Y95_SLICE_X5Y95_A2 = CLBLL_L_X4Y94_SLICE_X5Y94_DQ;
  assign CLBLL_L_X4Y95_SLICE_X5Y95_A3 = CLBLL_L_X4Y91_SLICE_X4Y91_AO6;
  assign CLBLL_L_X4Y95_SLICE_X5Y95_A4 = CLBLM_R_X3Y96_SLICE_X3Y96_AO6;
  assign CLBLL_L_X4Y95_SLICE_X5Y95_A5 = CLBLL_L_X4Y92_SLICE_X5Y92_CQ;
  assign CLBLL_L_X4Y95_SLICE_X5Y95_A6 = CLBLM_R_X3Y93_SLICE_X3Y93_DQ;
  assign CLBLL_L_X4Y95_SLICE_X5Y95_AX = CLBLL_L_X4Y95_SLICE_X5Y95_DO6;
  assign CLBLM_R_X5Y99_SLICE_X7Y99_D1 = CLBLL_L_X4Y97_SLICE_X4Y97_BQ;
  assign CLBLL_L_X4Y95_SLICE_X5Y95_B1 = CLBLL_L_X4Y93_SLICE_X4Y93_DQ;
  assign CLBLL_L_X4Y95_SLICE_X5Y95_B2 = CLBLL_L_X4Y94_SLICE_X4Y94_BQ;
  assign CLBLL_L_X4Y95_SLICE_X5Y95_B3 = CLBLL_L_X4Y91_SLICE_X4Y91_AO6;
  assign CLBLL_L_X4Y95_SLICE_X5Y95_B4 = CLBLM_R_X3Y96_SLICE_X3Y96_AO6;
  assign CLBLL_L_X4Y95_SLICE_X5Y95_B5 = CLBLM_R_X5Y94_SLICE_X6Y94_BQ;
  assign CLBLL_L_X4Y95_SLICE_X5Y95_B6 = CLBLL_L_X4Y92_SLICE_X4Y92_B5Q;
  assign CLBLM_R_X5Y99_SLICE_X7Y99_D2 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO1;
  assign CLBLM_R_X5Y99_SLICE_X7Y99_D3 = CLBLM_R_X5Y98_SLICE_X6Y98_DO6;
  assign CLBLM_R_X5Y99_SLICE_X7Y99_D4 = CLBLM_R_X5Y98_SLICE_X6Y98_BO6;
  assign CLBLL_L_X4Y95_SLICE_X5Y95_C1 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLL_L_X4Y95_SLICE_X5Y95_C2 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLL_L_X4Y95_SLICE_X5Y95_C3 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO6;
  assign CLBLL_L_X4Y95_SLICE_X5Y95_C4 = CLBLL_L_X4Y95_SLICE_X5Y95_F7AMUX_O;
  assign CLBLL_L_X4Y95_SLICE_X5Y95_C5 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLL_L_X4Y95_SLICE_X5Y95_C6 = CLBLL_L_X4Y91_SLICE_X4Y91_AO5;
  assign CLBLM_R_X5Y99_SLICE_X6Y99_A1 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLM_R_X5Y99_SLICE_X6Y99_A2 = CLBLM_R_X5Y99_SLICE_X7Y99_BO6;
  assign CLBLM_R_X5Y99_SLICE_X6Y99_A3 = CLBLL_L_X4Y98_SLICE_X5Y98_AO6;
  assign CLBLM_R_X5Y99_SLICE_X6Y99_A4 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X5Y99_SLICE_X6Y99_A5 = CLBLM_R_X7Y98_SLICE_X8Y98_F7AMUX_O;
  assign CLBLM_R_X5Y99_SLICE_X6Y99_A6 = CLBLM_R_X5Y99_SLICE_X6Y99_CO6;
  assign CLBLM_R_X5Y99_SLICE_X6Y99_B1 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLL_L_X4Y95_SLICE_X5Y95_D1 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLL_L_X4Y95_SLICE_X5Y95_D2 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLL_L_X4Y95_SLICE_X5Y95_D3 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO7;
  assign CLBLL_L_X4Y95_SLICE_X5Y95_D4 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLL_L_X4Y95_SLICE_X5Y95_D5 = 1'b1;
  assign CLBLL_L_X4Y95_SLICE_X5Y95_D6 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X5Y99_SLICE_X6Y99_B2 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X5Y99_SLICE_X6Y99_B3 = CLBLL_L_X4Y97_SLICE_X4Y97_BQ;
  assign CLBLM_R_X5Y99_SLICE_X6Y99_B4 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO1;
  assign CLBLM_R_X5Y99_SLICE_X6Y99_B5 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X5Y99_SLICE_X6Y99_B6 = CLBLM_R_X5Y95_SLICE_X6Y95_AQ;
  assign CLBLM_R_X5Y99_SLICE_X6Y99_C1 = CLBLL_L_X4Y97_SLICE_X4Y97_BQ;
  assign CLBLM_R_X5Y99_SLICE_X6Y99_C2 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO2;
  assign CLBLM_R_X5Y99_SLICE_X6Y99_C3 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X5Y99_SLICE_X6Y99_C4 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X5Y99_SLICE_X6Y99_C5 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X5Y99_SLICE_X6Y99_C6 = CLBLM_R_X5Y95_SLICE_X6Y95_AQ;
  assign CLBLM_R_X5Y99_SLICE_X6Y99_CE = CLBLM_R_X7Y99_SLICE_X9Y99_DO6;
  assign CLBLM_R_X5Y99_SLICE_X6Y99_D1 = 1'b1;
  assign CLBLM_R_X5Y99_SLICE_X6Y99_D2 = 1'b1;
  assign CLBLM_R_X5Y99_SLICE_X6Y99_D3 = 1'b1;
  assign CLBLM_R_X5Y99_SLICE_X6Y99_D4 = 1'b1;
  assign CLBLM_R_X5Y99_SLICE_X6Y99_D5 = 1'b1;
  assign CLBLM_R_X5Y99_SLICE_X6Y99_D6 = 1'b1;
  assign CLBLM_R_X5Y99_SLICE_X6Y99_SR = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y98_SLICE_X9Y98_B2 = CLBLM_L_X8Y98_SLICE_X10Y98_CO6;
  assign CLBLM_R_X7Y98_SLICE_X9Y98_B5 = CLBLM_R_X5Y95_SLICE_X6Y95_AQ;
  assign CLBLL_L_X4Y97_SLICE_X5Y97_B1 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO5;
  assign CLBLL_L_X4Y97_SLICE_X5Y97_B2 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLL_L_X4Y97_SLICE_X5Y97_B3 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLL_L_X4Y97_SLICE_X5Y97_B4 = CLBLM_R_X5Y95_SLICE_X6Y95_AQ;
  assign CLBLL_L_X4Y97_SLICE_X5Y97_C1 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLL_L_X4Y97_SLICE_X5Y97_C2 = CLBLM_R_X5Y97_SLICE_X7Y97_AO5;
  assign CLBLL_L_X4Y97_SLICE_X5Y97_C3 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLL_L_X4Y96_SLICE_X4Y96_A1 = CLBLM_R_X3Y98_SLICE_X3Y98_AO6;
  assign CLBLL_L_X4Y96_SLICE_X4Y96_A2 = CLBLL_L_X4Y98_SLICE_X4Y98_AO6;
  assign CLBLL_L_X4Y96_SLICE_X4Y96_A3 = CLBLL_L_X4Y97_SLICE_X4Y97_CO6;
  assign CLBLL_L_X4Y96_SLICE_X4Y96_A4 = CLBLL_L_X4Y96_SLICE_X4Y96_BO6;
  assign CLBLL_L_X4Y96_SLICE_X4Y96_A5 = CLBLL_L_X4Y97_SLICE_X4Y97_AO6;
  assign CLBLL_L_X4Y96_SLICE_X4Y96_A6 = CLBLM_R_X3Y96_SLICE_X2Y96_DO6;
  assign CLBLL_L_X4Y96_SLICE_X4Y96_B1 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO4;
  assign CLBLL_L_X4Y96_SLICE_X4Y96_B2 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLL_L_X4Y96_SLICE_X4Y96_B3 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLL_L_X4Y96_SLICE_X4Y96_B4 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLL_L_X4Y96_SLICE_X4Y96_B5 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLL_L_X4Y96_SLICE_X4Y96_B6 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLL_L_X4Y96_SLICE_X4Y96_C1 = CLBLL_L_X4Y97_SLICE_X4Y97_AO6;
  assign CLBLL_L_X4Y96_SLICE_X4Y96_C2 = CLBLL_L_X4Y96_SLICE_X5Y96_CO6;
  assign CLBLL_L_X4Y96_SLICE_X4Y96_C3 = CLBLM_R_X3Y96_SLICE_X2Y96_BO6;
  assign CLBLL_L_X4Y96_SLICE_X4Y96_C4 = CLBLL_L_X4Y98_SLICE_X4Y98_AO6;
  assign CLBLL_L_X4Y96_SLICE_X4Y96_C5 = CLBLL_L_X4Y97_SLICE_X4Y97_CO6;
  assign CLBLL_L_X4Y96_SLICE_X4Y96_C6 = CLBLM_R_X3Y98_SLICE_X3Y98_AO6;
  assign CLBLL_L_X4Y96_SLICE_X4Y96_D1 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO14;
  assign CLBLL_L_X4Y96_SLICE_X4Y96_D2 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO10;
  assign CLBLL_L_X4Y96_SLICE_X4Y96_D3 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO15;
  assign CLBLL_L_X4Y96_SLICE_X4Y96_D4 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO13;
  assign CLBLL_L_X4Y96_SLICE_X4Y96_D5 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO12;
  assign CLBLL_L_X4Y96_SLICE_X4Y96_D6 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO11;
  assign CLBLM_R_X3Y90_SLICE_X3Y90_A1 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X3Y90_A2 = 1'b1;
  assign CLBLL_L_X4Y96_SLICE_X5Y96_A1 = CLBLL_L_X4Y98_SLICE_X4Y98_AO6;
  assign CLBLL_L_X4Y96_SLICE_X5Y96_A2 = CLBLM_R_X3Y96_SLICE_X2Y96_AO6;
  assign CLBLL_L_X4Y96_SLICE_X5Y96_A3 = CLBLL_L_X4Y97_SLICE_X4Y97_AO6;
  assign CLBLM_R_X3Y90_SLICE_X3Y90_A6 = 1'b1;
  assign CLBLL_L_X4Y96_SLICE_X5Y96_A4 = CLBLL_L_X4Y96_SLICE_X5Y96_BO6;
  assign CLBLL_L_X4Y96_SLICE_X5Y96_A5 = CLBLL_L_X4Y97_SLICE_X4Y97_CO6;
  assign CLBLM_R_X3Y90_SLICE_X3Y90_AX = CLBLL_L_X4Y92_SLICE_X4Y92_AO5;
  assign CLBLL_L_X4Y96_SLICE_X5Y96_A6 = CLBLM_R_X3Y98_SLICE_X3Y98_AO6;
  assign CLBLM_R_X3Y90_SLICE_X3Y90_B1 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X3Y90_B2 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X3Y90_B3 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X3Y90_B4 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X3Y90_B5 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X3Y90_B6 = 1'b1;
  assign CLBLL_L_X4Y96_SLICE_X5Y96_B1 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLL_L_X4Y96_SLICE_X5Y96_B2 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X3Y90_SLICE_X3Y90_C1 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X3Y90_C2 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X3Y90_C3 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X3Y90_C4 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X3Y90_C5 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X3Y90_C6 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X3Y90_CE = CLBLL_L_X2Y92_SLICE_X1Y92_AO6;
  assign CLBLL_L_X4Y96_SLICE_X5Y96_C1 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLL_L_X4Y96_SLICE_X5Y96_C4 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLL_L_X4Y96_SLICE_X5Y96_C5 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO6;
  assign CLBLL_L_X4Y96_SLICE_X5Y96_C6 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLM_R_X7Y93_SLICE_X9Y93_A1 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X3Y90_D1 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X3Y90_D2 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X3Y90_D3 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X3Y90_D4 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X3Y90_D5 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X3Y90_D6 = 1'b1;
  assign CLBLL_L_X4Y96_SLICE_X5Y96_D5 = 1'b1;
  assign CLBLL_L_X4Y96_SLICE_X5Y96_D6 = 1'b1;
  assign CLBLL_L_X4Y96_SLICE_X5Y96_D1 = 1'b1;
  assign CLBLL_L_X4Y96_SLICE_X5Y96_D2 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X2Y90_A1 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X2Y90_A2 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X2Y90_A3 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X2Y90_A4 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X2Y90_A5 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X2Y90_A6 = 1'b1;
  assign CLBLM_R_X7Y93_SLICE_X9Y93_A4 = 1'b1;
  assign CLBLM_R_X7Y93_SLICE_X9Y93_A5 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X2Y90_AX = CLBLL_L_X4Y92_SLICE_X4Y92_AO6;
  assign CLBLM_R_X7Y93_SLICE_X9Y93_A6 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X2Y90_B1 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X2Y90_B2 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X2Y90_B3 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X2Y90_B4 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X2Y90_B5 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X2Y90_B6 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X2Y90_C1 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X2Y90_C2 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X2Y90_C3 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X2Y90_C4 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X2Y90_C5 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X2Y90_C6 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X2Y90_CE = CLBLL_L_X2Y93_SLICE_X1Y93_DO6;
  assign CLBLM_R_X7Y98_SLICE_X8Y98_B3 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X7Y98_SLICE_X8Y98_B4 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X7Y98_SLICE_X8Y98_B5 = CLBLL_L_X4Y97_SLICE_X4Y97_BQ;
  assign CLBLM_R_X7Y93_SLICE_X9Y93_B1 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X2Y90_D1 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X2Y90_D2 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X2Y90_D3 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X2Y90_D4 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X2Y90_D5 = 1'b1;
  assign CLBLM_R_X3Y90_SLICE_X2Y90_D6 = 1'b1;
  assign CLBLM_R_X7Y93_SLICE_X9Y93_B2 = 1'b1;
  assign CLBLM_R_X7Y93_SLICE_X9Y93_B3 = 1'b1;
  assign CLBLM_R_X7Y98_SLICE_X8Y98_B6 = CLBLM_R_X5Y95_SLICE_X6Y95_AQ;
  assign CLBLM_R_X7Y93_SLICE_X9Y93_B4 = 1'b1;
  assign CLBLM_R_X7Y93_SLICE_X9Y93_B5 = 1'b1;
  assign CLBLM_R_X7Y93_SLICE_X9Y93_B6 = 1'b1;
  assign CLBLM_R_X7Y93_SLICE_X9Y93_C1 = 1'b1;
  assign CLBLM_R_X7Y93_SLICE_X9Y93_C2 = 1'b1;
  assign CLBLM_R_X7Y93_SLICE_X9Y93_C3 = 1'b1;
  assign CLBLM_R_X7Y93_SLICE_X9Y93_C4 = 1'b1;
  assign CLBLM_R_X7Y93_SLICE_X9Y93_C5 = 1'b1;
  assign CLBLM_R_X7Y93_SLICE_X9Y93_C6 = 1'b1;
  assign CLBLL_L_X2Y95_SLICE_X1Y95_DX = 1'b0;
  assign CLBLM_R_X7Y93_SLICE_X9Y93_D1 = 1'b1;
  assign CLBLM_R_X7Y93_SLICE_X9Y93_D2 = 1'b1;
  assign CLBLM_R_X7Y93_SLICE_X9Y93_D3 = 1'b1;
  assign CLBLM_R_X7Y93_SLICE_X9Y93_D4 = 1'b1;
  assign CLBLM_R_X7Y93_SLICE_X9Y93_D5 = 1'b1;
  assign CLBLM_R_X7Y93_SLICE_X9Y93_D6 = 1'b1;
  assign CLBLL_L_X4Y97_SLICE_X4Y97_A1 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLL_L_X4Y97_SLICE_X4Y97_A2 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLL_L_X4Y97_SLICE_X4Y97_A3 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLL_L_X4Y97_SLICE_X4Y97_A4 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLL_L_X4Y97_SLICE_X4Y97_A5 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLL_L_X4Y97_SLICE_X4Y97_A6 = 1'b1;
  assign CLBLL_L_X4Y97_SLICE_X4Y97_B1 = CLBLL_L_X2Y97_SLICE_X1Y97_DO6;
  assign CLBLL_L_X4Y97_SLICE_X4Y97_B2 = CLBLL_L_X4Y97_SLICE_X4Y97_BQ;
  assign CLBLL_L_X4Y97_SLICE_X4Y97_B3 = 1'b1;
  assign CLBLL_L_X4Y97_SLICE_X4Y97_B4 = CLBLL_L_X2Y97_SLICE_X0Y97_DO6;
  assign CLBLL_L_X4Y97_SLICE_X4Y97_B5 = 1'b1;
  assign CLBLL_L_X4Y97_SLICE_X4Y97_B6 = CLBLL_L_X4Y97_SLICE_X4Y97_AO5;
  assign CLBLL_L_X4Y97_SLICE_X4Y97_C1 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLL_L_X4Y97_SLICE_X4Y97_C2 = CLBLL_L_X4Y97_SLICE_X5Y97_AO6;
  assign CLBLL_L_X4Y97_SLICE_X4Y97_C3 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLL_L_X4Y97_SLICE_X4Y97_C4 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO6;
  assign CLBLL_L_X4Y97_SLICE_X4Y97_C5 = CLBLL_L_X4Y97_SLICE_X4Y97_DO6;
  assign CLBLL_L_X4Y97_SLICE_X4Y97_C6 = CLBLM_R_X3Y96_SLICE_X3Y96_AO5;
  assign CLBLM_R_X7Y93_SLICE_X8Y93_A1 = CLBLM_R_X7Y93_SLICE_X8Y93_DO6;
  assign CLBLL_L_X4Y97_SLICE_X4Y97_D1 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO11;
  assign CLBLL_L_X4Y97_SLICE_X4Y97_D2 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO15;
  assign CLBLL_L_X4Y97_SLICE_X4Y97_D3 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO13;
  assign CLBLL_L_X4Y97_SLICE_X4Y97_D4 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO6;
  assign CLBLL_L_X4Y97_SLICE_X4Y97_D5 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO12;
  assign CLBLL_L_X4Y97_SLICE_X4Y97_D6 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO14;
  assign CLBLM_R_X7Y93_SLICE_X8Y93_A2 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X7Y93_SLICE_X8Y93_A3 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLL_L_X4Y97_SLICE_X4Y97_SR = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y93_SLICE_X8Y93_A4 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X7Y93_SLICE_X8Y93_A5 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLM_R_X7Y93_SLICE_X8Y93_A6 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLL_L_X4Y97_SLICE_X5Y97_A1 = CLBLM_R_X5Y95_SLICE_X6Y95_AQ;
  assign CLBLL_L_X4Y97_SLICE_X5Y97_A2 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLL_L_X4Y97_SLICE_X5Y97_A3 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLL_L_X4Y97_SLICE_X5Y97_A4 = CLBLL_L_X4Y97_SLICE_X4Y97_BQ;
  assign CLBLM_R_X3Y91_SLICE_X3Y91_A2 = CLBLM_R_X3Y92_SLICE_X3Y92_BQ;
  assign CLBLM_R_X3Y91_SLICE_X3Y91_A3 = CLBLL_L_X4Y91_SLICE_X5Y91_F7AMUX_O;
  assign CLBLM_R_X3Y91_SLICE_X3Y91_A4 = CLBLL_L_X4Y91_SLICE_X5Y91_BQ;
  assign CLBLM_R_X3Y91_SLICE_X3Y91_A5 = CLBLM_R_X5Y93_SLICE_X6Y93_F7AMUX_O;
  assign CLBLM_R_X3Y91_SLICE_X3Y91_A6 = CLBLM_R_X3Y91_SLICE_X3Y91_DQ;
  assign CLBLL_L_X4Y97_SLICE_X5Y97_A5 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLL_L_X4Y97_SLICE_X5Y97_A6 = 1'b1;
  assign CLBLM_R_X3Y91_SLICE_X3Y91_AX = CLBLL_L_X2Y93_SLICE_X0Y93_F7AMUX_O;
  assign CLBLM_R_X3Y91_SLICE_X3Y91_A1 = CLBLM_R_X3Y91_SLICE_X2Y91_DQ;
  assign CLBLM_R_X3Y91_SLICE_X3Y91_B1 = CLBLL_L_X4Y91_SLICE_X5Y91_F7AMUX_O;
  assign CLBLM_R_X3Y91_SLICE_X3Y91_B2 = CLBLL_L_X4Y92_SLICE_X4Y92_DQ;
  assign CLBLM_R_X3Y91_SLICE_X3Y91_B3 = CLBLM_R_X3Y90_SLICE_X3Y90_AQ;
  assign CLBLM_R_X3Y91_SLICE_X3Y91_B4 = CLBLM_R_X5Y92_SLICE_X6Y92_BQ;
  assign CLBLM_R_X3Y91_SLICE_X3Y91_B5 = CLBLM_R_X5Y93_SLICE_X6Y93_F7AMUX_O;
  assign CLBLM_R_X3Y91_SLICE_X3Y91_B6 = CLBLL_L_X4Y91_SLICE_X4Y91_BQ;
  assign CLBLL_L_X4Y97_SLICE_X5Y97_B5 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLL_L_X4Y97_SLICE_X5Y97_B6 = CLBLL_L_X4Y97_SLICE_X5Y97_CO6;
  assign CLBLM_R_X3Y91_SLICE_X3Y91_BX = CLBLL_L_X4Y92_SLICE_X4Y92_AO6;
  assign CLBLM_R_X3Y91_SLICE_X3Y91_C1 = CLBLL_L_X4Y91_SLICE_X5Y91_BQ;
  assign CLBLM_R_X3Y91_SLICE_X3Y91_C2 = CLBLM_R_X3Y96_SLICE_X3Y96_AO6;
  assign CLBLM_R_X3Y91_SLICE_X3Y91_C3 = CLBLM_R_X3Y91_SLICE_X3Y91_DQ;
  assign CLBLM_R_X3Y91_SLICE_X3Y91_C4 = CLBLL_L_X4Y91_SLICE_X4Y91_AO6;
  assign CLBLM_R_X3Y91_SLICE_X3Y91_C5 = CLBLM_R_X3Y91_SLICE_X2Y91_DQ;
  assign CLBLM_R_X3Y91_SLICE_X3Y91_C6 = CLBLM_R_X3Y92_SLICE_X3Y92_BQ;
  assign CLBLM_R_X3Y91_SLICE_X3Y91_CE = CLBLM_R_X3Y93_SLICE_X3Y93_CO6;
  assign CLBLL_L_X4Y97_SLICE_X5Y97_C6 = CLBLL_L_X4Y97_SLICE_X4Y97_BQ;
  assign CLBLL_L_X4Y97_SLICE_X5Y97_C4 = CLBLM_R_X5Y97_SLICE_X6Y97_BO6;
  assign CLBLL_L_X4Y97_SLICE_X5Y97_C5 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO5;
  assign CLBLL_L_X4Y97_SLICE_X5Y97_D1 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLM_R_X3Y91_SLICE_X3Y91_CX = CLBLL_L_X4Y95_SLICE_X5Y95_DO6;
  assign CLBLL_L_X4Y97_SLICE_X5Y97_D2 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X3Y91_SLICE_X3Y91_D1 = CLBLM_R_X3Y90_SLICE_X3Y90_AQ;
  assign CLBLM_R_X3Y91_SLICE_X3Y91_D2 = CLBLL_L_X4Y91_SLICE_X4Y91_BQ;
  assign CLBLM_R_X3Y91_SLICE_X3Y91_D3 = CLBLL_L_X4Y92_SLICE_X4Y92_DQ;
  assign CLBLM_R_X3Y91_SLICE_X3Y91_D4 = CLBLM_R_X3Y96_SLICE_X3Y96_AO6;
  assign CLBLM_R_X3Y91_SLICE_X3Y91_D5 = CLBLM_R_X5Y92_SLICE_X6Y92_BQ;
  assign CLBLM_R_X3Y91_SLICE_X3Y91_D6 = CLBLL_L_X4Y91_SLICE_X4Y91_AO6;
  assign CLBLL_L_X4Y97_SLICE_X5Y97_D3 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLM_R_X3Y91_SLICE_X3Y91_DX = CLBLL_L_X4Y92_SLICE_X4Y92_AO5;
  assign CLBLL_L_X4Y97_SLICE_X5Y97_D4 = CLBLL_L_X4Y97_SLICE_X5Y97_AO5;
  assign CLBLL_L_X4Y97_SLICE_X5Y97_D5 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLL_L_X4Y97_SLICE_X5Y97_D6 = 1'b1;
  assign CLBLM_R_X7Y93_SLICE_X8Y93_B6 = CLBLM_R_X7Y93_SLICE_X8Y93_CO6;
  assign CLBLM_R_X3Y91_SLICE_X2Y91_A1 = CLBLL_L_X2Y91_SLICE_X0Y91_AQ;
  assign CLBLM_R_X3Y91_SLICE_X2Y91_A2 = CLBLM_R_X3Y91_SLICE_X2Y91_BQ;
  assign CLBLM_R_X3Y91_SLICE_X2Y91_A3 = CLBLM_R_X5Y93_SLICE_X6Y93_F7AMUX_O;
  assign CLBLM_R_X3Y91_SLICE_X2Y91_A4 = CLBLM_R_X3Y91_SLICE_X3Y91_BQ;
  assign CLBLM_R_X3Y91_SLICE_X2Y91_A5 = CLBLL_L_X4Y91_SLICE_X5Y91_F7AMUX_O;
  assign CLBLM_R_X3Y91_SLICE_X2Y91_A6 = CLBLM_R_X3Y90_SLICE_X2Y90_AQ;
  assign CLBLM_R_X3Y91_SLICE_X2Y91_AX = CLBLL_L_X2Y93_SLICE_X0Y93_F7AMUX_O;
  assign CLBLM_R_X7Y87_SLICE_X8Y87_C3 = 1'b1;
  assign CLBLM_R_X3Y91_SLICE_X2Y91_B1 = CLBLL_L_X4Y91_SLICE_X5Y91_F7AMUX_O;
  assign CLBLM_R_X3Y91_SLICE_X2Y91_B2 = CLBLM_R_X5Y93_SLICE_X6Y93_F7AMUX_O;
  assign CLBLM_R_X3Y91_SLICE_X2Y91_B3 = CLBLL_L_X2Y90_SLICE_X1Y90_AQ;
  assign CLBLM_R_X3Y91_SLICE_X2Y91_B4 = CLBLL_L_X2Y92_SLICE_X1Y92_BQ;
  assign CLBLM_R_X3Y91_SLICE_X2Y91_B5 = CLBLL_L_X2Y91_SLICE_X1Y91_BQ;
  assign CLBLM_R_X3Y91_SLICE_X2Y91_B6 = CLBLM_R_X5Y92_SLICE_X6Y92_AQ;
  assign CLBLM_R_X3Y91_SLICE_X2Y91_BX = CLBLL_L_X4Y92_SLICE_X4Y92_AO6;
  assign CLBLM_R_X3Y91_SLICE_X2Y91_C1 = CLBLL_L_X4Y91_SLICE_X4Y91_AO6;
  assign CLBLM_R_X3Y91_SLICE_X2Y91_C2 = CLBLM_R_X3Y96_SLICE_X3Y96_AO6;
  assign CLBLM_R_X3Y91_SLICE_X2Y91_C3 = CLBLL_L_X2Y91_SLICE_X0Y91_AQ;
  assign CLBLM_R_X3Y91_SLICE_X2Y91_C4 = CLBLM_R_X3Y90_SLICE_X2Y90_AQ;
  assign CLBLM_R_X3Y91_SLICE_X2Y91_C5 = CLBLM_R_X3Y91_SLICE_X2Y91_BQ;
  assign CLBLM_R_X3Y91_SLICE_X2Y91_C6 = CLBLM_R_X3Y91_SLICE_X3Y91_BQ;
  assign CLBLM_R_X3Y91_SLICE_X2Y91_CE = CLBLM_R_X3Y93_SLICE_X3Y93_BO6;
  assign CLBLM_R_X7Y93_SLICE_X8Y93_C2 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO15;
  assign CLBLM_R_X7Y93_SLICE_X8Y93_C3 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLM_R_X3Y91_SLICE_X2Y91_CX = CLBLL_L_X4Y95_SLICE_X5Y95_DO6;
  assign CLBLM_R_X7Y93_SLICE_X8Y93_C4 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO13;
  assign CLBLM_R_X3Y91_SLICE_X2Y91_D1 = CLBLL_L_X2Y91_SLICE_X1Y91_BQ;
  assign CLBLM_R_X3Y91_SLICE_X2Y91_D2 = CLBLM_R_X3Y96_SLICE_X3Y96_AO6;
  assign CLBLM_R_X3Y91_SLICE_X2Y91_D3 = CLBLL_L_X2Y90_SLICE_X1Y90_AQ;
  assign CLBLM_R_X3Y91_SLICE_X2Y91_D4 = CLBLM_R_X5Y92_SLICE_X6Y92_AQ;
  assign CLBLM_R_X3Y91_SLICE_X2Y91_D5 = CLBLL_L_X4Y91_SLICE_X4Y91_AO6;
  assign CLBLM_R_X3Y91_SLICE_X2Y91_D6 = CLBLL_L_X2Y92_SLICE_X1Y92_BQ;
  assign CLBLM_R_X7Y93_SLICE_X8Y93_C5 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO12;
  assign CLBLM_R_X7Y93_SLICE_X8Y93_C6 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO14;
  assign CLBLM_R_X3Y91_SLICE_X2Y91_DX = CLBLL_L_X4Y92_SLICE_X4Y92_AO5;
  assign CLBLM_R_X7Y93_SLICE_X8Y93_CE = CLBLM_R_X7Y94_SLICE_X8Y94_CO6;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y95_SLICE_X6Y95_A4 = CLBLM_R_X5Y95_SLICE_X6Y95_BO6;
  assign CLBLM_R_X7Y93_SLICE_X8Y93_D1 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO11;
  assign CLBLL_L_X4Y98_SLICE_X4Y98_A1 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLL_L_X4Y98_SLICE_X4Y98_A2 = CLBLM_R_X3Y96_SLICE_X3Y96_AO5;
  assign CLBLL_L_X4Y98_SLICE_X4Y98_A3 = CLBLL_L_X4Y97_SLICE_X5Y97_AO6;
  assign CLBLL_L_X4Y98_SLICE_X4Y98_A4 = CLBLL_L_X4Y98_SLICE_X4Y98_BO6;
  assign CLBLL_L_X4Y98_SLICE_X4Y98_A5 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLL_L_X4Y98_SLICE_X4Y98_A6 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO5;
  assign CLBLM_R_X7Y88_SLICE_X8Y88_A4 = 1'b1;
  assign CLBLM_R_X7Y88_SLICE_X8Y88_A5 = 1'b1;
  assign CLBLL_L_X4Y98_SLICE_X4Y98_B1 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO13;
  assign CLBLL_L_X4Y98_SLICE_X4Y98_B2 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO11;
  assign CLBLL_L_X4Y98_SLICE_X4Y98_B3 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO14;
  assign CLBLL_L_X4Y98_SLICE_X4Y98_B4 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO5;
  assign CLBLL_L_X4Y98_SLICE_X4Y98_B5 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO12;
  assign CLBLL_L_X4Y98_SLICE_X4Y98_B6 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO15;
  assign CLBLM_R_X7Y88_SLICE_X8Y88_A6 = 1'b1;
  assign CLBLL_L_X4Y98_SLICE_X4Y98_C1 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO12;
  assign CLBLL_L_X4Y98_SLICE_X4Y98_C2 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO13;
  assign CLBLL_L_X4Y98_SLICE_X4Y98_C3 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO15;
  assign CLBLL_L_X4Y98_SLICE_X4Y98_C4 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO14;
  assign CLBLL_L_X4Y98_SLICE_X4Y98_C5 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO11;
  assign CLBLL_L_X4Y98_SLICE_X4Y98_C6 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO1;
  assign CLBLM_R_X5Y95_SLICE_X6Y95_C6 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO11;
  assign CLBLM_R_X5Y90_SLICE_X7Y90_C3 = 1'b1;
  assign CLBLL_L_X4Y98_SLICE_X4Y98_D1 = CLBLL_L_X4Y97_SLICE_X5Y97_AO6;
  assign CLBLL_L_X4Y98_SLICE_X4Y98_D2 = CLBLM_R_X3Y96_SLICE_X3Y96_AO5;
  assign CLBLL_L_X4Y98_SLICE_X4Y98_D3 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLL_L_X4Y98_SLICE_X4Y98_D4 = CLBLL_L_X4Y98_SLICE_X4Y98_CO6;
  assign CLBLL_L_X4Y98_SLICE_X4Y98_D5 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLL_L_X4Y98_SLICE_X4Y98_D6 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO1;
  assign CLBLM_R_X5Y90_SLICE_X7Y90_CE = CLBLM_R_X5Y90_SLICE_X7Y90_AO6;
  assign CLBLM_R_X7Y88_SLICE_X8Y88_B6 = CLBLM_R_X7Y91_SLICE_X8Y91_AQ;
  assign CLBLL_L_X4Y98_SLICE_X5Y98_A1 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLL_L_X4Y98_SLICE_X5Y98_A2 = CLBLM_R_X5Y95_SLICE_X6Y95_AQ;
  assign CLBLL_L_X4Y98_SLICE_X5Y98_A3 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLL_L_X4Y98_SLICE_X5Y98_A4 = CLBLM_R_X7Y94_SLICE_X9Y94_BQ;
  assign CLBLL_L_X4Y98_SLICE_X5Y98_A5 = CLBLM_R_X5Y98_SLICE_X7Y98_BO6;
  assign CLBLL_L_X4Y98_SLICE_X5Y98_A6 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO2;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRL0 = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRL1 = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRARDADDRL2 = CLBLM_R_X5Y90_SLICE_X7Y90_AQ;
  assign CLBLM_R_X3Y92_SLICE_X3Y92_A3 = 1'b1;
  assign CLBLM_R_X3Y92_SLICE_X3Y92_A4 = 1'b1;
  assign CLBLM_R_X3Y92_SLICE_X3Y92_A5 = 1'b1;
  assign CLBLM_R_X3Y92_SLICE_X3Y92_A6 = 1'b1;
  assign CLBLL_L_X4Y98_SLICE_X5Y98_B1 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLL_L_X4Y98_SLICE_X5Y98_B2 = CLBLM_R_X7Y94_SLICE_X9Y94_AQ;
  assign CLBLL_L_X4Y98_SLICE_X5Y98_B3 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign CLBLL_L_X4Y98_SLICE_X5Y98_B4 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO1;
  assign CLBLM_R_X3Y92_SLICE_X3Y92_B1 = 1'b1;
  assign CLBLM_R_X3Y92_SLICE_X3Y92_B2 = 1'b1;
  assign CLBLM_R_X3Y92_SLICE_X3Y92_B3 = 1'b1;
  assign CLBLM_R_X3Y92_SLICE_X3Y92_B4 = 1'b1;
  assign CLBLM_R_X3Y92_SLICE_X3Y92_B5 = 1'b1;
  assign CLBLM_R_X3Y92_SLICE_X3Y92_B6 = 1'b1;
  assign CLBLL_L_X4Y98_SLICE_X5Y98_B6 = CLBLM_R_X7Y93_SLICE_X8Y93_BQ;
  assign CLBLM_R_X3Y92_SLICE_X3Y92_BX = CLBLL_L_X4Y92_SLICE_X4Y92_AO5;
  assign CLBLL_L_X4Y98_SLICE_X5Y98_C1 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO14;
  assign CLBLM_R_X3Y92_SLICE_X3Y92_C1 = 1'b1;
  assign CLBLM_R_X3Y92_SLICE_X3Y92_C2 = 1'b1;
  assign CLBLM_R_X3Y92_SLICE_X3Y92_C3 = 1'b1;
  assign CLBLM_R_X3Y92_SLICE_X3Y92_C4 = 1'b1;
  assign CLBLL_L_X4Y98_SLICE_X5Y98_C4 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO13;
  assign CLBLL_L_X4Y98_SLICE_X5Y98_C5 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO12;
  assign CLBLL_L_X4Y98_SLICE_X5Y98_C6 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO11;
  assign CLBLL_L_X4Y98_SLICE_X5Y98_D1 = CLBLL_L_X4Y97_SLICE_X5Y97_AO6;
  assign CLBLL_L_X4Y98_SLICE_X5Y98_D2 = CLBLM_R_X3Y96_SLICE_X3Y96_AO5;
  assign CLBLL_L_X4Y98_SLICE_X5Y98_D3 = CLBLM_R_X7Y94_SLICE_X8Y94_AQ;
  assign CLBLL_L_X4Y98_SLICE_X5Y98_D4 = CLBLL_L_X4Y98_SLICE_X5Y98_CO6;
  assign CLBLL_L_X4Y98_SLICE_X5Y98_D5 = BRAM_L_X6Y95_RAMB36_X0Y19_DOADO4;
  assign CLBLL_L_X4Y98_SLICE_X5Y98_D6 = CLBLM_R_X7Y93_SLICE_X8Y93_AQ;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRL4 = CLBLM_R_X7Y90_SLICE_X9Y90_CQ;
  assign CLBLM_R_X3Y92_SLICE_X3Y92_D1 = 1'b1;
  assign CLBLM_R_X3Y92_SLICE_X3Y92_D2 = 1'b1;
  assign CLBLM_R_X3Y92_SLICE_X3Y92_D3 = 1'b1;
  assign CLBLM_R_X3Y92_SLICE_X3Y92_D4 = 1'b1;
  assign CLBLM_R_X3Y92_SLICE_X3Y92_D5 = 1'b1;
  assign CLBLM_R_X3Y92_SLICE_X3Y92_D6 = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRL7 = CLBLM_R_X7Y91_SLICE_X8Y91_AQ;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRL9 = CLBLM_L_X8Y89_SLICE_X10Y89_A5Q;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRL10 = CLBLM_R_X7Y89_SLICE_X9Y89_AQ;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRL11 = CLBLM_R_X7Y89_SLICE_X9Y89_BQ;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRL14 = CLBLM_R_X7Y89_SLICE_X8Y89_B5Q;
  assign CLBLM_R_X3Y92_SLICE_X2Y92_A1 = CLBLM_R_X3Y93_SLICE_X2Y93_CQ;
  assign CLBLM_R_X3Y92_SLICE_X2Y92_A2 = CLBLM_R_X3Y92_SLICE_X2Y92_DQ;
  assign CLBLM_R_X3Y92_SLICE_X2Y92_A3 = CLBLM_R_X5Y93_SLICE_X6Y93_F7AMUX_O;
  assign CLBLM_R_X3Y92_SLICE_X2Y92_A4 = CLBLL_L_X4Y91_SLICE_X5Y91_F7AMUX_O;
  assign CLBLM_R_X3Y92_SLICE_X2Y92_A5 = CLBLL_L_X2Y92_SLICE_X0Y92_AQ;
  assign CLBLM_R_X3Y92_SLICE_X2Y92_A6 = CLBLM_R_X3Y92_SLICE_X3Y92_CQ;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRU3 = CLBLM_R_X7Y90_SLICE_X9Y90_BQ;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRU4 = CLBLM_R_X7Y90_SLICE_X9Y90_CQ;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRU5 = CLBLM_R_X7Y91_SLICE_X9Y91_AQ;
  assign CLBLM_R_X3Y92_SLICE_X2Y92_AX = CLBLL_L_X2Y93_SLICE_X0Y93_F7AMUX_O;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_ADDRBWRADDRU7 = CLBLM_R_X7Y91_SLICE_X8Y91_AQ;
  assign CLBLM_R_X3Y92_SLICE_X3Y92_AX = CLBLM_R_X3Y94_SLICE_X2Y94_DO5;
  assign CLBLM_R_X3Y92_SLICE_X2Y92_B1 = CLBLL_L_X2Y94_SLICE_X1Y94_DQ;
  assign CLBLM_R_X3Y92_SLICE_X2Y92_B2 = CLBLL_L_X2Y92_SLICE_X1Y92_CQ;
  assign CLBLM_R_X3Y92_SLICE_X2Y92_B3 = CLBLM_R_X3Y94_SLICE_X2Y94_CQ;
  assign CLBLM_R_X3Y92_SLICE_X2Y92_B4 = CLBLL_L_X2Y91_SLICE_X1Y91_CQ;
  assign CLBLM_R_X3Y92_SLICE_X2Y92_B6 = CLBLL_L_X4Y91_SLICE_X5Y91_F7AMUX_O;
  assign CLBLM_R_X3Y92_SLICE_X2Y92_B5 = CLBLM_R_X5Y93_SLICE_X6Y93_F7AMUX_O;
  assign CLBLM_R_X3Y92_SLICE_X2Y92_BX = CLBLM_R_X3Y94_SLICE_X2Y94_DO6;
  assign CLBLM_R_X3Y92_SLICE_X2Y92_C1 = CLBLL_L_X2Y92_SLICE_X0Y92_AQ;
  assign CLBLM_R_X3Y92_SLICE_X2Y92_C2 = CLBLM_R_X3Y96_SLICE_X3Y96_AO6;
  assign CLBLM_R_X3Y92_SLICE_X2Y92_C3 = CLBLM_R_X3Y92_SLICE_X2Y92_DQ;
  assign CLBLM_R_X3Y92_SLICE_X2Y92_C4 = CLBLM_R_X3Y92_SLICE_X3Y92_CQ;
  assign CLBLM_R_X3Y92_SLICE_X2Y92_C5 = CLBLM_R_X3Y93_SLICE_X2Y93_CQ;
  assign CLBLM_R_X3Y92_SLICE_X2Y92_C6 = CLBLL_L_X4Y91_SLICE_X4Y91_AO6;
  assign CLBLM_R_X3Y92_SLICE_X2Y92_CE = CLBLM_R_X3Y93_SLICE_X3Y93_CO6;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIADI0 = CLBLM_R_X5Y93_SLICE_X7Y93_BQ;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIADI2 = CLBLM_R_X5Y91_SLICE_X6Y91_AQ;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIADI4 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIADI6 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIADI8 = 1'b0;
  assign CLBLM_R_X3Y92_SLICE_X2Y92_CX = CLBLL_L_X4Y95_SLICE_X5Y95_DO6;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIADI12 = 1'b0;
  assign CLBLM_R_X3Y92_SLICE_X2Y92_D1 = CLBLL_L_X4Y91_SLICE_X4Y91_AO6;
  assign CLBLM_R_X3Y92_SLICE_X2Y92_D2 = CLBLM_R_X3Y96_SLICE_X3Y96_AO6;
  assign CLBLM_R_X3Y92_SLICE_X2Y92_D3 = CLBLL_L_X2Y92_SLICE_X1Y92_CQ;
  assign CLBLM_R_X3Y92_SLICE_X2Y92_D4 = CLBLM_R_X3Y94_SLICE_X2Y94_CQ;
  assign CLBLM_R_X3Y92_SLICE_X2Y92_D5 = CLBLL_L_X2Y94_SLICE_X1Y94_DQ;
  assign CLBLM_R_X3Y92_SLICE_X2Y92_D6 = CLBLL_L_X2Y91_SLICE_X1Y91_CQ;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIADI26 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIADI28 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIADI30 = 1'b0;
  assign CLBLM_R_X3Y92_SLICE_X2Y92_DX = CLBLL_L_X4Y94_SLICE_X4Y94_CO5;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIADI3 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIADI5 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIADI7 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIADI9 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIADI29 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIADI13 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIADI15 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIADI17 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIADI19 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIADI23 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIADI25 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIADI27 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIADI31 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI0 = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI2 = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI4 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI6 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI8 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI10 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI12 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI14 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI16 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI18 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI20 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI22 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI24 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI26 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI28 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI30 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI1 = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI3 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI5 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI7 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI9 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI11 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI13 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI15 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI17 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI19 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI21 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI23 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI25 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI27 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI29 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIBDI31 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIPADIP0 = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIPADIP2 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIPADIP1 = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIPADIP3 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIPBDIP0 = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIPBDIP2 = 1'b0;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIPBDIP1 = 1'b1;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_DIPBDIP3 = 1'b0;
  assign CLBLM_R_X3Y92_SLICE_X3Y92_C6 = 1'b1;
  assign CLBLM_R_X3Y92_SLICE_X3Y92_CE = CLBLL_L_X2Y93_SLICE_X1Y93_DO6;
  assign CLBLM_R_X3Y92_SLICE_X3Y92_CX = CLBLL_L_X4Y94_SLICE_X4Y94_CO5;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X7Y93_SLICE_X8Y93_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLL_L_X4Y92_SLICE_X5Y92_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X5Y96_SLICE_X6Y96_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLL_L_X2Y91_SLICE_X1Y91_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X3Y99_SLICE_X2Y99_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X5Y90_SLICE_X7Y90_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_CLKARDCLKL = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign BRAM_L_X6Y95_RAMB36_X0Y19_CLKARDCLKU = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X3Y93_SLICE_X3Y93_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X5Y90_SLICE_X6Y90_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X3Y93_SLICE_X2Y93_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLL_L_X4Y93_SLICE_X4Y93_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X7Y94_SLICE_X9Y94_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLL_L_X2Y92_SLICE_X0Y92_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X7Y94_SLICE_X8Y94_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLL_L_X4Y93_SLICE_X5Y93_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLL_L_X2Y92_SLICE_X1Y92_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X5Y97_SLICE_X6Y97_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLL_L_X2Y99_SLICE_X0Y99_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLL_L_X2Y99_SLICE_X1Y99_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X3Y94_SLICE_X3Y94_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X7Y88_SLICE_X8Y88_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X5Y91_SLICE_X6Y91_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X3Y94_SLICE_X2Y94_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLL_L_X4Y94_SLICE_X4Y94_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLL_L_X2Y93_SLICE_X0Y93_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLL_L_X4Y94_SLICE_X5Y94_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLL_L_X2Y93_SLICE_X1Y93_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X5Y98_SLICE_X6Y98_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X5Y92_SLICE_X6Y92_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLL_L_X4Y95_SLICE_X4Y95_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X7Y96_SLICE_X9Y96_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X5Y99_SLICE_X7Y99_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X7Y96_SLICE_X8Y96_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLL_L_X2Y94_SLICE_X1Y94_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X5Y99_SLICE_X6Y99_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X5Y93_SLICE_X7Y93_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X5Y93_SLICE_X6Y93_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X3Y96_SLICE_X2Y96_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X7Y97_SLICE_X9Y97_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_L_X8Y97_SLICE_X11Y97_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X3Y90_SLICE_X3Y90_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X7Y97_SLICE_X8Y97_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_L_X8Y97_SLICE_X10Y97_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X3Y90_SLICE_X2Y90_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X5Y94_SLICE_X6Y94_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLL_L_X4Y90_SLICE_X5Y90_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X3Y97_SLICE_X2Y97_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLL_L_X4Y97_SLICE_X4Y97_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X7Y98_SLICE_X9Y98_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X3Y91_SLICE_X3Y91_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X3Y91_SLICE_X2Y91_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLL_L_X4Y91_SLICE_X4Y91_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLL_L_X4Y91_SLICE_X5Y91_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X5Y95_SLICE_X6Y95_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLL_L_X2Y90_SLICE_X1Y90_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X7Y99_SLICE_X9Y99_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X3Y92_SLICE_X3Y92_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X7Y99_SLICE_X8Y99_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_CLKARDCLKL = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_CLKARDCLKU = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_CLKBWRCLKL = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign BRAM_L_X6Y90_RAMB36_X0Y18_CLKBWRCLKU = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X3Y92_SLICE_X2Y92_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLL_L_X4Y92_SLICE_X4Y92_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLL_L_X2Y91_SLICE_X0Y91_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X5Y96_SLICE_X7Y96_CLK = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
endmodule
