// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 12 2017 08:25:46

// File Generated:     Jan 24 2019 12:17:51

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "atahost" view "INTERFACE"

module atahost (
    wb_dat_o,
    dd_pad_i,
    da_pad_o,
    wb_sel_i,
    wb_dat_i,
    wb_adr_i,
    dd_pad_o,
    wb_we_i,
    wb_stb_i,
    wb_rty_o,
    wb_rst_i,
    wb_inta_o,
    wb_err_o,
    wb_cyc_i,
    wb_clk_i,
    wb_ack_o,
    resetn_pad_o,
    iordy_pad_i,
    intrq_pad_i,
    dmarq_pad_i,
    dmackn_pad_o,
    diown_pad_o,
    diorn_pad_o,
    dd_padoe_o,
    cs1n_pad_o,
    cs0n_pad_o,
    arst_i,
    DMA_req,
    DMA_Ack);

    output [31:0] wb_dat_o;
    input [15:0] dd_pad_i;
    output [2:0] da_pad_o;
    input [3:0] wb_sel_i;
    input [31:0] wb_dat_i;
    input [6:2] wb_adr_i;
    output [15:0] dd_pad_o;
    input wb_we_i;
    input wb_stb_i;
    output wb_rty_o;
    input wb_rst_i;
    output wb_inta_o;
    output wb_err_o;
    input wb_cyc_i;
    input wb_clk_i;
    output wb_ack_o;
    output resetn_pad_o;
    input iordy_pad_i;
    input intrq_pad_i;
    input dmarq_pad_i;
    output dmackn_pad_o;
    output diown_pad_o;
    output diorn_pad_o;
    output dd_padoe_o;
    output cs1n_pad_o;
    output cs0n_pad_o;
    input arst_i;
    output DMA_req;
    input DMA_Ack;

    wire N__55912;
    wire N__55911;
    wire N__55910;
    wire N__55901;
    wire N__55900;
    wire N__55899;
    wire N__55892;
    wire N__55891;
    wire N__55890;
    wire N__55883;
    wire N__55882;
    wire N__55881;
    wire N__55874;
    wire N__55873;
    wire N__55872;
    wire N__55865;
    wire N__55864;
    wire N__55863;
    wire N__55856;
    wire N__55855;
    wire N__55854;
    wire N__55847;
    wire N__55846;
    wire N__55845;
    wire N__55838;
    wire N__55837;
    wire N__55836;
    wire N__55829;
    wire N__55828;
    wire N__55827;
    wire N__55820;
    wire N__55819;
    wire N__55818;
    wire N__55811;
    wire N__55810;
    wire N__55809;
    wire N__55802;
    wire N__55801;
    wire N__55800;
    wire N__55793;
    wire N__55792;
    wire N__55791;
    wire N__55784;
    wire N__55783;
    wire N__55782;
    wire N__55775;
    wire N__55774;
    wire N__55773;
    wire N__55766;
    wire N__55765;
    wire N__55764;
    wire N__55757;
    wire N__55756;
    wire N__55755;
    wire N__55748;
    wire N__55747;
    wire N__55746;
    wire N__55739;
    wire N__55738;
    wire N__55737;
    wire N__55730;
    wire N__55729;
    wire N__55728;
    wire N__55721;
    wire N__55720;
    wire N__55719;
    wire N__55712;
    wire N__55711;
    wire N__55710;
    wire N__55703;
    wire N__55702;
    wire N__55701;
    wire N__55694;
    wire N__55693;
    wire N__55692;
    wire N__55685;
    wire N__55684;
    wire N__55683;
    wire N__55676;
    wire N__55675;
    wire N__55674;
    wire N__55667;
    wire N__55666;
    wire N__55665;
    wire N__55658;
    wire N__55657;
    wire N__55656;
    wire N__55649;
    wire N__55648;
    wire N__55647;
    wire N__55640;
    wire N__55639;
    wire N__55638;
    wire N__55631;
    wire N__55630;
    wire N__55629;
    wire N__55622;
    wire N__55621;
    wire N__55620;
    wire N__55613;
    wire N__55612;
    wire N__55611;
    wire N__55604;
    wire N__55603;
    wire N__55602;
    wire N__55595;
    wire N__55594;
    wire N__55593;
    wire N__55586;
    wire N__55585;
    wire N__55584;
    wire N__55577;
    wire N__55576;
    wire N__55575;
    wire N__55568;
    wire N__55567;
    wire N__55566;
    wire N__55559;
    wire N__55558;
    wire N__55557;
    wire N__55550;
    wire N__55549;
    wire N__55548;
    wire N__55541;
    wire N__55540;
    wire N__55539;
    wire N__55532;
    wire N__55531;
    wire N__55530;
    wire N__55523;
    wire N__55522;
    wire N__55521;
    wire N__55514;
    wire N__55513;
    wire N__55512;
    wire N__55505;
    wire N__55504;
    wire N__55503;
    wire N__55496;
    wire N__55495;
    wire N__55494;
    wire N__55487;
    wire N__55486;
    wire N__55485;
    wire N__55478;
    wire N__55477;
    wire N__55476;
    wire N__55469;
    wire N__55468;
    wire N__55467;
    wire N__55460;
    wire N__55459;
    wire N__55458;
    wire N__55451;
    wire N__55450;
    wire N__55449;
    wire N__55442;
    wire N__55441;
    wire N__55440;
    wire N__55433;
    wire N__55432;
    wire N__55431;
    wire N__55424;
    wire N__55423;
    wire N__55422;
    wire N__55415;
    wire N__55414;
    wire N__55413;
    wire N__55406;
    wire N__55405;
    wire N__55404;
    wire N__55397;
    wire N__55396;
    wire N__55395;
    wire N__55388;
    wire N__55387;
    wire N__55386;
    wire N__55379;
    wire N__55378;
    wire N__55377;
    wire N__55370;
    wire N__55369;
    wire N__55368;
    wire N__55361;
    wire N__55360;
    wire N__55359;
    wire N__55352;
    wire N__55351;
    wire N__55350;
    wire N__55343;
    wire N__55342;
    wire N__55341;
    wire N__55334;
    wire N__55333;
    wire N__55332;
    wire N__55325;
    wire N__55324;
    wire N__55323;
    wire N__55316;
    wire N__55315;
    wire N__55314;
    wire N__55307;
    wire N__55306;
    wire N__55305;
    wire N__55298;
    wire N__55297;
    wire N__55296;
    wire N__55289;
    wire N__55288;
    wire N__55287;
    wire N__55280;
    wire N__55279;
    wire N__55278;
    wire N__55271;
    wire N__55270;
    wire N__55269;
    wire N__55262;
    wire N__55261;
    wire N__55260;
    wire N__55253;
    wire N__55252;
    wire N__55251;
    wire N__55244;
    wire N__55243;
    wire N__55242;
    wire N__55235;
    wire N__55234;
    wire N__55233;
    wire N__55226;
    wire N__55225;
    wire N__55224;
    wire N__55217;
    wire N__55216;
    wire N__55215;
    wire N__55208;
    wire N__55207;
    wire N__55206;
    wire N__55199;
    wire N__55198;
    wire N__55197;
    wire N__55190;
    wire N__55189;
    wire N__55188;
    wire N__55181;
    wire N__55180;
    wire N__55179;
    wire N__55172;
    wire N__55171;
    wire N__55170;
    wire N__55163;
    wire N__55162;
    wire N__55161;
    wire N__55154;
    wire N__55153;
    wire N__55152;
    wire N__55145;
    wire N__55144;
    wire N__55143;
    wire N__55136;
    wire N__55135;
    wire N__55134;
    wire N__55127;
    wire N__55126;
    wire N__55125;
    wire N__55118;
    wire N__55117;
    wire N__55116;
    wire N__55109;
    wire N__55108;
    wire N__55107;
    wire N__55100;
    wire N__55099;
    wire N__55098;
    wire N__55091;
    wire N__55090;
    wire N__55089;
    wire N__55082;
    wire N__55081;
    wire N__55080;
    wire N__55073;
    wire N__55072;
    wire N__55071;
    wire N__55064;
    wire N__55063;
    wire N__55062;
    wire N__55055;
    wire N__55054;
    wire N__55053;
    wire N__55046;
    wire N__55045;
    wire N__55044;
    wire N__55037;
    wire N__55036;
    wire N__55035;
    wire N__55028;
    wire N__55027;
    wire N__55026;
    wire N__55019;
    wire N__55018;
    wire N__55017;
    wire N__55010;
    wire N__55009;
    wire N__55008;
    wire N__55001;
    wire N__55000;
    wire N__54999;
    wire N__54992;
    wire N__54991;
    wire N__54990;
    wire N__54983;
    wire N__54982;
    wire N__54981;
    wire N__54974;
    wire N__54973;
    wire N__54972;
    wire N__54965;
    wire N__54964;
    wire N__54963;
    wire N__54956;
    wire N__54955;
    wire N__54954;
    wire N__54947;
    wire N__54946;
    wire N__54945;
    wire N__54938;
    wire N__54937;
    wire N__54936;
    wire N__54929;
    wire N__54928;
    wire N__54927;
    wire N__54920;
    wire N__54919;
    wire N__54918;
    wire N__54911;
    wire N__54910;
    wire N__54909;
    wire N__54902;
    wire N__54901;
    wire N__54900;
    wire N__54893;
    wire N__54892;
    wire N__54891;
    wire N__54884;
    wire N__54883;
    wire N__54882;
    wire N__54875;
    wire N__54874;
    wire N__54873;
    wire N__54866;
    wire N__54865;
    wire N__54864;
    wire N__54857;
    wire N__54856;
    wire N__54855;
    wire N__54848;
    wire N__54847;
    wire N__54846;
    wire N__54839;
    wire N__54838;
    wire N__54837;
    wire N__54830;
    wire N__54829;
    wire N__54828;
    wire N__54821;
    wire N__54820;
    wire N__54819;
    wire N__54812;
    wire N__54811;
    wire N__54810;
    wire N__54803;
    wire N__54802;
    wire N__54801;
    wire N__54794;
    wire N__54793;
    wire N__54792;
    wire N__54785;
    wire N__54784;
    wire N__54783;
    wire N__54776;
    wire N__54775;
    wire N__54774;
    wire N__54767;
    wire N__54766;
    wire N__54765;
    wire N__54758;
    wire N__54757;
    wire N__54756;
    wire N__54749;
    wire N__54748;
    wire N__54747;
    wire N__54730;
    wire N__54727;
    wire N__54724;
    wire N__54721;
    wire N__54718;
    wire N__54717;
    wire N__54716;
    wire N__54715;
    wire N__54714;
    wire N__54713;
    wire N__54712;
    wire N__54709;
    wire N__54708;
    wire N__54707;
    wire N__54706;
    wire N__54705;
    wire N__54704;
    wire N__54701;
    wire N__54698;
    wire N__54693;
    wire N__54690;
    wire N__54689;
    wire N__54688;
    wire N__54687;
    wire N__54686;
    wire N__54679;
    wire N__54676;
    wire N__54675;
    wire N__54674;
    wire N__54673;
    wire N__54670;
    wire N__54667;
    wire N__54664;
    wire N__54661;
    wire N__54658;
    wire N__54655;
    wire N__54652;
    wire N__54643;
    wire N__54638;
    wire N__54635;
    wire N__54634;
    wire N__54631;
    wire N__54630;
    wire N__54629;
    wire N__54626;
    wire N__54621;
    wire N__54618;
    wire N__54613;
    wire N__54606;
    wire N__54601;
    wire N__54598;
    wire N__54595;
    wire N__54590;
    wire N__54589;
    wire N__54588;
    wire N__54587;
    wire N__54584;
    wire N__54575;
    wire N__54570;
    wire N__54565;
    wire N__54562;
    wire N__54559;
    wire N__54556;
    wire N__54541;
    wire N__54538;
    wire N__54535;
    wire N__54532;
    wire N__54529;
    wire N__54526;
    wire N__54523;
    wire N__54522;
    wire N__54519;
    wire N__54516;
    wire N__54513;
    wire N__54510;
    wire N__54507;
    wire N__54504;
    wire N__54501;
    wire N__54498;
    wire N__54493;
    wire N__54490;
    wire N__54487;
    wire N__54484;
    wire N__54481;
    wire N__54478;
    wire N__54475;
    wire N__54472;
    wire N__54469;
    wire N__54468;
    wire N__54467;
    wire N__54466;
    wire N__54465;
    wire N__54462;
    wire N__54461;
    wire N__54460;
    wire N__54459;
    wire N__54456;
    wire N__54455;
    wire N__54452;
    wire N__54449;
    wire N__54446;
    wire N__54443;
    wire N__54440;
    wire N__54437;
    wire N__54434;
    wire N__54431;
    wire N__54428;
    wire N__54423;
    wire N__54420;
    wire N__54411;
    wire N__54408;
    wire N__54405;
    wire N__54402;
    wire N__54399;
    wire N__54396;
    wire N__54393;
    wire N__54390;
    wire N__54387;
    wire N__54384;
    wire N__54381;
    wire N__54376;
    wire N__54369;
    wire N__54366;
    wire N__54363;
    wire N__54358;
    wire N__54357;
    wire N__54354;
    wire N__54351;
    wire N__54348;
    wire N__54345;
    wire N__54342;
    wire N__54339;
    wire N__54334;
    wire N__54333;
    wire N__54332;
    wire N__54331;
    wire N__54330;
    wire N__54329;
    wire N__54328;
    wire N__54327;
    wire N__54326;
    wire N__54325;
    wire N__54324;
    wire N__54323;
    wire N__54322;
    wire N__54321;
    wire N__54320;
    wire N__54319;
    wire N__54318;
    wire N__54317;
    wire N__54316;
    wire N__54315;
    wire N__54314;
    wire N__54313;
    wire N__54312;
    wire N__54311;
    wire N__54310;
    wire N__54309;
    wire N__54308;
    wire N__54307;
    wire N__54306;
    wire N__54305;
    wire N__54304;
    wire N__54303;
    wire N__54302;
    wire N__54301;
    wire N__54300;
    wire N__54299;
    wire N__54298;
    wire N__54297;
    wire N__54296;
    wire N__54295;
    wire N__54294;
    wire N__54293;
    wire N__54292;
    wire N__54291;
    wire N__54290;
    wire N__54289;
    wire N__54288;
    wire N__54287;
    wire N__54286;
    wire N__54285;
    wire N__54284;
    wire N__54283;
    wire N__54282;
    wire N__54281;
    wire N__54280;
    wire N__54279;
    wire N__54278;
    wire N__54277;
    wire N__54276;
    wire N__54275;
    wire N__54274;
    wire N__54273;
    wire N__54272;
    wire N__54271;
    wire N__54270;
    wire N__54269;
    wire N__54268;
    wire N__54267;
    wire N__54266;
    wire N__54265;
    wire N__54264;
    wire N__54263;
    wire N__54262;
    wire N__54261;
    wire N__54260;
    wire N__54259;
    wire N__54258;
    wire N__54257;
    wire N__54256;
    wire N__54255;
    wire N__54254;
    wire N__54253;
    wire N__54252;
    wire N__54251;
    wire N__54250;
    wire N__54249;
    wire N__54248;
    wire N__54247;
    wire N__54246;
    wire N__54245;
    wire N__54244;
    wire N__54243;
    wire N__54242;
    wire N__54241;
    wire N__54240;
    wire N__54239;
    wire N__54238;
    wire N__54237;
    wire N__54236;
    wire N__54235;
    wire N__54234;
    wire N__54233;
    wire N__54232;
    wire N__54231;
    wire N__54230;
    wire N__54229;
    wire N__54228;
    wire N__54227;
    wire N__54226;
    wire N__54225;
    wire N__54224;
    wire N__54223;
    wire N__54222;
    wire N__54221;
    wire N__54220;
    wire N__54219;
    wire N__54218;
    wire N__54217;
    wire N__54216;
    wire N__54215;
    wire N__54214;
    wire N__54213;
    wire N__54212;
    wire N__54211;
    wire N__54210;
    wire N__54209;
    wire N__54208;
    wire N__54207;
    wire N__54206;
    wire N__54205;
    wire N__54204;
    wire N__54203;
    wire N__54202;
    wire N__54201;
    wire N__54200;
    wire N__54199;
    wire N__54198;
    wire N__54197;
    wire N__54196;
    wire N__54195;
    wire N__54194;
    wire N__54193;
    wire N__54192;
    wire N__54191;
    wire N__54190;
    wire N__54189;
    wire N__54188;
    wire N__54187;
    wire N__54186;
    wire N__54185;
    wire N__54184;
    wire N__54183;
    wire N__54182;
    wire N__54181;
    wire N__54180;
    wire N__54179;
    wire N__54178;
    wire N__54177;
    wire N__54176;
    wire N__54175;
    wire N__54174;
    wire N__54173;
    wire N__54172;
    wire N__54171;
    wire N__54170;
    wire N__54169;
    wire N__54168;
    wire N__54167;
    wire N__54166;
    wire N__54165;
    wire N__54164;
    wire N__54163;
    wire N__54162;
    wire N__54161;
    wire N__54160;
    wire N__54159;
    wire N__54158;
    wire N__54157;
    wire N__54156;
    wire N__54155;
    wire N__54154;
    wire N__54153;
    wire N__54152;
    wire N__54151;
    wire N__54150;
    wire N__54149;
    wire N__54148;
    wire N__54147;
    wire N__54146;
    wire N__54145;
    wire N__54144;
    wire N__54143;
    wire N__54142;
    wire N__54141;
    wire N__54140;
    wire N__54139;
    wire N__54138;
    wire N__54137;
    wire N__54136;
    wire N__54135;
    wire N__54134;
    wire N__54133;
    wire N__54132;
    wire N__54131;
    wire N__54130;
    wire N__54129;
    wire N__54128;
    wire N__54127;
    wire N__54126;
    wire N__54125;
    wire N__54124;
    wire N__54123;
    wire N__54122;
    wire N__54121;
    wire N__54120;
    wire N__54119;
    wire N__54118;
    wire N__54117;
    wire N__54116;
    wire N__54115;
    wire N__54114;
    wire N__54113;
    wire N__54112;
    wire N__54111;
    wire N__54110;
    wire N__53659;
    wire N__53656;
    wire N__53653;
    wire N__53652;
    wire N__53651;
    wire N__53648;
    wire N__53647;
    wire N__53646;
    wire N__53645;
    wire N__53644;
    wire N__53643;
    wire N__53642;
    wire N__53641;
    wire N__53638;
    wire N__53635;
    wire N__53634;
    wire N__53631;
    wire N__53628;
    wire N__53625;
    wire N__53622;
    wire N__53619;
    wire N__53616;
    wire N__53615;
    wire N__53614;
    wire N__53611;
    wire N__53610;
    wire N__53607;
    wire N__53606;
    wire N__53601;
    wire N__53598;
    wire N__53591;
    wire N__53588;
    wire N__53587;
    wire N__53582;
    wire N__53579;
    wire N__53576;
    wire N__53575;
    wire N__53572;
    wire N__53569;
    wire N__53566;
    wire N__53565;
    wire N__53562;
    wire N__53561;
    wire N__53560;
    wire N__53555;
    wire N__53550;
    wire N__53549;
    wire N__53546;
    wire N__53539;
    wire N__53536;
    wire N__53531;
    wire N__53530;
    wire N__53527;
    wire N__53524;
    wire N__53521;
    wire N__53518;
    wire N__53515;
    wire N__53514;
    wire N__53513;
    wire N__53510;
    wire N__53507;
    wire N__53504;
    wire N__53501;
    wire N__53496;
    wire N__53493;
    wire N__53490;
    wire N__53487;
    wire N__53484;
    wire N__53477;
    wire N__53474;
    wire N__53471;
    wire N__53464;
    wire N__53459;
    wire N__53454;
    wire N__53447;
    wire N__53444;
    wire N__53441;
    wire N__53438;
    wire N__53433;
    wire N__53430;
    wire N__53425;
    wire N__53422;
    wire N__53413;
    wire N__53412;
    wire N__53411;
    wire N__53410;
    wire N__53409;
    wire N__53408;
    wire N__53407;
    wire N__53406;
    wire N__53405;
    wire N__53404;
    wire N__53403;
    wire N__53402;
    wire N__53401;
    wire N__53400;
    wire N__53399;
    wire N__53398;
    wire N__53397;
    wire N__53396;
    wire N__53395;
    wire N__53394;
    wire N__53393;
    wire N__53392;
    wire N__53391;
    wire N__53390;
    wire N__53389;
    wire N__53388;
    wire N__53387;
    wire N__53386;
    wire N__53385;
    wire N__53384;
    wire N__53383;
    wire N__53382;
    wire N__53381;
    wire N__53380;
    wire N__53379;
    wire N__53378;
    wire N__53377;
    wire N__53376;
    wire N__53375;
    wire N__53374;
    wire N__53373;
    wire N__53372;
    wire N__53371;
    wire N__53370;
    wire N__53369;
    wire N__53368;
    wire N__53367;
    wire N__53366;
    wire N__53365;
    wire N__53364;
    wire N__53363;
    wire N__53362;
    wire N__53361;
    wire N__53360;
    wire N__53359;
    wire N__53358;
    wire N__53357;
    wire N__53356;
    wire N__53355;
    wire N__53354;
    wire N__53353;
    wire N__53352;
    wire N__53351;
    wire N__53350;
    wire N__53349;
    wire N__53348;
    wire N__53347;
    wire N__53346;
    wire N__53345;
    wire N__53344;
    wire N__53343;
    wire N__53342;
    wire N__53341;
    wire N__53340;
    wire N__53339;
    wire N__53338;
    wire N__53337;
    wire N__53336;
    wire N__53335;
    wire N__53334;
    wire N__53333;
    wire N__53332;
    wire N__53331;
    wire N__53330;
    wire N__53329;
    wire N__53328;
    wire N__53327;
    wire N__53326;
    wire N__53325;
    wire N__53324;
    wire N__53323;
    wire N__53322;
    wire N__53321;
    wire N__53320;
    wire N__53319;
    wire N__53318;
    wire N__53317;
    wire N__53316;
    wire N__53315;
    wire N__53314;
    wire N__53313;
    wire N__53312;
    wire N__53311;
    wire N__53310;
    wire N__53309;
    wire N__53308;
    wire N__53307;
    wire N__53306;
    wire N__53305;
    wire N__53086;
    wire N__53083;
    wire N__53080;
    wire N__53079;
    wire N__53078;
    wire N__53077;
    wire N__53074;
    wire N__53071;
    wire N__53070;
    wire N__53069;
    wire N__53068;
    wire N__53067;
    wire N__53066;
    wire N__53065;
    wire N__53062;
    wire N__53059;
    wire N__53058;
    wire N__53057;
    wire N__53056;
    wire N__53047;
    wire N__53044;
    wire N__53041;
    wire N__53038;
    wire N__53031;
    wire N__53028;
    wire N__53025;
    wire N__53024;
    wire N__53023;
    wire N__53020;
    wire N__53019;
    wire N__53016;
    wire N__53015;
    wire N__53012;
    wire N__53007;
    wire N__53006;
    wire N__53003;
    wire N__53000;
    wire N__52991;
    wire N__52988;
    wire N__52985;
    wire N__52982;
    wire N__52979;
    wire N__52976;
    wire N__52973;
    wire N__52964;
    wire N__52959;
    wire N__52956;
    wire N__52951;
    wire N__52948;
    wire N__52945;
    wire N__52942;
    wire N__52939;
    wire N__52934;
    wire N__52931;
    wire N__52928;
    wire N__52925;
    wire N__52922;
    wire N__52917;
    wire N__52912;
    wire N__52911;
    wire N__52910;
    wire N__52909;
    wire N__52908;
    wire N__52907;
    wire N__52904;
    wire N__52893;
    wire N__52888;
    wire N__52887;
    wire N__52886;
    wire N__52883;
    wire N__52880;
    wire N__52877;
    wire N__52874;
    wire N__52869;
    wire N__52864;
    wire N__52861;
    wire N__52860;
    wire N__52857;
    wire N__52854;
    wire N__52851;
    wire N__52848;
    wire N__52845;
    wire N__52842;
    wire N__52839;
    wire N__52836;
    wire N__52831;
    wire N__52828;
    wire N__52827;
    wire N__52824;
    wire N__52821;
    wire N__52818;
    wire N__52815;
    wire N__52812;
    wire N__52809;
    wire N__52804;
    wire N__52801;
    wire N__52798;
    wire N__52795;
    wire N__52792;
    wire N__52789;
    wire N__52788;
    wire N__52787;
    wire N__52784;
    wire N__52783;
    wire N__52782;
    wire N__52781;
    wire N__52780;
    wire N__52779;
    wire N__52778;
    wire N__52775;
    wire N__52774;
    wire N__52773;
    wire N__52772;
    wire N__52771;
    wire N__52770;
    wire N__52769;
    wire N__52768;
    wire N__52767;
    wire N__52764;
    wire N__52763;
    wire N__52762;
    wire N__52761;
    wire N__52758;
    wire N__52751;
    wire N__52742;
    wire N__52739;
    wire N__52736;
    wire N__52733;
    wire N__52732;
    wire N__52729;
    wire N__52726;
    wire N__52723;
    wire N__52720;
    wire N__52717;
    wire N__52714;
    wire N__52711;
    wire N__52710;
    wire N__52709;
    wire N__52708;
    wire N__52707;
    wire N__52704;
    wire N__52701;
    wire N__52700;
    wire N__52699;
    wire N__52698;
    wire N__52697;
    wire N__52696;
    wire N__52695;
    wire N__52694;
    wire N__52693;
    wire N__52692;
    wire N__52685;
    wire N__52680;
    wire N__52677;
    wire N__52670;
    wire N__52667;
    wire N__52664;
    wire N__52661;
    wire N__52656;
    wire N__52653;
    wire N__52652;
    wire N__52651;
    wire N__52648;
    wire N__52647;
    wire N__52646;
    wire N__52645;
    wire N__52644;
    wire N__52643;
    wire N__52642;
    wire N__52641;
    wire N__52640;
    wire N__52639;
    wire N__52638;
    wire N__52637;
    wire N__52636;
    wire N__52635;
    wire N__52632;
    wire N__52631;
    wire N__52630;
    wire N__52629;
    wire N__52628;
    wire N__52627;
    wire N__52624;
    wire N__52623;
    wire N__52618;
    wire N__52615;
    wire N__52612;
    wire N__52611;
    wire N__52610;
    wire N__52609;
    wire N__52608;
    wire N__52607;
    wire N__52606;
    wire N__52603;
    wire N__52602;
    wire N__52601;
    wire N__52598;
    wire N__52595;
    wire N__52592;
    wire N__52589;
    wire N__52588;
    wire N__52585;
    wire N__52582;
    wire N__52581;
    wire N__52580;
    wire N__52579;
    wire N__52578;
    wire N__52577;
    wire N__52576;
    wire N__52575;
    wire N__52574;
    wire N__52573;
    wire N__52560;
    wire N__52553;
    wire N__52550;
    wire N__52547;
    wire N__52544;
    wire N__52537;
    wire N__52526;
    wire N__52519;
    wire N__52518;
    wire N__52517;
    wire N__52516;
    wire N__52515;
    wire N__52514;
    wire N__52513;
    wire N__52512;
    wire N__52511;
    wire N__52510;
    wire N__52509;
    wire N__52508;
    wire N__52507;
    wire N__52506;
    wire N__52505;
    wire N__52504;
    wire N__52503;
    wire N__52502;
    wire N__52501;
    wire N__52498;
    wire N__52495;
    wire N__52494;
    wire N__52493;
    wire N__52490;
    wire N__52485;
    wire N__52482;
    wire N__52479;
    wire N__52476;
    wire N__52473;
    wire N__52472;
    wire N__52471;
    wire N__52470;
    wire N__52469;
    wire N__52468;
    wire N__52467;
    wire N__52464;
    wire N__52463;
    wire N__52462;
    wire N__52461;
    wire N__52460;
    wire N__52459;
    wire N__52456;
    wire N__52451;
    wire N__52450;
    wire N__52449;
    wire N__52446;
    wire N__52445;
    wire N__52444;
    wire N__52441;
    wire N__52440;
    wire N__52437;
    wire N__52436;
    wire N__52433;
    wire N__52430;
    wire N__52427;
    wire N__52426;
    wire N__52425;
    wire N__52424;
    wire N__52423;
    wire N__52422;
    wire N__52417;
    wire N__52414;
    wire N__52405;
    wire N__52396;
    wire N__52393;
    wire N__52390;
    wire N__52387;
    wire N__52384;
    wire N__52381;
    wire N__52378;
    wire N__52375;
    wire N__52372;
    wire N__52369;
    wire N__52354;
    wire N__52337;
    wire N__52322;
    wire N__52319;
    wire N__52312;
    wire N__52309;
    wire N__52308;
    wire N__52307;
    wire N__52306;
    wire N__52305;
    wire N__52302;
    wire N__52301;
    wire N__52298;
    wire N__52297;
    wire N__52292;
    wire N__52287;
    wire N__52282;
    wire N__52275;
    wire N__52264;
    wire N__52263;
    wire N__52262;
    wire N__52259;
    wire N__52256;
    wire N__52255;
    wire N__52254;
    wire N__52253;
    wire N__52252;
    wire N__52249;
    wire N__52246;
    wire N__52245;
    wire N__52244;
    wire N__52243;
    wire N__52242;
    wire N__52241;
    wire N__52236;
    wire N__52233;
    wire N__52230;
    wire N__52227;
    wire N__52218;
    wire N__52213;
    wire N__52206;
    wire N__52205;
    wire N__52204;
    wire N__52201;
    wire N__52200;
    wire N__52199;
    wire N__52198;
    wire N__52197;
    wire N__52196;
    wire N__52195;
    wire N__52194;
    wire N__52187;
    wire N__52186;
    wire N__52183;
    wire N__52182;
    wire N__52181;
    wire N__52180;
    wire N__52179;
    wire N__52178;
    wire N__52169;
    wire N__52160;
    wire N__52151;
    wire N__52136;
    wire N__52133;
    wire N__52130;
    wire N__52127;
    wire N__52124;
    wire N__52119;
    wire N__52116;
    wire N__52115;
    wire N__52114;
    wire N__52113;
    wire N__52112;
    wire N__52111;
    wire N__52110;
    wire N__52107;
    wire N__52106;
    wire N__52105;
    wire N__52100;
    wire N__52093;
    wire N__52088;
    wire N__52081;
    wire N__52078;
    wire N__52069;
    wire N__52066;
    wire N__52063;
    wire N__52060;
    wire N__52059;
    wire N__52058;
    wire N__52055;
    wire N__52052;
    wire N__52051;
    wire N__52046;
    wire N__52039;
    wire N__52034;
    wire N__52031;
    wire N__52026;
    wire N__52021;
    wire N__52018;
    wire N__52015;
    wire N__52012;
    wire N__52011;
    wire N__52008;
    wire N__52007;
    wire N__52004;
    wire N__52003;
    wire N__52000;
    wire N__51991;
    wire N__51988;
    wire N__51987;
    wire N__51986;
    wire N__51983;
    wire N__51982;
    wire N__51979;
    wire N__51974;
    wire N__51969;
    wire N__51962;
    wire N__51959;
    wire N__51954;
    wire N__51951;
    wire N__51950;
    wire N__51949;
    wire N__51948;
    wire N__51947;
    wire N__51946;
    wire N__51943;
    wire N__51942;
    wire N__51941;
    wire N__51940;
    wire N__51939;
    wire N__51938;
    wire N__51935;
    wire N__51934;
    wire N__51933;
    wire N__51932;
    wire N__51929;
    wire N__51928;
    wire N__51925;
    wire N__51924;
    wire N__51923;
    wire N__51922;
    wire N__51919;
    wire N__51918;
    wire N__51917;
    wire N__51914;
    wire N__51911;
    wire N__51908;
    wire N__51907;
    wire N__51900;
    wire N__51893;
    wire N__51890;
    wire N__51887;
    wire N__51884;
    wire N__51881;
    wire N__51880;
    wire N__51879;
    wire N__51878;
    wire N__51877;
    wire N__51876;
    wire N__51875;
    wire N__51874;
    wire N__51873;
    wire N__51872;
    wire N__51871;
    wire N__51870;
    wire N__51869;
    wire N__51868;
    wire N__51867;
    wire N__51864;
    wire N__51863;
    wire N__51862;
    wire N__51859;
    wire N__51856;
    wire N__51855;
    wire N__51854;
    wire N__51853;
    wire N__51852;
    wire N__51851;
    wire N__51850;
    wire N__51849;
    wire N__51848;
    wire N__51845;
    wire N__51844;
    wire N__51843;
    wire N__51842;
    wire N__51841;
    wire N__51840;
    wire N__51839;
    wire N__51826;
    wire N__51819;
    wire N__51810;
    wire N__51809;
    wire N__51808;
    wire N__51807;
    wire N__51806;
    wire N__51803;
    wire N__51802;
    wire N__51797;
    wire N__51784;
    wire N__51783;
    wire N__51782;
    wire N__51773;
    wire N__51768;
    wire N__51761;
    wire N__51758;
    wire N__51755;
    wire N__51754;
    wire N__51751;
    wire N__51748;
    wire N__51745;
    wire N__51742;
    wire N__51725;
    wire N__51724;
    wire N__51723;
    wire N__51722;
    wire N__51721;
    wire N__51720;
    wire N__51719;
    wire N__51718;
    wire N__51717;
    wire N__51716;
    wire N__51715;
    wire N__51714;
    wire N__51713;
    wire N__51712;
    wire N__51697;
    wire N__51696;
    wire N__51689;
    wire N__51686;
    wire N__51685;
    wire N__51684;
    wire N__51683;
    wire N__51678;
    wire N__51675;
    wire N__51670;
    wire N__51667;
    wire N__51654;
    wire N__51639;
    wire N__51638;
    wire N__51637;
    wire N__51636;
    wire N__51635;
    wire N__51634;
    wire N__51633;
    wire N__51632;
    wire N__51631;
    wire N__51628;
    wire N__51627;
    wire N__51626;
    wire N__51623;
    wire N__51622;
    wire N__51621;
    wire N__51618;
    wire N__51615;
    wire N__51614;
    wire N__51613;
    wire N__51612;
    wire N__51611;
    wire N__51610;
    wire N__51607;
    wire N__51604;
    wire N__51601;
    wire N__51598;
    wire N__51595;
    wire N__51594;
    wire N__51591;
    wire N__51588;
    wire N__51585;
    wire N__51584;
    wire N__51569;
    wire N__51566;
    wire N__51565;
    wire N__51564;
    wire N__51561;
    wire N__51560;
    wire N__51553;
    wire N__51552;
    wire N__51551;
    wire N__51550;
    wire N__51549;
    wire N__51548;
    wire N__51547;
    wire N__51546;
    wire N__51545;
    wire N__51544;
    wire N__51543;
    wire N__51542;
    wire N__51541;
    wire N__51532;
    wire N__51529;
    wire N__51526;
    wire N__51521;
    wire N__51516;
    wire N__51511;
    wire N__51504;
    wire N__51501;
    wire N__51500;
    wire N__51489;
    wire N__51474;
    wire N__51471;
    wire N__51460;
    wire N__51459;
    wire N__51458;
    wire N__51457;
    wire N__51454;
    wire N__51451;
    wire N__51446;
    wire N__51443;
    wire N__51440;
    wire N__51437;
    wire N__51436;
    wire N__51433;
    wire N__51428;
    wire N__51421;
    wire N__51408;
    wire N__51397;
    wire N__51394;
    wire N__51391;
    wire N__51388;
    wire N__51383;
    wire N__51380;
    wire N__51377;
    wire N__51374;
    wire N__51373;
    wire N__51370;
    wire N__51367;
    wire N__51366;
    wire N__51365;
    wire N__51364;
    wire N__51363;
    wire N__51358;
    wire N__51349;
    wire N__51340;
    wire N__51337;
    wire N__51334;
    wire N__51325;
    wire N__51322;
    wire N__51315;
    wire N__51312;
    wire N__51311;
    wire N__51310;
    wire N__51309;
    wire N__51308;
    wire N__51307;
    wire N__51306;
    wire N__51305;
    wire N__51304;
    wire N__51303;
    wire N__51302;
    wire N__51301;
    wire N__51300;
    wire N__51299;
    wire N__51298;
    wire N__51283;
    wire N__51280;
    wire N__51279;
    wire N__51278;
    wire N__51277;
    wire N__51276;
    wire N__51275;
    wire N__51274;
    wire N__51273;
    wire N__51272;
    wire N__51271;
    wire N__51270;
    wire N__51269;
    wire N__51268;
    wire N__51267;
    wire N__51266;
    wire N__51265;
    wire N__51264;
    wire N__51261;
    wire N__51256;
    wire N__51251;
    wire N__51244;
    wire N__51241;
    wire N__51232;
    wire N__51229;
    wire N__51226;
    wire N__51223;
    wire N__51218;
    wire N__51213;
    wire N__51212;
    wire N__51207;
    wire N__51204;
    wire N__51203;
    wire N__51202;
    wire N__51191;
    wire N__51184;
    wire N__51175;
    wire N__51172;
    wire N__51167;
    wire N__51164;
    wire N__51161;
    wire N__51158;
    wire N__51155;
    wire N__51152;
    wire N__51141;
    wire N__51138;
    wire N__51133;
    wire N__51130;
    wire N__51117;
    wire N__51114;
    wire N__51101;
    wire N__51096;
    wire N__51081;
    wire N__51074;
    wire N__51063;
    wire N__51060;
    wire N__51055;
    wire N__51050;
    wire N__51039;
    wire N__51034;
    wire N__51031;
    wire N__51026;
    wire N__51023;
    wire N__51020;
    wire N__51017;
    wire N__51014;
    wire N__50999;
    wire N__50998;
    wire N__50997;
    wire N__50992;
    wire N__50987;
    wire N__50968;
    wire N__50961;
    wire N__50958;
    wire N__50949;
    wire N__50942;
    wire N__50939;
    wire N__50936;
    wire N__50933;
    wire N__50928;
    wire N__50925;
    wire N__50920;
    wire N__50917;
    wire N__50914;
    wire N__50911;
    wire N__50906;
    wire N__50903;
    wire N__50900;
    wire N__50897;
    wire N__50892;
    wire N__50887;
    wire N__50882;
    wire N__50879;
    wire N__50872;
    wire N__50869;
    wire N__50868;
    wire N__50865;
    wire N__50864;
    wire N__50863;
    wire N__50860;
    wire N__50857;
    wire N__50854;
    wire N__50851;
    wire N__50850;
    wire N__50847;
    wire N__50842;
    wire N__50839;
    wire N__50838;
    wire N__50835;
    wire N__50832;
    wire N__50831;
    wire N__50826;
    wire N__50823;
    wire N__50822;
    wire N__50819;
    wire N__50816;
    wire N__50813;
    wire N__50810;
    wire N__50807;
    wire N__50804;
    wire N__50801;
    wire N__50796;
    wire N__50793;
    wire N__50790;
    wire N__50787;
    wire N__50784;
    wire N__50781;
    wire N__50774;
    wire N__50767;
    wire N__50766;
    wire N__50765;
    wire N__50762;
    wire N__50761;
    wire N__50758;
    wire N__50757;
    wire N__50752;
    wire N__50751;
    wire N__50750;
    wire N__50749;
    wire N__50748;
    wire N__50747;
    wire N__50744;
    wire N__50741;
    wire N__50738;
    wire N__50735;
    wire N__50726;
    wire N__50725;
    wire N__50724;
    wire N__50721;
    wire N__50720;
    wire N__50719;
    wire N__50718;
    wire N__50717;
    wire N__50716;
    wire N__50713;
    wire N__50708;
    wire N__50703;
    wire N__50702;
    wire N__50699;
    wire N__50696;
    wire N__50693;
    wire N__50690;
    wire N__50687;
    wire N__50682;
    wire N__50679;
    wire N__50678;
    wire N__50677;
    wire N__50676;
    wire N__50673;
    wire N__50670;
    wire N__50667;
    wire N__50664;
    wire N__50663;
    wire N__50660;
    wire N__50651;
    wire N__50646;
    wire N__50643;
    wire N__50640;
    wire N__50637;
    wire N__50632;
    wire N__50629;
    wire N__50626;
    wire N__50623;
    wire N__50614;
    wire N__50611;
    wire N__50608;
    wire N__50593;
    wire N__50590;
    wire N__50587;
    wire N__50584;
    wire N__50581;
    wire N__50578;
    wire N__50577;
    wire N__50576;
    wire N__50575;
    wire N__50574;
    wire N__50573;
    wire N__50570;
    wire N__50563;
    wire N__50562;
    wire N__50561;
    wire N__50560;
    wire N__50559;
    wire N__50558;
    wire N__50557;
    wire N__50554;
    wire N__50551;
    wire N__50548;
    wire N__50545;
    wire N__50542;
    wire N__50531;
    wire N__50526;
    wire N__50525;
    wire N__50522;
    wire N__50519;
    wire N__50514;
    wire N__50511;
    wire N__50508;
    wire N__50505;
    wire N__50500;
    wire N__50497;
    wire N__50494;
    wire N__50491;
    wire N__50488;
    wire N__50485;
    wire N__50482;
    wire N__50477;
    wire N__50472;
    wire N__50467;
    wire N__50466;
    wire N__50465;
    wire N__50464;
    wire N__50463;
    wire N__50460;
    wire N__50459;
    wire N__50458;
    wire N__50457;
    wire N__50454;
    wire N__50451;
    wire N__50448;
    wire N__50445;
    wire N__50444;
    wire N__50443;
    wire N__50442;
    wire N__50439;
    wire N__50436;
    wire N__50433;
    wire N__50430;
    wire N__50427;
    wire N__50422;
    wire N__50419;
    wire N__50416;
    wire N__50413;
    wire N__50410;
    wire N__50409;
    wire N__50408;
    wire N__50401;
    wire N__50398;
    wire N__50393;
    wire N__50388;
    wire N__50385;
    wire N__50378;
    wire N__50377;
    wire N__50374;
    wire N__50371;
    wire N__50370;
    wire N__50369;
    wire N__50360;
    wire N__50357;
    wire N__50354;
    wire N__50351;
    wire N__50348;
    wire N__50345;
    wire N__50342;
    wire N__50339;
    wire N__50336;
    wire N__50331;
    wire N__50328;
    wire N__50323;
    wire N__50318;
    wire N__50315;
    wire N__50310;
    wire N__50307;
    wire N__50304;
    wire N__50301;
    wire N__50298;
    wire N__50293;
    wire N__50292;
    wire N__50291;
    wire N__50290;
    wire N__50289;
    wire N__50288;
    wire N__50285;
    wire N__50284;
    wire N__50273;
    wire N__50270;
    wire N__50267;
    wire N__50264;
    wire N__50261;
    wire N__50258;
    wire N__50257;
    wire N__50254;
    wire N__50251;
    wire N__50248;
    wire N__50245;
    wire N__50242;
    wire N__50237;
    wire N__50234;
    wire N__50227;
    wire N__50224;
    wire N__50221;
    wire N__50218;
    wire N__50215;
    wire N__50212;
    wire N__50209;
    wire N__50208;
    wire N__50207;
    wire N__50206;
    wire N__50205;
    wire N__50202;
    wire N__50199;
    wire N__50198;
    wire N__50195;
    wire N__50194;
    wire N__50193;
    wire N__50190;
    wire N__50189;
    wire N__50188;
    wire N__50185;
    wire N__50180;
    wire N__50179;
    wire N__50176;
    wire N__50175;
    wire N__50174;
    wire N__50173;
    wire N__50172;
    wire N__50171;
    wire N__50170;
    wire N__50169;
    wire N__50168;
    wire N__50167;
    wire N__50166;
    wire N__50165;
    wire N__50162;
    wire N__50157;
    wire N__50154;
    wire N__50153;
    wire N__50152;
    wire N__50147;
    wire N__50142;
    wire N__50141;
    wire N__50140;
    wire N__50139;
    wire N__50138;
    wire N__50137;
    wire N__50136;
    wire N__50135;
    wire N__50134;
    wire N__50131;
    wire N__50128;
    wire N__50125;
    wire N__50120;
    wire N__50115;
    wire N__50114;
    wire N__50113;
    wire N__50112;
    wire N__50111;
    wire N__50106;
    wire N__50101;
    wire N__50096;
    wire N__50089;
    wire N__50084;
    wire N__50081;
    wire N__50078;
    wire N__50075;
    wire N__50070;
    wire N__50065;
    wire N__50064;
    wire N__50061;
    wire N__50060;
    wire N__50059;
    wire N__50058;
    wire N__50053;
    wire N__50052;
    wire N__50049;
    wire N__50040;
    wire N__50039;
    wire N__50038;
    wire N__50037;
    wire N__50036;
    wire N__50033;
    wire N__50030;
    wire N__50027;
    wire N__50024;
    wire N__50021;
    wire N__50020;
    wire N__50019;
    wire N__50018;
    wire N__50017;
    wire N__50016;
    wire N__50015;
    wire N__50014;
    wire N__50013;
    wire N__50012;
    wire N__50003;
    wire N__49996;
    wire N__49991;
    wire N__49984;
    wire N__49979;
    wire N__49978;
    wire N__49977;
    wire N__49974;
    wire N__49971;
    wire N__49966;
    wire N__49961;
    wire N__49956;
    wire N__49953;
    wire N__49944;
    wire N__49939;
    wire N__49938;
    wire N__49937;
    wire N__49934;
    wire N__49929;
    wire N__49924;
    wire N__49919;
    wire N__49918;
    wire N__49917;
    wire N__49916;
    wire N__49915;
    wire N__49912;
    wire N__49905;
    wire N__49902;
    wire N__49897;
    wire N__49892;
    wire N__49885;
    wire N__49878;
    wire N__49873;
    wire N__49864;
    wire N__49859;
    wire N__49854;
    wire N__49853;
    wire N__49852;
    wire N__49851;
    wire N__49848;
    wire N__49841;
    wire N__49836;
    wire N__49835;
    wire N__49834;
    wire N__49829;
    wire N__49824;
    wire N__49821;
    wire N__49814;
    wire N__49811;
    wire N__49806;
    wire N__49803;
    wire N__49802;
    wire N__49801;
    wire N__49798;
    wire N__49797;
    wire N__49794;
    wire N__49787;
    wire N__49784;
    wire N__49781;
    wire N__49778;
    wire N__49775;
    wire N__49768;
    wire N__49763;
    wire N__49750;
    wire N__49747;
    wire N__49744;
    wire N__49741;
    wire N__49738;
    wire N__49735;
    wire N__49732;
    wire N__49729;
    wire N__49726;
    wire N__49723;
    wire N__49720;
    wire N__49717;
    wire N__49716;
    wire N__49713;
    wire N__49710;
    wire N__49707;
    wire N__49702;
    wire N__49701;
    wire N__49700;
    wire N__49699;
    wire N__49698;
    wire N__49697;
    wire N__49696;
    wire N__49695;
    wire N__49694;
    wire N__49693;
    wire N__49692;
    wire N__49691;
    wire N__49690;
    wire N__49663;
    wire N__49660;
    wire N__49657;
    wire N__49654;
    wire N__49651;
    wire N__49648;
    wire N__49645;
    wire N__49644;
    wire N__49641;
    wire N__49638;
    wire N__49637;
    wire N__49634;
    wire N__49631;
    wire N__49628;
    wire N__49625;
    wire N__49624;
    wire N__49623;
    wire N__49620;
    wire N__49617;
    wire N__49614;
    wire N__49611;
    wire N__49608;
    wire N__49607;
    wire N__49606;
    wire N__49601;
    wire N__49596;
    wire N__49593;
    wire N__49590;
    wire N__49587;
    wire N__49576;
    wire N__49573;
    wire N__49570;
    wire N__49567;
    wire N__49564;
    wire N__49561;
    wire N__49558;
    wire N__49555;
    wire N__49552;
    wire N__49549;
    wire N__49546;
    wire N__49545;
    wire N__49544;
    wire N__49541;
    wire N__49538;
    wire N__49535;
    wire N__49534;
    wire N__49533;
    wire N__49530;
    wire N__49527;
    wire N__49526;
    wire N__49523;
    wire N__49520;
    wire N__49517;
    wire N__49512;
    wire N__49509;
    wire N__49502;
    wire N__49501;
    wire N__49500;
    wire N__49497;
    wire N__49494;
    wire N__49493;
    wire N__49490;
    wire N__49485;
    wire N__49480;
    wire N__49477;
    wire N__49472;
    wire N__49469;
    wire N__49466;
    wire N__49465;
    wire N__49462;
    wire N__49457;
    wire N__49454;
    wire N__49451;
    wire N__49448;
    wire N__49445;
    wire N__49442;
    wire N__49439;
    wire N__49436;
    wire N__49431;
    wire N__49428;
    wire N__49425;
    wire N__49422;
    wire N__49417;
    wire N__49416;
    wire N__49413;
    wire N__49410;
    wire N__49407;
    wire N__49404;
    wire N__49401;
    wire N__49398;
    wire N__49395;
    wire N__49392;
    wire N__49389;
    wire N__49384;
    wire N__49383;
    wire N__49382;
    wire N__49381;
    wire N__49380;
    wire N__49379;
    wire N__49378;
    wire N__49377;
    wire N__49376;
    wire N__49375;
    wire N__49354;
    wire N__49351;
    wire N__49348;
    wire N__49345;
    wire N__49344;
    wire N__49343;
    wire N__49342;
    wire N__49339;
    wire N__49336;
    wire N__49335;
    wire N__49332;
    wire N__49329;
    wire N__49326;
    wire N__49323;
    wire N__49320;
    wire N__49315;
    wire N__49314;
    wire N__49311;
    wire N__49306;
    wire N__49303;
    wire N__49300;
    wire N__49297;
    wire N__49294;
    wire N__49289;
    wire N__49288;
    wire N__49285;
    wire N__49282;
    wire N__49279;
    wire N__49276;
    wire N__49273;
    wire N__49266;
    wire N__49263;
    wire N__49260;
    wire N__49255;
    wire N__49252;
    wire N__49249;
    wire N__49246;
    wire N__49243;
    wire N__49242;
    wire N__49239;
    wire N__49236;
    wire N__49233;
    wire N__49230;
    wire N__49227;
    wire N__49224;
    wire N__49219;
    wire N__49218;
    wire N__49215;
    wire N__49212;
    wire N__49209;
    wire N__49206;
    wire N__49203;
    wire N__49200;
    wire N__49195;
    wire N__49192;
    wire N__49189;
    wire N__49186;
    wire N__49183;
    wire N__49180;
    wire N__49177;
    wire N__49174;
    wire N__49171;
    wire N__49168;
    wire N__49165;
    wire N__49162;
    wire N__49159;
    wire N__49158;
    wire N__49155;
    wire N__49152;
    wire N__49149;
    wire N__49146;
    wire N__49143;
    wire N__49140;
    wire N__49137;
    wire N__49134;
    wire N__49129;
    wire N__49126;
    wire N__49123;
    wire N__49120;
    wire N__49117;
    wire N__49114;
    wire N__49111;
    wire N__49108;
    wire N__49105;
    wire N__49102;
    wire N__49099;
    wire N__49096;
    wire N__49093;
    wire N__49090;
    wire N__49087;
    wire N__49084;
    wire N__49081;
    wire N__49078;
    wire N__49075;
    wire N__49072;
    wire N__49069;
    wire N__49066;
    wire N__49063;
    wire N__49060;
    wire N__49057;
    wire N__49054;
    wire N__49051;
    wire N__49048;
    wire N__49045;
    wire N__49042;
    wire N__49039;
    wire N__49036;
    wire N__49033;
    wire N__49030;
    wire N__49027;
    wire N__49024;
    wire N__49021;
    wire N__49018;
    wire N__49015;
    wire N__49012;
    wire N__49009;
    wire N__49006;
    wire N__49003;
    wire N__49000;
    wire N__48997;
    wire N__48994;
    wire N__48991;
    wire N__48988;
    wire N__48987;
    wire N__48986;
    wire N__48985;
    wire N__48982;
    wire N__48979;
    wire N__48976;
    wire N__48975;
    wire N__48972;
    wire N__48971;
    wire N__48970;
    wire N__48969;
    wire N__48968;
    wire N__48967;
    wire N__48964;
    wire N__48959;
    wire N__48958;
    wire N__48955;
    wire N__48952;
    wire N__48949;
    wire N__48946;
    wire N__48945;
    wire N__48944;
    wire N__48941;
    wire N__48940;
    wire N__48939;
    wire N__48938;
    wire N__48937;
    wire N__48934;
    wire N__48931;
    wire N__48930;
    wire N__48929;
    wire N__48924;
    wire N__48921;
    wire N__48918;
    wire N__48911;
    wire N__48910;
    wire N__48907;
    wire N__48904;
    wire N__48901;
    wire N__48898;
    wire N__48895;
    wire N__48892;
    wire N__48891;
    wire N__48890;
    wire N__48889;
    wire N__48886;
    wire N__48883;
    wire N__48880;
    wire N__48877;
    wire N__48874;
    wire N__48869;
    wire N__48868;
    wire N__48865;
    wire N__48862;
    wire N__48859;
    wire N__48858;
    wire N__48851;
    wire N__48846;
    wire N__48843;
    wire N__48840;
    wire N__48837;
    wire N__48834;
    wire N__48833;
    wire N__48832;
    wire N__48831;
    wire N__48830;
    wire N__48829;
    wire N__48826;
    wire N__48817;
    wire N__48814;
    wire N__48813;
    wire N__48810;
    wire N__48807;
    wire N__48804;
    wire N__48801;
    wire N__48798;
    wire N__48785;
    wire N__48782;
    wire N__48779;
    wire N__48776;
    wire N__48773;
    wire N__48770;
    wire N__48769;
    wire N__48768;
    wire N__48763;
    wire N__48760;
    wire N__48757;
    wire N__48754;
    wire N__48745;
    wire N__48736;
    wire N__48733;
    wire N__48730;
    wire N__48725;
    wire N__48722;
    wire N__48719;
    wire N__48716;
    wire N__48713;
    wire N__48710;
    wire N__48709;
    wire N__48708;
    wire N__48707;
    wire N__48706;
    wire N__48705;
    wire N__48702;
    wire N__48695;
    wire N__48688;
    wire N__48683;
    wire N__48678;
    wire N__48671;
    wire N__48666;
    wire N__48655;
    wire N__48652;
    wire N__48649;
    wire N__48646;
    wire N__48643;
    wire N__48640;
    wire N__48637;
    wire N__48634;
    wire N__48631;
    wire N__48628;
    wire N__48625;
    wire N__48622;
    wire N__48619;
    wire N__48616;
    wire N__48613;
    wire N__48610;
    wire N__48607;
    wire N__48604;
    wire N__48601;
    wire N__48600;
    wire N__48599;
    wire N__48598;
    wire N__48597;
    wire N__48594;
    wire N__48591;
    wire N__48588;
    wire N__48587;
    wire N__48584;
    wire N__48583;
    wire N__48582;
    wire N__48579;
    wire N__48578;
    wire N__48577;
    wire N__48574;
    wire N__48571;
    wire N__48570;
    wire N__48567;
    wire N__48566;
    wire N__48565;
    wire N__48562;
    wire N__48559;
    wire N__48556;
    wire N__48553;
    wire N__48550;
    wire N__48549;
    wire N__48548;
    wire N__48545;
    wire N__48544;
    wire N__48541;
    wire N__48540;
    wire N__48535;
    wire N__48532;
    wire N__48531;
    wire N__48528;
    wire N__48525;
    wire N__48522;
    wire N__48521;
    wire N__48518;
    wire N__48515;
    wire N__48512;
    wire N__48507;
    wire N__48504;
    wire N__48501;
    wire N__48498;
    wire N__48495;
    wire N__48492;
    wire N__48489;
    wire N__48484;
    wire N__48481;
    wire N__48480;
    wire N__48473;
    wire N__48470;
    wire N__48469;
    wire N__48468;
    wire N__48465;
    wire N__48456;
    wire N__48453;
    wire N__48440;
    wire N__48437;
    wire N__48436;
    wire N__48433;
    wire N__48430;
    wire N__48427;
    wire N__48424;
    wire N__48417;
    wire N__48412;
    wire N__48409;
    wire N__48394;
    wire N__48391;
    wire N__48388;
    wire N__48385;
    wire N__48384;
    wire N__48381;
    wire N__48378;
    wire N__48375;
    wire N__48372;
    wire N__48367;
    wire N__48364;
    wire N__48361;
    wire N__48358;
    wire N__48355;
    wire N__48352;
    wire N__48349;
    wire N__48346;
    wire N__48343;
    wire N__48340;
    wire N__48337;
    wire N__48334;
    wire N__48333;
    wire N__48332;
    wire N__48331;
    wire N__48330;
    wire N__48329;
    wire N__48328;
    wire N__48327;
    wire N__48326;
    wire N__48325;
    wire N__48324;
    wire N__48321;
    wire N__48318;
    wire N__48315;
    wire N__48312;
    wire N__48311;
    wire N__48308;
    wire N__48305;
    wire N__48302;
    wire N__48299;
    wire N__48296;
    wire N__48293;
    wire N__48290;
    wire N__48289;
    wire N__48284;
    wire N__48283;
    wire N__48280;
    wire N__48279;
    wire N__48278;
    wire N__48277;
    wire N__48276;
    wire N__48275;
    wire N__48272;
    wire N__48269;
    wire N__48266;
    wire N__48263;
    wire N__48258;
    wire N__48255;
    wire N__48254;
    wire N__48253;
    wire N__48250;
    wire N__48247;
    wire N__48244;
    wire N__48241;
    wire N__48238;
    wire N__48237;
    wire N__48234;
    wire N__48223;
    wire N__48218;
    wire N__48215;
    wire N__48208;
    wire N__48205;
    wire N__48202;
    wire N__48197;
    wire N__48194;
    wire N__48189;
    wire N__48186;
    wire N__48181;
    wire N__48176;
    wire N__48173;
    wire N__48170;
    wire N__48167;
    wire N__48158;
    wire N__48145;
    wire N__48144;
    wire N__48141;
    wire N__48138;
    wire N__48135;
    wire N__48134;
    wire N__48133;
    wire N__48132;
    wire N__48129;
    wire N__48128;
    wire N__48127;
    wire N__48126;
    wire N__48125;
    wire N__48124;
    wire N__48121;
    wire N__48120;
    wire N__48115;
    wire N__48114;
    wire N__48113;
    wire N__48112;
    wire N__48111;
    wire N__48110;
    wire N__48107;
    wire N__48106;
    wire N__48103;
    wire N__48092;
    wire N__48089;
    wire N__48086;
    wire N__48085;
    wire N__48082;
    wire N__48075;
    wire N__48072;
    wire N__48069;
    wire N__48066;
    wire N__48065;
    wire N__48062;
    wire N__48061;
    wire N__48060;
    wire N__48055;
    wire N__48050;
    wire N__48047;
    wire N__48042;
    wire N__48037;
    wire N__48034;
    wire N__48031;
    wire N__48028;
    wire N__48027;
    wire N__48024;
    wire N__48021;
    wire N__48020;
    wire N__48019;
    wire N__48018;
    wire N__48015;
    wire N__48010;
    wire N__48003;
    wire N__47998;
    wire N__47995;
    wire N__47992;
    wire N__47989;
    wire N__47984;
    wire N__47981;
    wire N__47962;
    wire N__47959;
    wire N__47956;
    wire N__47955;
    wire N__47952;
    wire N__47949;
    wire N__47946;
    wire N__47943;
    wire N__47938;
    wire N__47935;
    wire N__47932;
    wire N__47929;
    wire N__47926;
    wire N__47923;
    wire N__47920;
    wire N__47919;
    wire N__47916;
    wire N__47913;
    wire N__47908;
    wire N__47905;
    wire N__47902;
    wire N__47899;
    wire N__47896;
    wire N__47893;
    wire N__47890;
    wire N__47887;
    wire N__47884;
    wire N__47883;
    wire N__47880;
    wire N__47877;
    wire N__47874;
    wire N__47871;
    wire N__47868;
    wire N__47865;
    wire N__47862;
    wire N__47857;
    wire N__47854;
    wire N__47851;
    wire N__47848;
    wire N__47845;
    wire N__47842;
    wire N__47839;
    wire N__47838;
    wire N__47835;
    wire N__47832;
    wire N__47831;
    wire N__47826;
    wire N__47823;
    wire N__47822;
    wire N__47821;
    wire N__47816;
    wire N__47813;
    wire N__47810;
    wire N__47807;
    wire N__47804;
    wire N__47801;
    wire N__47796;
    wire N__47795;
    wire N__47794;
    wire N__47791;
    wire N__47788;
    wire N__47785;
    wire N__47782;
    wire N__47779;
    wire N__47776;
    wire N__47773;
    wire N__47770;
    wire N__47767;
    wire N__47762;
    wire N__47759;
    wire N__47752;
    wire N__47749;
    wire N__47746;
    wire N__47743;
    wire N__47740;
    wire N__47737;
    wire N__47736;
    wire N__47735;
    wire N__47732;
    wire N__47731;
    wire N__47728;
    wire N__47727;
    wire N__47724;
    wire N__47721;
    wire N__47720;
    wire N__47719;
    wire N__47716;
    wire N__47715;
    wire N__47712;
    wire N__47709;
    wire N__47708;
    wire N__47707;
    wire N__47706;
    wire N__47705;
    wire N__47704;
    wire N__47703;
    wire N__47702;
    wire N__47701;
    wire N__47700;
    wire N__47697;
    wire N__47694;
    wire N__47685;
    wire N__47682;
    wire N__47679;
    wire N__47674;
    wire N__47667;
    wire N__47660;
    wire N__47657;
    wire N__47654;
    wire N__47653;
    wire N__47650;
    wire N__47647;
    wire N__47644;
    wire N__47635;
    wire N__47634;
    wire N__47631;
    wire N__47628;
    wire N__47625;
    wire N__47620;
    wire N__47615;
    wire N__47612;
    wire N__47605;
    wire N__47598;
    wire N__47595;
    wire N__47592;
    wire N__47589;
    wire N__47586;
    wire N__47581;
    wire N__47578;
    wire N__47575;
    wire N__47572;
    wire N__47569;
    wire N__47566;
    wire N__47563;
    wire N__47560;
    wire N__47557;
    wire N__47554;
    wire N__47551;
    wire N__47548;
    wire N__47545;
    wire N__47542;
    wire N__47539;
    wire N__47536;
    wire N__47533;
    wire N__47530;
    wire N__47527;
    wire N__47524;
    wire N__47521;
    wire N__47518;
    wire N__47517;
    wire N__47516;
    wire N__47513;
    wire N__47512;
    wire N__47511;
    wire N__47510;
    wire N__47505;
    wire N__47498;
    wire N__47497;
    wire N__47494;
    wire N__47493;
    wire N__47488;
    wire N__47487;
    wire N__47484;
    wire N__47483;
    wire N__47482;
    wire N__47481;
    wire N__47478;
    wire N__47475;
    wire N__47472;
    wire N__47469;
    wire N__47468;
    wire N__47467;
    wire N__47464;
    wire N__47461;
    wire N__47458;
    wire N__47455;
    wire N__47454;
    wire N__47453;
    wire N__47450;
    wire N__47447;
    wire N__47442;
    wire N__47439;
    wire N__47436;
    wire N__47435;
    wire N__47432;
    wire N__47429;
    wire N__47424;
    wire N__47423;
    wire N__47420;
    wire N__47417;
    wire N__47416;
    wire N__47411;
    wire N__47406;
    wire N__47405;
    wire N__47402;
    wire N__47399;
    wire N__47398;
    wire N__47395;
    wire N__47392;
    wire N__47389;
    wire N__47386;
    wire N__47383;
    wire N__47380;
    wire N__47377;
    wire N__47376;
    wire N__47375;
    wire N__47374;
    wire N__47373;
    wire N__47370;
    wire N__47367;
    wire N__47364;
    wire N__47361;
    wire N__47358;
    wire N__47355;
    wire N__47348;
    wire N__47345;
    wire N__47340;
    wire N__47335;
    wire N__47332;
    wire N__47327;
    wire N__47320;
    wire N__47313;
    wire N__47310;
    wire N__47299;
    wire N__47296;
    wire N__47293;
    wire N__47290;
    wire N__47285;
    wire N__47282;
    wire N__47279;
    wire N__47276;
    wire N__47273;
    wire N__47268;
    wire N__47263;
    wire N__47262;
    wire N__47259;
    wire N__47256;
    wire N__47255;
    wire N__47254;
    wire N__47253;
    wire N__47250;
    wire N__47249;
    wire N__47246;
    wire N__47245;
    wire N__47242;
    wire N__47239;
    wire N__47238;
    wire N__47235;
    wire N__47232;
    wire N__47229;
    wire N__47228;
    wire N__47225;
    wire N__47224;
    wire N__47221;
    wire N__47220;
    wire N__47217;
    wire N__47214;
    wire N__47213;
    wire N__47210;
    wire N__47209;
    wire N__47206;
    wire N__47201;
    wire N__47198;
    wire N__47197;
    wire N__47196;
    wire N__47193;
    wire N__47190;
    wire N__47187;
    wire N__47184;
    wire N__47183;
    wire N__47182;
    wire N__47181;
    wire N__47178;
    wire N__47175;
    wire N__47172;
    wire N__47169;
    wire N__47168;
    wire N__47167;
    wire N__47164;
    wire N__47157;
    wire N__47152;
    wire N__47149;
    wire N__47146;
    wire N__47145;
    wire N__47144;
    wire N__47139;
    wire N__47136;
    wire N__47133;
    wire N__47130;
    wire N__47121;
    wire N__47118;
    wire N__47115;
    wire N__47112;
    wire N__47111;
    wire N__47106;
    wire N__47101;
    wire N__47098;
    wire N__47095;
    wire N__47090;
    wire N__47085;
    wire N__47078;
    wire N__47075;
    wire N__47072;
    wire N__47071;
    wire N__47070;
    wire N__47061;
    wire N__47050;
    wire N__47047;
    wire N__47044;
    wire N__47035;
    wire N__47032;
    wire N__47029;
    wire N__47026;
    wire N__47023;
    wire N__47020;
    wire N__47017;
    wire N__47014;
    wire N__47011;
    wire N__47010;
    wire N__47007;
    wire N__47004;
    wire N__46999;
    wire N__46996;
    wire N__46993;
    wire N__46990;
    wire N__46987;
    wire N__46984;
    wire N__46983;
    wire N__46980;
    wire N__46979;
    wire N__46978;
    wire N__46975;
    wire N__46972;
    wire N__46969;
    wire N__46966;
    wire N__46963;
    wire N__46962;
    wire N__46961;
    wire N__46960;
    wire N__46955;
    wire N__46952;
    wire N__46951;
    wire N__46948;
    wire N__46941;
    wire N__46940;
    wire N__46939;
    wire N__46938;
    wire N__46937;
    wire N__46936;
    wire N__46931;
    wire N__46928;
    wire N__46923;
    wire N__46920;
    wire N__46917;
    wire N__46912;
    wire N__46909;
    wire N__46908;
    wire N__46907;
    wire N__46906;
    wire N__46905;
    wire N__46904;
    wire N__46899;
    wire N__46894;
    wire N__46891;
    wire N__46890;
    wire N__46889;
    wire N__46888;
    wire N__46883;
    wire N__46880;
    wire N__46877;
    wire N__46874;
    wire N__46871;
    wire N__46868;
    wire N__46867;
    wire N__46866;
    wire N__46865;
    wire N__46864;
    wire N__46861;
    wire N__46856;
    wire N__46853;
    wire N__46850;
    wire N__46847;
    wire N__46840;
    wire N__46833;
    wire N__46830;
    wire N__46827;
    wire N__46824;
    wire N__46821;
    wire N__46798;
    wire N__46797;
    wire N__46794;
    wire N__46791;
    wire N__46788;
    wire N__46785;
    wire N__46782;
    wire N__46779;
    wire N__46776;
    wire N__46771;
    wire N__46768;
    wire N__46767;
    wire N__46764;
    wire N__46761;
    wire N__46758;
    wire N__46755;
    wire N__46752;
    wire N__46749;
    wire N__46744;
    wire N__46741;
    wire N__46738;
    wire N__46735;
    wire N__46734;
    wire N__46733;
    wire N__46732;
    wire N__46731;
    wire N__46730;
    wire N__46729;
    wire N__46726;
    wire N__46719;
    wire N__46714;
    wire N__46711;
    wire N__46702;
    wire N__46701;
    wire N__46698;
    wire N__46695;
    wire N__46692;
    wire N__46689;
    wire N__46686;
    wire N__46683;
    wire N__46680;
    wire N__46675;
    wire N__46672;
    wire N__46669;
    wire N__46666;
    wire N__46663;
    wire N__46660;
    wire N__46657;
    wire N__46654;
    wire N__46651;
    wire N__46648;
    wire N__46645;
    wire N__46642;
    wire N__46639;
    wire N__46638;
    wire N__46635;
    wire N__46632;
    wire N__46627;
    wire N__46624;
    wire N__46623;
    wire N__46620;
    wire N__46617;
    wire N__46614;
    wire N__46611;
    wire N__46606;
    wire N__46603;
    wire N__46602;
    wire N__46601;
    wire N__46598;
    wire N__46595;
    wire N__46594;
    wire N__46593;
    wire N__46590;
    wire N__46589;
    wire N__46586;
    wire N__46583;
    wire N__46580;
    wire N__46577;
    wire N__46574;
    wire N__46571;
    wire N__46568;
    wire N__46567;
    wire N__46566;
    wire N__46559;
    wire N__46554;
    wire N__46551;
    wire N__46546;
    wire N__46541;
    wire N__46536;
    wire N__46535;
    wire N__46532;
    wire N__46529;
    wire N__46526;
    wire N__46519;
    wire N__46518;
    wire N__46515;
    wire N__46512;
    wire N__46509;
    wire N__46506;
    wire N__46503;
    wire N__46500;
    wire N__46495;
    wire N__46492;
    wire N__46489;
    wire N__46486;
    wire N__46483;
    wire N__46480;
    wire N__46477;
    wire N__46474;
    wire N__46471;
    wire N__46468;
    wire N__46465;
    wire N__46462;
    wire N__46459;
    wire N__46456;
    wire N__46453;
    wire N__46450;
    wire N__46447;
    wire N__46444;
    wire N__46441;
    wire N__46438;
    wire N__46435;
    wire N__46432;
    wire N__46429;
    wire N__46426;
    wire N__46423;
    wire N__46420;
    wire N__46417;
    wire N__46416;
    wire N__46415;
    wire N__46414;
    wire N__46413;
    wire N__46412;
    wire N__46409;
    wire N__46402;
    wire N__46399;
    wire N__46396;
    wire N__46387;
    wire N__46384;
    wire N__46381;
    wire N__46378;
    wire N__46375;
    wire N__46372;
    wire N__46369;
    wire N__46366;
    wire N__46363;
    wire N__46360;
    wire N__46357;
    wire N__46354;
    wire N__46351;
    wire N__46348;
    wire N__46345;
    wire N__46342;
    wire N__46339;
    wire N__46336;
    wire N__46333;
    wire N__46330;
    wire N__46327;
    wire N__46324;
    wire N__46321;
    wire N__46318;
    wire N__46315;
    wire N__46312;
    wire N__46309;
    wire N__46306;
    wire N__46303;
    wire N__46302;
    wire N__46299;
    wire N__46296;
    wire N__46291;
    wire N__46290;
    wire N__46289;
    wire N__46288;
    wire N__46285;
    wire N__46282;
    wire N__46279;
    wire N__46276;
    wire N__46273;
    wire N__46272;
    wire N__46271;
    wire N__46266;
    wire N__46265;
    wire N__46264;
    wire N__46261;
    wire N__46258;
    wire N__46255;
    wire N__46252;
    wire N__46249;
    wire N__46246;
    wire N__46243;
    wire N__46240;
    wire N__46233;
    wire N__46228;
    wire N__46225;
    wire N__46222;
    wire N__46219;
    wire N__46216;
    wire N__46213;
    wire N__46210;
    wire N__46207;
    wire N__46204;
    wire N__46201;
    wire N__46196;
    wire N__46193;
    wire N__46190;
    wire N__46187;
    wire N__46184;
    wire N__46177;
    wire N__46174;
    wire N__46173;
    wire N__46170;
    wire N__46167;
    wire N__46164;
    wire N__46161;
    wire N__46156;
    wire N__46153;
    wire N__46150;
    wire N__46149;
    wire N__46146;
    wire N__46143;
    wire N__46140;
    wire N__46137;
    wire N__46132;
    wire N__46131;
    wire N__46128;
    wire N__46125;
    wire N__46124;
    wire N__46123;
    wire N__46118;
    wire N__46115;
    wire N__46112;
    wire N__46111;
    wire N__46106;
    wire N__46105;
    wire N__46102;
    wire N__46099;
    wire N__46096;
    wire N__46093;
    wire N__46090;
    wire N__46087;
    wire N__46084;
    wire N__46081;
    wire N__46076;
    wire N__46073;
    wire N__46070;
    wire N__46067;
    wire N__46060;
    wire N__46057;
    wire N__46054;
    wire N__46051;
    wire N__46048;
    wire N__46045;
    wire N__46042;
    wire N__46039;
    wire N__46036;
    wire N__46033;
    wire N__46030;
    wire N__46027;
    wire N__46024;
    wire N__46021;
    wire N__46018;
    wire N__46017;
    wire N__46014;
    wire N__46011;
    wire N__46008;
    wire N__46005;
    wire N__46000;
    wire N__45997;
    wire N__45994;
    wire N__45991;
    wire N__45988;
    wire N__45985;
    wire N__45982;
    wire N__45979;
    wire N__45976;
    wire N__45975;
    wire N__45974;
    wire N__45971;
    wire N__45966;
    wire N__45963;
    wire N__45960;
    wire N__45955;
    wire N__45952;
    wire N__45949;
    wire N__45946;
    wire N__45943;
    wire N__45940;
    wire N__45937;
    wire N__45936;
    wire N__45933;
    wire N__45932;
    wire N__45931;
    wire N__45928;
    wire N__45927;
    wire N__45926;
    wire N__45925;
    wire N__45922;
    wire N__45919;
    wire N__45916;
    wire N__45913;
    wire N__45910;
    wire N__45909;
    wire N__45908;
    wire N__45907;
    wire N__45904;
    wire N__45903;
    wire N__45900;
    wire N__45899;
    wire N__45896;
    wire N__45893;
    wire N__45890;
    wire N__45885;
    wire N__45882;
    wire N__45881;
    wire N__45880;
    wire N__45877;
    wire N__45874;
    wire N__45873;
    wire N__45870;
    wire N__45867;
    wire N__45864;
    wire N__45861;
    wire N__45856;
    wire N__45853;
    wire N__45848;
    wire N__45845;
    wire N__45842;
    wire N__45839;
    wire N__45836;
    wire N__45833;
    wire N__45830;
    wire N__45823;
    wire N__45820;
    wire N__45817;
    wire N__45814;
    wire N__45811;
    wire N__45808;
    wire N__45805;
    wire N__45802;
    wire N__45797;
    wire N__45794;
    wire N__45791;
    wire N__45788;
    wire N__45785;
    wire N__45782;
    wire N__45775;
    wire N__45770;
    wire N__45763;
    wire N__45754;
    wire N__45751;
    wire N__45750;
    wire N__45747;
    wire N__45744;
    wire N__45741;
    wire N__45738;
    wire N__45735;
    wire N__45732;
    wire N__45727;
    wire N__45724;
    wire N__45721;
    wire N__45718;
    wire N__45715;
    wire N__45712;
    wire N__45709;
    wire N__45706;
    wire N__45703;
    wire N__45702;
    wire N__45701;
    wire N__45700;
    wire N__45699;
    wire N__45698;
    wire N__45697;
    wire N__45696;
    wire N__45695;
    wire N__45694;
    wire N__45693;
    wire N__45692;
    wire N__45691;
    wire N__45690;
    wire N__45689;
    wire N__45688;
    wire N__45687;
    wire N__45686;
    wire N__45685;
    wire N__45684;
    wire N__45683;
    wire N__45682;
    wire N__45681;
    wire N__45680;
    wire N__45677;
    wire N__45676;
    wire N__45675;
    wire N__45674;
    wire N__45673;
    wire N__45670;
    wire N__45669;
    wire N__45668;
    wire N__45667;
    wire N__45664;
    wire N__45663;
    wire N__45662;
    wire N__45661;
    wire N__45660;
    wire N__45659;
    wire N__45658;
    wire N__45657;
    wire N__45656;
    wire N__45655;
    wire N__45654;
    wire N__45653;
    wire N__45652;
    wire N__45651;
    wire N__45650;
    wire N__45645;
    wire N__45638;
    wire N__45637;
    wire N__45636;
    wire N__45635;
    wire N__45634;
    wire N__45633;
    wire N__45632;
    wire N__45625;
    wire N__45620;
    wire N__45619;
    wire N__45618;
    wire N__45617;
    wire N__45616;
    wire N__45615;
    wire N__45610;
    wire N__45607;
    wire N__45604;
    wire N__45595;
    wire N__45588;
    wire N__45583;
    wire N__45576;
    wire N__45573;
    wire N__45566;
    wire N__45563;
    wire N__45560;
    wire N__45553;
    wire N__45552;
    wire N__45551;
    wire N__45550;
    wire N__45549;
    wire N__45546;
    wire N__45539;
    wire N__45532;
    wire N__45525;
    wire N__45520;
    wire N__45515;
    wire N__45514;
    wire N__45513;
    wire N__45512;
    wire N__45511;
    wire N__45510;
    wire N__45509;
    wire N__45508;
    wire N__45507;
    wire N__45506;
    wire N__45505;
    wire N__45496;
    wire N__45495;
    wire N__45494;
    wire N__45493;
    wire N__45492;
    wire N__45489;
    wire N__45486;
    wire N__45481;
    wire N__45474;
    wire N__45467;
    wire N__45466;
    wire N__45465;
    wire N__45464;
    wire N__45463;
    wire N__45462;
    wire N__45461;
    wire N__45458;
    wire N__45453;
    wire N__45440;
    wire N__45437;
    wire N__45434;
    wire N__45431;
    wire N__45430;
    wire N__45427;
    wire N__45426;
    wire N__45425;
    wire N__45424;
    wire N__45423;
    wire N__45422;
    wire N__45421;
    wire N__45420;
    wire N__45419;
    wire N__45418;
    wire N__45417;
    wire N__45408;
    wire N__45403;
    wire N__45394;
    wire N__45381;
    wire N__45378;
    wire N__45369;
    wire N__45360;
    wire N__45357;
    wire N__45350;
    wire N__45347;
    wire N__45344;
    wire N__45341;
    wire N__45340;
    wire N__45339;
    wire N__45338;
    wire N__45337;
    wire N__45334;
    wire N__45325;
    wire N__45318;
    wire N__45311;
    wire N__45302;
    wire N__45295;
    wire N__45294;
    wire N__45285;
    wire N__45280;
    wire N__45273;
    wire N__45268;
    wire N__45265;
    wire N__45262;
    wire N__45259;
    wire N__45254;
    wire N__45253;
    wire N__45250;
    wire N__45247;
    wire N__45244;
    wire N__45237;
    wire N__45234;
    wire N__45231;
    wire N__45228;
    wire N__45219;
    wire N__45214;
    wire N__45211;
    wire N__45210;
    wire N__45203;
    wire N__45198;
    wire N__45191;
    wire N__45188;
    wire N__45183;
    wire N__45182;
    wire N__45181;
    wire N__45178;
    wire N__45175;
    wire N__45172;
    wire N__45169;
    wire N__45166;
    wire N__45163;
    wire N__45160;
    wire N__45145;
    wire N__45142;
    wire N__45141;
    wire N__45138;
    wire N__45135;
    wire N__45134;
    wire N__45133;
    wire N__45130;
    wire N__45127;
    wire N__45124;
    wire N__45121;
    wire N__45118;
    wire N__45117;
    wire N__45114;
    wire N__45111;
    wire N__45108;
    wire N__45105;
    wire N__45102;
    wire N__45099;
    wire N__45096;
    wire N__45093;
    wire N__45088;
    wire N__45083;
    wire N__45080;
    wire N__45077;
    wire N__45074;
    wire N__45071;
    wire N__45068;
    wire N__45063;
    wire N__45060;
    wire N__45055;
    wire N__45052;
    wire N__45049;
    wire N__45048;
    wire N__45047;
    wire N__45046;
    wire N__45043;
    wire N__45040;
    wire N__45037;
    wire N__45034;
    wire N__45031;
    wire N__45030;
    wire N__45029;
    wire N__45026;
    wire N__45025;
    wire N__45020;
    wire N__45017;
    wire N__45014;
    wire N__45011;
    wire N__45008;
    wire N__45005;
    wire N__44996;
    wire N__44995;
    wire N__44990;
    wire N__44987;
    wire N__44984;
    wire N__44981;
    wire N__44976;
    wire N__44973;
    wire N__44970;
    wire N__44965;
    wire N__44962;
    wire N__44959;
    wire N__44956;
    wire N__44953;
    wire N__44950;
    wire N__44949;
    wire N__44946;
    wire N__44943;
    wire N__44938;
    wire N__44937;
    wire N__44936;
    wire N__44935;
    wire N__44932;
    wire N__44929;
    wire N__44928;
    wire N__44927;
    wire N__44924;
    wire N__44921;
    wire N__44918;
    wire N__44915;
    wire N__44912;
    wire N__44911;
    wire N__44908;
    wire N__44905;
    wire N__44904;
    wire N__44901;
    wire N__44894;
    wire N__44891;
    wire N__44886;
    wire N__44883;
    wire N__44880;
    wire N__44877;
    wire N__44874;
    wire N__44871;
    wire N__44868;
    wire N__44861;
    wire N__44856;
    wire N__44853;
    wire N__44850;
    wire N__44847;
    wire N__44842;
    wire N__44839;
    wire N__44838;
    wire N__44835;
    wire N__44832;
    wire N__44831;
    wire N__44826;
    wire N__44823;
    wire N__44820;
    wire N__44819;
    wire N__44818;
    wire N__44815;
    wire N__44812;
    wire N__44809;
    wire N__44806;
    wire N__44803;
    wire N__44798;
    wire N__44795;
    wire N__44792;
    wire N__44789;
    wire N__44786;
    wire N__44783;
    wire N__44780;
    wire N__44773;
    wire N__44770;
    wire N__44767;
    wire N__44764;
    wire N__44761;
    wire N__44758;
    wire N__44755;
    wire N__44752;
    wire N__44749;
    wire N__44746;
    wire N__44743;
    wire N__44740;
    wire N__44737;
    wire N__44734;
    wire N__44731;
    wire N__44730;
    wire N__44727;
    wire N__44724;
    wire N__44719;
    wire N__44716;
    wire N__44713;
    wire N__44710;
    wire N__44707;
    wire N__44704;
    wire N__44701;
    wire N__44698;
    wire N__44695;
    wire N__44692;
    wire N__44691;
    wire N__44688;
    wire N__44685;
    wire N__44682;
    wire N__44679;
    wire N__44674;
    wire N__44673;
    wire N__44670;
    wire N__44667;
    wire N__44664;
    wire N__44661;
    wire N__44658;
    wire N__44655;
    wire N__44650;
    wire N__44647;
    wire N__44644;
    wire N__44641;
    wire N__44638;
    wire N__44635;
    wire N__44632;
    wire N__44629;
    wire N__44626;
    wire N__44623;
    wire N__44620;
    wire N__44617;
    wire N__44614;
    wire N__44611;
    wire N__44608;
    wire N__44605;
    wire N__44602;
    wire N__44599;
    wire N__44596;
    wire N__44593;
    wire N__44590;
    wire N__44587;
    wire N__44584;
    wire N__44581;
    wire N__44578;
    wire N__44575;
    wire N__44572;
    wire N__44571;
    wire N__44570;
    wire N__44567;
    wire N__44562;
    wire N__44559;
    wire N__44556;
    wire N__44553;
    wire N__44550;
    wire N__44545;
    wire N__44542;
    wire N__44539;
    wire N__44536;
    wire N__44533;
    wire N__44530;
    wire N__44527;
    wire N__44524;
    wire N__44521;
    wire N__44518;
    wire N__44515;
    wire N__44512;
    wire N__44509;
    wire N__44506;
    wire N__44503;
    wire N__44500;
    wire N__44497;
    wire N__44494;
    wire N__44491;
    wire N__44488;
    wire N__44485;
    wire N__44482;
    wire N__44481;
    wire N__44480;
    wire N__44477;
    wire N__44472;
    wire N__44469;
    wire N__44466;
    wire N__44461;
    wire N__44458;
    wire N__44455;
    wire N__44452;
    wire N__44449;
    wire N__44446;
    wire N__44443;
    wire N__44440;
    wire N__44437;
    wire N__44434;
    wire N__44431;
    wire N__44428;
    wire N__44425;
    wire N__44422;
    wire N__44419;
    wire N__44416;
    wire N__44415;
    wire N__44412;
    wire N__44409;
    wire N__44406;
    wire N__44403;
    wire N__44400;
    wire N__44397;
    wire N__44394;
    wire N__44391;
    wire N__44386;
    wire N__44383;
    wire N__44380;
    wire N__44377;
    wire N__44374;
    wire N__44371;
    wire N__44368;
    wire N__44365;
    wire N__44362;
    wire N__44359;
    wire N__44356;
    wire N__44353;
    wire N__44350;
    wire N__44347;
    wire N__44344;
    wire N__44341;
    wire N__44338;
    wire N__44337;
    wire N__44334;
    wire N__44331;
    wire N__44328;
    wire N__44325;
    wire N__44322;
    wire N__44319;
    wire N__44316;
    wire N__44313;
    wire N__44308;
    wire N__44305;
    wire N__44302;
    wire N__44301;
    wire N__44298;
    wire N__44295;
    wire N__44292;
    wire N__44289;
    wire N__44284;
    wire N__44281;
    wire N__44280;
    wire N__44277;
    wire N__44274;
    wire N__44271;
    wire N__44268;
    wire N__44263;
    wire N__44260;
    wire N__44257;
    wire N__44254;
    wire N__44251;
    wire N__44248;
    wire N__44245;
    wire N__44242;
    wire N__44239;
    wire N__44238;
    wire N__44237;
    wire N__44234;
    wire N__44231;
    wire N__44230;
    wire N__44227;
    wire N__44222;
    wire N__44219;
    wire N__44218;
    wire N__44215;
    wire N__44210;
    wire N__44207;
    wire N__44206;
    wire N__44205;
    wire N__44202;
    wire N__44199;
    wire N__44196;
    wire N__44193;
    wire N__44190;
    wire N__44187;
    wire N__44182;
    wire N__44179;
    wire N__44176;
    wire N__44171;
    wire N__44166;
    wire N__44161;
    wire N__44158;
    wire N__44155;
    wire N__44152;
    wire N__44149;
    wire N__44146;
    wire N__44143;
    wire N__44140;
    wire N__44139;
    wire N__44136;
    wire N__44133;
    wire N__44128;
    wire N__44125;
    wire N__44122;
    wire N__44121;
    wire N__44118;
    wire N__44115;
    wire N__44112;
    wire N__44109;
    wire N__44106;
    wire N__44103;
    wire N__44100;
    wire N__44095;
    wire N__44094;
    wire N__44091;
    wire N__44088;
    wire N__44085;
    wire N__44082;
    wire N__44079;
    wire N__44076;
    wire N__44071;
    wire N__44068;
    wire N__44065;
    wire N__44062;
    wire N__44061;
    wire N__44060;
    wire N__44059;
    wire N__44058;
    wire N__44055;
    wire N__44052;
    wire N__44049;
    wire N__44046;
    wire N__44043;
    wire N__44036;
    wire N__44035;
    wire N__44032;
    wire N__44029;
    wire N__44028;
    wire N__44025;
    wire N__44022;
    wire N__44019;
    wire N__44016;
    wire N__44015;
    wire N__44012;
    wire N__44007;
    wire N__44006;
    wire N__44003;
    wire N__44000;
    wire N__43997;
    wire N__43994;
    wire N__43991;
    wire N__43988;
    wire N__43983;
    wire N__43980;
    wire N__43977;
    wire N__43972;
    wire N__43967;
    wire N__43964;
    wire N__43961;
    wire N__43954;
    wire N__43951;
    wire N__43948;
    wire N__43945;
    wire N__43944;
    wire N__43941;
    wire N__43938;
    wire N__43933;
    wire N__43930;
    wire N__43927;
    wire N__43924;
    wire N__43921;
    wire N__43918;
    wire N__43915;
    wire N__43912;
    wire N__43909;
    wire N__43906;
    wire N__43903;
    wire N__43900;
    wire N__43897;
    wire N__43894;
    wire N__43891;
    wire N__43888;
    wire N__43887;
    wire N__43884;
    wire N__43881;
    wire N__43878;
    wire N__43875;
    wire N__43872;
    wire N__43869;
    wire N__43866;
    wire N__43863;
    wire N__43860;
    wire N__43855;
    wire N__43854;
    wire N__43851;
    wire N__43848;
    wire N__43845;
    wire N__43842;
    wire N__43839;
    wire N__43836;
    wire N__43833;
    wire N__43830;
    wire N__43825;
    wire N__43822;
    wire N__43819;
    wire N__43818;
    wire N__43815;
    wire N__43812;
    wire N__43809;
    wire N__43806;
    wire N__43803;
    wire N__43798;
    wire N__43795;
    wire N__43792;
    wire N__43789;
    wire N__43786;
    wire N__43783;
    wire N__43780;
    wire N__43779;
    wire N__43776;
    wire N__43773;
    wire N__43768;
    wire N__43765;
    wire N__43762;
    wire N__43759;
    wire N__43756;
    wire N__43753;
    wire N__43752;
    wire N__43749;
    wire N__43746;
    wire N__43741;
    wire N__43738;
    wire N__43735;
    wire N__43732;
    wire N__43729;
    wire N__43726;
    wire N__43723;
    wire N__43720;
    wire N__43717;
    wire N__43714;
    wire N__43711;
    wire N__43708;
    wire N__43705;
    wire N__43702;
    wire N__43701;
    wire N__43700;
    wire N__43699;
    wire N__43696;
    wire N__43693;
    wire N__43690;
    wire N__43687;
    wire N__43682;
    wire N__43677;
    wire N__43676;
    wire N__43673;
    wire N__43672;
    wire N__43671;
    wire N__43668;
    wire N__43665;
    wire N__43662;
    wire N__43659;
    wire N__43656;
    wire N__43653;
    wire N__43650;
    wire N__43643;
    wire N__43640;
    wire N__43639;
    wire N__43634;
    wire N__43631;
    wire N__43628;
    wire N__43627;
    wire N__43624;
    wire N__43619;
    wire N__43616;
    wire N__43613;
    wire N__43610;
    wire N__43607;
    wire N__43604;
    wire N__43599;
    wire N__43594;
    wire N__43591;
    wire N__43588;
    wire N__43585;
    wire N__43584;
    wire N__43581;
    wire N__43578;
    wire N__43575;
    wire N__43572;
    wire N__43567;
    wire N__43564;
    wire N__43561;
    wire N__43560;
    wire N__43557;
    wire N__43554;
    wire N__43551;
    wire N__43548;
    wire N__43543;
    wire N__43540;
    wire N__43537;
    wire N__43536;
    wire N__43533;
    wire N__43530;
    wire N__43527;
    wire N__43524;
    wire N__43519;
    wire N__43516;
    wire N__43513;
    wire N__43510;
    wire N__43509;
    wire N__43506;
    wire N__43503;
    wire N__43500;
    wire N__43497;
    wire N__43494;
    wire N__43491;
    wire N__43486;
    wire N__43485;
    wire N__43482;
    wire N__43479;
    wire N__43476;
    wire N__43473;
    wire N__43468;
    wire N__43465;
    wire N__43462;
    wire N__43459;
    wire N__43456;
    wire N__43453;
    wire N__43450;
    wire N__43447;
    wire N__43444;
    wire N__43441;
    wire N__43438;
    wire N__43435;
    wire N__43432;
    wire N__43429;
    wire N__43426;
    wire N__43423;
    wire N__43420;
    wire N__43417;
    wire N__43414;
    wire N__43411;
    wire N__43408;
    wire N__43405;
    wire N__43402;
    wire N__43399;
    wire N__43396;
    wire N__43393;
    wire N__43390;
    wire N__43387;
    wire N__43384;
    wire N__43381;
    wire N__43380;
    wire N__43379;
    wire N__43376;
    wire N__43371;
    wire N__43368;
    wire N__43365;
    wire N__43362;
    wire N__43359;
    wire N__43356;
    wire N__43353;
    wire N__43350;
    wire N__43347;
    wire N__43342;
    wire N__43339;
    wire N__43336;
    wire N__43333;
    wire N__43330;
    wire N__43327;
    wire N__43324;
    wire N__43321;
    wire N__43318;
    wire N__43315;
    wire N__43312;
    wire N__43309;
    wire N__43306;
    wire N__43303;
    wire N__43300;
    wire N__43297;
    wire N__43294;
    wire N__43291;
    wire N__43290;
    wire N__43287;
    wire N__43286;
    wire N__43285;
    wire N__43282;
    wire N__43279;
    wire N__43276;
    wire N__43273;
    wire N__43270;
    wire N__43261;
    wire N__43258;
    wire N__43255;
    wire N__43252;
    wire N__43249;
    wire N__43246;
    wire N__43243;
    wire N__43240;
    wire N__43237;
    wire N__43236;
    wire N__43233;
    wire N__43232;
    wire N__43231;
    wire N__43230;
    wire N__43229;
    wire N__43226;
    wire N__43225;
    wire N__43220;
    wire N__43217;
    wire N__43212;
    wire N__43207;
    wire N__43206;
    wire N__43205;
    wire N__43204;
    wire N__43203;
    wire N__43202;
    wire N__43199;
    wire N__43194;
    wire N__43191;
    wire N__43186;
    wire N__43183;
    wire N__43178;
    wire N__43177;
    wire N__43176;
    wire N__43173;
    wire N__43170;
    wire N__43165;
    wire N__43160;
    wire N__43157;
    wire N__43154;
    wire N__43141;
    wire N__43140;
    wire N__43139;
    wire N__43138;
    wire N__43137;
    wire N__43136;
    wire N__43135;
    wire N__43134;
    wire N__43131;
    wire N__43126;
    wire N__43121;
    wire N__43118;
    wire N__43117;
    wire N__43114;
    wire N__43109;
    wire N__43108;
    wire N__43103;
    wire N__43098;
    wire N__43097;
    wire N__43096;
    wire N__43095;
    wire N__43094;
    wire N__43089;
    wire N__43086;
    wire N__43081;
    wire N__43078;
    wire N__43075;
    wire N__43074;
    wire N__43071;
    wire N__43068;
    wire N__43065;
    wire N__43056;
    wire N__43053;
    wire N__43050;
    wire N__43039;
    wire N__43038;
    wire N__43037;
    wire N__43036;
    wire N__43035;
    wire N__43034;
    wire N__43033;
    wire N__43032;
    wire N__43031;
    wire N__43030;
    wire N__43029;
    wire N__43028;
    wire N__43027;
    wire N__43026;
    wire N__43025;
    wire N__43024;
    wire N__43023;
    wire N__43022;
    wire N__43021;
    wire N__43020;
    wire N__43019;
    wire N__43018;
    wire N__43017;
    wire N__43016;
    wire N__43015;
    wire N__43014;
    wire N__43013;
    wire N__43012;
    wire N__43011;
    wire N__43010;
    wire N__43009;
    wire N__43008;
    wire N__43007;
    wire N__43006;
    wire N__42997;
    wire N__42988;
    wire N__42987;
    wire N__42986;
    wire N__42985;
    wire N__42984;
    wire N__42983;
    wire N__42982;
    wire N__42981;
    wire N__42980;
    wire N__42979;
    wire N__42978;
    wire N__42977;
    wire N__42976;
    wire N__42975;
    wire N__42974;
    wire N__42973;
    wire N__42972;
    wire N__42971;
    wire N__42970;
    wire N__42969;
    wire N__42968;
    wire N__42967;
    wire N__42966;
    wire N__42965;
    wire N__42964;
    wire N__42963;
    wire N__42962;
    wire N__42961;
    wire N__42960;
    wire N__42959;
    wire N__42958;
    wire N__42957;
    wire N__42956;
    wire N__42955;
    wire N__42954;
    wire N__42953;
    wire N__42952;
    wire N__42951;
    wire N__42950;
    wire N__42949;
    wire N__42948;
    wire N__42947;
    wire N__42946;
    wire N__42945;
    wire N__42944;
    wire N__42943;
    wire N__42942;
    wire N__42941;
    wire N__42940;
    wire N__42939;
    wire N__42938;
    wire N__42937;
    wire N__42936;
    wire N__42935;
    wire N__42934;
    wire N__42933;
    wire N__42932;
    wire N__42931;
    wire N__42930;
    wire N__42929;
    wire N__42928;
    wire N__42927;
    wire N__42926;
    wire N__42925;
    wire N__42918;
    wire N__42915;
    wire N__42910;
    wire N__42909;
    wire N__42908;
    wire N__42907;
    wire N__42906;
    wire N__42905;
    wire N__42904;
    wire N__42903;
    wire N__42902;
    wire N__42901;
    wire N__42900;
    wire N__42899;
    wire N__42898;
    wire N__42897;
    wire N__42896;
    wire N__42893;
    wire N__42876;
    wire N__42859;
    wire N__42856;
    wire N__42855;
    wire N__42854;
    wire N__42853;
    wire N__42852;
    wire N__42851;
    wire N__42850;
    wire N__42849;
    wire N__42848;
    wire N__42847;
    wire N__42846;
    wire N__42845;
    wire N__42844;
    wire N__42843;
    wire N__42842;
    wire N__42839;
    wire N__42836;
    wire N__42835;
    wire N__42834;
    wire N__42833;
    wire N__42832;
    wire N__42831;
    wire N__42830;
    wire N__42825;
    wire N__42818;
    wire N__42817;
    wire N__42816;
    wire N__42813;
    wire N__42812;
    wire N__42811;
    wire N__42810;
    wire N__42809;
    wire N__42808;
    wire N__42807;
    wire N__42790;
    wire N__42785;
    wire N__42784;
    wire N__42777;
    wire N__42768;
    wire N__42767;
    wire N__42764;
    wire N__42763;
    wire N__42762;
    wire N__42761;
    wire N__42760;
    wire N__42759;
    wire N__42758;
    wire N__42757;
    wire N__42756;
    wire N__42753;
    wire N__42750;
    wire N__42747;
    wire N__42746;
    wire N__42743;
    wire N__42742;
    wire N__42741;
    wire N__42740;
    wire N__42739;
    wire N__42738;
    wire N__42737;
    wire N__42736;
    wire N__42735;
    wire N__42734;
    wire N__42733;
    wire N__42732;
    wire N__42731;
    wire N__42730;
    wire N__42729;
    wire N__42728;
    wire N__42727;
    wire N__42726;
    wire N__42725;
    wire N__42724;
    wire N__42723;
    wire N__42722;
    wire N__42721;
    wire N__42720;
    wire N__42719;
    wire N__42716;
    wire N__42713;
    wire N__42712;
    wire N__42711;
    wire N__42710;
    wire N__42709;
    wire N__42708;
    wire N__42707;
    wire N__42706;
    wire N__42705;
    wire N__42704;
    wire N__42703;
    wire N__42694;
    wire N__42677;
    wire N__42664;
    wire N__42655;
    wire N__42644;
    wire N__42627;
    wire N__42620;
    wire N__42615;
    wire N__42610;
    wire N__42601;
    wire N__42592;
    wire N__42587;
    wire N__42586;
    wire N__42585;
    wire N__42584;
    wire N__42583;
    wire N__42582;
    wire N__42581;
    wire N__42580;
    wire N__42579;
    wire N__42570;
    wire N__42561;
    wire N__42544;
    wire N__42539;
    wire N__42530;
    wire N__42525;
    wire N__42520;
    wire N__42515;
    wire N__42510;
    wire N__42509;
    wire N__42508;
    wire N__42507;
    wire N__42506;
    wire N__42505;
    wire N__42504;
    wire N__42503;
    wire N__42502;
    wire N__42501;
    wire N__42500;
    wire N__42499;
    wire N__42498;
    wire N__42497;
    wire N__42496;
    wire N__42495;
    wire N__42494;
    wire N__42493;
    wire N__42492;
    wire N__42491;
    wire N__42490;
    wire N__42489;
    wire N__42488;
    wire N__42487;
    wire N__42486;
    wire N__42485;
    wire N__42484;
    wire N__42483;
    wire N__42482;
    wire N__42481;
    wire N__42480;
    wire N__42479;
    wire N__42478;
    wire N__42477;
    wire N__42474;
    wire N__42461;
    wire N__42456;
    wire N__42453;
    wire N__42448;
    wire N__42445;
    wire N__42440;
    wire N__42435;
    wire N__42424;
    wire N__42421;
    wire N__42414;
    wire N__42411;
    wire N__42400;
    wire N__42399;
    wire N__42398;
    wire N__42397;
    wire N__42396;
    wire N__42395;
    wire N__42394;
    wire N__42393;
    wire N__42392;
    wire N__42391;
    wire N__42390;
    wire N__42389;
    wire N__42388;
    wire N__42387;
    wire N__42386;
    wire N__42385;
    wire N__42384;
    wire N__42383;
    wire N__42382;
    wire N__42381;
    wire N__42380;
    wire N__42379;
    wire N__42378;
    wire N__42377;
    wire N__42376;
    wire N__42375;
    wire N__42374;
    wire N__42373;
    wire N__42372;
    wire N__42371;
    wire N__42370;
    wire N__42369;
    wire N__42368;
    wire N__42367;
    wire N__42366;
    wire N__42365;
    wire N__42364;
    wire N__42363;
    wire N__42362;
    wire N__42361;
    wire N__42360;
    wire N__42359;
    wire N__42358;
    wire N__42357;
    wire N__42356;
    wire N__42355;
    wire N__42354;
    wire N__42353;
    wire N__42352;
    wire N__42351;
    wire N__42350;
    wire N__42349;
    wire N__42348;
    wire N__42347;
    wire N__42346;
    wire N__42345;
    wire N__42334;
    wire N__42323;
    wire N__42314;
    wire N__42303;
    wire N__42300;
    wire N__42297;
    wire N__42292;
    wire N__42275;
    wire N__42272;
    wire N__42269;
    wire N__42260;
    wire N__42251;
    wire N__42246;
    wire N__42245;
    wire N__42244;
    wire N__42243;
    wire N__42242;
    wire N__42241;
    wire N__42240;
    wire N__42239;
    wire N__42238;
    wire N__42221;
    wire N__42216;
    wire N__42209;
    wire N__42200;
    wire N__42183;
    wire N__42174;
    wire N__42159;
    wire N__42142;
    wire N__42129;
    wire N__42120;
    wire N__42115;
    wire N__42112;
    wire N__42105;
    wire N__42098;
    wire N__42081;
    wire N__42064;
    wire N__42049;
    wire N__42032;
    wire N__42015;
    wire N__41998;
    wire N__41981;
    wire N__41976;
    wire N__41971;
    wire N__41964;
    wire N__41951;
    wire N__41934;
    wire N__41925;
    wire N__41922;
    wire N__41909;
    wire N__41902;
    wire N__41869;
    wire N__41866;
    wire N__41863;
    wire N__41860;
    wire N__41859;
    wire N__41856;
    wire N__41855;
    wire N__41854;
    wire N__41853;
    wire N__41850;
    wire N__41849;
    wire N__41846;
    wire N__41843;
    wire N__41840;
    wire N__41837;
    wire N__41834;
    wire N__41833;
    wire N__41830;
    wire N__41827;
    wire N__41822;
    wire N__41819;
    wire N__41818;
    wire N__41815;
    wire N__41812;
    wire N__41809;
    wire N__41802;
    wire N__41799;
    wire N__41798;
    wire N__41795;
    wire N__41792;
    wire N__41785;
    wire N__41782;
    wire N__41777;
    wire N__41774;
    wire N__41771;
    wire N__41764;
    wire N__41761;
    wire N__41758;
    wire N__41755;
    wire N__41752;
    wire N__41749;
    wire N__41746;
    wire N__41743;
    wire N__41740;
    wire N__41739;
    wire N__41738;
    wire N__41737;
    wire N__41734;
    wire N__41733;
    wire N__41732;
    wire N__41731;
    wire N__41730;
    wire N__41725;
    wire N__41722;
    wire N__41719;
    wire N__41714;
    wire N__41709;
    wire N__41704;
    wire N__41703;
    wire N__41702;
    wire N__41701;
    wire N__41696;
    wire N__41693;
    wire N__41690;
    wire N__41685;
    wire N__41684;
    wire N__41683;
    wire N__41682;
    wire N__41681;
    wire N__41678;
    wire N__41675;
    wire N__41672;
    wire N__41667;
    wire N__41662;
    wire N__41657;
    wire N__41644;
    wire N__41643;
    wire N__41642;
    wire N__41641;
    wire N__41638;
    wire N__41633;
    wire N__41630;
    wire N__41629;
    wire N__41628;
    wire N__41627;
    wire N__41626;
    wire N__41625;
    wire N__41618;
    wire N__41615;
    wire N__41612;
    wire N__41609;
    wire N__41606;
    wire N__41603;
    wire N__41602;
    wire N__41595;
    wire N__41590;
    wire N__41585;
    wire N__41584;
    wire N__41583;
    wire N__41582;
    wire N__41581;
    wire N__41578;
    wire N__41575;
    wire N__41572;
    wire N__41569;
    wire N__41566;
    wire N__41563;
    wire N__41560;
    wire N__41545;
    wire N__41542;
    wire N__41539;
    wire N__41536;
    wire N__41535;
    wire N__41534;
    wire N__41531;
    wire N__41528;
    wire N__41525;
    wire N__41522;
    wire N__41521;
    wire N__41520;
    wire N__41519;
    wire N__41518;
    wire N__41515;
    wire N__41514;
    wire N__41513;
    wire N__41512;
    wire N__41511;
    wire N__41510;
    wire N__41509;
    wire N__41506;
    wire N__41503;
    wire N__41500;
    wire N__41497;
    wire N__41492;
    wire N__41489;
    wire N__41486;
    wire N__41485;
    wire N__41484;
    wire N__41481;
    wire N__41476;
    wire N__41471;
    wire N__41462;
    wire N__41459;
    wire N__41454;
    wire N__41451;
    wire N__41448;
    wire N__41445;
    wire N__41442;
    wire N__41435;
    wire N__41432;
    wire N__41419;
    wire N__41418;
    wire N__41417;
    wire N__41414;
    wire N__41413;
    wire N__41412;
    wire N__41411;
    wire N__41410;
    wire N__41409;
    wire N__41406;
    wire N__41403;
    wire N__41402;
    wire N__41399;
    wire N__41396;
    wire N__41393;
    wire N__41390;
    wire N__41387;
    wire N__41384;
    wire N__41383;
    wire N__41382;
    wire N__41379;
    wire N__41376;
    wire N__41373;
    wire N__41372;
    wire N__41371;
    wire N__41362;
    wire N__41357;
    wire N__41354;
    wire N__41351;
    wire N__41350;
    wire N__41345;
    wire N__41342;
    wire N__41339;
    wire N__41336;
    wire N__41327;
    wire N__41324;
    wire N__41311;
    wire N__41308;
    wire N__41305;
    wire N__41302;
    wire N__41299;
    wire N__41298;
    wire N__41297;
    wire N__41296;
    wire N__41295;
    wire N__41292;
    wire N__41289;
    wire N__41288;
    wire N__41285;
    wire N__41282;
    wire N__41279;
    wire N__41276;
    wire N__41273;
    wire N__41270;
    wire N__41269;
    wire N__41268;
    wire N__41265;
    wire N__41262;
    wire N__41253;
    wire N__41250;
    wire N__41247;
    wire N__41246;
    wire N__41243;
    wire N__41238;
    wire N__41235;
    wire N__41232;
    wire N__41229;
    wire N__41226;
    wire N__41223;
    wire N__41220;
    wire N__41217;
    wire N__41214;
    wire N__41203;
    wire N__41200;
    wire N__41197;
    wire N__41194;
    wire N__41191;
    wire N__41188;
    wire N__41185;
    wire N__41182;
    wire N__41179;
    wire N__41176;
    wire N__41173;
    wire N__41170;
    wire N__41167;
    wire N__41164;
    wire N__41161;
    wire N__41160;
    wire N__41157;
    wire N__41154;
    wire N__41149;
    wire N__41146;
    wire N__41143;
    wire N__41140;
    wire N__41137;
    wire N__41134;
    wire N__41131;
    wire N__41128;
    wire N__41125;
    wire N__41122;
    wire N__41119;
    wire N__41116;
    wire N__41113;
    wire N__41110;
    wire N__41107;
    wire N__41104;
    wire N__41101;
    wire N__41098;
    wire N__41095;
    wire N__41092;
    wire N__41089;
    wire N__41086;
    wire N__41083;
    wire N__41080;
    wire N__41077;
    wire N__41074;
    wire N__41071;
    wire N__41068;
    wire N__41065;
    wire N__41062;
    wire N__41059;
    wire N__41056;
    wire N__41053;
    wire N__41050;
    wire N__41047;
    wire N__41044;
    wire N__41041;
    wire N__41038;
    wire N__41035;
    wire N__41034;
    wire N__41031;
    wire N__41028;
    wire N__41023;
    wire N__41020;
    wire N__41019;
    wire N__41018;
    wire N__41015;
    wire N__41012;
    wire N__41009;
    wire N__41006;
    wire N__41001;
    wire N__41000;
    wire N__40995;
    wire N__40994;
    wire N__40991;
    wire N__40988;
    wire N__40985;
    wire N__40982;
    wire N__40977;
    wire N__40974;
    wire N__40971;
    wire N__40968;
    wire N__40965;
    wire N__40960;
    wire N__40957;
    wire N__40954;
    wire N__40951;
    wire N__40948;
    wire N__40945;
    wire N__40942;
    wire N__40939;
    wire N__40936;
    wire N__40933;
    wire N__40930;
    wire N__40927;
    wire N__40924;
    wire N__40921;
    wire N__40918;
    wire N__40915;
    wire N__40912;
    wire N__40909;
    wire N__40906;
    wire N__40903;
    wire N__40900;
    wire N__40897;
    wire N__40894;
    wire N__40891;
    wire N__40888;
    wire N__40885;
    wire N__40882;
    wire N__40879;
    wire N__40876;
    wire N__40873;
    wire N__40872;
    wire N__40871;
    wire N__40868;
    wire N__40867;
    wire N__40864;
    wire N__40861;
    wire N__40858;
    wire N__40855;
    wire N__40854;
    wire N__40851;
    wire N__40848;
    wire N__40843;
    wire N__40840;
    wire N__40839;
    wire N__40834;
    wire N__40831;
    wire N__40828;
    wire N__40825;
    wire N__40822;
    wire N__40819;
    wire N__40816;
    wire N__40813;
    wire N__40812;
    wire N__40807;
    wire N__40802;
    wire N__40799;
    wire N__40792;
    wire N__40789;
    wire N__40786;
    wire N__40783;
    wire N__40780;
    wire N__40777;
    wire N__40774;
    wire N__40771;
    wire N__40768;
    wire N__40765;
    wire N__40762;
    wire N__40761;
    wire N__40758;
    wire N__40755;
    wire N__40750;
    wire N__40747;
    wire N__40746;
    wire N__40743;
    wire N__40740;
    wire N__40735;
    wire N__40732;
    wire N__40729;
    wire N__40726;
    wire N__40725;
    wire N__40722;
    wire N__40719;
    wire N__40716;
    wire N__40713;
    wire N__40708;
    wire N__40705;
    wire N__40702;
    wire N__40701;
    wire N__40698;
    wire N__40695;
    wire N__40692;
    wire N__40687;
    wire N__40684;
    wire N__40683;
    wire N__40682;
    wire N__40679;
    wire N__40674;
    wire N__40671;
    wire N__40668;
    wire N__40663;
    wire N__40660;
    wire N__40657;
    wire N__40654;
    wire N__40651;
    wire N__40648;
    wire N__40645;
    wire N__40642;
    wire N__40639;
    wire N__40636;
    wire N__40633;
    wire N__40630;
    wire N__40627;
    wire N__40624;
    wire N__40623;
    wire N__40620;
    wire N__40619;
    wire N__40616;
    wire N__40613;
    wire N__40610;
    wire N__40607;
    wire N__40604;
    wire N__40601;
    wire N__40598;
    wire N__40593;
    wire N__40588;
    wire N__40585;
    wire N__40582;
    wire N__40579;
    wire N__40578;
    wire N__40575;
    wire N__40572;
    wire N__40567;
    wire N__40564;
    wire N__40561;
    wire N__40558;
    wire N__40557;
    wire N__40554;
    wire N__40551;
    wire N__40548;
    wire N__40545;
    wire N__40542;
    wire N__40537;
    wire N__40534;
    wire N__40531;
    wire N__40528;
    wire N__40527;
    wire N__40526;
    wire N__40523;
    wire N__40520;
    wire N__40519;
    wire N__40516;
    wire N__40511;
    wire N__40508;
    wire N__40505;
    wire N__40504;
    wire N__40497;
    wire N__40494;
    wire N__40489;
    wire N__40488;
    wire N__40487;
    wire N__40484;
    wire N__40481;
    wire N__40478;
    wire N__40475;
    wire N__40472;
    wire N__40469;
    wire N__40466;
    wire N__40463;
    wire N__40460;
    wire N__40453;
    wire N__40450;
    wire N__40447;
    wire N__40444;
    wire N__40441;
    wire N__40438;
    wire N__40435;
    wire N__40434;
    wire N__40431;
    wire N__40428;
    wire N__40425;
    wire N__40422;
    wire N__40419;
    wire N__40416;
    wire N__40411;
    wire N__40408;
    wire N__40405;
    wire N__40402;
    wire N__40399;
    wire N__40398;
    wire N__40395;
    wire N__40392;
    wire N__40389;
    wire N__40384;
    wire N__40381;
    wire N__40378;
    wire N__40375;
    wire N__40372;
    wire N__40369;
    wire N__40366;
    wire N__40363;
    wire N__40362;
    wire N__40359;
    wire N__40356;
    wire N__40353;
    wire N__40348;
    wire N__40345;
    wire N__40342;
    wire N__40341;
    wire N__40338;
    wire N__40335;
    wire N__40332;
    wire N__40329;
    wire N__40326;
    wire N__40323;
    wire N__40318;
    wire N__40315;
    wire N__40312;
    wire N__40309;
    wire N__40306;
    wire N__40305;
    wire N__40302;
    wire N__40299;
    wire N__40296;
    wire N__40293;
    wire N__40288;
    wire N__40285;
    wire N__40282;
    wire N__40279;
    wire N__40276;
    wire N__40275;
    wire N__40272;
    wire N__40269;
    wire N__40264;
    wire N__40261;
    wire N__40260;
    wire N__40257;
    wire N__40254;
    wire N__40251;
    wire N__40248;
    wire N__40243;
    wire N__40240;
    wire N__40239;
    wire N__40236;
    wire N__40233;
    wire N__40230;
    wire N__40227;
    wire N__40224;
    wire N__40221;
    wire N__40218;
    wire N__40213;
    wire N__40210;
    wire N__40207;
    wire N__40204;
    wire N__40201;
    wire N__40198;
    wire N__40197;
    wire N__40194;
    wire N__40191;
    wire N__40186;
    wire N__40185;
    wire N__40182;
    wire N__40179;
    wire N__40174;
    wire N__40173;
    wire N__40172;
    wire N__40169;
    wire N__40168;
    wire N__40167;
    wire N__40166;
    wire N__40163;
    wire N__40160;
    wire N__40157;
    wire N__40154;
    wire N__40151;
    wire N__40148;
    wire N__40145;
    wire N__40142;
    wire N__40135;
    wire N__40132;
    wire N__40129;
    wire N__40128;
    wire N__40123;
    wire N__40122;
    wire N__40119;
    wire N__40116;
    wire N__40113;
    wire N__40110;
    wire N__40107;
    wire N__40100;
    wire N__40097;
    wire N__40094;
    wire N__40091;
    wire N__40088;
    wire N__40085;
    wire N__40082;
    wire N__40079;
    wire N__40076;
    wire N__40069;
    wire N__40066;
    wire N__40063;
    wire N__40060;
    wire N__40057;
    wire N__40056;
    wire N__40053;
    wire N__40050;
    wire N__40045;
    wire N__40042;
    wire N__40039;
    wire N__40036;
    wire N__40033;
    wire N__40030;
    wire N__40027;
    wire N__40024;
    wire N__40021;
    wire N__40018;
    wire N__40015;
    wire N__40012;
    wire N__40009;
    wire N__40006;
    wire N__40003;
    wire N__40000;
    wire N__39997;
    wire N__39994;
    wire N__39993;
    wire N__39990;
    wire N__39987;
    wire N__39984;
    wire N__39981;
    wire N__39976;
    wire N__39973;
    wire N__39970;
    wire N__39967;
    wire N__39964;
    wire N__39963;
    wire N__39960;
    wire N__39957;
    wire N__39952;
    wire N__39949;
    wire N__39948;
    wire N__39945;
    wire N__39942;
    wire N__39939;
    wire N__39936;
    wire N__39933;
    wire N__39928;
    wire N__39925;
    wire N__39922;
    wire N__39921;
    wire N__39920;
    wire N__39917;
    wire N__39914;
    wire N__39911;
    wire N__39908;
    wire N__39907;
    wire N__39904;
    wire N__39901;
    wire N__39898;
    wire N__39895;
    wire N__39892;
    wire N__39889;
    wire N__39884;
    wire N__39883;
    wire N__39880;
    wire N__39879;
    wire N__39878;
    wire N__39875;
    wire N__39872;
    wire N__39869;
    wire N__39866;
    wire N__39863;
    wire N__39860;
    wire N__39857;
    wire N__39852;
    wire N__39847;
    wire N__39844;
    wire N__39841;
    wire N__39838;
    wire N__39835;
    wire N__39832;
    wire N__39829;
    wire N__39826;
    wire N__39821;
    wire N__39818;
    wire N__39815;
    wire N__39812;
    wire N__39805;
    wire N__39802;
    wire N__39799;
    wire N__39796;
    wire N__39793;
    wire N__39790;
    wire N__39787;
    wire N__39784;
    wire N__39781;
    wire N__39778;
    wire N__39775;
    wire N__39772;
    wire N__39769;
    wire N__39766;
    wire N__39763;
    wire N__39760;
    wire N__39757;
    wire N__39754;
    wire N__39753;
    wire N__39750;
    wire N__39747;
    wire N__39742;
    wire N__39741;
    wire N__39740;
    wire N__39737;
    wire N__39736;
    wire N__39733;
    wire N__39730;
    wire N__39727;
    wire N__39724;
    wire N__39723;
    wire N__39720;
    wire N__39717;
    wire N__39714;
    wire N__39711;
    wire N__39708;
    wire N__39705;
    wire N__39702;
    wire N__39697;
    wire N__39694;
    wire N__39693;
    wire N__39690;
    wire N__39685;
    wire N__39682;
    wire N__39679;
    wire N__39676;
    wire N__39671;
    wire N__39668;
    wire N__39661;
    wire N__39658;
    wire N__39657;
    wire N__39654;
    wire N__39651;
    wire N__39650;
    wire N__39649;
    wire N__39644;
    wire N__39641;
    wire N__39640;
    wire N__39637;
    wire N__39632;
    wire N__39629;
    wire N__39628;
    wire N__39625;
    wire N__39624;
    wire N__39621;
    wire N__39618;
    wire N__39615;
    wire N__39614;
    wire N__39611;
    wire N__39608;
    wire N__39607;
    wire N__39604;
    wire N__39601;
    wire N__39598;
    wire N__39595;
    wire N__39592;
    wire N__39589;
    wire N__39586;
    wire N__39583;
    wire N__39576;
    wire N__39569;
    wire N__39566;
    wire N__39563;
    wire N__39560;
    wire N__39553;
    wire N__39552;
    wire N__39547;
    wire N__39544;
    wire N__39543;
    wire N__39542;
    wire N__39539;
    wire N__39536;
    wire N__39533;
    wire N__39532;
    wire N__39529;
    wire N__39526;
    wire N__39523;
    wire N__39520;
    wire N__39517;
    wire N__39512;
    wire N__39509;
    wire N__39506;
    wire N__39503;
    wire N__39500;
    wire N__39495;
    wire N__39492;
    wire N__39487;
    wire N__39484;
    wire N__39481;
    wire N__39480;
    wire N__39477;
    wire N__39476;
    wire N__39475;
    wire N__39472;
    wire N__39471;
    wire N__39468;
    wire N__39465;
    wire N__39462;
    wire N__39459;
    wire N__39456;
    wire N__39455;
    wire N__39450;
    wire N__39449;
    wire N__39446;
    wire N__39443;
    wire N__39440;
    wire N__39437;
    wire N__39434;
    wire N__39431;
    wire N__39430;
    wire N__39427;
    wire N__39422;
    wire N__39421;
    wire N__39418;
    wire N__39415;
    wire N__39412;
    wire N__39409;
    wire N__39406;
    wire N__39403;
    wire N__39400;
    wire N__39397;
    wire N__39390;
    wire N__39387;
    wire N__39382;
    wire N__39377;
    wire N__39372;
    wire N__39369;
    wire N__39366;
    wire N__39363;
    wire N__39358;
    wire N__39355;
    wire N__39354;
    wire N__39353;
    wire N__39352;
    wire N__39349;
    wire N__39346;
    wire N__39345;
    wire N__39342;
    wire N__39341;
    wire N__39338;
    wire N__39337;
    wire N__39334;
    wire N__39331;
    wire N__39328;
    wire N__39325;
    wire N__39322;
    wire N__39319;
    wire N__39316;
    wire N__39309;
    wire N__39308;
    wire N__39305;
    wire N__39302;
    wire N__39299;
    wire N__39296;
    wire N__39295;
    wire N__39292;
    wire N__39289;
    wire N__39286;
    wire N__39279;
    wire N__39276;
    wire N__39273;
    wire N__39270;
    wire N__39263;
    wire N__39258;
    wire N__39255;
    wire N__39252;
    wire N__39249;
    wire N__39246;
    wire N__39241;
    wire N__39238;
    wire N__39237;
    wire N__39234;
    wire N__39231;
    wire N__39228;
    wire N__39225;
    wire N__39222;
    wire N__39219;
    wire N__39216;
    wire N__39213;
    wire N__39208;
    wire N__39207;
    wire N__39206;
    wire N__39205;
    wire N__39202;
    wire N__39201;
    wire N__39198;
    wire N__39195;
    wire N__39192;
    wire N__39189;
    wire N__39188;
    wire N__39185;
    wire N__39180;
    wire N__39177;
    wire N__39174;
    wire N__39171;
    wire N__39168;
    wire N__39165;
    wire N__39162;
    wire N__39159;
    wire N__39156;
    wire N__39155;
    wire N__39154;
    wire N__39151;
    wire N__39148;
    wire N__39145;
    wire N__39140;
    wire N__39137;
    wire N__39134;
    wire N__39121;
    wire N__39120;
    wire N__39117;
    wire N__39114;
    wire N__39111;
    wire N__39106;
    wire N__39103;
    wire N__39100;
    wire N__39097;
    wire N__39094;
    wire N__39091;
    wire N__39088;
    wire N__39085;
    wire N__39082;
    wire N__39079;
    wire N__39076;
    wire N__39073;
    wire N__39070;
    wire N__39067;
    wire N__39064;
    wire N__39061;
    wire N__39058;
    wire N__39055;
    wire N__39052;
    wire N__39049;
    wire N__39046;
    wire N__39043;
    wire N__39040;
    wire N__39037;
    wire N__39034;
    wire N__39031;
    wire N__39028;
    wire N__39025;
    wire N__39022;
    wire N__39019;
    wire N__39016;
    wire N__39013;
    wire N__39010;
    wire N__39007;
    wire N__39004;
    wire N__39001;
    wire N__38998;
    wire N__38995;
    wire N__38992;
    wire N__38989;
    wire N__38986;
    wire N__38983;
    wire N__38980;
    wire N__38977;
    wire N__38974;
    wire N__38971;
    wire N__38968;
    wire N__38965;
    wire N__38962;
    wire N__38959;
    wire N__38956;
    wire N__38953;
    wire N__38950;
    wire N__38947;
    wire N__38944;
    wire N__38941;
    wire N__38938;
    wire N__38935;
    wire N__38932;
    wire N__38929;
    wire N__38928;
    wire N__38925;
    wire N__38922;
    wire N__38917;
    wire N__38914;
    wire N__38911;
    wire N__38908;
    wire N__38905;
    wire N__38902;
    wire N__38899;
    wire N__38896;
    wire N__38893;
    wire N__38890;
    wire N__38887;
    wire N__38884;
    wire N__38881;
    wire N__38878;
    wire N__38875;
    wire N__38872;
    wire N__38869;
    wire N__38866;
    wire N__38863;
    wire N__38860;
    wire N__38857;
    wire N__38856;
    wire N__38855;
    wire N__38852;
    wire N__38851;
    wire N__38850;
    wire N__38849;
    wire N__38846;
    wire N__38845;
    wire N__38842;
    wire N__38841;
    wire N__38840;
    wire N__38839;
    wire N__38834;
    wire N__38831;
    wire N__38830;
    wire N__38829;
    wire N__38826;
    wire N__38821;
    wire N__38816;
    wire N__38811;
    wire N__38808;
    wire N__38805;
    wire N__38804;
    wire N__38803;
    wire N__38802;
    wire N__38797;
    wire N__38792;
    wire N__38789;
    wire N__38786;
    wire N__38781;
    wire N__38778;
    wire N__38773;
    wire N__38768;
    wire N__38765;
    wire N__38760;
    wire N__38749;
    wire N__38746;
    wire N__38745;
    wire N__38744;
    wire N__38743;
    wire N__38742;
    wire N__38741;
    wire N__38740;
    wire N__38739;
    wire N__38736;
    wire N__38731;
    wire N__38728;
    wire N__38725;
    wire N__38722;
    wire N__38717;
    wire N__38716;
    wire N__38715;
    wire N__38710;
    wire N__38707;
    wire N__38702;
    wire N__38699;
    wire N__38694;
    wire N__38693;
    wire N__38692;
    wire N__38691;
    wire N__38690;
    wire N__38687;
    wire N__38682;
    wire N__38677;
    wire N__38674;
    wire N__38671;
    wire N__38668;
    wire N__38665;
    wire N__38650;
    wire N__38647;
    wire N__38644;
    wire N__38641;
    wire N__38638;
    wire N__38635;
    wire N__38632;
    wire N__38629;
    wire N__38628;
    wire N__38627;
    wire N__38626;
    wire N__38625;
    wire N__38624;
    wire N__38623;
    wire N__38620;
    wire N__38619;
    wire N__38618;
    wire N__38615;
    wire N__38610;
    wire N__38609;
    wire N__38606;
    wire N__38601;
    wire N__38598;
    wire N__38595;
    wire N__38592;
    wire N__38587;
    wire N__38586;
    wire N__38585;
    wire N__38584;
    wire N__38583;
    wire N__38580;
    wire N__38577;
    wire N__38574;
    wire N__38565;
    wire N__38560;
    wire N__38555;
    wire N__38552;
    wire N__38549;
    wire N__38544;
    wire N__38533;
    wire N__38532;
    wire N__38531;
    wire N__38530;
    wire N__38529;
    wire N__38528;
    wire N__38527;
    wire N__38526;
    wire N__38523;
    wire N__38520;
    wire N__38517;
    wire N__38514;
    wire N__38509;
    wire N__38508;
    wire N__38505;
    wire N__38502;
    wire N__38495;
    wire N__38492;
    wire N__38489;
    wire N__38486;
    wire N__38485;
    wire N__38484;
    wire N__38483;
    wire N__38478;
    wire N__38473;
    wire N__38468;
    wire N__38465;
    wire N__38462;
    wire N__38461;
    wire N__38460;
    wire N__38459;
    wire N__38456;
    wire N__38453;
    wire N__38448;
    wire N__38445;
    wire N__38440;
    wire N__38437;
    wire N__38434;
    wire N__38419;
    wire N__38416;
    wire N__38413;
    wire N__38410;
    wire N__38407;
    wire N__38404;
    wire N__38401;
    wire N__38398;
    wire N__38395;
    wire N__38392;
    wire N__38391;
    wire N__38390;
    wire N__38387;
    wire N__38382;
    wire N__38379;
    wire N__38376;
    wire N__38373;
    wire N__38370;
    wire N__38367;
    wire N__38364;
    wire N__38359;
    wire N__38356;
    wire N__38353;
    wire N__38350;
    wire N__38347;
    wire N__38344;
    wire N__38341;
    wire N__38340;
    wire N__38339;
    wire N__38336;
    wire N__38335;
    wire N__38330;
    wire N__38327;
    wire N__38326;
    wire N__38323;
    wire N__38320;
    wire N__38317;
    wire N__38314;
    wire N__38311;
    wire N__38308;
    wire N__38299;
    wire N__38296;
    wire N__38293;
    wire N__38290;
    wire N__38287;
    wire N__38284;
    wire N__38281;
    wire N__38278;
    wire N__38275;
    wire N__38272;
    wire N__38269;
    wire N__38266;
    wire N__38263;
    wire N__38260;
    wire N__38257;
    wire N__38254;
    wire N__38251;
    wire N__38248;
    wire N__38245;
    wire N__38242;
    wire N__38239;
    wire N__38236;
    wire N__38233;
    wire N__38230;
    wire N__38227;
    wire N__38224;
    wire N__38221;
    wire N__38218;
    wire N__38215;
    wire N__38212;
    wire N__38209;
    wire N__38206;
    wire N__38203;
    wire N__38200;
    wire N__38197;
    wire N__38194;
    wire N__38191;
    wire N__38188;
    wire N__38185;
    wire N__38184;
    wire N__38183;
    wire N__38182;
    wire N__38179;
    wire N__38176;
    wire N__38173;
    wire N__38170;
    wire N__38165;
    wire N__38162;
    wire N__38159;
    wire N__38156;
    wire N__38153;
    wire N__38150;
    wire N__38149;
    wire N__38146;
    wire N__38143;
    wire N__38140;
    wire N__38137;
    wire N__38134;
    wire N__38129;
    wire N__38126;
    wire N__38123;
    wire N__38118;
    wire N__38113;
    wire N__38110;
    wire N__38107;
    wire N__38104;
    wire N__38101;
    wire N__38098;
    wire N__38095;
    wire N__38092;
    wire N__38089;
    wire N__38086;
    wire N__38083;
    wire N__38080;
    wire N__38077;
    wire N__38076;
    wire N__38073;
    wire N__38070;
    wire N__38069;
    wire N__38066;
    wire N__38063;
    wire N__38060;
    wire N__38057;
    wire N__38056;
    wire N__38051;
    wire N__38048;
    wire N__38047;
    wire N__38044;
    wire N__38041;
    wire N__38038;
    wire N__38035;
    wire N__38032;
    wire N__38029;
    wire N__38024;
    wire N__38021;
    wire N__38018;
    wire N__38015;
    wire N__38008;
    wire N__38005;
    wire N__38002;
    wire N__37999;
    wire N__37996;
    wire N__37993;
    wire N__37990;
    wire N__37987;
    wire N__37984;
    wire N__37981;
    wire N__37978;
    wire N__37975;
    wire N__37972;
    wire N__37969;
    wire N__37966;
    wire N__37963;
    wire N__37960;
    wire N__37957;
    wire N__37954;
    wire N__37951;
    wire N__37948;
    wire N__37945;
    wire N__37942;
    wire N__37939;
    wire N__37936;
    wire N__37933;
    wire N__37930;
    wire N__37927;
    wire N__37924;
    wire N__37921;
    wire N__37918;
    wire N__37915;
    wire N__37912;
    wire N__37911;
    wire N__37908;
    wire N__37905;
    wire N__37902;
    wire N__37899;
    wire N__37894;
    wire N__37891;
    wire N__37888;
    wire N__37885;
    wire N__37882;
    wire N__37879;
    wire N__37876;
    wire N__37873;
    wire N__37870;
    wire N__37867;
    wire N__37864;
    wire N__37861;
    wire N__37858;
    wire N__37855;
    wire N__37854;
    wire N__37851;
    wire N__37848;
    wire N__37845;
    wire N__37842;
    wire N__37839;
    wire N__37836;
    wire N__37833;
    wire N__37828;
    wire N__37827;
    wire N__37824;
    wire N__37821;
    wire N__37818;
    wire N__37815;
    wire N__37812;
    wire N__37809;
    wire N__37804;
    wire N__37801;
    wire N__37800;
    wire N__37797;
    wire N__37794;
    wire N__37791;
    wire N__37788;
    wire N__37783;
    wire N__37780;
    wire N__37779;
    wire N__37776;
    wire N__37773;
    wire N__37770;
    wire N__37767;
    wire N__37762;
    wire N__37759;
    wire N__37756;
    wire N__37753;
    wire N__37750;
    wire N__37749;
    wire N__37746;
    wire N__37743;
    wire N__37740;
    wire N__37735;
    wire N__37732;
    wire N__37729;
    wire N__37726;
    wire N__37723;
    wire N__37720;
    wire N__37717;
    wire N__37716;
    wire N__37715;
    wire N__37714;
    wire N__37711;
    wire N__37708;
    wire N__37707;
    wire N__37704;
    wire N__37701;
    wire N__37696;
    wire N__37693;
    wire N__37688;
    wire N__37687;
    wire N__37684;
    wire N__37681;
    wire N__37678;
    wire N__37675;
    wire N__37674;
    wire N__37669;
    wire N__37666;
    wire N__37663;
    wire N__37660;
    wire N__37657;
    wire N__37650;
    wire N__37647;
    wire N__37644;
    wire N__37641;
    wire N__37638;
    wire N__37633;
    wire N__37630;
    wire N__37627;
    wire N__37624;
    wire N__37621;
    wire N__37620;
    wire N__37617;
    wire N__37614;
    wire N__37611;
    wire N__37608;
    wire N__37605;
    wire N__37602;
    wire N__37597;
    wire N__37594;
    wire N__37591;
    wire N__37588;
    wire N__37585;
    wire N__37582;
    wire N__37579;
    wire N__37578;
    wire N__37575;
    wire N__37572;
    wire N__37569;
    wire N__37564;
    wire N__37561;
    wire N__37558;
    wire N__37555;
    wire N__37552;
    wire N__37549;
    wire N__37546;
    wire N__37543;
    wire N__37542;
    wire N__37539;
    wire N__37536;
    wire N__37533;
    wire N__37528;
    wire N__37525;
    wire N__37524;
    wire N__37521;
    wire N__37518;
    wire N__37515;
    wire N__37512;
    wire N__37507;
    wire N__37504;
    wire N__37501;
    wire N__37500;
    wire N__37497;
    wire N__37494;
    wire N__37491;
    wire N__37486;
    wire N__37483;
    wire N__37480;
    wire N__37477;
    wire N__37474;
    wire N__37471;
    wire N__37468;
    wire N__37465;
    wire N__37464;
    wire N__37461;
    wire N__37458;
    wire N__37455;
    wire N__37452;
    wire N__37449;
    wire N__37444;
    wire N__37441;
    wire N__37440;
    wire N__37437;
    wire N__37434;
    wire N__37431;
    wire N__37426;
    wire N__37423;
    wire N__37420;
    wire N__37417;
    wire N__37414;
    wire N__37413;
    wire N__37410;
    wire N__37407;
    wire N__37404;
    wire N__37399;
    wire N__37398;
    wire N__37395;
    wire N__37392;
    wire N__37389;
    wire N__37386;
    wire N__37381;
    wire N__37378;
    wire N__37377;
    wire N__37374;
    wire N__37371;
    wire N__37370;
    wire N__37369;
    wire N__37368;
    wire N__37365;
    wire N__37364;
    wire N__37363;
    wire N__37360;
    wire N__37357;
    wire N__37354;
    wire N__37351;
    wire N__37348;
    wire N__37345;
    wire N__37342;
    wire N__37341;
    wire N__37338;
    wire N__37333;
    wire N__37330;
    wire N__37327;
    wire N__37322;
    wire N__37319;
    wire N__37318;
    wire N__37313;
    wire N__37310;
    wire N__37303;
    wire N__37300;
    wire N__37297;
    wire N__37292;
    wire N__37289;
    wire N__37284;
    wire N__37281;
    wire N__37278;
    wire N__37273;
    wire N__37270;
    wire N__37269;
    wire N__37266;
    wire N__37263;
    wire N__37260;
    wire N__37257;
    wire N__37254;
    wire N__37251;
    wire N__37246;
    wire N__37245;
    wire N__37242;
    wire N__37241;
    wire N__37238;
    wire N__37237;
    wire N__37234;
    wire N__37233;
    wire N__37230;
    wire N__37227;
    wire N__37226;
    wire N__37225;
    wire N__37222;
    wire N__37221;
    wire N__37218;
    wire N__37215;
    wire N__37212;
    wire N__37209;
    wire N__37206;
    wire N__37203;
    wire N__37200;
    wire N__37197;
    wire N__37194;
    wire N__37191;
    wire N__37190;
    wire N__37187;
    wire N__37182;
    wire N__37179;
    wire N__37176;
    wire N__37173;
    wire N__37168;
    wire N__37165;
    wire N__37162;
    wire N__37159;
    wire N__37152;
    wire N__37147;
    wire N__37144;
    wire N__37139;
    wire N__37136;
    wire N__37131;
    wire N__37128;
    wire N__37123;
    wire N__37120;
    wire N__37117;
    wire N__37114;
    wire N__37111;
    wire N__37108;
    wire N__37105;
    wire N__37102;
    wire N__37099;
    wire N__37096;
    wire N__37095;
    wire N__37092;
    wire N__37089;
    wire N__37086;
    wire N__37083;
    wire N__37080;
    wire N__37079;
    wire N__37076;
    wire N__37073;
    wire N__37070;
    wire N__37063;
    wire N__37060;
    wire N__37059;
    wire N__37056;
    wire N__37053;
    wire N__37050;
    wire N__37047;
    wire N__37042;
    wire N__37041;
    wire N__37038;
    wire N__37035;
    wire N__37032;
    wire N__37029;
    wire N__37026;
    wire N__37023;
    wire N__37018;
    wire N__37017;
    wire N__37014;
    wire N__37011;
    wire N__37008;
    wire N__37005;
    wire N__37002;
    wire N__36999;
    wire N__36994;
    wire N__36991;
    wire N__36990;
    wire N__36989;
    wire N__36986;
    wire N__36985;
    wire N__36982;
    wire N__36981;
    wire N__36978;
    wire N__36975;
    wire N__36972;
    wire N__36971;
    wire N__36968;
    wire N__36965;
    wire N__36962;
    wire N__36961;
    wire N__36958;
    wire N__36955;
    wire N__36952;
    wire N__36951;
    wire N__36948;
    wire N__36945;
    wire N__36942;
    wire N__36939;
    wire N__36938;
    wire N__36935;
    wire N__36930;
    wire N__36927;
    wire N__36922;
    wire N__36917;
    wire N__36914;
    wire N__36905;
    wire N__36900;
    wire N__36897;
    wire N__36894;
    wire N__36891;
    wire N__36888;
    wire N__36883;
    wire N__36880;
    wire N__36879;
    wire N__36876;
    wire N__36873;
    wire N__36870;
    wire N__36867;
    wire N__36864;
    wire N__36861;
    wire N__36856;
    wire N__36853;
    wire N__36852;
    wire N__36849;
    wire N__36846;
    wire N__36843;
    wire N__36840;
    wire N__36837;
    wire N__36834;
    wire N__36829;
    wire N__36826;
    wire N__36823;
    wire N__36822;
    wire N__36819;
    wire N__36816;
    wire N__36811;
    wire N__36808;
    wire N__36805;
    wire N__36802;
    wire N__36799;
    wire N__36798;
    wire N__36795;
    wire N__36792;
    wire N__36787;
    wire N__36784;
    wire N__36783;
    wire N__36782;
    wire N__36781;
    wire N__36780;
    wire N__36779;
    wire N__36778;
    wire N__36777;
    wire N__36776;
    wire N__36775;
    wire N__36774;
    wire N__36773;
    wire N__36772;
    wire N__36771;
    wire N__36768;
    wire N__36765;
    wire N__36760;
    wire N__36755;
    wire N__36752;
    wire N__36749;
    wire N__36746;
    wire N__36743;
    wire N__36742;
    wire N__36741;
    wire N__36740;
    wire N__36731;
    wire N__36730;
    wire N__36727;
    wire N__36720;
    wire N__36715;
    wire N__36710;
    wire N__36707;
    wire N__36702;
    wire N__36699;
    wire N__36698;
    wire N__36695;
    wire N__36694;
    wire N__36691;
    wire N__36688;
    wire N__36685;
    wire N__36678;
    wire N__36675;
    wire N__36672;
    wire N__36669;
    wire N__36668;
    wire N__36665;
    wire N__36664;
    wire N__36663;
    wire N__36662;
    wire N__36659;
    wire N__36656;
    wire N__36653;
    wire N__36650;
    wire N__36645;
    wire N__36642;
    wire N__36639;
    wire N__36630;
    wire N__36613;
    wire N__36610;
    wire N__36609;
    wire N__36606;
    wire N__36603;
    wire N__36600;
    wire N__36597;
    wire N__36594;
    wire N__36589;
    wire N__36586;
    wire N__36583;
    wire N__36580;
    wire N__36577;
    wire N__36574;
    wire N__36571;
    wire N__36570;
    wire N__36567;
    wire N__36564;
    wire N__36561;
    wire N__36558;
    wire N__36553;
    wire N__36552;
    wire N__36551;
    wire N__36550;
    wire N__36549;
    wire N__36544;
    wire N__36539;
    wire N__36538;
    wire N__36537;
    wire N__36536;
    wire N__36535;
    wire N__36534;
    wire N__36531;
    wire N__36530;
    wire N__36529;
    wire N__36526;
    wire N__36523;
    wire N__36520;
    wire N__36517;
    wire N__36512;
    wire N__36509;
    wire N__36504;
    wire N__36503;
    wire N__36500;
    wire N__36499;
    wire N__36498;
    wire N__36495;
    wire N__36488;
    wire N__36485;
    wire N__36482;
    wire N__36479;
    wire N__36474;
    wire N__36471;
    wire N__36468;
    wire N__36465;
    wire N__36460;
    wire N__36453;
    wire N__36448;
    wire N__36439;
    wire N__36438;
    wire N__36437;
    wire N__36436;
    wire N__36435;
    wire N__36432;
    wire N__36431;
    wire N__36428;
    wire N__36427;
    wire N__36426;
    wire N__36421;
    wire N__36418;
    wire N__36413;
    wire N__36412;
    wire N__36411;
    wire N__36410;
    wire N__36409;
    wire N__36404;
    wire N__36403;
    wire N__36402;
    wire N__36399;
    wire N__36396;
    wire N__36393;
    wire N__36390;
    wire N__36385;
    wire N__36380;
    wire N__36377;
    wire N__36374;
    wire N__36371;
    wire N__36366;
    wire N__36361;
    wire N__36354;
    wire N__36347;
    wire N__36344;
    wire N__36341;
    wire N__36338;
    wire N__36331;
    wire N__36328;
    wire N__36327;
    wire N__36326;
    wire N__36325;
    wire N__36324;
    wire N__36323;
    wire N__36322;
    wire N__36321;
    wire N__36318;
    wire N__36301;
    wire N__36298;
    wire N__36295;
    wire N__36292;
    wire N__36291;
    wire N__36290;
    wire N__36289;
    wire N__36288;
    wire N__36287;
    wire N__36286;
    wire N__36285;
    wire N__36284;
    wire N__36283;
    wire N__36282;
    wire N__36279;
    wire N__36276;
    wire N__36273;
    wire N__36258;
    wire N__36257;
    wire N__36256;
    wire N__36255;
    wire N__36254;
    wire N__36253;
    wire N__36252;
    wire N__36251;
    wire N__36248;
    wire N__36245;
    wire N__36242;
    wire N__36241;
    wire N__36238;
    wire N__36235;
    wire N__36232;
    wire N__36231;
    wire N__36230;
    wire N__36229;
    wire N__36228;
    wire N__36227;
    wire N__36218;
    wire N__36217;
    wire N__36216;
    wire N__36213;
    wire N__36210;
    wire N__36209;
    wire N__36208;
    wire N__36205;
    wire N__36202;
    wire N__36199;
    wire N__36196;
    wire N__36191;
    wire N__36188;
    wire N__36177;
    wire N__36174;
    wire N__36171;
    wire N__36170;
    wire N__36167;
    wire N__36164;
    wire N__36161;
    wire N__36158;
    wire N__36155;
    wire N__36152;
    wire N__36145;
    wire N__36138;
    wire N__36133;
    wire N__36128;
    wire N__36125;
    wire N__36120;
    wire N__36103;
    wire N__36100;
    wire N__36097;
    wire N__36094;
    wire N__36091;
    wire N__36090;
    wire N__36087;
    wire N__36084;
    wire N__36081;
    wire N__36078;
    wire N__36075;
    wire N__36072;
    wire N__36067;
    wire N__36064;
    wire N__36063;
    wire N__36060;
    wire N__36057;
    wire N__36054;
    wire N__36051;
    wire N__36048;
    wire N__36043;
    wire N__36042;
    wire N__36039;
    wire N__36036;
    wire N__36033;
    wire N__36030;
    wire N__36027;
    wire N__36022;
    wire N__36019;
    wire N__36018;
    wire N__36017;
    wire N__36014;
    wire N__36011;
    wire N__36010;
    wire N__36007;
    wire N__36004;
    wire N__36001;
    wire N__35998;
    wire N__35995;
    wire N__35994;
    wire N__35991;
    wire N__35986;
    wire N__35985;
    wire N__35982;
    wire N__35979;
    wire N__35974;
    wire N__35971;
    wire N__35966;
    wire N__35965;
    wire N__35960;
    wire N__35957;
    wire N__35954;
    wire N__35953;
    wire N__35952;
    wire N__35949;
    wire N__35944;
    wire N__35941;
    wire N__35938;
    wire N__35935;
    wire N__35932;
    wire N__35927;
    wire N__35924;
    wire N__35921;
    wire N__35918;
    wire N__35911;
    wire N__35908;
    wire N__35905;
    wire N__35902;
    wire N__35901;
    wire N__35900;
    wire N__35899;
    wire N__35896;
    wire N__35893;
    wire N__35892;
    wire N__35891;
    wire N__35890;
    wire N__35887;
    wire N__35884;
    wire N__35879;
    wire N__35878;
    wire N__35875;
    wire N__35872;
    wire N__35869;
    wire N__35866;
    wire N__35863;
    wire N__35860;
    wire N__35857;
    wire N__35852;
    wire N__35849;
    wire N__35846;
    wire N__35843;
    wire N__35840;
    wire N__35837;
    wire N__35834;
    wire N__35827;
    wire N__35824;
    wire N__35815;
    wire N__35812;
    wire N__35809;
    wire N__35806;
    wire N__35803;
    wire N__35800;
    wire N__35797;
    wire N__35794;
    wire N__35791;
    wire N__35788;
    wire N__35785;
    wire N__35782;
    wire N__35779;
    wire N__35776;
    wire N__35773;
    wire N__35770;
    wire N__35767;
    wire N__35764;
    wire N__35761;
    wire N__35758;
    wire N__35755;
    wire N__35752;
    wire N__35749;
    wire N__35746;
    wire N__35743;
    wire N__35740;
    wire N__35737;
    wire N__35734;
    wire N__35731;
    wire N__35728;
    wire N__35725;
    wire N__35722;
    wire N__35719;
    wire N__35716;
    wire N__35713;
    wire N__35710;
    wire N__35707;
    wire N__35704;
    wire N__35701;
    wire N__35698;
    wire N__35695;
    wire N__35692;
    wire N__35689;
    wire N__35686;
    wire N__35683;
    wire N__35680;
    wire N__35677;
    wire N__35674;
    wire N__35671;
    wire N__35670;
    wire N__35669;
    wire N__35668;
    wire N__35667;
    wire N__35666;
    wire N__35665;
    wire N__35664;
    wire N__35661;
    wire N__35658;
    wire N__35655;
    wire N__35654;
    wire N__35653;
    wire N__35648;
    wire N__35645;
    wire N__35642;
    wire N__35639;
    wire N__35638;
    wire N__35637;
    wire N__35634;
    wire N__35629;
    wire N__35626;
    wire N__35623;
    wire N__35620;
    wire N__35617;
    wire N__35614;
    wire N__35609;
    wire N__35606;
    wire N__35605;
    wire N__35604;
    wire N__35603;
    wire N__35594;
    wire N__35591;
    wire N__35584;
    wire N__35579;
    wire N__35576;
    wire N__35573;
    wire N__35560;
    wire N__35559;
    wire N__35558;
    wire N__35557;
    wire N__35556;
    wire N__35553;
    wire N__35552;
    wire N__35551;
    wire N__35550;
    wire N__35549;
    wire N__35548;
    wire N__35547;
    wire N__35542;
    wire N__35537;
    wire N__35534;
    wire N__35531;
    wire N__35526;
    wire N__35521;
    wire N__35518;
    wire N__35517;
    wire N__35514;
    wire N__35511;
    wire N__35504;
    wire N__35501;
    wire N__35496;
    wire N__35495;
    wire N__35494;
    wire N__35491;
    wire N__35482;
    wire N__35477;
    wire N__35474;
    wire N__35471;
    wire N__35468;
    wire N__35461;
    wire N__35458;
    wire N__35455;
    wire N__35452;
    wire N__35449;
    wire N__35446;
    wire N__35443;
    wire N__35442;
    wire N__35441;
    wire N__35440;
    wire N__35439;
    wire N__35438;
    wire N__35437;
    wire N__35434;
    wire N__35431;
    wire N__35428;
    wire N__35427;
    wire N__35426;
    wire N__35421;
    wire N__35420;
    wire N__35419;
    wire N__35416;
    wire N__35413;
    wire N__35410;
    wire N__35407;
    wire N__35402;
    wire N__35399;
    wire N__35398;
    wire N__35395;
    wire N__35390;
    wire N__35379;
    wire N__35376;
    wire N__35375;
    wire N__35374;
    wire N__35373;
    wire N__35370;
    wire N__35365;
    wire N__35360;
    wire N__35357;
    wire N__35352;
    wire N__35341;
    wire N__35340;
    wire N__35339;
    wire N__35338;
    wire N__35337;
    wire N__35336;
    wire N__35335;
    wire N__35332;
    wire N__35329;
    wire N__35324;
    wire N__35323;
    wire N__35320;
    wire N__35317;
    wire N__35314;
    wire N__35313;
    wire N__35312;
    wire N__35311;
    wire N__35310;
    wire N__35307;
    wire N__35304;
    wire N__35301;
    wire N__35298;
    wire N__35297;
    wire N__35296;
    wire N__35291;
    wire N__35286;
    wire N__35283;
    wire N__35280;
    wire N__35277;
    wire N__35272;
    wire N__35269;
    wire N__35266;
    wire N__35263;
    wire N__35260;
    wire N__35249;
    wire N__35236;
    wire N__35233;
    wire N__35230;
    wire N__35227;
    wire N__35224;
    wire N__35221;
    wire N__35218;
    wire N__35215;
    wire N__35212;
    wire N__35209;
    wire N__35206;
    wire N__35203;
    wire N__35200;
    wire N__35197;
    wire N__35194;
    wire N__35191;
    wire N__35188;
    wire N__35185;
    wire N__35182;
    wire N__35179;
    wire N__35176;
    wire N__35173;
    wire N__35170;
    wire N__35167;
    wire N__35164;
    wire N__35161;
    wire N__35158;
    wire N__35157;
    wire N__35154;
    wire N__35151;
    wire N__35146;
    wire N__35143;
    wire N__35142;
    wire N__35139;
    wire N__35136;
    wire N__35133;
    wire N__35130;
    wire N__35127;
    wire N__35124;
    wire N__35119;
    wire N__35116;
    wire N__35113;
    wire N__35110;
    wire N__35107;
    wire N__35104;
    wire N__35101;
    wire N__35098;
    wire N__35095;
    wire N__35092;
    wire N__35089;
    wire N__35086;
    wire N__35083;
    wire N__35080;
    wire N__35077;
    wire N__35074;
    wire N__35071;
    wire N__35068;
    wire N__35065;
    wire N__35062;
    wire N__35059;
    wire N__35056;
    wire N__35053;
    wire N__35050;
    wire N__35047;
    wire N__35044;
    wire N__35043;
    wire N__35040;
    wire N__35037;
    wire N__35036;
    wire N__35033;
    wire N__35030;
    wire N__35027;
    wire N__35022;
    wire N__35021;
    wire N__35020;
    wire N__35017;
    wire N__35014;
    wire N__35011;
    wire N__35008;
    wire N__35005;
    wire N__35002;
    wire N__34999;
    wire N__34996;
    wire N__34989;
    wire N__34986;
    wire N__34981;
    wire N__34978;
    wire N__34975;
    wire N__34972;
    wire N__34971;
    wire N__34968;
    wire N__34965;
    wire N__34962;
    wire N__34959;
    wire N__34956;
    wire N__34951;
    wire N__34948;
    wire N__34945;
    wire N__34942;
    wire N__34939;
    wire N__34936;
    wire N__34933;
    wire N__34930;
    wire N__34927;
    wire N__34924;
    wire N__34921;
    wire N__34918;
    wire N__34915;
    wire N__34912;
    wire N__34911;
    wire N__34910;
    wire N__34905;
    wire N__34902;
    wire N__34899;
    wire N__34896;
    wire N__34893;
    wire N__34890;
    wire N__34887;
    wire N__34884;
    wire N__34879;
    wire N__34876;
    wire N__34873;
    wire N__34870;
    wire N__34867;
    wire N__34864;
    wire N__34861;
    wire N__34858;
    wire N__34855;
    wire N__34852;
    wire N__34849;
    wire N__34846;
    wire N__34843;
    wire N__34840;
    wire N__34837;
    wire N__34834;
    wire N__34833;
    wire N__34830;
    wire N__34827;
    wire N__34822;
    wire N__34819;
    wire N__34816;
    wire N__34815;
    wire N__34812;
    wire N__34809;
    wire N__34804;
    wire N__34803;
    wire N__34800;
    wire N__34797;
    wire N__34792;
    wire N__34789;
    wire N__34788;
    wire N__34787;
    wire N__34784;
    wire N__34781;
    wire N__34780;
    wire N__34777;
    wire N__34772;
    wire N__34769;
    wire N__34766;
    wire N__34761;
    wire N__34758;
    wire N__34755;
    wire N__34752;
    wire N__34749;
    wire N__34744;
    wire N__34741;
    wire N__34738;
    wire N__34735;
    wire N__34732;
    wire N__34729;
    wire N__34726;
    wire N__34723;
    wire N__34720;
    wire N__34717;
    wire N__34714;
    wire N__34711;
    wire N__34708;
    wire N__34705;
    wire N__34704;
    wire N__34703;
    wire N__34700;
    wire N__34699;
    wire N__34698;
    wire N__34695;
    wire N__34692;
    wire N__34689;
    wire N__34688;
    wire N__34687;
    wire N__34684;
    wire N__34681;
    wire N__34676;
    wire N__34673;
    wire N__34670;
    wire N__34667;
    wire N__34666;
    wire N__34663;
    wire N__34658;
    wire N__34653;
    wire N__34650;
    wire N__34647;
    wire N__34646;
    wire N__34643;
    wire N__34640;
    wire N__34637;
    wire N__34632;
    wire N__34629;
    wire N__34624;
    wire N__34621;
    wire N__34616;
    wire N__34613;
    wire N__34608;
    wire N__34605;
    wire N__34602;
    wire N__34597;
    wire N__34594;
    wire N__34591;
    wire N__34588;
    wire N__34587;
    wire N__34584;
    wire N__34581;
    wire N__34576;
    wire N__34573;
    wire N__34570;
    wire N__34569;
    wire N__34568;
    wire N__34565;
    wire N__34562;
    wire N__34559;
    wire N__34554;
    wire N__34551;
    wire N__34550;
    wire N__34549;
    wire N__34546;
    wire N__34543;
    wire N__34542;
    wire N__34541;
    wire N__34538;
    wire N__34535;
    wire N__34530;
    wire N__34527;
    wire N__34524;
    wire N__34523;
    wire N__34522;
    wire N__34519;
    wire N__34516;
    wire N__34513;
    wire N__34508;
    wire N__34505;
    wire N__34502;
    wire N__34497;
    wire N__34492;
    wire N__34489;
    wire N__34486;
    wire N__34483;
    wire N__34480;
    wire N__34477;
    wire N__34474;
    wire N__34471;
    wire N__34468;
    wire N__34463;
    wire N__34460;
    wire N__34457;
    wire N__34454;
    wire N__34447;
    wire N__34444;
    wire N__34441;
    wire N__34440;
    wire N__34437;
    wire N__34434;
    wire N__34431;
    wire N__34426;
    wire N__34423;
    wire N__34420;
    wire N__34417;
    wire N__34414;
    wire N__34411;
    wire N__34408;
    wire N__34405;
    wire N__34402;
    wire N__34399;
    wire N__34398;
    wire N__34395;
    wire N__34392;
    wire N__34389;
    wire N__34384;
    wire N__34381;
    wire N__34378;
    wire N__34375;
    wire N__34372;
    wire N__34369;
    wire N__34368;
    wire N__34365;
    wire N__34362;
    wire N__34359;
    wire N__34358;
    wire N__34355;
    wire N__34352;
    wire N__34349;
    wire N__34346;
    wire N__34341;
    wire N__34338;
    wire N__34337;
    wire N__34334;
    wire N__34333;
    wire N__34330;
    wire N__34327;
    wire N__34324;
    wire N__34321;
    wire N__34318;
    wire N__34315;
    wire N__34312;
    wire N__34309;
    wire N__34304;
    wire N__34299;
    wire N__34294;
    wire N__34291;
    wire N__34290;
    wire N__34287;
    wire N__34284;
    wire N__34281;
    wire N__34276;
    wire N__34273;
    wire N__34272;
    wire N__34271;
    wire N__34268;
    wire N__34265;
    wire N__34264;
    wire N__34261;
    wire N__34258;
    wire N__34255;
    wire N__34252;
    wire N__34249;
    wire N__34244;
    wire N__34243;
    wire N__34242;
    wire N__34241;
    wire N__34238;
    wire N__34237;
    wire N__34236;
    wire N__34233;
    wire N__34230;
    wire N__34227;
    wire N__34224;
    wire N__34221;
    wire N__34218;
    wire N__34215;
    wire N__34212;
    wire N__34209;
    wire N__34204;
    wire N__34201;
    wire N__34198;
    wire N__34195;
    wire N__34192;
    wire N__34189;
    wire N__34186;
    wire N__34183;
    wire N__34178;
    wire N__34175;
    wire N__34170;
    wire N__34165;
    wire N__34162;
    wire N__34157;
    wire N__34154;
    wire N__34151;
    wire N__34148;
    wire N__34141;
    wire N__34138;
    wire N__34137;
    wire N__34134;
    wire N__34131;
    wire N__34128;
    wire N__34125;
    wire N__34122;
    wire N__34119;
    wire N__34116;
    wire N__34111;
    wire N__34108;
    wire N__34105;
    wire N__34102;
    wire N__34099;
    wire N__34096;
    wire N__34093;
    wire N__34090;
    wire N__34087;
    wire N__34084;
    wire N__34081;
    wire N__34078;
    wire N__34075;
    wire N__34072;
    wire N__34069;
    wire N__34066;
    wire N__34063;
    wire N__34060;
    wire N__34057;
    wire N__34054;
    wire N__34051;
    wire N__34048;
    wire N__34045;
    wire N__34042;
    wire N__34039;
    wire N__34036;
    wire N__34033;
    wire N__34030;
    wire N__34027;
    wire N__34026;
    wire N__34025;
    wire N__34022;
    wire N__34017;
    wire N__34014;
    wire N__34011;
    wire N__34008;
    wire N__34005;
    wire N__34002;
    wire N__33999;
    wire N__33994;
    wire N__33991;
    wire N__33988;
    wire N__33985;
    wire N__33982;
    wire N__33981;
    wire N__33978;
    wire N__33975;
    wire N__33972;
    wire N__33969;
    wire N__33964;
    wire N__33961;
    wire N__33960;
    wire N__33957;
    wire N__33954;
    wire N__33951;
    wire N__33948;
    wire N__33945;
    wire N__33942;
    wire N__33937;
    wire N__33936;
    wire N__33933;
    wire N__33930;
    wire N__33927;
    wire N__33924;
    wire N__33921;
    wire N__33916;
    wire N__33913;
    wire N__33910;
    wire N__33907;
    wire N__33904;
    wire N__33901;
    wire N__33898;
    wire N__33895;
    wire N__33892;
    wire N__33889;
    wire N__33886;
    wire N__33883;
    wire N__33880;
    wire N__33877;
    wire N__33874;
    wire N__33871;
    wire N__33868;
    wire N__33865;
    wire N__33864;
    wire N__33863;
    wire N__33862;
    wire N__33861;
    wire N__33860;
    wire N__33859;
    wire N__33856;
    wire N__33855;
    wire N__33854;
    wire N__33853;
    wire N__33850;
    wire N__33847;
    wire N__33842;
    wire N__33837;
    wire N__33832;
    wire N__33831;
    wire N__33830;
    wire N__33825;
    wire N__33824;
    wire N__33821;
    wire N__33816;
    wire N__33813;
    wire N__33810;
    wire N__33805;
    wire N__33802;
    wire N__33801;
    wire N__33800;
    wire N__33797;
    wire N__33792;
    wire N__33787;
    wire N__33784;
    wire N__33781;
    wire N__33778;
    wire N__33775;
    wire N__33760;
    wire N__33759;
    wire N__33758;
    wire N__33757;
    wire N__33756;
    wire N__33755;
    wire N__33750;
    wire N__33745;
    wire N__33742;
    wire N__33741;
    wire N__33738;
    wire N__33737;
    wire N__33736;
    wire N__33735;
    wire N__33730;
    wire N__33729;
    wire N__33728;
    wire N__33723;
    wire N__33718;
    wire N__33713;
    wire N__33712;
    wire N__33709;
    wire N__33706;
    wire N__33703;
    wire N__33700;
    wire N__33697;
    wire N__33696;
    wire N__33693;
    wire N__33690;
    wire N__33687;
    wire N__33682;
    wire N__33677;
    wire N__33674;
    wire N__33669;
    wire N__33658;
    wire N__33655;
    wire N__33652;
    wire N__33649;
    wire N__33646;
    wire N__33643;
    wire N__33640;
    wire N__33637;
    wire N__33634;
    wire N__33631;
    wire N__33628;
    wire N__33625;
    wire N__33622;
    wire N__33619;
    wire N__33616;
    wire N__33613;
    wire N__33610;
    wire N__33607;
    wire N__33604;
    wire N__33601;
    wire N__33600;
    wire N__33599;
    wire N__33598;
    wire N__33595;
    wire N__33594;
    wire N__33593;
    wire N__33592;
    wire N__33591;
    wire N__33588;
    wire N__33585;
    wire N__33582;
    wire N__33579;
    wire N__33576;
    wire N__33575;
    wire N__33572;
    wire N__33571;
    wire N__33566;
    wire N__33563;
    wire N__33562;
    wire N__33561;
    wire N__33560;
    wire N__33555;
    wire N__33552;
    wire N__33549;
    wire N__33546;
    wire N__33543;
    wire N__33540;
    wire N__33537;
    wire N__33534;
    wire N__33531;
    wire N__33530;
    wire N__33525;
    wire N__33524;
    wire N__33521;
    wire N__33518;
    wire N__33515;
    wire N__33508;
    wire N__33501;
    wire N__33498;
    wire N__33495;
    wire N__33492;
    wire N__33489;
    wire N__33482;
    wire N__33477;
    wire N__33474;
    wire N__33463;
    wire N__33462;
    wire N__33461;
    wire N__33460;
    wire N__33459;
    wire N__33458;
    wire N__33457;
    wire N__33456;
    wire N__33455;
    wire N__33454;
    wire N__33451;
    wire N__33450;
    wire N__33447;
    wire N__33444;
    wire N__33441;
    wire N__33440;
    wire N__33437;
    wire N__33434;
    wire N__33431;
    wire N__33426;
    wire N__33425;
    wire N__33424;
    wire N__33421;
    wire N__33416;
    wire N__33413;
    wire N__33410;
    wire N__33407;
    wire N__33404;
    wire N__33399;
    wire N__33394;
    wire N__33391;
    wire N__33388;
    wire N__33385;
    wire N__33380;
    wire N__33377;
    wire N__33368;
    wire N__33363;
    wire N__33360;
    wire N__33355;
    wire N__33352;
    wire N__33343;
    wire N__33340;
    wire N__33337;
    wire N__33334;
    wire N__33331;
    wire N__33328;
    wire N__33325;
    wire N__33322;
    wire N__33319;
    wire N__33316;
    wire N__33313;
    wire N__33310;
    wire N__33307;
    wire N__33304;
    wire N__33301;
    wire N__33298;
    wire N__33295;
    wire N__33292;
    wire N__33289;
    wire N__33286;
    wire N__33283;
    wire N__33280;
    wire N__33277;
    wire N__33274;
    wire N__33271;
    wire N__33268;
    wire N__33265;
    wire N__33262;
    wire N__33261;
    wire N__33260;
    wire N__33257;
    wire N__33256;
    wire N__33253;
    wire N__33250;
    wire N__33247;
    wire N__33244;
    wire N__33241;
    wire N__33238;
    wire N__33235;
    wire N__33232;
    wire N__33229;
    wire N__33226;
    wire N__33217;
    wire N__33214;
    wire N__33211;
    wire N__33208;
    wire N__33205;
    wire N__33202;
    wire N__33199;
    wire N__33196;
    wire N__33193;
    wire N__33190;
    wire N__33187;
    wire N__33184;
    wire N__33181;
    wire N__33178;
    wire N__33175;
    wire N__33172;
    wire N__33169;
    wire N__33166;
    wire N__33163;
    wire N__33160;
    wire N__33157;
    wire N__33154;
    wire N__33151;
    wire N__33148;
    wire N__33145;
    wire N__33142;
    wire N__33139;
    wire N__33136;
    wire N__33133;
    wire N__33130;
    wire N__33127;
    wire N__33124;
    wire N__33123;
    wire N__33118;
    wire N__33115;
    wire N__33112;
    wire N__33111;
    wire N__33108;
    wire N__33105;
    wire N__33102;
    wire N__33099;
    wire N__33096;
    wire N__33093;
    wire N__33088;
    wire N__33085;
    wire N__33082;
    wire N__33079;
    wire N__33076;
    wire N__33075;
    wire N__33074;
    wire N__33073;
    wire N__33072;
    wire N__33069;
    wire N__33068;
    wire N__33063;
    wire N__33062;
    wire N__33061;
    wire N__33056;
    wire N__33055;
    wire N__33054;
    wire N__33049;
    wire N__33046;
    wire N__33041;
    wire N__33040;
    wire N__33039;
    wire N__33036;
    wire N__33031;
    wire N__33030;
    wire N__33029;
    wire N__33028;
    wire N__33025;
    wire N__33020;
    wire N__33015;
    wire N__33010;
    wire N__33005;
    wire N__33002;
    wire N__32999;
    wire N__32994;
    wire N__32989;
    wire N__32980;
    wire N__32979;
    wire N__32978;
    wire N__32977;
    wire N__32974;
    wire N__32973;
    wire N__32970;
    wire N__32969;
    wire N__32968;
    wire N__32967;
    wire N__32964;
    wire N__32963;
    wire N__32960;
    wire N__32959;
    wire N__32954;
    wire N__32949;
    wire N__32946;
    wire N__32945;
    wire N__32944;
    wire N__32941;
    wire N__32940;
    wire N__32935;
    wire N__32930;
    wire N__32927;
    wire N__32926;
    wire N__32923;
    wire N__32918;
    wire N__32915;
    wire N__32910;
    wire N__32903;
    wire N__32900;
    wire N__32895;
    wire N__32890;
    wire N__32885;
    wire N__32882;
    wire N__32879;
    wire N__32876;
    wire N__32873;
    wire N__32866;
    wire N__32865;
    wire N__32860;
    wire N__32857;
    wire N__32854;
    wire N__32851;
    wire N__32850;
    wire N__32847;
    wire N__32844;
    wire N__32839;
    wire N__32836;
    wire N__32833;
    wire N__32830;
    wire N__32827;
    wire N__32826;
    wire N__32825;
    wire N__32824;
    wire N__32823;
    wire N__32822;
    wire N__32821;
    wire N__32820;
    wire N__32819;
    wire N__32816;
    wire N__32813;
    wire N__32810;
    wire N__32807;
    wire N__32806;
    wire N__32805;
    wire N__32802;
    wire N__32799;
    wire N__32796;
    wire N__32795;
    wire N__32790;
    wire N__32789;
    wire N__32786;
    wire N__32779;
    wire N__32774;
    wire N__32767;
    wire N__32764;
    wire N__32763;
    wire N__32762;
    wire N__32759;
    wire N__32756;
    wire N__32749;
    wire N__32746;
    wire N__32741;
    wire N__32738;
    wire N__32733;
    wire N__32730;
    wire N__32725;
    wire N__32716;
    wire N__32715;
    wire N__32714;
    wire N__32713;
    wire N__32712;
    wire N__32711;
    wire N__32708;
    wire N__32707;
    wire N__32706;
    wire N__32701;
    wire N__32698;
    wire N__32693;
    wire N__32692;
    wire N__32687;
    wire N__32684;
    wire N__32683;
    wire N__32682;
    wire N__32681;
    wire N__32676;
    wire N__32673;
    wire N__32670;
    wire N__32667;
    wire N__32664;
    wire N__32661;
    wire N__32658;
    wire N__32655;
    wire N__32652;
    wire N__32647;
    wire N__32640;
    wire N__32635;
    wire N__32634;
    wire N__32633;
    wire N__32630;
    wire N__32623;
    wire N__32618;
    wire N__32611;
    wire N__32610;
    wire N__32609;
    wire N__32608;
    wire N__32607;
    wire N__32602;
    wire N__32601;
    wire N__32600;
    wire N__32599;
    wire N__32598;
    wire N__32597;
    wire N__32594;
    wire N__32591;
    wire N__32590;
    wire N__32589;
    wire N__32586;
    wire N__32585;
    wire N__32584;
    wire N__32581;
    wire N__32576;
    wire N__32571;
    wire N__32568;
    wire N__32563;
    wire N__32558;
    wire N__32553;
    wire N__32550;
    wire N__32549;
    wire N__32544;
    wire N__32541;
    wire N__32538;
    wire N__32535;
    wire N__32532;
    wire N__32527;
    wire N__32524;
    wire N__32521;
    wire N__32516;
    wire N__32511;
    wire N__32508;
    wire N__32497;
    wire N__32496;
    wire N__32493;
    wire N__32492;
    wire N__32491;
    wire N__32490;
    wire N__32489;
    wire N__32486;
    wire N__32485;
    wire N__32480;
    wire N__32479;
    wire N__32478;
    wire N__32477;
    wire N__32474;
    wire N__32473;
    wire N__32468;
    wire N__32463;
    wire N__32460;
    wire N__32457;
    wire N__32454;
    wire N__32451;
    wire N__32446;
    wire N__32445;
    wire N__32444;
    wire N__32443;
    wire N__32440;
    wire N__32437;
    wire N__32428;
    wire N__32425;
    wire N__32420;
    wire N__32417;
    wire N__32414;
    wire N__32409;
    wire N__32406;
    wire N__32401;
    wire N__32392;
    wire N__32391;
    wire N__32386;
    wire N__32383;
    wire N__32382;
    wire N__32379;
    wire N__32376;
    wire N__32371;
    wire N__32368;
    wire N__32365;
    wire N__32362;
    wire N__32359;
    wire N__32356;
    wire N__32355;
    wire N__32352;
    wire N__32349;
    wire N__32346;
    wire N__32343;
    wire N__32340;
    wire N__32337;
    wire N__32336;
    wire N__32333;
    wire N__32330;
    wire N__32327;
    wire N__32324;
    wire N__32319;
    wire N__32316;
    wire N__32313;
    wire N__32310;
    wire N__32307;
    wire N__32302;
    wire N__32299;
    wire N__32298;
    wire N__32297;
    wire N__32294;
    wire N__32291;
    wire N__32288;
    wire N__32285;
    wire N__32282;
    wire N__32279;
    wire N__32276;
    wire N__32273;
    wire N__32270;
    wire N__32267;
    wire N__32262;
    wire N__32257;
    wire N__32254;
    wire N__32251;
    wire N__32248;
    wire N__32245;
    wire N__32242;
    wire N__32239;
    wire N__32236;
    wire N__32233;
    wire N__32230;
    wire N__32227;
    wire N__32224;
    wire N__32221;
    wire N__32218;
    wire N__32215;
    wire N__32214;
    wire N__32213;
    wire N__32212;
    wire N__32211;
    wire N__32208;
    wire N__32207;
    wire N__32206;
    wire N__32201;
    wire N__32198;
    wire N__32195;
    wire N__32194;
    wire N__32189;
    wire N__32186;
    wire N__32185;
    wire N__32184;
    wire N__32179;
    wire N__32174;
    wire N__32173;
    wire N__32168;
    wire N__32165;
    wire N__32164;
    wire N__32163;
    wire N__32162;
    wire N__32159;
    wire N__32154;
    wire N__32151;
    wire N__32146;
    wire N__32141;
    wire N__32140;
    wire N__32137;
    wire N__32134;
    wire N__32131;
    wire N__32128;
    wire N__32123;
    wire N__32120;
    wire N__32107;
    wire N__32104;
    wire N__32103;
    wire N__32102;
    wire N__32097;
    wire N__32096;
    wire N__32093;
    wire N__32092;
    wire N__32089;
    wire N__32088;
    wire N__32087;
    wire N__32084;
    wire N__32083;
    wire N__32082;
    wire N__32081;
    wire N__32076;
    wire N__32075;
    wire N__32074;
    wire N__32071;
    wire N__32066;
    wire N__32063;
    wire N__32060;
    wire N__32059;
    wire N__32056;
    wire N__32053;
    wire N__32050;
    wire N__32049;
    wire N__32046;
    wire N__32043;
    wire N__32040;
    wire N__32035;
    wire N__32030;
    wire N__32023;
    wire N__32020;
    wire N__32017;
    wire N__32014;
    wire N__32011;
    wire N__32008;
    wire N__32003;
    wire N__31990;
    wire N__31987;
    wire N__31984;
    wire N__31981;
    wire N__31978;
    wire N__31975;
    wire N__31972;
    wire N__31969;
    wire N__31966;
    wire N__31963;
    wire N__31960;
    wire N__31957;
    wire N__31954;
    wire N__31951;
    wire N__31948;
    wire N__31945;
    wire N__31942;
    wire N__31939;
    wire N__31936;
    wire N__31933;
    wire N__31930;
    wire N__31927;
    wire N__31924;
    wire N__31921;
    wire N__31918;
    wire N__31915;
    wire N__31912;
    wire N__31909;
    wire N__31906;
    wire N__31903;
    wire N__31900;
    wire N__31899;
    wire N__31896;
    wire N__31893;
    wire N__31890;
    wire N__31887;
    wire N__31884;
    wire N__31881;
    wire N__31876;
    wire N__31873;
    wire N__31870;
    wire N__31867;
    wire N__31864;
    wire N__31863;
    wire N__31862;
    wire N__31859;
    wire N__31854;
    wire N__31849;
    wire N__31846;
    wire N__31843;
    wire N__31840;
    wire N__31837;
    wire N__31834;
    wire N__31831;
    wire N__31828;
    wire N__31825;
    wire N__31822;
    wire N__31819;
    wire N__31816;
    wire N__31813;
    wire N__31810;
    wire N__31807;
    wire N__31804;
    wire N__31801;
    wire N__31798;
    wire N__31795;
    wire N__31792;
    wire N__31789;
    wire N__31786;
    wire N__31783;
    wire N__31780;
    wire N__31777;
    wire N__31774;
    wire N__31771;
    wire N__31768;
    wire N__31765;
    wire N__31762;
    wire N__31761;
    wire N__31758;
    wire N__31755;
    wire N__31752;
    wire N__31749;
    wire N__31746;
    wire N__31743;
    wire N__31740;
    wire N__31735;
    wire N__31732;
    wire N__31731;
    wire N__31728;
    wire N__31725;
    wire N__31720;
    wire N__31717;
    wire N__31714;
    wire N__31711;
    wire N__31708;
    wire N__31705;
    wire N__31702;
    wire N__31701;
    wire N__31698;
    wire N__31695;
    wire N__31690;
    wire N__31687;
    wire N__31684;
    wire N__31683;
    wire N__31680;
    wire N__31677;
    wire N__31674;
    wire N__31671;
    wire N__31668;
    wire N__31663;
    wire N__31660;
    wire N__31657;
    wire N__31654;
    wire N__31651;
    wire N__31648;
    wire N__31647;
    wire N__31644;
    wire N__31641;
    wire N__31638;
    wire N__31635;
    wire N__31630;
    wire N__31627;
    wire N__31624;
    wire N__31621;
    wire N__31618;
    wire N__31615;
    wire N__31612;
    wire N__31609;
    wire N__31606;
    wire N__31603;
    wire N__31600;
    wire N__31597;
    wire N__31594;
    wire N__31591;
    wire N__31588;
    wire N__31585;
    wire N__31582;
    wire N__31579;
    wire N__31576;
    wire N__31573;
    wire N__31570;
    wire N__31567;
    wire N__31564;
    wire N__31561;
    wire N__31560;
    wire N__31557;
    wire N__31554;
    wire N__31551;
    wire N__31548;
    wire N__31545;
    wire N__31540;
    wire N__31537;
    wire N__31534;
    wire N__31533;
    wire N__31530;
    wire N__31527;
    wire N__31524;
    wire N__31521;
    wire N__31516;
    wire N__31513;
    wire N__31510;
    wire N__31507;
    wire N__31506;
    wire N__31503;
    wire N__31500;
    wire N__31497;
    wire N__31494;
    wire N__31491;
    wire N__31488;
    wire N__31483;
    wire N__31482;
    wire N__31479;
    wire N__31476;
    wire N__31473;
    wire N__31470;
    wire N__31467;
    wire N__31462;
    wire N__31459;
    wire N__31456;
    wire N__31453;
    wire N__31450;
    wire N__31447;
    wire N__31444;
    wire N__31443;
    wire N__31442;
    wire N__31439;
    wire N__31436;
    wire N__31433;
    wire N__31430;
    wire N__31429;
    wire N__31426;
    wire N__31425;
    wire N__31422;
    wire N__31419;
    wire N__31416;
    wire N__31413;
    wire N__31410;
    wire N__31407;
    wire N__31396;
    wire N__31395;
    wire N__31392;
    wire N__31389;
    wire N__31386;
    wire N__31383;
    wire N__31380;
    wire N__31375;
    wire N__31372;
    wire N__31369;
    wire N__31366;
    wire N__31365;
    wire N__31362;
    wire N__31359;
    wire N__31356;
    wire N__31353;
    wire N__31348;
    wire N__31345;
    wire N__31342;
    wire N__31339;
    wire N__31336;
    wire N__31333;
    wire N__31330;
    wire N__31327;
    wire N__31326;
    wire N__31323;
    wire N__31320;
    wire N__31317;
    wire N__31314;
    wire N__31311;
    wire N__31306;
    wire N__31303;
    wire N__31302;
    wire N__31299;
    wire N__31296;
    wire N__31293;
    wire N__31288;
    wire N__31287;
    wire N__31284;
    wire N__31281;
    wire N__31278;
    wire N__31275;
    wire N__31272;
    wire N__31269;
    wire N__31266;
    wire N__31261;
    wire N__31258;
    wire N__31255;
    wire N__31252;
    wire N__31249;
    wire N__31246;
    wire N__31243;
    wire N__31240;
    wire N__31237;
    wire N__31234;
    wire N__31231;
    wire N__31228;
    wire N__31225;
    wire N__31222;
    wire N__31219;
    wire N__31216;
    wire N__31213;
    wire N__31210;
    wire N__31207;
    wire N__31206;
    wire N__31203;
    wire N__31200;
    wire N__31197;
    wire N__31194;
    wire N__31191;
    wire N__31188;
    wire N__31185;
    wire N__31180;
    wire N__31177;
    wire N__31176;
    wire N__31173;
    wire N__31170;
    wire N__31167;
    wire N__31164;
    wire N__31161;
    wire N__31158;
    wire N__31153;
    wire N__31150;
    wire N__31147;
    wire N__31144;
    wire N__31141;
    wire N__31138;
    wire N__31135;
    wire N__31132;
    wire N__31129;
    wire N__31126;
    wire N__31123;
    wire N__31120;
    wire N__31117;
    wire N__31114;
    wire N__31111;
    wire N__31108;
    wire N__31105;
    wire N__31102;
    wire N__31099;
    wire N__31096;
    wire N__31093;
    wire N__31090;
    wire N__31087;
    wire N__31084;
    wire N__31081;
    wire N__31078;
    wire N__31075;
    wire N__31072;
    wire N__31069;
    wire N__31066;
    wire N__31063;
    wire N__31060;
    wire N__31057;
    wire N__31054;
    wire N__31051;
    wire N__31048;
    wire N__31045;
    wire N__31042;
    wire N__31039;
    wire N__31036;
    wire N__31033;
    wire N__31030;
    wire N__31027;
    wire N__31024;
    wire N__31021;
    wire N__31018;
    wire N__31017;
    wire N__31014;
    wire N__31011;
    wire N__31010;
    wire N__31009;
    wire N__31008;
    wire N__31007;
    wire N__31006;
    wire N__31005;
    wire N__31004;
    wire N__31003;
    wire N__31002;
    wire N__31001;
    wire N__30996;
    wire N__30993;
    wire N__30990;
    wire N__30985;
    wire N__30980;
    wire N__30979;
    wire N__30976;
    wire N__30973;
    wire N__30968;
    wire N__30959;
    wire N__30956;
    wire N__30955;
    wire N__30954;
    wire N__30951;
    wire N__30946;
    wire N__30943;
    wire N__30938;
    wire N__30933;
    wire N__30922;
    wire N__30921;
    wire N__30918;
    wire N__30915;
    wire N__30914;
    wire N__30913;
    wire N__30912;
    wire N__30911;
    wire N__30906;
    wire N__30901;
    wire N__30900;
    wire N__30899;
    wire N__30896;
    wire N__30893;
    wire N__30892;
    wire N__30891;
    wire N__30890;
    wire N__30889;
    wire N__30884;
    wire N__30879;
    wire N__30874;
    wire N__30869;
    wire N__30866;
    wire N__30863;
    wire N__30862;
    wire N__30861;
    wire N__30858;
    wire N__30855;
    wire N__30852;
    wire N__30849;
    wire N__30844;
    wire N__30841;
    wire N__30838;
    wire N__30823;
    wire N__30820;
    wire N__30817;
    wire N__30814;
    wire N__30813;
    wire N__30812;
    wire N__30809;
    wire N__30808;
    wire N__30807;
    wire N__30806;
    wire N__30803;
    wire N__30800;
    wire N__30797;
    wire N__30794;
    wire N__30791;
    wire N__30788;
    wire N__30787;
    wire N__30784;
    wire N__30781;
    wire N__30776;
    wire N__30773;
    wire N__30770;
    wire N__30767;
    wire N__30766;
    wire N__30761;
    wire N__30758;
    wire N__30755;
    wire N__30750;
    wire N__30747;
    wire N__30744;
    wire N__30739;
    wire N__30736;
    wire N__30733;
    wire N__30724;
    wire N__30721;
    wire N__30718;
    wire N__30715;
    wire N__30712;
    wire N__30709;
    wire N__30706;
    wire N__30703;
    wire N__30700;
    wire N__30697;
    wire N__30694;
    wire N__30691;
    wire N__30688;
    wire N__30685;
    wire N__30682;
    wire N__30679;
    wire N__30676;
    wire N__30673;
    wire N__30670;
    wire N__30667;
    wire N__30664;
    wire N__30661;
    wire N__30658;
    wire N__30655;
    wire N__30652;
    wire N__30649;
    wire N__30646;
    wire N__30643;
    wire N__30640;
    wire N__30637;
    wire N__30634;
    wire N__30631;
    wire N__30628;
    wire N__30625;
    wire N__30622;
    wire N__30619;
    wire N__30616;
    wire N__30613;
    wire N__30610;
    wire N__30607;
    wire N__30604;
    wire N__30601;
    wire N__30598;
    wire N__30595;
    wire N__30592;
    wire N__30589;
    wire N__30586;
    wire N__30583;
    wire N__30580;
    wire N__30577;
    wire N__30574;
    wire N__30571;
    wire N__30568;
    wire N__30565;
    wire N__30562;
    wire N__30559;
    wire N__30556;
    wire N__30553;
    wire N__30550;
    wire N__30547;
    wire N__30544;
    wire N__30541;
    wire N__30538;
    wire N__30535;
    wire N__30532;
    wire N__30529;
    wire N__30526;
    wire N__30523;
    wire N__30520;
    wire N__30517;
    wire N__30514;
    wire N__30511;
    wire N__30508;
    wire N__30505;
    wire N__30502;
    wire N__30499;
    wire N__30498;
    wire N__30495;
    wire N__30494;
    wire N__30493;
    wire N__30492;
    wire N__30491;
    wire N__30488;
    wire N__30487;
    wire N__30486;
    wire N__30481;
    wire N__30480;
    wire N__30479;
    wire N__30474;
    wire N__30473;
    wire N__30472;
    wire N__30469;
    wire N__30464;
    wire N__30461;
    wire N__30460;
    wire N__30457;
    wire N__30454;
    wire N__30451;
    wire N__30448;
    wire N__30445;
    wire N__30442;
    wire N__30439;
    wire N__30434;
    wire N__30433;
    wire N__30432;
    wire N__30429;
    wire N__30426;
    wire N__30423;
    wire N__30420;
    wire N__30417;
    wire N__30412;
    wire N__30407;
    wire N__30404;
    wire N__30401;
    wire N__30398;
    wire N__30393;
    wire N__30390;
    wire N__30381;
    wire N__30378;
    wire N__30367;
    wire N__30364;
    wire N__30363;
    wire N__30362;
    wire N__30361;
    wire N__30360;
    wire N__30359;
    wire N__30358;
    wire N__30353;
    wire N__30348;
    wire N__30343;
    wire N__30340;
    wire N__30339;
    wire N__30338;
    wire N__30337;
    wire N__30336;
    wire N__30335;
    wire N__30332;
    wire N__30327;
    wire N__30324;
    wire N__30321;
    wire N__30318;
    wire N__30315;
    wire N__30310;
    wire N__30309;
    wire N__30306;
    wire N__30299;
    wire N__30296;
    wire N__30293;
    wire N__30290;
    wire N__30287;
    wire N__30286;
    wire N__30283;
    wire N__30280;
    wire N__30275;
    wire N__30272;
    wire N__30269;
    wire N__30266;
    wire N__30263;
    wire N__30260;
    wire N__30253;
    wire N__30250;
    wire N__30241;
    wire N__30238;
    wire N__30235;
    wire N__30232;
    wire N__30229;
    wire N__30226;
    wire N__30223;
    wire N__30220;
    wire N__30217;
    wire N__30214;
    wire N__30211;
    wire N__30208;
    wire N__30205;
    wire N__30202;
    wire N__30199;
    wire N__30196;
    wire N__30193;
    wire N__30190;
    wire N__30187;
    wire N__30184;
    wire N__30181;
    wire N__30178;
    wire N__30175;
    wire N__30172;
    wire N__30169;
    wire N__30166;
    wire N__30163;
    wire N__30160;
    wire N__30157;
    wire N__30154;
    wire N__30151;
    wire N__30148;
    wire N__30145;
    wire N__30142;
    wire N__30139;
    wire N__30136;
    wire N__30133;
    wire N__30130;
    wire N__30127;
    wire N__30124;
    wire N__30121;
    wire N__30118;
    wire N__30115;
    wire N__30112;
    wire N__30109;
    wire N__30106;
    wire N__30103;
    wire N__30100;
    wire N__30097;
    wire N__30094;
    wire N__30091;
    wire N__30088;
    wire N__30085;
    wire N__30082;
    wire N__30079;
    wire N__30076;
    wire N__30073;
    wire N__30070;
    wire N__30067;
    wire N__30064;
    wire N__30061;
    wire N__30058;
    wire N__30055;
    wire N__30052;
    wire N__30049;
    wire N__30046;
    wire N__30043;
    wire N__30040;
    wire N__30037;
    wire N__30034;
    wire N__30031;
    wire N__30028;
    wire N__30025;
    wire N__30022;
    wire N__30019;
    wire N__30016;
    wire N__30013;
    wire N__30010;
    wire N__30007;
    wire N__30004;
    wire N__30001;
    wire N__29998;
    wire N__29995;
    wire N__29992;
    wire N__29989;
    wire N__29986;
    wire N__29983;
    wire N__29980;
    wire N__29977;
    wire N__29974;
    wire N__29971;
    wire N__29968;
    wire N__29965;
    wire N__29962;
    wire N__29959;
    wire N__29956;
    wire N__29953;
    wire N__29950;
    wire N__29947;
    wire N__29944;
    wire N__29941;
    wire N__29938;
    wire N__29935;
    wire N__29932;
    wire N__29929;
    wire N__29926;
    wire N__29923;
    wire N__29920;
    wire N__29917;
    wire N__29914;
    wire N__29911;
    wire N__29908;
    wire N__29905;
    wire N__29902;
    wire N__29899;
    wire N__29896;
    wire N__29893;
    wire N__29890;
    wire N__29887;
    wire N__29884;
    wire N__29881;
    wire N__29878;
    wire N__29875;
    wire N__29872;
    wire N__29869;
    wire N__29868;
    wire N__29865;
    wire N__29862;
    wire N__29859;
    wire N__29856;
    wire N__29853;
    wire N__29848;
    wire N__29845;
    wire N__29842;
    wire N__29839;
    wire N__29836;
    wire N__29833;
    wire N__29830;
    wire N__29827;
    wire N__29824;
    wire N__29821;
    wire N__29818;
    wire N__29815;
    wire N__29812;
    wire N__29811;
    wire N__29810;
    wire N__29807;
    wire N__29802;
    wire N__29799;
    wire N__29796;
    wire N__29793;
    wire N__29790;
    wire N__29785;
    wire N__29782;
    wire N__29779;
    wire N__29776;
    wire N__29773;
    wire N__29770;
    wire N__29767;
    wire N__29764;
    wire N__29761;
    wire N__29758;
    wire N__29755;
    wire N__29752;
    wire N__29749;
    wire N__29746;
    wire N__29743;
    wire N__29740;
    wire N__29737;
    wire N__29734;
    wire N__29731;
    wire N__29728;
    wire N__29725;
    wire N__29722;
    wire N__29719;
    wire N__29716;
    wire N__29713;
    wire N__29710;
    wire N__29707;
    wire N__29704;
    wire N__29701;
    wire N__29698;
    wire N__29695;
    wire N__29692;
    wire N__29689;
    wire N__29686;
    wire N__29683;
    wire N__29682;
    wire N__29679;
    wire N__29676;
    wire N__29671;
    wire N__29668;
    wire N__29665;
    wire N__29662;
    wire N__29659;
    wire N__29656;
    wire N__29653;
    wire N__29650;
    wire N__29647;
    wire N__29644;
    wire N__29641;
    wire N__29638;
    wire N__29635;
    wire N__29634;
    wire N__29631;
    wire N__29628;
    wire N__29623;
    wire N__29620;
    wire N__29619;
    wire N__29616;
    wire N__29613;
    wire N__29610;
    wire N__29607;
    wire N__29604;
    wire N__29599;
    wire N__29596;
    wire N__29595;
    wire N__29592;
    wire N__29589;
    wire N__29584;
    wire N__29581;
    wire N__29580;
    wire N__29577;
    wire N__29574;
    wire N__29571;
    wire N__29568;
    wire N__29563;
    wire N__29562;
    wire N__29559;
    wire N__29556;
    wire N__29553;
    wire N__29550;
    wire N__29545;
    wire N__29542;
    wire N__29539;
    wire N__29536;
    wire N__29533;
    wire N__29530;
    wire N__29527;
    wire N__29524;
    wire N__29521;
    wire N__29518;
    wire N__29515;
    wire N__29512;
    wire N__29509;
    wire N__29506;
    wire N__29503;
    wire N__29500;
    wire N__29497;
    wire N__29494;
    wire N__29491;
    wire N__29488;
    wire N__29485;
    wire N__29482;
    wire N__29479;
    wire N__29476;
    wire N__29473;
    wire N__29470;
    wire N__29467;
    wire N__29464;
    wire N__29463;
    wire N__29462;
    wire N__29461;
    wire N__29460;
    wire N__29459;
    wire N__29458;
    wire N__29457;
    wire N__29456;
    wire N__29453;
    wire N__29452;
    wire N__29451;
    wire N__29450;
    wire N__29449;
    wire N__29448;
    wire N__29447;
    wire N__29446;
    wire N__29445;
    wire N__29442;
    wire N__29441;
    wire N__29440;
    wire N__29439;
    wire N__29438;
    wire N__29437;
    wire N__29436;
    wire N__29429;
    wire N__29420;
    wire N__29415;
    wire N__29412;
    wire N__29411;
    wire N__29410;
    wire N__29407;
    wire N__29406;
    wire N__29403;
    wire N__29402;
    wire N__29399;
    wire N__29396;
    wire N__29393;
    wire N__29390;
    wire N__29389;
    wire N__29388;
    wire N__29381;
    wire N__29380;
    wire N__29377;
    wire N__29376;
    wire N__29373;
    wire N__29370;
    wire N__29367;
    wire N__29366;
    wire N__29365;
    wire N__29362;
    wire N__29359;
    wire N__29356;
    wire N__29353;
    wire N__29340;
    wire N__29329;
    wire N__29326;
    wire N__29323;
    wire N__29316;
    wire N__29307;
    wire N__29304;
    wire N__29281;
    wire N__29280;
    wire N__29279;
    wire N__29278;
    wire N__29277;
    wire N__29276;
    wire N__29271;
    wire N__29270;
    wire N__29269;
    wire N__29268;
    wire N__29267;
    wire N__29258;
    wire N__29257;
    wire N__29256;
    wire N__29255;
    wire N__29254;
    wire N__29253;
    wire N__29252;
    wire N__29249;
    wire N__29248;
    wire N__29247;
    wire N__29246;
    wire N__29245;
    wire N__29244;
    wire N__29243;
    wire N__29234;
    wire N__29231;
    wire N__29228;
    wire N__29225;
    wire N__29216;
    wire N__29215;
    wire N__29214;
    wire N__29213;
    wire N__29212;
    wire N__29211;
    wire N__29210;
    wire N__29209;
    wire N__29208;
    wire N__29207;
    wire N__29206;
    wire N__29203;
    wire N__29194;
    wire N__29189;
    wire N__29186;
    wire N__29181;
    wire N__29176;
    wire N__29167;
    wire N__29154;
    wire N__29137;
    wire N__29134;
    wire N__29131;
    wire N__29128;
    wire N__29125;
    wire N__29122;
    wire N__29119;
    wire N__29116;
    wire N__29113;
    wire N__29110;
    wire N__29107;
    wire N__29104;
    wire N__29101;
    wire N__29098;
    wire N__29097;
    wire N__29096;
    wire N__29095;
    wire N__29094;
    wire N__29093;
    wire N__29092;
    wire N__29091;
    wire N__29090;
    wire N__29085;
    wire N__29072;
    wire N__29071;
    wire N__29070;
    wire N__29069;
    wire N__29068;
    wire N__29067;
    wire N__29066;
    wire N__29063;
    wire N__29062;
    wire N__29061;
    wire N__29056;
    wire N__29051;
    wire N__29042;
    wire N__29041;
    wire N__29040;
    wire N__29039;
    wire N__29038;
    wire N__29037;
    wire N__29036;
    wire N__29035;
    wire N__29034;
    wire N__29033;
    wire N__29032;
    wire N__29031;
    wire N__29030;
    wire N__29029;
    wire N__29028;
    wire N__29027;
    wire N__29024;
    wire N__29019;
    wire N__29016;
    wire N__29011;
    wire N__29002;
    wire N__28993;
    wire N__28986;
    wire N__28977;
    wire N__28960;
    wire N__28957;
    wire N__28954;
    wire N__28951;
    wire N__28948;
    wire N__28945;
    wire N__28944;
    wire N__28943;
    wire N__28942;
    wire N__28939;
    wire N__28934;
    wire N__28931;
    wire N__28924;
    wire N__28921;
    wire N__28920;
    wire N__28917;
    wire N__28914;
    wire N__28913;
    wire N__28908;
    wire N__28905;
    wire N__28900;
    wire N__28897;
    wire N__28894;
    wire N__28891;
    wire N__28888;
    wire N__28885;
    wire N__28884;
    wire N__28881;
    wire N__28878;
    wire N__28873;
    wire N__28870;
    wire N__28867;
    wire N__28864;
    wire N__28861;
    wire N__28858;
    wire N__28857;
    wire N__28854;
    wire N__28851;
    wire N__28850;
    wire N__28847;
    wire N__28844;
    wire N__28841;
    wire N__28834;
    wire N__28831;
    wire N__28828;
    wire N__28825;
    wire N__28822;
    wire N__28821;
    wire N__28818;
    wire N__28815;
    wire N__28814;
    wire N__28811;
    wire N__28808;
    wire N__28805;
    wire N__28798;
    wire N__28795;
    wire N__28792;
    wire N__28789;
    wire N__28786;
    wire N__28783;
    wire N__28782;
    wire N__28779;
    wire N__28776;
    wire N__28771;
    wire N__28768;
    wire N__28765;
    wire N__28762;
    wire N__28759;
    wire N__28756;
    wire N__28753;
    wire N__28750;
    wire N__28747;
    wire N__28744;
    wire N__28743;
    wire N__28740;
    wire N__28737;
    wire N__28732;
    wire N__28731;
    wire N__28730;
    wire N__28729;
    wire N__28728;
    wire N__28727;
    wire N__28724;
    wire N__28721;
    wire N__28718;
    wire N__28715;
    wire N__28712;
    wire N__28709;
    wire N__28708;
    wire N__28707;
    wire N__28706;
    wire N__28705;
    wire N__28704;
    wire N__28703;
    wire N__28702;
    wire N__28701;
    wire N__28700;
    wire N__28699;
    wire N__28692;
    wire N__28685;
    wire N__28684;
    wire N__28683;
    wire N__28682;
    wire N__28679;
    wire N__28674;
    wire N__28671;
    wire N__28668;
    wire N__28665;
    wire N__28662;
    wire N__28659;
    wire N__28656;
    wire N__28653;
    wire N__28652;
    wire N__28651;
    wire N__28650;
    wire N__28649;
    wire N__28648;
    wire N__28647;
    wire N__28642;
    wire N__28641;
    wire N__28638;
    wire N__28637;
    wire N__28634;
    wire N__28633;
    wire N__28630;
    wire N__28627;
    wire N__28624;
    wire N__28617;
    wire N__28614;
    wire N__28607;
    wire N__28604;
    wire N__28601;
    wire N__28598;
    wire N__28595;
    wire N__28592;
    wire N__28589;
    wire N__28586;
    wire N__28585;
    wire N__28584;
    wire N__28583;
    wire N__28582;
    wire N__28581;
    wire N__28580;
    wire N__28579;
    wire N__28578;
    wire N__28577;
    wire N__28576;
    wire N__28575;
    wire N__28562;
    wire N__28557;
    wire N__28554;
    wire N__28549;
    wire N__28542;
    wire N__28535;
    wire N__28532;
    wire N__28527;
    wire N__28524;
    wire N__28523;
    wire N__28520;
    wire N__28519;
    wire N__28516;
    wire N__28515;
    wire N__28512;
    wire N__28511;
    wire N__28510;
    wire N__28509;
    wire N__28508;
    wire N__28507;
    wire N__28504;
    wire N__28501;
    wire N__28500;
    wire N__28497;
    wire N__28494;
    wire N__28491;
    wire N__28488;
    wire N__28477;
    wire N__28470;
    wire N__28457;
    wire N__28454;
    wire N__28451;
    wire N__28448;
    wire N__28447;
    wire N__28444;
    wire N__28441;
    wire N__28432;
    wire N__28427;
    wire N__28426;
    wire N__28425;
    wire N__28424;
    wire N__28423;
    wire N__28418;
    wire N__28415;
    wire N__28412;
    wire N__28407;
    wire N__28398;
    wire N__28393;
    wire N__28390;
    wire N__28383;
    wire N__28366;
    wire N__28363;
    wire N__28360;
    wire N__28357;
    wire N__28354;
    wire N__28351;
    wire N__28348;
    wire N__28345;
    wire N__28344;
    wire N__28341;
    wire N__28338;
    wire N__28333;
    wire N__28330;
    wire N__28327;
    wire N__28324;
    wire N__28321;
    wire N__28318;
    wire N__28315;
    wire N__28312;
    wire N__28309;
    wire N__28306;
    wire N__28303;
    wire N__28300;
    wire N__28297;
    wire N__28294;
    wire N__28293;
    wire N__28292;
    wire N__28291;
    wire N__28290;
    wire N__28289;
    wire N__28286;
    wire N__28283;
    wire N__28280;
    wire N__28277;
    wire N__28274;
    wire N__28271;
    wire N__28264;
    wire N__28261;
    wire N__28260;
    wire N__28257;
    wire N__28254;
    wire N__28251;
    wire N__28248;
    wire N__28245;
    wire N__28240;
    wire N__28233;
    wire N__28230;
    wire N__28227;
    wire N__28222;
    wire N__28219;
    wire N__28216;
    wire N__28213;
    wire N__28210;
    wire N__28207;
    wire N__28204;
    wire N__28201;
    wire N__28198;
    wire N__28195;
    wire N__28192;
    wire N__28189;
    wire N__28186;
    wire N__28183;
    wire N__28180;
    wire N__28177;
    wire N__28174;
    wire N__28171;
    wire N__28168;
    wire N__28165;
    wire N__28162;
    wire N__28159;
    wire N__28156;
    wire N__28153;
    wire N__28150;
    wire N__28147;
    wire N__28146;
    wire N__28145;
    wire N__28142;
    wire N__28139;
    wire N__28138;
    wire N__28137;
    wire N__28134;
    wire N__28129;
    wire N__28126;
    wire N__28123;
    wire N__28120;
    wire N__28115;
    wire N__28112;
    wire N__28107;
    wire N__28104;
    wire N__28101;
    wire N__28098;
    wire N__28093;
    wire N__28090;
    wire N__28087;
    wire N__28084;
    wire N__28081;
    wire N__28078;
    wire N__28075;
    wire N__28072;
    wire N__28069;
    wire N__28066;
    wire N__28063;
    wire N__28060;
    wire N__28057;
    wire N__28054;
    wire N__28051;
    wire N__28048;
    wire N__28045;
    wire N__28042;
    wire N__28039;
    wire N__28036;
    wire N__28033;
    wire N__28030;
    wire N__28027;
    wire N__28024;
    wire N__28021;
    wire N__28018;
    wire N__28015;
    wire N__28012;
    wire N__28009;
    wire N__28006;
    wire N__28003;
    wire N__28000;
    wire N__27997;
    wire N__27994;
    wire N__27991;
    wire N__27988;
    wire N__27985;
    wire N__27982;
    wire N__27979;
    wire N__27976;
    wire N__27973;
    wire N__27970;
    wire N__27967;
    wire N__27964;
    wire N__27961;
    wire N__27958;
    wire N__27955;
    wire N__27952;
    wire N__27949;
    wire N__27946;
    wire N__27943;
    wire N__27940;
    wire N__27937;
    wire N__27934;
    wire N__27931;
    wire N__27928;
    wire N__27925;
    wire N__27922;
    wire N__27919;
    wire N__27916;
    wire N__27913;
    wire N__27910;
    wire N__27907;
    wire N__27904;
    wire N__27901;
    wire N__27898;
    wire N__27895;
    wire N__27892;
    wire N__27889;
    wire N__27886;
    wire N__27883;
    wire N__27880;
    wire N__27877;
    wire N__27874;
    wire N__27871;
    wire N__27868;
    wire N__27865;
    wire N__27862;
    wire N__27859;
    wire N__27856;
    wire N__27855;
    wire N__27852;
    wire N__27849;
    wire N__27846;
    wire N__27843;
    wire N__27838;
    wire N__27835;
    wire N__27832;
    wire N__27831;
    wire N__27828;
    wire N__27825;
    wire N__27822;
    wire N__27819;
    wire N__27814;
    wire N__27811;
    wire N__27808;
    wire N__27807;
    wire N__27804;
    wire N__27801;
    wire N__27796;
    wire N__27793;
    wire N__27792;
    wire N__27789;
    wire N__27786;
    wire N__27783;
    wire N__27780;
    wire N__27775;
    wire N__27772;
    wire N__27771;
    wire N__27768;
    wire N__27765;
    wire N__27762;
    wire N__27759;
    wire N__27756;
    wire N__27753;
    wire N__27750;
    wire N__27745;
    wire N__27744;
    wire N__27743;
    wire N__27742;
    wire N__27739;
    wire N__27738;
    wire N__27733;
    wire N__27730;
    wire N__27727;
    wire N__27724;
    wire N__27719;
    wire N__27716;
    wire N__27713;
    wire N__27708;
    wire N__27705;
    wire N__27702;
    wire N__27697;
    wire N__27694;
    wire N__27691;
    wire N__27690;
    wire N__27687;
    wire N__27684;
    wire N__27683;
    wire N__27678;
    wire N__27675;
    wire N__27672;
    wire N__27669;
    wire N__27666;
    wire N__27663;
    wire N__27658;
    wire N__27655;
    wire N__27652;
    wire N__27651;
    wire N__27648;
    wire N__27645;
    wire N__27642;
    wire N__27639;
    wire N__27634;
    wire N__27631;
    wire N__27628;
    wire N__27625;
    wire N__27622;
    wire N__27619;
    wire N__27616;
    wire N__27613;
    wire N__27610;
    wire N__27607;
    wire N__27604;
    wire N__27601;
    wire N__27598;
    wire N__27595;
    wire N__27592;
    wire N__27589;
    wire N__27586;
    wire N__27583;
    wire N__27580;
    wire N__27577;
    wire N__27574;
    wire N__27571;
    wire N__27568;
    wire N__27565;
    wire N__27562;
    wire N__27559;
    wire N__27556;
    wire N__27553;
    wire N__27550;
    wire N__27547;
    wire N__27544;
    wire N__27541;
    wire N__27538;
    wire N__27535;
    wire N__27532;
    wire N__27529;
    wire N__27526;
    wire N__27523;
    wire N__27520;
    wire N__27517;
    wire N__27514;
    wire N__27511;
    wire N__27508;
    wire N__27505;
    wire N__27502;
    wire N__27499;
    wire N__27496;
    wire N__27493;
    wire N__27490;
    wire N__27487;
    wire N__27484;
    wire N__27481;
    wire N__27478;
    wire N__27475;
    wire N__27472;
    wire N__27469;
    wire N__27466;
    wire N__27463;
    wire N__27460;
    wire N__27457;
    wire N__27454;
    wire N__27451;
    wire N__27448;
    wire N__27445;
    wire N__27442;
    wire N__27439;
    wire N__27436;
    wire N__27433;
    wire N__27430;
    wire N__27427;
    wire N__27424;
    wire N__27423;
    wire N__27420;
    wire N__27417;
    wire N__27414;
    wire N__27411;
    wire N__27408;
    wire N__27405;
    wire N__27402;
    wire N__27399;
    wire N__27394;
    wire N__27391;
    wire N__27388;
    wire N__27385;
    wire N__27382;
    wire N__27379;
    wire N__27376;
    wire N__27373;
    wire N__27370;
    wire N__27367;
    wire N__27364;
    wire N__27363;
    wire N__27360;
    wire N__27357;
    wire N__27352;
    wire N__27349;
    wire N__27346;
    wire N__27343;
    wire N__27340;
    wire N__27337;
    wire N__27334;
    wire N__27331;
    wire N__27328;
    wire N__27325;
    wire N__27322;
    wire N__27319;
    wire N__27316;
    wire N__27313;
    wire N__27310;
    wire N__27307;
    wire N__27304;
    wire N__27301;
    wire N__27298;
    wire N__27295;
    wire N__27292;
    wire N__27289;
    wire N__27286;
    wire N__27283;
    wire N__27280;
    wire N__27277;
    wire N__27274;
    wire N__27271;
    wire N__27268;
    wire N__27265;
    wire N__27262;
    wire N__27259;
    wire N__27256;
    wire N__27253;
    wire N__27250;
    wire N__27247;
    wire N__27244;
    wire N__27241;
    wire N__27238;
    wire N__27235;
    wire N__27232;
    wire N__27229;
    wire N__27226;
    wire N__27223;
    wire N__27220;
    wire N__27217;
    wire N__27214;
    wire N__27211;
    wire N__27208;
    wire N__27205;
    wire N__27202;
    wire N__27199;
    wire N__27196;
    wire N__27193;
    wire N__27190;
    wire N__27187;
    wire N__27184;
    wire N__27181;
    wire N__27178;
    wire N__27175;
    wire N__27172;
    wire N__27169;
    wire N__27166;
    wire N__27163;
    wire N__27160;
    wire N__27157;
    wire N__27154;
    wire N__27151;
    wire N__27148;
    wire N__27145;
    wire N__27142;
    wire N__27139;
    wire N__27136;
    wire N__27133;
    wire N__27130;
    wire N__27127;
    wire N__27124;
    wire N__27121;
    wire N__27118;
    wire N__27115;
    wire N__27112;
    wire N__27109;
    wire N__27106;
    wire N__27103;
    wire N__27100;
    wire N__27097;
    wire N__27094;
    wire N__27091;
    wire N__27088;
    wire N__27085;
    wire N__27082;
    wire N__27079;
    wire N__27076;
    wire N__27073;
    wire N__27070;
    wire N__27067;
    wire N__27064;
    wire N__27061;
    wire N__27058;
    wire N__27055;
    wire N__27052;
    wire N__27049;
    wire N__27046;
    wire N__27043;
    wire N__27040;
    wire N__27037;
    wire N__27034;
    wire N__27031;
    wire N__27028;
    wire N__27025;
    wire N__27022;
    wire N__27019;
    wire N__27016;
    wire N__27013;
    wire N__27010;
    wire N__27007;
    wire N__27006;
    wire N__27003;
    wire N__27000;
    wire N__26995;
    wire N__26992;
    wire N__26991;
    wire N__26990;
    wire N__26987;
    wire N__26982;
    wire N__26977;
    wire N__26974;
    wire N__26971;
    wire N__26968;
    wire N__26965;
    wire N__26962;
    wire N__26959;
    wire N__26956;
    wire N__26953;
    wire N__26950;
    wire N__26947;
    wire N__26944;
    wire N__26941;
    wire N__26938;
    wire N__26935;
    wire N__26932;
    wire N__26929;
    wire N__26928;
    wire N__26927;
    wire N__26926;
    wire N__26925;
    wire N__26922;
    wire N__26921;
    wire N__26920;
    wire N__26919;
    wire N__26918;
    wire N__26917;
    wire N__26914;
    wire N__26911;
    wire N__26908;
    wire N__26905;
    wire N__26904;
    wire N__26903;
    wire N__26900;
    wire N__26897;
    wire N__26896;
    wire N__26895;
    wire N__26894;
    wire N__26893;
    wire N__26892;
    wire N__26891;
    wire N__26890;
    wire N__26889;
    wire N__26888;
    wire N__26879;
    wire N__26878;
    wire N__26877;
    wire N__26876;
    wire N__26867;
    wire N__26862;
    wire N__26857;
    wire N__26856;
    wire N__26855;
    wire N__26854;
    wire N__26853;
    wire N__26850;
    wire N__26841;
    wire N__26832;
    wire N__26829;
    wire N__26822;
    wire N__26819;
    wire N__26814;
    wire N__26805;
    wire N__26802;
    wire N__26795;
    wire N__26794;
    wire N__26793;
    wire N__26792;
    wire N__26791;
    wire N__26790;
    wire N__26785;
    wire N__26776;
    wire N__26769;
    wire N__26764;
    wire N__26755;
    wire N__26752;
    wire N__26749;
    wire N__26746;
    wire N__26743;
    wire N__26740;
    wire N__26737;
    wire N__26734;
    wire N__26731;
    wire N__26728;
    wire N__26725;
    wire N__26722;
    wire N__26719;
    wire N__26716;
    wire N__26713;
    wire N__26710;
    wire N__26707;
    wire N__26704;
    wire N__26701;
    wire N__26698;
    wire N__26695;
    wire N__26692;
    wire N__26689;
    wire N__26686;
    wire N__26683;
    wire N__26680;
    wire N__26679;
    wire N__26678;
    wire N__26677;
    wire N__26674;
    wire N__26671;
    wire N__26668;
    wire N__26665;
    wire N__26656;
    wire N__26653;
    wire N__26650;
    wire N__26647;
    wire N__26644;
    wire N__26641;
    wire N__26638;
    wire N__26635;
    wire N__26632;
    wire N__26629;
    wire N__26626;
    wire N__26623;
    wire N__26620;
    wire N__26617;
    wire N__26614;
    wire N__26611;
    wire N__26608;
    wire N__26605;
    wire N__26602;
    wire N__26599;
    wire N__26596;
    wire N__26593;
    wire N__26590;
    wire N__26587;
    wire N__26584;
    wire N__26581;
    wire N__26578;
    wire N__26575;
    wire N__26574;
    wire N__26571;
    wire N__26568;
    wire N__26563;
    wire N__26560;
    wire N__26557;
    wire N__26554;
    wire N__26551;
    wire N__26548;
    wire N__26545;
    wire N__26542;
    wire N__26539;
    wire N__26536;
    wire N__26533;
    wire N__26530;
    wire N__26527;
    wire N__26524;
    wire N__26521;
    wire N__26518;
    wire N__26515;
    wire N__26512;
    wire N__26509;
    wire N__26506;
    wire N__26503;
    wire N__26500;
    wire N__26497;
    wire N__26494;
    wire N__26493;
    wire N__26490;
    wire N__26487;
    wire N__26482;
    wire N__26479;
    wire N__26476;
    wire N__26473;
    wire N__26472;
    wire N__26471;
    wire N__26470;
    wire N__26469;
    wire N__26468;
    wire N__26455;
    wire N__26452;
    wire N__26451;
    wire N__26450;
    wire N__26447;
    wire N__26442;
    wire N__26437;
    wire N__26434;
    wire N__26431;
    wire N__26428;
    wire N__26427;
    wire N__26424;
    wire N__26421;
    wire N__26416;
    wire N__26415;
    wire N__26412;
    wire N__26409;
    wire N__26404;
    wire N__26403;
    wire N__26400;
    wire N__26399;
    wire N__26396;
    wire N__26391;
    wire N__26386;
    wire N__26383;
    wire N__26380;
    wire N__26377;
    wire N__26374;
    wire N__26371;
    wire N__26368;
    wire N__26365;
    wire N__26364;
    wire N__26361;
    wire N__26360;
    wire N__26357;
    wire N__26354;
    wire N__26351;
    wire N__26348;
    wire N__26345;
    wire N__26344;
    wire N__26341;
    wire N__26336;
    wire N__26333;
    wire N__26326;
    wire N__26323;
    wire N__26320;
    wire N__26317;
    wire N__26314;
    wire N__26311;
    wire N__26308;
    wire N__26307;
    wire N__26304;
    wire N__26301;
    wire N__26298;
    wire N__26297;
    wire N__26296;
    wire N__26295;
    wire N__26292;
    wire N__26289;
    wire N__26282;
    wire N__26275;
    wire N__26274;
    wire N__26273;
    wire N__26268;
    wire N__26265;
    wire N__26262;
    wire N__26257;
    wire N__26254;
    wire N__26253;
    wire N__26252;
    wire N__26249;
    wire N__26246;
    wire N__26243;
    wire N__26240;
    wire N__26233;
    wire N__26232;
    wire N__26227;
    wire N__26226;
    wire N__26223;
    wire N__26220;
    wire N__26219;
    wire N__26216;
    wire N__26211;
    wire N__26206;
    wire N__26203;
    wire N__26200;
    wire N__26197;
    wire N__26194;
    wire N__26191;
    wire N__26188;
    wire N__26185;
    wire N__26182;
    wire N__26179;
    wire N__26176;
    wire N__26173;
    wire N__26170;
    wire N__26167;
    wire N__26164;
    wire N__26161;
    wire N__26158;
    wire N__26155;
    wire N__26152;
    wire N__26149;
    wire N__26146;
    wire N__26143;
    wire N__26140;
    wire N__26137;
    wire N__26134;
    wire N__26131;
    wire N__26128;
    wire N__26125;
    wire N__26122;
    wire N__26119;
    wire N__26116;
    wire N__26113;
    wire N__26110;
    wire N__26107;
    wire N__26104;
    wire N__26101;
    wire N__26098;
    wire N__26095;
    wire N__26092;
    wire N__26089;
    wire N__26086;
    wire N__26083;
    wire N__26080;
    wire N__26079;
    wire N__26078;
    wire N__26075;
    wire N__26070;
    wire N__26069;
    wire N__26068;
    wire N__26065;
    wire N__26062;
    wire N__26057;
    wire N__26056;
    wire N__26053;
    wire N__26048;
    wire N__26045;
    wire N__26038;
    wire N__26035;
    wire N__26032;
    wire N__26029;
    wire N__26026;
    wire N__26023;
    wire N__26020;
    wire N__26017;
    wire N__26014;
    wire N__26011;
    wire N__26008;
    wire N__26005;
    wire N__26002;
    wire N__25999;
    wire N__25998;
    wire N__25995;
    wire N__25992;
    wire N__25989;
    wire N__25986;
    wire N__25981;
    wire N__25978;
    wire N__25975;
    wire N__25972;
    wire N__25969;
    wire N__25966;
    wire N__25963;
    wire N__25960;
    wire N__25957;
    wire N__25954;
    wire N__25951;
    wire N__25948;
    wire N__25945;
    wire N__25942;
    wire N__25939;
    wire N__25936;
    wire N__25933;
    wire N__25930;
    wire N__25927;
    wire N__25924;
    wire N__25921;
    wire N__25918;
    wire N__25915;
    wire N__25912;
    wire N__25909;
    wire N__25906;
    wire N__25903;
    wire N__25900;
    wire N__25897;
    wire N__25894;
    wire N__25891;
    wire N__25888;
    wire N__25885;
    wire N__25882;
    wire N__25881;
    wire N__25878;
    wire N__25875;
    wire N__25872;
    wire N__25869;
    wire N__25866;
    wire N__25861;
    wire N__25858;
    wire N__25855;
    wire N__25852;
    wire N__25849;
    wire N__25846;
    wire N__25845;
    wire N__25842;
    wire N__25839;
    wire N__25836;
    wire N__25833;
    wire N__25830;
    wire N__25827;
    wire N__25822;
    wire N__25819;
    wire N__25816;
    wire N__25813;
    wire N__25810;
    wire N__25807;
    wire N__25804;
    wire N__25803;
    wire N__25800;
    wire N__25797;
    wire N__25794;
    wire N__25791;
    wire N__25788;
    wire N__25783;
    wire N__25780;
    wire N__25777;
    wire N__25774;
    wire N__25771;
    wire N__25768;
    wire N__25765;
    wire N__25762;
    wire N__25761;
    wire N__25758;
    wire N__25755;
    wire N__25750;
    wire N__25747;
    wire N__25744;
    wire N__25741;
    wire N__25738;
    wire N__25735;
    wire N__25732;
    wire N__25729;
    wire N__25728;
    wire N__25725;
    wire N__25722;
    wire N__25719;
    wire N__25716;
    wire N__25713;
    wire N__25708;
    wire N__25705;
    wire N__25702;
    wire N__25699;
    wire N__25696;
    wire N__25693;
    wire N__25690;
    wire N__25687;
    wire N__25684;
    wire N__25681;
    wire N__25678;
    wire N__25675;
    wire N__25674;
    wire N__25671;
    wire N__25668;
    wire N__25665;
    wire N__25662;
    wire N__25659;
    wire N__25654;
    wire N__25651;
    wire N__25648;
    wire N__25647;
    wire N__25644;
    wire N__25641;
    wire N__25638;
    wire N__25635;
    wire N__25630;
    wire N__25629;
    wire N__25626;
    wire N__25625;
    wire N__25624;
    wire N__25623;
    wire N__25622;
    wire N__25621;
    wire N__25620;
    wire N__25619;
    wire N__25618;
    wire N__25615;
    wire N__25614;
    wire N__25613;
    wire N__25612;
    wire N__25611;
    wire N__25610;
    wire N__25609;
    wire N__25608;
    wire N__25607;
    wire N__25604;
    wire N__25597;
    wire N__25594;
    wire N__25589;
    wire N__25586;
    wire N__25585;
    wire N__25574;
    wire N__25573;
    wire N__25572;
    wire N__25571;
    wire N__25570;
    wire N__25569;
    wire N__25568;
    wire N__25567;
    wire N__25564;
    wire N__25563;
    wire N__25562;
    wire N__25561;
    wire N__25558;
    wire N__25555;
    wire N__25552;
    wire N__25551;
    wire N__25550;
    wire N__25549;
    wire N__25546;
    wire N__25543;
    wire N__25540;
    wire N__25537;
    wire N__25534;
    wire N__25531;
    wire N__25530;
    wire N__25529;
    wire N__25528;
    wire N__25527;
    wire N__25524;
    wire N__25521;
    wire N__25506;
    wire N__25489;
    wire N__25486;
    wire N__25483;
    wire N__25480;
    wire N__25477;
    wire N__25472;
    wire N__25467;
    wire N__25462;
    wire N__25455;
    wire N__25452;
    wire N__25445;
    wire N__25442;
    wire N__25439;
    wire N__25432;
    wire N__25423;
    wire N__25414;
    wire N__25411;
    wire N__25408;
    wire N__25405;
    wire N__25402;
    wire N__25399;
    wire N__25396;
    wire N__25395;
    wire N__25392;
    wire N__25391;
    wire N__25388;
    wire N__25385;
    wire N__25382;
    wire N__25381;
    wire N__25378;
    wire N__25373;
    wire N__25370;
    wire N__25367;
    wire N__25364;
    wire N__25361;
    wire N__25354;
    wire N__25351;
    wire N__25348;
    wire N__25345;
    wire N__25342;
    wire N__25339;
    wire N__25336;
    wire N__25333;
    wire N__25330;
    wire N__25327;
    wire N__25324;
    wire N__25321;
    wire N__25318;
    wire N__25317;
    wire N__25314;
    wire N__25311;
    wire N__25306;
    wire N__25303;
    wire N__25300;
    wire N__25297;
    wire N__25294;
    wire N__25291;
    wire N__25288;
    wire N__25285;
    wire N__25282;
    wire N__25279;
    wire N__25276;
    wire N__25273;
    wire N__25270;
    wire N__25267;
    wire N__25264;
    wire N__25261;
    wire N__25258;
    wire N__25255;
    wire N__25252;
    wire N__25249;
    wire N__25246;
    wire N__25243;
    wire N__25240;
    wire N__25237;
    wire N__25234;
    wire N__25231;
    wire N__25230;
    wire N__25225;
    wire N__25222;
    wire N__25221;
    wire N__25218;
    wire N__25215;
    wire N__25212;
    wire N__25209;
    wire N__25204;
    wire N__25201;
    wire N__25198;
    wire N__25195;
    wire N__25192;
    wire N__25189;
    wire N__25186;
    wire N__25183;
    wire N__25180;
    wire N__25177;
    wire N__25174;
    wire N__25171;
    wire N__25168;
    wire N__25165;
    wire N__25162;
    wire N__25159;
    wire N__25156;
    wire N__25153;
    wire N__25150;
    wire N__25147;
    wire N__25144;
    wire N__25141;
    wire N__25138;
    wire N__25135;
    wire N__25132;
    wire N__25129;
    wire N__25126;
    wire N__25123;
    wire N__25120;
    wire N__25117;
    wire N__25114;
    wire N__25111;
    wire N__25108;
    wire N__25105;
    wire N__25102;
    wire N__25099;
    wire N__25096;
    wire N__25093;
    wire N__25090;
    wire N__25087;
    wire N__25086;
    wire N__25085;
    wire N__25082;
    wire N__25079;
    wire N__25076;
    wire N__25073;
    wire N__25070;
    wire N__25067;
    wire N__25064;
    wire N__25061;
    wire N__25054;
    wire N__25051;
    wire N__25048;
    wire N__25047;
    wire N__25044;
    wire N__25041;
    wire N__25038;
    wire N__25035;
    wire N__25030;
    wire N__25027;
    wire N__25026;
    wire N__25023;
    wire N__25020;
    wire N__25015;
    wire N__25012;
    wire N__25009;
    wire N__25006;
    wire N__25003;
    wire N__25000;
    wire N__24997;
    wire N__24994;
    wire N__24991;
    wire N__24988;
    wire N__24987;
    wire N__24984;
    wire N__24981;
    wire N__24976;
    wire N__24973;
    wire N__24972;
    wire N__24971;
    wire N__24968;
    wire N__24965;
    wire N__24964;
    wire N__24961;
    wire N__24954;
    wire N__24953;
    wire N__24950;
    wire N__24947;
    wire N__24944;
    wire N__24939;
    wire N__24936;
    wire N__24931;
    wire N__24928;
    wire N__24925;
    wire N__24924;
    wire N__24921;
    wire N__24918;
    wire N__24913;
    wire N__24910;
    wire N__24907;
    wire N__24904;
    wire N__24901;
    wire N__24898;
    wire N__24895;
    wire N__24894;
    wire N__24891;
    wire N__24888;
    wire N__24885;
    wire N__24884;
    wire N__24883;
    wire N__24882;
    wire N__24879;
    wire N__24876;
    wire N__24873;
    wire N__24870;
    wire N__24867;
    wire N__24864;
    wire N__24859;
    wire N__24856;
    wire N__24853;
    wire N__24848;
    wire N__24845;
    wire N__24842;
    wire N__24835;
    wire N__24832;
    wire N__24829;
    wire N__24828;
    wire N__24827;
    wire N__24826;
    wire N__24825;
    wire N__24824;
    wire N__24823;
    wire N__24822;
    wire N__24819;
    wire N__24806;
    wire N__24803;
    wire N__24796;
    wire N__24793;
    wire N__24790;
    wire N__24787;
    wire N__24784;
    wire N__24783;
    wire N__24780;
    wire N__24777;
    wire N__24774;
    wire N__24771;
    wire N__24768;
    wire N__24763;
    wire N__24760;
    wire N__24759;
    wire N__24756;
    wire N__24753;
    wire N__24752;
    wire N__24749;
    wire N__24746;
    wire N__24743;
    wire N__24740;
    wire N__24735;
    wire N__24732;
    wire N__24729;
    wire N__24724;
    wire N__24723;
    wire N__24720;
    wire N__24717;
    wire N__24716;
    wire N__24715;
    wire N__24712;
    wire N__24709;
    wire N__24706;
    wire N__24703;
    wire N__24698;
    wire N__24691;
    wire N__24688;
    wire N__24685;
    wire N__24682;
    wire N__24679;
    wire N__24676;
    wire N__24673;
    wire N__24670;
    wire N__24669;
    wire N__24666;
    wire N__24663;
    wire N__24660;
    wire N__24657;
    wire N__24652;
    wire N__24649;
    wire N__24646;
    wire N__24643;
    wire N__24640;
    wire N__24637;
    wire N__24634;
    wire N__24631;
    wire N__24628;
    wire N__24625;
    wire N__24622;
    wire N__24619;
    wire N__24616;
    wire N__24613;
    wire N__24610;
    wire N__24607;
    wire N__24604;
    wire N__24603;
    wire N__24600;
    wire N__24599;
    wire N__24596;
    wire N__24593;
    wire N__24590;
    wire N__24589;
    wire N__24588;
    wire N__24587;
    wire N__24584;
    wire N__24579;
    wire N__24572;
    wire N__24565;
    wire N__24562;
    wire N__24561;
    wire N__24560;
    wire N__24557;
    wire N__24554;
    wire N__24551;
    wire N__24548;
    wire N__24547;
    wire N__24546;
    wire N__24543;
    wire N__24540;
    wire N__24537;
    wire N__24534;
    wire N__24531;
    wire N__24520;
    wire N__24517;
    wire N__24516;
    wire N__24515;
    wire N__24512;
    wire N__24511;
    wire N__24506;
    wire N__24505;
    wire N__24504;
    wire N__24503;
    wire N__24502;
    wire N__24499;
    wire N__24496;
    wire N__24493;
    wire N__24484;
    wire N__24475;
    wire N__24472;
    wire N__24469;
    wire N__24466;
    wire N__24463;
    wire N__24460;
    wire N__24457;
    wire N__24454;
    wire N__24451;
    wire N__24448;
    wire N__24447;
    wire N__24446;
    wire N__24445;
    wire N__24442;
    wire N__24439;
    wire N__24436;
    wire N__24433;
    wire N__24430;
    wire N__24427;
    wire N__24424;
    wire N__24421;
    wire N__24418;
    wire N__24413;
    wire N__24406;
    wire N__24405;
    wire N__24404;
    wire N__24403;
    wire N__24400;
    wire N__24397;
    wire N__24394;
    wire N__24391;
    wire N__24388;
    wire N__24385;
    wire N__24382;
    wire N__24379;
    wire N__24376;
    wire N__24371;
    wire N__24364;
    wire N__24361;
    wire N__24358;
    wire N__24355;
    wire N__24352;
    wire N__24349;
    wire N__24346;
    wire N__24343;
    wire N__24340;
    wire N__24337;
    wire N__24334;
    wire N__24331;
    wire N__24328;
    wire N__24325;
    wire N__24322;
    wire N__24321;
    wire N__24320;
    wire N__24317;
    wire N__24310;
    wire N__24309;
    wire N__24308;
    wire N__24307;
    wire N__24306;
    wire N__24305;
    wire N__24304;
    wire N__24303;
    wire N__24302;
    wire N__24301;
    wire N__24300;
    wire N__24297;
    wire N__24284;
    wire N__24275;
    wire N__24272;
    wire N__24269;
    wire N__24262;
    wire N__24261;
    wire N__24260;
    wire N__24259;
    wire N__24258;
    wire N__24257;
    wire N__24256;
    wire N__24253;
    wire N__24252;
    wire N__24251;
    wire N__24248;
    wire N__24247;
    wire N__24244;
    wire N__24243;
    wire N__24240;
    wire N__24239;
    wire N__24236;
    wire N__24233;
    wire N__24222;
    wire N__24209;
    wire N__24206;
    wire N__24203;
    wire N__24200;
    wire N__24197;
    wire N__24192;
    wire N__24187;
    wire N__24184;
    wire N__24183;
    wire N__24182;
    wire N__24181;
    wire N__24178;
    wire N__24175;
    wire N__24174;
    wire N__24173;
    wire N__24170;
    wire N__24169;
    wire N__24168;
    wire N__24165;
    wire N__24152;
    wire N__24149;
    wire N__24148;
    wire N__24147;
    wire N__24146;
    wire N__24141;
    wire N__24132;
    wire N__24127;
    wire N__24126;
    wire N__24125;
    wire N__24124;
    wire N__24123;
    wire N__24122;
    wire N__24109;
    wire N__24108;
    wire N__24107;
    wire N__24106;
    wire N__24103;
    wire N__24100;
    wire N__24095;
    wire N__24088;
    wire N__24085;
    wire N__24082;
    wire N__24079;
    wire N__24076;
    wire N__24073;
    wire N__24070;
    wire N__24067;
    wire N__24064;
    wire N__24061;
    wire N__24058;
    wire N__24055;
    wire N__24052;
    wire N__24049;
    wire N__24046;
    wire N__24043;
    wire N__24040;
    wire N__24039;
    wire N__24036;
    wire N__24033;
    wire N__24030;
    wire N__24025;
    wire N__24022;
    wire N__24019;
    wire N__24016;
    wire N__24013;
    wire N__24010;
    wire N__24007;
    wire N__24006;
    wire N__24003;
    wire N__24000;
    wire N__23997;
    wire N__23994;
    wire N__23991;
    wire N__23986;
    wire N__23983;
    wire N__23980;
    wire N__23977;
    wire N__23974;
    wire N__23971;
    wire N__23968;
    wire N__23965;
    wire N__23962;
    wire N__23959;
    wire N__23956;
    wire N__23955;
    wire N__23952;
    wire N__23949;
    wire N__23944;
    wire N__23941;
    wire N__23938;
    wire N__23935;
    wire N__23932;
    wire N__23929;
    wire N__23926;
    wire N__23923;
    wire N__23922;
    wire N__23919;
    wire N__23916;
    wire N__23913;
    wire N__23910;
    wire N__23907;
    wire N__23904;
    wire N__23899;
    wire N__23896;
    wire N__23893;
    wire N__23890;
    wire N__23887;
    wire N__23884;
    wire N__23881;
    wire N__23878;
    wire N__23877;
    wire N__23876;
    wire N__23875;
    wire N__23874;
    wire N__23873;
    wire N__23872;
    wire N__23871;
    wire N__23870;
    wire N__23869;
    wire N__23868;
    wire N__23867;
    wire N__23866;
    wire N__23865;
    wire N__23864;
    wire N__23863;
    wire N__23862;
    wire N__23861;
    wire N__23860;
    wire N__23859;
    wire N__23858;
    wire N__23841;
    wire N__23840;
    wire N__23839;
    wire N__23838;
    wire N__23837;
    wire N__23836;
    wire N__23835;
    wire N__23834;
    wire N__23833;
    wire N__23832;
    wire N__23831;
    wire N__23830;
    wire N__23829;
    wire N__23828;
    wire N__23827;
    wire N__23826;
    wire N__23825;
    wire N__23824;
    wire N__23813;
    wire N__23796;
    wire N__23793;
    wire N__23776;
    wire N__23759;
    wire N__23756;
    wire N__23755;
    wire N__23754;
    wire N__23753;
    wire N__23752;
    wire N__23749;
    wire N__23746;
    wire N__23739;
    wire N__23736;
    wire N__23727;
    wire N__23716;
    wire N__23715;
    wire N__23714;
    wire N__23713;
    wire N__23706;
    wire N__23703;
    wire N__23700;
    wire N__23697;
    wire N__23694;
    wire N__23689;
    wire N__23686;
    wire N__23683;
    wire N__23680;
    wire N__23677;
    wire N__23674;
    wire N__23671;
    wire N__23668;
    wire N__23665;
    wire N__23662;
    wire N__23661;
    wire N__23660;
    wire N__23659;
    wire N__23658;
    wire N__23657;
    wire N__23656;
    wire N__23655;
    wire N__23654;
    wire N__23653;
    wire N__23652;
    wire N__23651;
    wire N__23650;
    wire N__23643;
    wire N__23638;
    wire N__23635;
    wire N__23632;
    wire N__23629;
    wire N__23626;
    wire N__23619;
    wire N__23616;
    wire N__23611;
    wire N__23608;
    wire N__23603;
    wire N__23598;
    wire N__23595;
    wire N__23592;
    wire N__23585;
    wire N__23578;
    wire N__23575;
    wire N__23574;
    wire N__23569;
    wire N__23566;
    wire N__23563;
    wire N__23560;
    wire N__23557;
    wire N__23554;
    wire N__23551;
    wire N__23548;
    wire N__23545;
    wire N__23542;
    wire N__23539;
    wire N__23536;
    wire N__23533;
    wire N__23530;
    wire N__23527;
    wire N__23526;
    wire N__23525;
    wire N__23524;
    wire N__23521;
    wire N__23518;
    wire N__23515;
    wire N__23514;
    wire N__23513;
    wire N__23512;
    wire N__23511;
    wire N__23510;
    wire N__23507;
    wire N__23504;
    wire N__23501;
    wire N__23492;
    wire N__23487;
    wire N__23484;
    wire N__23477;
    wire N__23470;
    wire N__23469;
    wire N__23464;
    wire N__23461;
    wire N__23458;
    wire N__23455;
    wire N__23454;
    wire N__23451;
    wire N__23450;
    wire N__23447;
    wire N__23440;
    wire N__23439;
    wire N__23436;
    wire N__23433;
    wire N__23430;
    wire N__23425;
    wire N__23424;
    wire N__23421;
    wire N__23418;
    wire N__23415;
    wire N__23412;
    wire N__23407;
    wire N__23404;
    wire N__23401;
    wire N__23398;
    wire N__23395;
    wire N__23392;
    wire N__23389;
    wire N__23386;
    wire N__23383;
    wire N__23380;
    wire N__23377;
    wire N__23374;
    wire N__23371;
    wire N__23368;
    wire N__23367;
    wire N__23366;
    wire N__23363;
    wire N__23362;
    wire N__23359;
    wire N__23350;
    wire N__23347;
    wire N__23346;
    wire N__23343;
    wire N__23340;
    wire N__23335;
    wire N__23332;
    wire N__23329;
    wire N__23328;
    wire N__23325;
    wire N__23322;
    wire N__23317;
    wire N__23314;
    wire N__23311;
    wire N__23308;
    wire N__23307;
    wire N__23304;
    wire N__23301;
    wire N__23296;
    wire N__23293;
    wire N__23290;
    wire N__23287;
    wire N__23284;
    wire N__23281;
    wire N__23280;
    wire N__23277;
    wire N__23274;
    wire N__23271;
    wire N__23268;
    wire N__23265;
    wire N__23262;
    wire N__23257;
    wire N__23256;
    wire N__23253;
    wire N__23252;
    wire N__23251;
    wire N__23248;
    wire N__23245;
    wire N__23242;
    wire N__23239;
    wire N__23238;
    wire N__23237;
    wire N__23234;
    wire N__23231;
    wire N__23228;
    wire N__23223;
    wire N__23220;
    wire N__23211;
    wire N__23206;
    wire N__23205;
    wire N__23200;
    wire N__23199;
    wire N__23196;
    wire N__23193;
    wire N__23188;
    wire N__23185;
    wire N__23182;
    wire N__23179;
    wire N__23176;
    wire N__23173;
    wire N__23170;
    wire N__23167;
    wire N__23166;
    wire N__23163;
    wire N__23160;
    wire N__23155;
    wire N__23152;
    wire N__23151;
    wire N__23146;
    wire N__23145;
    wire N__23142;
    wire N__23139;
    wire N__23136;
    wire N__23131;
    wire N__23130;
    wire N__23127;
    wire N__23124;
    wire N__23119;
    wire N__23116;
    wire N__23113;
    wire N__23110;
    wire N__23109;
    wire N__23106;
    wire N__23103;
    wire N__23098;
    wire N__23095;
    wire N__23092;
    wire N__23089;
    wire N__23088;
    wire N__23085;
    wire N__23082;
    wire N__23077;
    wire N__23074;
    wire N__23071;
    wire N__23068;
    wire N__23067;
    wire N__23064;
    wire N__23061;
    wire N__23056;
    wire N__23053;
    wire N__23050;
    wire N__23047;
    wire N__23046;
    wire N__23043;
    wire N__23040;
    wire N__23035;
    wire N__23032;
    wire N__23029;
    wire N__23026;
    wire N__23025;
    wire N__23022;
    wire N__23019;
    wire N__23014;
    wire N__23011;
    wire N__23008;
    wire N__23005;
    wire N__23002;
    wire N__22999;
    wire N__22996;
    wire N__22993;
    wire N__22990;
    wire N__22987;
    wire N__22984;
    wire N__22981;
    wire N__22978;
    wire N__22975;
    wire N__22972;
    wire N__22969;
    wire N__22966;
    wire N__22963;
    wire N__22960;
    wire N__22957;
    wire N__22954;
    wire N__22951;
    wire N__22948;
    wire N__22945;
    wire N__22942;
    wire N__22939;
    wire N__22936;
    wire N__22933;
    wire N__22930;
    wire N__22927;
    wire N__22924;
    wire N__22921;
    wire N__22918;
    wire N__22915;
    wire N__22912;
    wire N__22909;
    wire N__22906;
    wire N__22903;
    wire N__22900;
    wire N__22897;
    wire N__22894;
    wire N__22891;
    wire N__22888;
    wire N__22885;
    wire N__22882;
    wire N__22879;
    wire N__22876;
    wire N__22873;
    wire N__22870;
    wire N__22867;
    wire N__22864;
    wire N__22861;
    wire N__22858;
    wire N__22855;
    wire N__22852;
    wire N__22849;
    wire N__22846;
    wire N__22843;
    wire N__22840;
    wire N__22837;
    wire N__22834;
    wire N__22831;
    wire N__22828;
    wire N__22825;
    wire N__22822;
    wire N__22819;
    wire N__22818;
    wire N__22815;
    wire N__22812;
    wire N__22809;
    wire N__22806;
    wire N__22803;
    wire N__22800;
    wire N__22795;
    wire N__22792;
    wire N__22789;
    wire N__22786;
    wire N__22783;
    wire N__22780;
    wire N__22777;
    wire N__22774;
    wire N__22771;
    wire N__22770;
    wire N__22767;
    wire N__22764;
    wire N__22759;
    wire N__22756;
    wire N__22753;
    wire N__22750;
    wire N__22747;
    wire N__22744;
    wire N__22741;
    wire N__22738;
    wire N__22735;
    wire N__22732;
    wire N__22729;
    wire N__22726;
    wire N__22723;
    wire N__22720;
    wire N__22719;
    wire N__22716;
    wire N__22713;
    wire N__22708;
    wire N__22705;
    wire N__22702;
    wire N__22699;
    wire N__22696;
    wire N__22693;
    wire N__22690;
    wire N__22687;
    wire N__22686;
    wire N__22683;
    wire N__22680;
    wire N__22677;
    wire N__22674;
    wire N__22671;
    wire N__22668;
    wire N__22663;
    wire N__22660;
    wire N__22657;
    wire N__22654;
    wire N__22653;
    wire N__22650;
    wire N__22647;
    wire N__22642;
    wire N__22639;
    wire N__22636;
    wire N__22633;
    wire N__22630;
    wire N__22629;
    wire N__22626;
    wire N__22623;
    wire N__22620;
    wire N__22617;
    wire N__22614;
    wire N__22609;
    wire N__22608;
    wire N__22605;
    wire N__22602;
    wire N__22599;
    wire N__22594;
    wire N__22591;
    wire N__22588;
    wire N__22585;
    wire N__22582;
    wire N__22579;
    wire N__22576;
    wire N__22575;
    wire N__22572;
    wire N__22569;
    wire N__22566;
    wire N__22563;
    wire N__22558;
    wire N__22555;
    wire N__22552;
    wire N__22549;
    wire N__22546;
    wire N__22543;
    wire N__22540;
    wire N__22537;
    wire N__22534;
    wire N__22531;
    wire N__22528;
    wire N__22525;
    wire N__22522;
    wire N__22519;
    wire N__22516;
    wire N__22513;
    wire N__22510;
    wire N__22507;
    wire N__22504;
    wire N__22501;
    wire N__22498;
    wire N__22495;
    wire N__22494;
    wire N__22493;
    wire N__22490;
    wire N__22487;
    wire N__22484;
    wire N__22477;
    wire N__22474;
    wire N__22471;
    wire N__22470;
    wire N__22467;
    wire N__22464;
    wire N__22461;
    wire N__22458;
    wire N__22453;
    wire N__22450;
    wire N__22447;
    wire N__22446;
    wire N__22443;
    wire N__22440;
    wire N__22437;
    wire N__22434;
    wire N__22429;
    wire N__22426;
    wire N__22423;
    wire N__22420;
    wire N__22417;
    wire N__22414;
    wire N__22411;
    wire N__22410;
    wire N__22407;
    wire N__22404;
    wire N__22401;
    wire N__22398;
    wire N__22395;
    wire N__22392;
    wire N__22387;
    wire N__22384;
    wire N__22381;
    wire N__22380;
    wire N__22377;
    wire N__22374;
    wire N__22371;
    wire N__22368;
    wire N__22363;
    wire N__22360;
    wire N__22357;
    wire N__22354;
    wire N__22351;
    wire N__22350;
    wire N__22347;
    wire N__22344;
    wire N__22339;
    wire N__22336;
    wire N__22333;
    wire N__22330;
    wire N__22327;
    wire N__22324;
    wire N__22321;
    wire N__22320;
    wire N__22317;
    wire N__22314;
    wire N__22311;
    wire N__22308;
    wire N__22305;
    wire N__22302;
    wire N__22297;
    wire N__22294;
    wire N__22291;
    wire N__22288;
    wire N__22287;
    wire N__22284;
    wire N__22281;
    wire N__22276;
    wire N__22273;
    wire N__22270;
    wire N__22267;
    wire N__22264;
    wire N__22261;
    wire N__22258;
    wire N__22255;
    wire N__22252;
    wire N__22249;
    wire N__22246;
    wire N__22243;
    wire N__22242;
    wire N__22239;
    wire N__22236;
    wire N__22233;
    wire N__22228;
    wire N__22225;
    wire N__22222;
    wire N__22221;
    wire N__22220;
    wire N__22219;
    wire N__22218;
    wire N__22217;
    wire N__22216;
    wire N__22213;
    wire N__22200;
    wire N__22195;
    wire N__22192;
    wire N__22189;
    wire N__22186;
    wire N__22183;
    wire N__22180;
    wire N__22179;
    wire N__22176;
    wire N__22173;
    wire N__22168;
    wire N__22165;
    wire N__22162;
    wire N__22159;
    wire N__22158;
    wire N__22155;
    wire N__22152;
    wire N__22149;
    wire N__22146;
    wire N__22143;
    wire N__22140;
    wire N__22135;
    wire N__22134;
    wire N__22131;
    wire N__22128;
    wire N__22123;
    wire N__22120;
    wire N__22117;
    wire N__22114;
    wire N__22113;
    wire N__22110;
    wire N__22107;
    wire N__22102;
    wire N__22099;
    wire N__22096;
    wire N__22093;
    wire N__22090;
    wire N__22087;
    wire N__22086;
    wire N__22083;
    wire N__22080;
    wire N__22075;
    wire N__22072;
    wire N__22069;
    wire N__22066;
    wire N__22063;
    wire N__22062;
    wire N__22059;
    wire N__22056;
    wire N__22053;
    wire N__22048;
    wire N__22045;
    wire N__22042;
    wire N__22039;
    wire N__22036;
    wire N__22035;
    wire N__22032;
    wire N__22029;
    wire N__22026;
    wire N__22023;
    wire N__22020;
    wire N__22015;
    wire N__22012;
    wire N__22009;
    wire N__22006;
    wire N__22003;
    wire N__22000;
    wire N__21997;
    wire N__21994;
    wire N__21991;
    wire N__21988;
    wire N__21987;
    wire N__21984;
    wire N__21981;
    wire N__21978;
    wire N__21975;
    wire N__21970;
    wire N__21967;
    wire N__21964;
    wire N__21961;
    wire N__21960;
    wire N__21959;
    wire N__21956;
    wire N__21955;
    wire N__21952;
    wire N__21951;
    wire N__21950;
    wire N__21947;
    wire N__21944;
    wire N__21941;
    wire N__21940;
    wire N__21937;
    wire N__21934;
    wire N__21931;
    wire N__21928;
    wire N__21923;
    wire N__21920;
    wire N__21917;
    wire N__21914;
    wire N__21911;
    wire N__21906;
    wire N__21903;
    wire N__21896;
    wire N__21891;
    wire N__21886;
    wire N__21885;
    wire N__21880;
    wire N__21877;
    wire N__21874;
    wire N__21873;
    wire N__21870;
    wire N__21867;
    wire N__21862;
    wire N__21859;
    wire N__21856;
    wire N__21853;
    wire N__21852;
    wire N__21851;
    wire N__21850;
    wire N__21841;
    wire N__21840;
    wire N__21837;
    wire N__21834;
    wire N__21831;
    wire N__21828;
    wire N__21825;
    wire N__21822;
    wire N__21819;
    wire N__21816;
    wire N__21813;
    wire N__21810;
    wire N__21805;
    wire N__21804;
    wire N__21803;
    wire N__21800;
    wire N__21795;
    wire N__21792;
    wire N__21789;
    wire N__21786;
    wire N__21783;
    wire N__21780;
    wire N__21777;
    wire N__21774;
    wire N__21769;
    wire N__21766;
    wire N__21763;
    wire N__21760;
    wire N__21757;
    wire N__21754;
    wire N__21751;
    wire N__21748;
    wire N__21745;
    wire N__21742;
    wire N__21739;
    wire N__21736;
    wire N__21733;
    wire N__21730;
    wire N__21727;
    wire N__21724;
    wire N__21721;
    wire N__21718;
    wire N__21715;
    wire N__21712;
    wire N__21709;
    wire N__21706;
    wire N__21705;
    wire N__21702;
    wire N__21701;
    wire N__21694;
    wire N__21693;
    wire N__21690;
    wire N__21687;
    wire N__21682;
    wire N__21681;
    wire N__21678;
    wire N__21675;
    wire N__21670;
    wire N__21667;
    wire N__21664;
    wire N__21661;
    wire N__21658;
    wire N__21655;
    wire N__21652;
    wire N__21649;
    wire N__21646;
    wire N__21645;
    wire N__21644;
    wire N__21643;
    wire N__21638;
    wire N__21635;
    wire N__21632;
    wire N__21625;
    wire N__21622;
    wire N__21619;
    wire N__21616;
    wire N__21613;
    wire N__21610;
    wire N__21607;
    wire N__21604;
    wire N__21601;
    wire N__21598;
    wire N__21595;
    wire N__21592;
    wire N__21589;
    wire N__21586;
    wire N__21583;
    wire N__21580;
    wire N__21577;
    wire N__21574;
    wire N__21571;
    wire N__21568;
    wire N__21565;
    wire N__21562;
    wire N__21559;
    wire N__21556;
    wire N__21555;
    wire N__21552;
    wire N__21549;
    wire N__21548;
    wire N__21543;
    wire N__21540;
    wire N__21537;
    wire N__21532;
    wire N__21529;
    wire N__21526;
    wire N__21523;
    wire N__21522;
    wire N__21519;
    wire N__21516;
    wire N__21511;
    wire N__21508;
    wire N__21505;
    wire N__21502;
    wire N__21499;
    wire N__21498;
    wire N__21497;
    wire N__21494;
    wire N__21491;
    wire N__21490;
    wire N__21487;
    wire N__21484;
    wire N__21483;
    wire N__21482;
    wire N__21477;
    wire N__21472;
    wire N__21469;
    wire N__21466;
    wire N__21457;
    wire N__21456;
    wire N__21455;
    wire N__21450;
    wire N__21447;
    wire N__21442;
    wire N__21439;
    wire N__21436;
    wire N__21433;
    wire N__21430;
    wire N__21427;
    wire N__21426;
    wire N__21425;
    wire N__21424;
    wire N__21423;
    wire N__21420;
    wire N__21413;
    wire N__21410;
    wire N__21407;
    wire N__21404;
    wire N__21401;
    wire N__21394;
    wire N__21391;
    wire N__21388;
    wire N__21385;
    wire N__21382;
    wire N__21379;
    wire N__21376;
    wire N__21375;
    wire N__21370;
    wire N__21367;
    wire N__21366;
    wire N__21365;
    wire N__21362;
    wire N__21357;
    wire N__21352;
    wire N__21349;
    wire N__21346;
    wire N__21343;
    wire N__21340;
    wire N__21337;
    wire N__21334;
    wire N__21331;
    wire N__21328;
    wire N__21325;
    wire N__21322;
    wire N__21319;
    wire N__21316;
    wire N__21313;
    wire N__21310;
    wire N__21307;
    wire N__21304;
    wire N__21301;
    wire N__21298;
    wire N__21295;
    wire N__21292;
    wire N__21289;
    wire N__21286;
    wire N__21283;
    wire N__21280;
    wire N__21277;
    wire N__21274;
    wire N__21271;
    wire N__21268;
    wire N__21265;
    wire N__21262;
    wire N__21259;
    wire N__21256;
    wire N__21253;
    wire N__21250;
    wire N__21247;
    wire N__21244;
    wire N__21241;
    wire N__21238;
    wire N__21235;
    wire N__21232;
    wire N__21229;
    wire N__21226;
    wire N__21223;
    wire N__21220;
    wire N__21217;
    wire N__21214;
    wire N__21211;
    wire N__21208;
    wire N__21205;
    wire N__21202;
    wire N__21199;
    wire N__21196;
    wire N__21193;
    wire N__21190;
    wire N__21187;
    wire N__21184;
    wire N__21181;
    wire N__21178;
    wire N__21175;
    wire N__21172;
    wire N__21169;
    wire N__21166;
    wire N__21165;
    wire N__21164;
    wire N__21163;
    wire N__21154;
    wire N__21151;
    wire N__21148;
    wire N__21145;
    wire N__21142;
    wire N__21139;
    wire N__21138;
    wire N__21137;
    wire N__21136;
    wire N__21135;
    wire N__21134;
    wire N__21131;
    wire N__21130;
    wire N__21129;
    wire N__21122;
    wire N__21117;
    wire N__21114;
    wire N__21111;
    wire N__21108;
    wire N__21105;
    wire N__21100;
    wire N__21091;
    wire N__21088;
    wire N__21085;
    wire N__21082;
    wire N__21079;
    wire N__21078;
    wire N__21077;
    wire N__21076;
    wire N__21075;
    wire N__21074;
    wire N__21073;
    wire N__21072;
    wire N__21069;
    wire N__21068;
    wire N__21061;
    wire N__21052;
    wire N__21047;
    wire N__21042;
    wire N__21037;
    wire N__21036;
    wire N__21033;
    wire N__21030;
    wire N__21027;
    wire N__21022;
    wire N__21021;
    wire N__21016;
    wire N__21015;
    wire N__21014;
    wire N__21011;
    wire N__21008;
    wire N__21007;
    wire N__21004;
    wire N__21001;
    wire N__20996;
    wire N__20993;
    wire N__20986;
    wire N__20983;
    wire N__20980;
    wire N__20979;
    wire N__20976;
    wire N__20973;
    wire N__20968;
    wire N__20965;
    wire N__20962;
    wire N__20959;
    wire N__20956;
    wire N__20953;
    wire N__20950;
    wire N__20947;
    wire N__20944;
    wire N__20941;
    wire N__20940;
    wire N__20937;
    wire N__20934;
    wire N__20929;
    wire N__20926;
    wire N__20923;
    wire N__20922;
    wire N__20919;
    wire N__20916;
    wire N__20911;
    wire N__20908;
    wire N__20907;
    wire N__20902;
    wire N__20899;
    wire N__20896;
    wire N__20893;
    wire N__20890;
    wire N__20887;
    wire N__20884;
    wire N__20883;
    wire N__20880;
    wire N__20877;
    wire N__20874;
    wire N__20873;
    wire N__20870;
    wire N__20867;
    wire N__20864;
    wire N__20861;
    wire N__20856;
    wire N__20851;
    wire N__20850;
    wire N__20847;
    wire N__20844;
    wire N__20841;
    wire N__20838;
    wire N__20833;
    wire N__20830;
    wire N__20829;
    wire N__20826;
    wire N__20823;
    wire N__20820;
    wire N__20817;
    wire N__20812;
    wire N__20809;
    wire N__20806;
    wire N__20803;
    wire N__20802;
    wire N__20801;
    wire N__20798;
    wire N__20793;
    wire N__20788;
    wire N__20787;
    wire N__20786;
    wire N__20785;
    wire N__20776;
    wire N__20773;
    wire N__20770;
    wire N__20767;
    wire N__20764;
    wire N__20761;
    wire N__20758;
    wire N__20755;
    wire N__20752;
    wire N__20749;
    wire N__20748;
    wire N__20747;
    wire N__20744;
    wire N__20739;
    wire N__20734;
    wire N__20731;
    wire N__20728;
    wire N__20725;
    wire N__20722;
    wire N__20719;
    wire N__20716;
    wire N__20713;
    wire N__20710;
    wire N__20707;
    wire N__20704;
    wire N__20701;
    wire N__20698;
    wire N__20697;
    wire N__20696;
    wire N__20693;
    wire N__20688;
    wire N__20683;
    wire N__20680;
    wire N__20677;
    wire N__20674;
    wire N__20673;
    wire N__20672;
    wire N__20669;
    wire N__20666;
    wire N__20663;
    wire N__20660;
    wire N__20653;
    wire N__20650;
    wire N__20647;
    wire N__20646;
    wire N__20645;
    wire N__20644;
    wire N__20635;
    wire N__20632;
    wire N__20631;
    wire N__20630;
    wire N__20629;
    wire N__20620;
    wire N__20617;
    wire N__20614;
    wire N__20611;
    wire N__20608;
    wire N__20605;
    wire N__20602;
    wire N__20599;
    wire N__20596;
    wire N__20593;
    wire N__20590;
    wire N__20587;
    wire N__20584;
    wire N__20581;
    wire N__20578;
    wire N__20575;
    wire N__20572;
    wire N__20569;
    wire N__20566;
    wire N__20563;
    wire N__20560;
    wire N__20559;
    wire N__20558;
    wire N__20555;
    wire N__20552;
    wire N__20549;
    wire N__20546;
    wire N__20543;
    wire N__20536;
    wire N__20533;
    wire N__20530;
    wire N__20529;
    wire N__20528;
    wire N__20525;
    wire N__20522;
    wire N__20519;
    wire N__20512;
    wire N__20509;
    wire N__20506;
    wire N__20505;
    wire N__20502;
    wire N__20501;
    wire N__20498;
    wire N__20495;
    wire N__20492;
    wire N__20485;
    wire N__20482;
    wire N__20479;
    wire N__20478;
    wire N__20477;
    wire N__20474;
    wire N__20471;
    wire N__20468;
    wire N__20461;
    wire N__20458;
    wire N__20455;
    wire N__20454;
    wire N__20453;
    wire N__20450;
    wire N__20447;
    wire N__20444;
    wire N__20437;
    wire N__20434;
    wire N__20431;
    wire N__20430;
    wire N__20429;
    wire N__20426;
    wire N__20423;
    wire N__20420;
    wire N__20413;
    wire N__20410;
    wire N__20407;
    wire N__20404;
    wire N__20403;
    wire N__20402;
    wire N__20399;
    wire N__20396;
    wire N__20393;
    wire N__20386;
    wire N__20383;
    wire N__20382;
    wire N__20381;
    wire N__20380;
    wire N__20377;
    wire N__20370;
    wire N__20365;
    wire N__20362;
    wire N__20361;
    wire N__20358;
    wire N__20355;
    wire N__20352;
    wire N__20349;
    wire N__20348;
    wire N__20347;
    wire N__20342;
    wire N__20339;
    wire N__20336;
    wire N__20329;
    wire N__20326;
    wire N__20323;
    wire N__20320;
    wire N__20317;
    wire N__20314;
    wire N__20311;
    wire N__20308;
    wire N__20305;
    wire N__20302;
    wire N__20299;
    wire N__20296;
    wire N__20293;
    wire N__20290;
    wire N__20287;
    wire N__20284;
    wire N__20281;
    wire N__20278;
    wire N__20275;
    wire N__20272;
    wire N__20269;
    wire N__20266;
    wire N__20265;
    wire N__20264;
    wire N__20263;
    wire N__20260;
    wire N__20257;
    wire N__20252;
    wire N__20251;
    wire N__20250;
    wire N__20249;
    wire N__20246;
    wire N__20241;
    wire N__20234;
    wire N__20229;
    wire N__20224;
    wire N__20221;
    wire N__20218;
    wire N__20215;
    wire N__20212;
    wire N__20209;
    wire N__20206;
    wire N__20203;
    wire N__20200;
    wire N__20197;
    wire N__20196;
    wire N__20193;
    wire N__20190;
    wire N__20185;
    wire N__20182;
    wire N__20181;
    wire N__20176;
    wire N__20173;
    wire N__20170;
    wire N__20167;
    wire N__20164;
    wire N__20161;
    wire N__20158;
    wire N__20155;
    wire N__20152;
    wire N__20151;
    wire N__20146;
    wire N__20143;
    wire N__20140;
    wire N__20137;
    wire N__20134;
    wire N__20131;
    wire N__20128;
    wire N__20125;
    wire N__20122;
    wire N__20119;
    wire N__20116;
    wire N__20113;
    wire N__20110;
    wire N__20107;
    wire N__20106;
    wire N__20105;
    wire N__20102;
    wire N__20097;
    wire N__20094;
    wire N__20091;
    wire N__20086;
    wire N__20085;
    wire N__20082;
    wire N__20079;
    wire N__20078;
    wire N__20073;
    wire N__20070;
    wire N__20065;
    wire N__20062;
    wire N__20061;
    wire N__20060;
    wire N__20059;
    wire N__20054;
    wire N__20049;
    wire N__20044;
    wire N__20043;
    wire N__20042;
    wire N__20041;
    wire N__20034;
    wire N__20031;
    wire N__20026;
    wire N__20023;
    wire N__20022;
    wire N__20021;
    wire N__20020;
    wire N__20019;
    wire N__20018;
    wire N__20015;
    wire N__20010;
    wire N__20003;
    wire N__19996;
    wire N__19995;
    wire N__19992;
    wire N__19989;
    wire N__19984;
    wire N__19983;
    wire N__19982;
    wire N__19981;
    wire N__19978;
    wire N__19975;
    wire N__19972;
    wire N__19969;
    wire N__19966;
    wire N__19963;
    wire N__19954;
    wire N__19951;
    wire N__19948;
    wire N__19947;
    wire N__19944;
    wire N__19941;
    wire N__19938;
    wire N__19933;
    wire N__19930;
    wire N__19927;
    wire N__19926;
    wire N__19923;
    wire N__19920;
    wire N__19915;
    wire N__19914;
    wire N__19913;
    wire N__19908;
    wire N__19905;
    wire N__19900;
    wire N__19897;
    wire N__19894;
    wire N__19893;
    wire N__19890;
    wire N__19887;
    wire N__19882;
    wire N__19879;
    wire N__19876;
    wire N__19873;
    wire N__19870;
    wire N__19867;
    wire N__19864;
    wire N__19861;
    wire N__19860;
    wire N__19859;
    wire N__19856;
    wire N__19855;
    wire N__19854;
    wire N__19851;
    wire N__19848;
    wire N__19845;
    wire N__19840;
    wire N__19835;
    wire N__19828;
    wire N__19827;
    wire N__19826;
    wire N__19825;
    wire N__19824;
    wire N__19823;
    wire N__19822;
    wire N__19821;
    wire N__19808;
    wire N__19803;
    wire N__19798;
    wire N__19795;
    wire N__19792;
    wire N__19789;
    wire N__19786;
    wire N__19783;
    wire N__19782;
    wire N__19779;
    wire N__19776;
    wire N__19771;
    wire N__19770;
    wire N__19767;
    wire N__19764;
    wire N__19761;
    wire N__19756;
    wire N__19753;
    wire N__19750;
    wire N__19747;
    wire N__19744;
    wire N__19741;
    wire N__19738;
    wire N__19735;
    wire N__19734;
    wire N__19733;
    wire N__19730;
    wire N__19725;
    wire N__19720;
    wire N__19717;
    wire N__19714;
    wire N__19711;
    wire N__19710;
    wire N__19707;
    wire N__19704;
    wire N__19699;
    wire N__19696;
    wire N__19693;
    wire N__19692;
    wire N__19689;
    wire N__19686;
    wire N__19681;
    wire N__19678;
    wire N__19675;
    wire N__19672;
    wire N__19671;
    wire N__19668;
    wire N__19665;
    wire N__19660;
    wire N__19657;
    wire N__19656;
    wire N__19653;
    wire N__19650;
    wire N__19645;
    wire N__19642;
    wire N__19639;
    wire N__19636;
    wire N__19633;
    wire N__19630;
    wire N__19627;
    wire N__19624;
    wire N__19621;
    wire N__19618;
    wire N__19615;
    wire N__19612;
    wire N__19609;
    wire N__19606;
    wire N__19603;
    wire N__19600;
    wire N__19599;
    wire N__19596;
    wire N__19593;
    wire N__19588;
    wire N__19585;
    wire N__19582;
    wire N__19579;
    wire N__19576;
    wire N__19573;
    wire N__19570;
    wire N__19567;
    wire N__19564;
    wire N__19561;
    wire N__19558;
    wire N__19555;
    wire N__19552;
    wire N__19549;
    wire N__19546;
    wire N__19543;
    wire N__19540;
    wire N__19537;
    wire N__19534;
    wire N__19531;
    wire N__19528;
    wire N__19525;
    wire N__19522;
    wire N__19519;
    wire N__19516;
    wire N__19513;
    wire N__19510;
    wire N__19507;
    wire N__19504;
    wire N__19501;
    wire N__19498;
    wire N__19495;
    wire N__19492;
    wire N__19489;
    wire N__19488;
    wire N__19483;
    wire N__19480;
    wire N__19477;
    wire N__19476;
    wire N__19473;
    wire N__19470;
    wire N__19465;
    wire N__19464;
    wire N__19461;
    wire N__19458;
    wire N__19453;
    wire N__19450;
    wire N__19447;
    wire N__19444;
    wire N__19441;
    wire N__19440;
    wire N__19439;
    wire N__19438;
    wire N__19435;
    wire N__19430;
    wire N__19427;
    wire N__19420;
    wire N__19417;
    wire N__19414;
    wire N__19411;
    wire N__19408;
    wire N__19405;
    wire N__19402;
    wire N__19399;
    wire N__19398;
    wire N__19397;
    wire N__19394;
    wire N__19391;
    wire N__19388;
    wire N__19381;
    wire N__19378;
    wire N__19375;
    wire N__19372;
    wire N__19369;
    wire N__19366;
    wire N__19363;
    wire N__19360;
    wire N__19357;
    wire N__19354;
    wire N__19351;
    wire N__19350;
    wire N__19347;
    wire N__19344;
    wire N__19339;
    wire N__19336;
    wire N__19333;
    wire N__19330;
    wire N__19327;
    wire N__19324;
    wire N__19321;
    wire N__19318;
    wire N__19317;
    wire N__19314;
    wire N__19311;
    wire N__19306;
    wire N__19305;
    wire N__19302;
    wire N__19299;
    wire N__19296;
    wire N__19291;
    wire N__19290;
    wire N__19287;
    wire N__19284;
    wire N__19281;
    wire N__19278;
    wire N__19273;
    wire N__19272;
    wire N__19269;
    wire N__19266;
    wire N__19261;
    wire N__19258;
    wire N__19255;
    wire N__19252;
    wire N__19249;
    wire N__19246;
    wire N__19243;
    wire N__19240;
    wire N__19237;
    wire N__19236;
    wire N__19233;
    wire N__19230;
    wire N__19225;
    wire N__19222;
    wire N__19219;
    wire N__19216;
    wire N__19213;
    wire N__19212;
    wire N__19209;
    wire N__19206;
    wire N__19201;
    wire N__19198;
    wire N__19195;
    wire N__19192;
    wire N__19189;
    wire N__19186;
    wire N__19183;
    wire N__19180;
    wire N__19179;
    wire N__19176;
    wire N__19173;
    wire N__19168;
    wire N__19165;
    wire N__19162;
    wire N__19159;
    wire N__19156;
    wire N__19153;
    wire N__19150;
    wire N__19149;
    wire N__19146;
    wire N__19143;
    wire N__19138;
    wire N__19137;
    wire N__19136;
    wire N__19135;
    wire N__19134;
    wire N__19133;
    wire N__19132;
    wire N__19131;
    wire N__19120;
    wire N__19115;
    wire N__19112;
    wire N__19105;
    wire N__19102;
    wire N__19099;
    wire N__19096;
    wire N__19093;
    wire N__19090;
    wire N__19087;
    wire N__19086;
    wire N__19083;
    wire N__19080;
    wire N__19077;
    wire N__19072;
    wire N__19071;
    wire N__19070;
    wire N__19067;
    wire N__19064;
    wire N__19061;
    wire N__19058;
    wire N__19055;
    wire N__19052;
    wire N__19045;
    wire N__19042;
    wire N__19039;
    wire N__19036;
    wire N__19033;
    wire N__19030;
    wire N__19027;
    wire N__19024;
    wire N__19021;
    wire N__19020;
    wire N__19017;
    wire N__19014;
    wire N__19009;
    wire N__19006;
    wire N__19005;
    wire N__19002;
    wire N__18999;
    wire N__18994;
    wire N__18991;
    wire N__18990;
    wire N__18987;
    wire N__18984;
    wire N__18981;
    wire N__18978;
    wire N__18973;
    wire N__18970;
    wire N__18967;
    wire N__18964;
    wire N__18961;
    wire N__18958;
    wire N__18955;
    wire N__18952;
    wire N__18949;
    wire N__18948;
    wire N__18945;
    wire N__18942;
    wire N__18937;
    wire N__18934;
    wire N__18931;
    wire N__18928;
    wire N__18925;
    wire N__18922;
    wire N__18919;
    wire N__18916;
    wire N__18915;
    wire N__18912;
    wire N__18909;
    wire N__18904;
    wire N__18901;
    wire N__18898;
    wire N__18895;
    wire N__18892;
    wire N__18889;
    wire N__18888;
    wire N__18885;
    wire N__18882;
    wire N__18879;
    wire N__18876;
    wire N__18875;
    wire N__18872;
    wire N__18869;
    wire N__18866;
    wire N__18859;
    wire N__18858;
    wire N__18857;
    wire N__18856;
    wire N__18855;
    wire N__18854;
    wire N__18853;
    wire N__18852;
    wire N__18851;
    wire N__18850;
    wire N__18849;
    wire N__18848;
    wire N__18847;
    wire N__18846;
    wire N__18845;
    wire N__18828;
    wire N__18819;
    wire N__18812;
    wire N__18805;
    wire N__18802;
    wire N__18799;
    wire N__18796;
    wire N__18793;
    wire N__18790;
    wire N__18787;
    wire N__18786;
    wire N__18783;
    wire N__18780;
    wire N__18775;
    wire N__18772;
    wire N__18771;
    wire N__18768;
    wire N__18765;
    wire N__18762;
    wire N__18759;
    wire N__18756;
    wire N__18751;
    wire N__18748;
    wire N__18745;
    wire N__18742;
    wire N__18739;
    wire N__18736;
    wire N__18733;
    wire N__18730;
    wire N__18727;
    wire N__18724;
    wire N__18721;
    wire N__18718;
    wire N__18715;
    wire N__18712;
    wire N__18709;
    wire N__18706;
    wire N__18703;
    wire N__18700;
    wire N__18697;
    wire N__18694;
    wire N__18691;
    wire N__18688;
    wire N__18685;
    wire N__18682;
    wire N__18679;
    wire N__18676;
    wire N__18675;
    wire N__18672;
    wire N__18669;
    wire N__18664;
    wire N__18661;
    wire N__18658;
    wire N__18657;
    wire N__18654;
    wire N__18651;
    wire N__18648;
    wire N__18645;
    wire N__18642;
    wire N__18639;
    wire N__18636;
    wire N__18631;
    wire N__18628;
    wire N__18625;
    wire N__18622;
    wire N__18619;
    wire N__18616;
    wire N__18613;
    wire N__18610;
    wire N__18607;
    wire N__18604;
    wire N__18601;
    wire N__18598;
    wire N__18595;
    wire N__18592;
    wire N__18589;
    wire N__18586;
    wire N__18583;
    wire N__18580;
    wire N__18577;
    wire N__18574;
    wire N__18571;
    wire N__18568;
    wire N__18565;
    wire N__18562;
    wire N__18559;
    wire N__18556;
    wire N__18553;
    wire N__18550;
    wire N__18547;
    wire N__18544;
    wire N__18541;
    wire N__18538;
    wire N__18535;
    wire N__18532;
    wire N__18529;
    wire N__18526;
    wire N__18523;
    wire N__18520;
    wire N__18517;
    wire N__18514;
    wire N__18511;
    wire N__18508;
    wire N__18505;
    wire N__18504;
    wire N__18501;
    wire N__18498;
    wire N__18493;
    wire N__18490;
    wire N__18487;
    wire N__18484;
    wire N__18481;
    wire N__18478;
    wire N__18475;
    wire N__18472;
    wire N__18469;
    wire N__18466;
    wire N__18465;
    wire N__18462;
    wire N__18459;
    wire N__18454;
    wire N__18451;
    wire N__18448;
    wire N__18445;
    wire N__18442;
    wire N__18439;
    wire N__18436;
    wire N__18433;
    wire N__18430;
    wire N__18427;
    wire N__18424;
    wire N__18421;
    wire N__18418;
    wire N__18415;
    wire N__18414;
    wire N__18413;
    wire N__18410;
    wire N__18407;
    wire N__18402;
    wire N__18397;
    wire N__18394;
    wire N__18391;
    wire N__18390;
    wire N__18389;
    wire N__18386;
    wire N__18383;
    wire N__18380;
    wire N__18373;
    wire N__18370;
    wire N__18367;
    wire N__18364;
    wire N__18361;
    wire N__18358;
    wire N__18355;
    wire N__18352;
    wire N__18349;
    wire N__18346;
    wire N__18343;
    wire N__18340;
    wire N__18337;
    wire N__18334;
    wire N__18331;
    wire N__18328;
    wire N__18325;
    wire N__18322;
    wire N__18319;
    wire N__18316;
    wire N__18313;
    wire N__18310;
    wire N__18307;
    wire N__18304;
    wire N__18301;
    wire N__18298;
    wire N__18295;
    wire N__18292;
    wire N__18289;
    wire N__18286;
    wire N__18283;
    wire N__18280;
    wire N__18277;
    wire N__18274;
    wire N__18271;
    wire N__18268;
    wire N__18265;
    wire N__18262;
    wire N__18259;
    wire N__18256;
    wire N__18253;
    wire N__18250;
    wire N__18247;
    wire VCCG0;
    wire GNDG0;
    wire arst_i_c;
    wire arst_i_c_i;
    wire dmarq_pad_i_c;
    wire bfn_1_18_0_;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_cry_0 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_cry_1 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_cry_2 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_cry_3 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_cry_4 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_cry_5 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_cry_6 ;
    wire CONSTANT_ONE_NET_cascade_;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_s_0 ;
    wire \u1.cDMARQ ;
    wire intrq_pad_i_c;
    wire bfn_2_17_0_;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_cry_0 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_cry_1 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_cry_2 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_cry_3 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_cry_4 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_cry_5 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_cry_6 ;
    wire \u1.DMA_control.Teoc_7 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.val_c7_0_3_cascade_ ;
    wire \u1.Tdone_i_cascade_ ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNIDE5P1Z0Z_0 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.rciZ0 ;
    wire \u1.DMA_control.dTfw ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.QiZ0Z_0 ;
    wire bfn_2_21_0_;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_cry_0 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.QiZ0Z_2 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_s_2 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_cry_1 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_cry_2 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_cry_3 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_cry_4 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_cry_5 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.QiZ0Z_7 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_cry_6 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_s_7 ;
    wire \u1.DMA_control.Teoc_0 ;
    wire \u1.DMA_control.Teoc_2 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.N_2413_iZ0_cascade_ ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_s_0 ;
    wire \u1.DMA_control.Tm_2 ;
    wire bfn_2_24_0_;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_s_1 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_cry_0 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_s_2 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_cry_1 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_s_3 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_cry_2 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_s_4 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_cry_3 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_s_5 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_cry_4 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_s_6 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_cry_5 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_cry_6 ;
    wire wb_cyc_i_c;
    wire wb_stb_i_c;
    wire \u1.cINTRQ ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_s_0 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_s_1 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_s_2 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_s_3 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_s_4 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_s_5 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_s_6 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_s_7 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.val_c8_cascade_ ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.N_1545_cascade_ ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_s_1 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_s_6 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_s_7 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.val_c8_0_3 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_s_3 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.QiZ0Z_3 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.QiZ0Z_1 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNIPRNIZ0Z_0_cascade_ ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.QiZ0Z_6 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.val_c7_0_3 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_s_2 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.QiZ0Z_2 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_s_4 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.QiZ0Z_4 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_s_0 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.QiZ0Z_0 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.N_1545 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_s_5 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.QiZ0Z_5 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.N_290 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_1_sqmuxa_i_x0_0 ;
    wire \u1.DMA_control.Teoc_1 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_s_1 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.QiZ0Z_1 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_s_3 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.QiZ0Z_3 ;
    wire \u1.DMA_control.Teoc_4 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_s_4 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.QiZ0Z_4 ;
    wire \u1.DMA_control.Teoc_5 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_s_5 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.QiZ0Z_5 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_1_sqmuxa_i ;
    wire \u1.DMA_control.Teoc_6 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_s_6 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.QiZ0Z_6 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qie_0_iZ0 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.rd_dstrb ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.Tddone_i_cascade_ ;
    wire diown_pad_o_c;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.QiZ0Z_3 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.QiZ0Z_2 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.QiZ0Z_4 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.QiZ0Z_1 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.val_c8_a0_4_cascade_ ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.Tmdone_i_i_cascade_ ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.QiZ0Z_6 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.QiZ0Z_5 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.val_c8_a0_3 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.val_c8_a0_3_cascade_ ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.Qi_0 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.N_2415_i_xZ0Z1_cascade_ ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.val_c8_a0_4 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.DIOW_RNO_1_0 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.DIOW_RNOZ0Z_0 ;
    wire \u1.DMAdiow ;
    wire \u1.N_1395_cascade_ ;
    wire dd_padoe_o_c;
    wire \u1.N_1387_cascade_ ;
    wire \u1.PIOoe ;
    wire \u1.PIO_control.pong_d_9 ;
    wire \u1.N_1434_cascade_ ;
    wire dd_pad_o_c_9;
    wire \u1.N_1387 ;
    wire iordy_pad_i_c;
    wire \u1.cIORDY ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qilde_i_sxZ0 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.rci_3_i_a0_4_cascade_ ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qilde_i_sxZ0_cascade_ ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.N_1083 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.rci_3_i_a0_5 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.rci_3_i_a0_6 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.N_1377_cascade_ ;
    wire \u1.PIOdior ;
    wire diorn_pad_o_c;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.DIOR_RNOZ0Z_1 ;
    wire \u1.PIO_control.N_1450_cascade_ ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.DIOW_RNOZ0Z_1_cascade_ ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.N_1378_cascade_ ;
    wire \u1.PIOdiow ;
    wire bfn_4_20_0_;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_cry_0 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_cry_1 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_cry_2 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_cry_3 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_cry_4 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_cry_5 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_cry_6 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.val_c8_0_4 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_s_2 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.QiZ0Z_2 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_s_5 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.QiZ0Z_5 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_s_6 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.QiZ0Z_6 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_s_7 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.QiZ0Z_7 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_s_1 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.QiZ0Z_1 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.val_c8_0_3 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_s_3 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.QiZ0Z_3 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_s_0 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.Qi_0_0 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.N_2415_i ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_s_4 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.QiZ0Z_4 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qie_0_iZ0 ;
    wire \u1.DMA_control.iDMA_req_2_0_0_a2_0_2_cascade_ ;
    wire DMA_Ack_c;
    wire irq;
    wire \u0.dirq ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.DIOR_RNO_1_0 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.DIOR_RNOZ0Z_0 ;
    wire \u1.DMAdior ;
    wire \u1.DMA_control.igo ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.rci ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.Tmdone_i_i ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.Tddone_i ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.rci_0 ;
    wire \u1.Tfw ;
    wire \u1.DMA_control.iDMA_req_2_0_0_a2_1 ;
    wire \u1.DMA_control.N_1769 ;
    wire DMA_req_c;
    wire \u1.PIO_control.pong_d_2 ;
    wire \u1.N_1428_cascade_ ;
    wire dd_pad_o_c_2;
    wire \u1.PIO_control.pong_d_3 ;
    wire \u1.N_1449_cascade_ ;
    wire dd_pad_o_c_3;
    wire \u1.PIO_control.pong_d_15 ;
    wire \u1.PIO_control.pong_d_4 ;
    wire \u1.N_1436 ;
    wire dd_pad_o_c_15;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.Qi_6 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.Qi_5 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.Qi_7 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.Qi_2 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.Qi_4 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.Qi_3 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.val_c8_0_4_cascade_ ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.Qi_1 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.rci ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.val_c8_0_5_cascade_ ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.Qi_0 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.busy_3_i_0 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.N_1371_cascade_ ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.hold_goZ0 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.busyZ0 ;
    wire \u1.PIO_control.ping_d_9 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.val_c8_0_4_cascade_ ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_1_sqmuxa_i_xZ0Z0_cascade_ ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.val_c8_0_4 ;
    wire \u1.sIORDYZ0 ;
    wire da_pad_o_c_2;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.N_1358 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.N_1358_cascade_ ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.rciZ0 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.QiZ0Z_7 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.val_c7 ;
    wire \u1.N_1382 ;
    wire \u1.PIOdone_i_cascade_ ;
    wire \u1.N_1372 ;
    wire \u1.PIOgoZ0 ;
    wire N_468_cascade_;
    wire \u1.PIO_control.N_2409_cascade_ ;
    wire \u1.PIO_control.ping_valid_3_0_a2_0_1 ;
    wire \u1.PIO_control.pong_valid_3_0_a2_0_1 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.N_2138 ;
    wire \u1.PIO_control.iack_7_u_0_0_1_cascade_ ;
    wire \u1.PIO_control.iack_7_u_0_0_cascade_ ;
    wire \u1.PIO_control.pong_we ;
    wire \u1.PIO_control.ping_we ;
    wire \u1.PIO_control.N_1362 ;
    wire \u1.PIO_control.iack_7_u_0_a2_1_1 ;
    wire \u1.PIO_control.iack_7_u_0_a2_2_1 ;
    wire \u1.N_1359 ;
    wire \u1.PIO_control.rpp_2_i_0_cascade_ ;
    wire \u1.PIO_control.wpp ;
    wire \u1.PIO_control.pong_valid_3_0_a2_0 ;
    wire u1_PIO_control_gen_pingpong_pong_valid;
    wire \u1.PIO_control.dpong_valid ;
    wire \u1.DMAgoZ0 ;
    wire \u1.DMA_control.hgo_2_i_0_0 ;
    wire \u1.DMA_control.hgo ;
    wire \u1.DMA_control.gen_DMAbuf_Txbuf.N_319_g ;
    wire \u1.PIO_control.dping_valid_3 ;
    wire \u1.PIO_control.ping_d_15 ;
    wire \u1.PIO_control.ping_d_2 ;
    wire \u1.PIO_control.ping_d_3 ;
    wire \u1.PIO_control.ping_d_4 ;
    wire dd_pad_o_c_4;
    wire \u1.PIO_control.pong_d_5 ;
    wire \u1.PIO_control.ping_d_5 ;
    wire \u1.N_1430_cascade_ ;
    wire dd_pad_o_c_5;
    wire \u1.PIO_control.pong_d_6 ;
    wire \u1.PIO_control.ping_d_6 ;
    wire \u1.PIO_control.pong_d_8 ;
    wire \u1.PIO_control.ping_d_8 ;
    wire \u1.PIO_control.pong_d_7 ;
    wire \u1.PIO_control.ping_d_7 ;
    wire dd_pad_o_c_13;
    wire \u1.N_1431 ;
    wire dd_pad_o_c_6;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.val_c8_0_3 ;
    wire DMA_dmarq;
    wire \u1.c_state_RNIUC0A1Z0Z_1_cascade_ ;
    wire \u1.DMAtip_2_i_i_a2_0_1 ;
    wire \u1.DMAtip_2_i_i_a2_0_1_cascade_ ;
    wire dmackn_pad_o_c;
    wire \u1.N_2150 ;
    wire \u1.DMAtip_2_i_i_1 ;
    wire \u1.Tdone_i ;
    wire \u1.N_2150_cascade_ ;
    wire \u1.N_1874 ;
    wire \u1.DMA_control.Tm_0 ;
    wire DMAtip;
    wire u0_gen_bc_dec_store_pp_full;
    wire \u1.DMA_control.Td_2 ;
    wire \u1.DMA_control.Td_3 ;
    wire \u1.DMA_control.Td_4 ;
    wire \u1.DMA_control.Td_7 ;
    wire N_1369;
    wire u1_PIO_control_gen_pingpong_iack;
    wire \u0.N_1384_cascade_ ;
    wire \u0.ack_o_i_i_1_cascade_ ;
    wire N_410_i;
    wire N_1360;
    wire N_288_i;
    wire \u1.PIO_control.pong_d_10 ;
    wire \u1.DMA_control.Td_0 ;
    wire wb_we_i_c;
    wire wb_sel_i_c_3;
    wire N_1342;
    wire wb_sel_i_c_2;
    wire \u1.N_1435 ;
    wire dd_pad_o_c_10;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.N_2413_iZ0 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_s_7 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.QiZ0Z_7 ;
    wire \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qie_0_iZ0 ;
    wire \u1.DMA_control.TxbufQ_16 ;
    wire \u1.DMA_control.writeDlw_0 ;
    wire \u1.DMA_control.TxbufQ_17 ;
    wire \u1.DMA_control.writeDlw_1 ;
    wire \u1.DMA_control.TxbufQ_27 ;
    wire \u1.DMA_control.writeDlw_11 ;
    wire \u1.DMA_control.TxbufQ_28 ;
    wire \u1.DMA_control.writeDlw_12 ;
    wire \u1.DMA_control.TxbufQ_30 ;
    wire \u1.DMA_control.writeDlw_14 ;
    wire \u1.DMA_control.writeDfw_6_i_0_0 ;
    wire \u1.DMA_control.TxbufQ_8 ;
    wire \u1.DMA_control.dstrb ;
    wire \u1.DMA_control.writeDfw_6_i_0_1 ;
    wire \u1.DMA_control.TxbufQ_9 ;
    wire \u1.DMA_control.TxbufQ_2 ;
    wire \u1.DMAd_10 ;
    wire \u1.DMA_control.writeDfw_6_i_0_11 ;
    wire \u1.DMA_control.TxbufQ_3 ;
    wire \u1.DMA_control.TxbufQ_4 ;
    wire \u1.DMA_control.writeDfw_6_i_0_12 ;
    wire \u1.DMA_control.TxbufQ_5 ;
    wire \u1.DMAd_13 ;
    wire \u1.DMA_control.TxbufQ_6 ;
    wire \u1.DMA_control.writeDfw_6_i_m3_i_0_14 ;
    wire \u1.DMA_control.TxbufQ_21 ;
    wire \u1.DMA_control.writeDlw_5 ;
    wire \u1.DMA_control.writeDlw_6 ;
    wire \u1.DMA_control.TxbufQ_22 ;
    wire \u1.DMA_control.TxbufQ_14 ;
    wire \u1.DMA_control.writeDfw_6_i_0_6_cascade_ ;
    wire \u1.DMAd_6 ;
    wire \u1.DMA_control.writeDlw_7 ;
    wire \u1.DMA_control.TxbufQ_23 ;
    wire \u1.DMA_control.TxbufQ_15 ;
    wire \u1.DMA_control.writeDfw_6_i_0_7_cascade_ ;
    wire \u1.DMA_control.writeDlw_8 ;
    wire \u1.DMA_control.TxbufQ_24 ;
    wire \u1.DMA_control.TxbufQ_0 ;
    wire \u1.DMA_control.writeDfw_6_i_0_8_cascade_ ;
    wire \u1.DMA_control.TxbufQ_13 ;
    wire \u1.DMA_control.writeDfw_6_i_0_5 ;
    wire \u1.DMAd_5 ;
    wire \u1.PIO_control.pong_d_11 ;
    wire \u1.DMAd_11 ;
    wire \u1.N_1448_cascade_ ;
    wire dd_pad_o_c_11;
    wire \u1.PIO_control.pong_d_12 ;
    wire \u1.PIO_control.ping_d_12 ;
    wire \u1.PIO_control.pong_d_14 ;
    wire \u1.PIO_control.ping_d_14 ;
    wire \u1.PIO_control.pong_d_13 ;
    wire \u1.PIO_control.ping_d_13 ;
    wire \u1.N_1446 ;
    wire \u1.DMAd_12 ;
    wire \u1.N_1447 ;
    wire dd_pad_o_c_12;
    wire \u1.N_1445 ;
    wire \u1.DMAd_14 ;
    wire dd_pad_o_c_14;
    wire \u1.DMAd_8 ;
    wire \u1.N_1433 ;
    wire dd_pad_o_c_8;
    wire \u1.DMAd_7 ;
    wire \u1.N_1432 ;
    wire dd_pad_o_c_7;
    wire \u0.N_1384 ;
    wire wb_sel_i_c_1;
    wire \u0.un1_piosel ;
    wire wb_sel_i_c_0;
    wire N_284_i;
    wire bfn_7_17_0_;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.QiZ0Z_1 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_s_1 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_cry_0 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.QiZ0Z_2 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_s_2 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_cry_1 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.QiZ0Z_3 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_s_3 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_cry_2 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.QiZ0Z_4 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_s_4 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_cry_3 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.QiZ0Z_5 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_s_5 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_cry_4 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.QiZ0Z_6 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_s_6 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_cry_5 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_cry_6 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.N_1371 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.rci_0 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.T1done_i ;
    wire \u1.PIO_control.dsel_3_0_a2_0 ;
    wire \u1.PIO_control.N_2409 ;
    wire \u1.PIO_control.dsel ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.un1_ena_i_0_o3_sx_cascade_ ;
    wire N_1364;
    wire PIOq_10;
    wire N_1364_cascade_;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.un1_ena_i_0_o3_0_cascade_ ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.un1_ena_i_0_a2_sx ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.N_2092 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.drd_ptr_2 ;
    wire \u1.DMA_control.N_1346 ;
    wire \u1.DMA_control.gen_DMAbuf_Txbuf.N_1341 ;
    wire DMA_dev0_Td_0;
    wire DMA_dev1_Tm_0;
    wire da_pad_o_c_1;
    wire resetn_pad_o_c;
    wire u1_PIO_control_gen_pingpong_ping_valid;
    wire \u1.PIO_control.dping_valid ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.iQ_fast_3 ;
    wire DMActrl_dir;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.N_1385_i_cascade_ ;
    wire \u1.DMA_control.N_1326 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.iQ_fast_2 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_18 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_19 ;
    wire \u1.DMA_control.gen_DMAbuf_Txbuf.N_1602 ;
    wire \u1.DMA_control.gen_DMAbuf_Txbuf.N_1602_cascade_ ;
    wire \u1.DMA_control.gen_DMAbuf_Txbuf.N_319 ;
    wire \u1.DMA_control.writeDlw_13 ;
    wire \u1.DMA_control.TxbufQ_29 ;
    wire \u1.DMA_control.writeDfw_6_i_m2_i_0_13 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_6 ;
    wire \u1.DMA_control.TxbufQ_26 ;
    wire \u1.DMA_control.writeDlw_10 ;
    wire \u1.DMA_control.writeDfw_6_i_0_10 ;
    wire \u1.DMA_control.Td_5 ;
    wire \u1.DMA_control.TxbufQ_25 ;
    wire \u1.DMA_control.writeDlw_9 ;
    wire \u1.DMA_control.TxbufQ_1 ;
    wire \u1.DMA_control.writeDfw_6_i_0_9_cascade_ ;
    wire \u1.DMAd_9 ;
    wire \u1.DMA_control.wr_ptr_0 ;
    wire \u1.DMA_control.RxWrZ0 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.wr_ptr_1 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.wr_ptr_2 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_21 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_5 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_3 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_19 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNIA9TNZ0Z_6 ;
    wire mem_mem_ram6__RNIQPOD1_6_cascade_;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_6 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_18 ;
    wire \u1.DMA_control.Tm_1 ;
    wire \u1.PIO_control.PIO_access_control.T1Z0Z_0 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.hT2doneZ0 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.val_c8 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.iordy_done_0 ;
    wire \u1.PIO_control.PIO_access_control.T1Z0Z_2 ;
    wire \u1.PIO_control.PIO_access_control.T1Z0Z_4 ;
    wire \u1.c_stateZ0Z_0 ;
    wire \u1.c_stateZ0Z_1 ;
    wire \u1.c_state_ns_i_i_i_a2_1_1 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.N_1073 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_s_7 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.QiZ0Z_7 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.N_1071 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.rciZ0 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNI9LFIZ0Z_1_cascade_ ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.Qi_RNI7F9K_0 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.val_c8_0_4_0 ;
    wire \u1.PIO_control.PIO_access_control.it1_1_iv_0_0_4 ;
    wire \u1.PIO_control.pong_a_RNI914A1_0_cascade_ ;
    wire \u1.PIO_control.ping_a_RNIQNVQ_0 ;
    wire \u1.PIO_control.pong_we_1_sqmuxa ;
    wire \u1.PIO_control.ping_d_10 ;
    wire \u1.PIO_control.ping_d_11 ;
    wire \u1.PIO_control.ping_we_0_sqmuxa ;
    wire DMA_dev0_Td_5;
    wire \u1.N_1423 ;
    wire \u1.PIO_control.un3_idone_0_a2_0 ;
    wire \u1.N_1429 ;
    wire \u1.PIO_control.SelDev_e_1_cascade_ ;
    wire DMActrl_DMAen;
    wire \u0.dat_o_0_0_2_15_cascade_ ;
    wire DMA_dev0_Td_7;
    wire \u0.dat_o_0_0_3_15 ;
    wire \u0.dat_o_0_0_5_15_cascade_ ;
    wire wb_dat_o_c_15;
    wire mem_mem_ram6__RNIAVA71_15_cascade_;
    wire \u0.N_2029 ;
    wire iQ_RNIQGDM1_2;
    wire PIOq_15;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIEL7KZ0Z_19 ;
    wire iQ_RNIA1EM1_2_cascade_;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIA1VQZ0Z_19 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNII9GTZ0Z_19 ;
    wire mem_mem_ram6__RNIMBB71_19;
    wire \u0.CtrlRegZ0Z_19 ;
    wire \u0.dat_o_i_0_2_19_cascade_ ;
    wire \u0.N_1724 ;
    wire N_327_i;
    wire dd_pad_i_c_12;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_20 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_21 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_22 ;
    wire \u1.DMA_control.TxbufQ_12 ;
    wire \u1.DMAd_4 ;
    wire \u1.DMA_control.TxbufQ_18 ;
    wire \u1.DMA_control.writeDlw_2 ;
    wire \u1.DMA_control.TxbufQ_10 ;
    wire \u1.DMA_control.writeDfw_6_i_0_2_cascade_ ;
    wire \u1.DMAd_2 ;
    wire \u1.DMA_control.TxbufQ_19 ;
    wire \u1.DMA_control.writeDlw_3 ;
    wire \u1.DMA_control.TxbufQ_11 ;
    wire \u1.DMA_control.writeDfw_6_i_0_3_cascade_ ;
    wire \u1.DMAd_3 ;
    wire \u1.DMA_control.TxbufQ_20 ;
    wire \u1.DMA_control.writeDlw_4 ;
    wire \u1.DMA_control.writeDfw_6_i_0_4 ;
    wire \u1.DMA_control.writeDlw_15 ;
    wire \u1.DMA_control.TxbufQ_31 ;
    wire \u1.DMA_control.TxbufQ_7 ;
    wire \u1.DMA_control.TxRdZ0 ;
    wire \u1.DMA_control.writeDfw_6_i_m3_i_0_15_cascade_ ;
    wire \u1.DMAd_15 ;
    wire \u1.DMA_control.N_53 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_20 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_21 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_3 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_5 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_6 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_22 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_22 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_31 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_15 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI6D7KZ0Z_15 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_4 ;
    wire \u0.dat_o_0_0_3_13 ;
    wire \u0.dat_o_0_0_0_13 ;
    wire \u0.dat_o_0_0_2_13 ;
    wire wb_dat_o_c_13;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.Qi_0_0 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_s_0 ;
    wire \u0.int_3_i_0_0 ;
    wire PIO_dport1_T1_0;
    wire \u1.PIO_control.PIO_access_control.it1_1_iv_i_i_0_0 ;
    wire \u1.PIO_control.PIO_access_control.iteoc_1_iv_0_0_6_cascade_ ;
    wire \u1.PIO_control.PIO_access_control.TeocZ0Z_6 ;
    wire \u1.PIO_control.PIO_access_control.T1Z0Z_5 ;
    wire \u1.PIO_control.PIO_access_control.TeocZ0Z_7 ;
    wire \u1.PIO_control.PIO_access_control.it1_1_iv_i_i_0_3_cascade_ ;
    wire \u1.PIO_control.PIO_access_control.T1Z0Z_3 ;
    wire \u1.PIO_control.PIO_access_control.it1_1_iv_0_0_2 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_s_0 ;
    wire \u1.PIO_control.PIO_access_control.N_2110_cascade_ ;
    wire \u1.PIO_control.PIO_access_control.it1_1_iv_i_i_0_5 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_1_sqmuxa_i ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qie_0_iZ0 ;
    wire \u1.pong_a_0 ;
    wire \u1.ping_a_0 ;
    wire da_pad_o_c_0;
    wire \u1.PIO_control.N_1450 ;
    wire \u1.PIO_control.rpp_2_i_0 ;
    wire \u1.PIOdone_i ;
    wire \u1.PIO_control.ping_a_1 ;
    wire \u1.pong_a_2 ;
    wire \u1.ping_a_2 ;
    wire \u1.PIO_control.pong_a_1 ;
    wire \u1.PIO_control.PIO_access_control.it4_1_iv_i_i_o2_0_x0Z0Z_2_cascade_ ;
    wire \u1.PIO_control.PIO_access_control.it4_1_iv_i_i_o2_0_x1Z0Z_2 ;
    wire \u1.PIO_control.PIO_access_control.it4_1_iv_i_i_o2_0_2_cascade_ ;
    wire \u1.PIO_control.PIO_access_control.it4_1_iv_i_i_o3_x0Z0Z_2_cascade_ ;
    wire \u1.PIO_control.PIO_access_control.iiordyen_1_iv_i_i_0_cascade_ ;
    wire \u1.PIO_control.PIO_access_control.IORDYenZ0 ;
    wire \u1.PIO_control.PIO_access_control.it1_1_iv_i_i_0_1_cascade_ ;
    wire \u1.PIO_control.PIO_access_control.T1Z0Z_1 ;
    wire \u1.DMA_control.Td_1 ;
    wire \u1.PIO_control.PIO_access_control.it4_1_iv_i_i_o2_0_2 ;
    wire \u1.PIO_control.N_1315 ;
    wire \u1.PIO_control.PIO_access_control.N_2112_cascade_ ;
    wire \u1.PIO_control.PIO_access_control.iteoc_1_iv_i_i_0_7 ;
    wire \u1.PIO_control.PIO_access_control.it4_1_iv_i_i_0_2_cascade_ ;
    wire \u1.PIO_control.PIO_access_control.T4Z0Z_2 ;
    wire \u1.PIO_control.PIO_access_control.it4_1_iv_i_i_0_3_cascade_ ;
    wire \u1.PIO_control.PIO_access_control.T4Z0Z_3 ;
    wire \u1.PIO_control.PIO_access_control.it4_1_iv_0_0_4_cascade_ ;
    wire \u1.PIO_control.PIO_access_control.T4Z0Z_4 ;
    wire \u1.PIO_control.PIO_access_control.it4_1_iv_i_i_0_5_cascade_ ;
    wire \u1.PIO_control.PIO_access_control.T4Z0Z_5 ;
    wire \u1.DMAd_0 ;
    wire dd_pad_o_c_0;
    wire \u1.PIO_control.pong_a_3 ;
    wire \u1.PIO_control.ping_a_3 ;
    wire \u1.N_1425_cascade_ ;
    wire cs0n_pad_o_c;
    wire \u1.PIO_control.pong_d_0 ;
    wire \u1.PIO_control.ping_d_0 ;
    wire \u1.N_1426 ;
    wire \u1.rpp ;
    wire \u1.PIO_control.ping_d_1 ;
    wire \u1.PIO_control.pong_d_1 ;
    wire \u1.N_1427_cascade_ ;
    wire \u1.DMAd_1 ;
    wire dd_pad_o_c_1;
    wire \u1.N_1425 ;
    wire cs1n_pad_o_c;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_15 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_31 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI61KTZ0Z_31_cascade_ ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_31 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI2DBKZ0Z_31 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI4VG71Z0Z_31 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIIGLM1Z0Z_2_cascade_ ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_2 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_3 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_19 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_12 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_14 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_14 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_15 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIA1GTZ0Z_15 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_15 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_31 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_17 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_2 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_12 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_3 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_19 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_19 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_17 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_19 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_22 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_21 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_24 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_8 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_8 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_16 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_16 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_0 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_24 ;
    wire \u1.PIO_control.PIO_access_control.it1_1_iv_i_i_0_6_cascade_ ;
    wire \u1.PIO_control.PIO_access_control.T1Z0Z_6 ;
    wire PIO_dport1_T2_4;
    wire \u1.PIO_control.PIO_access_control.T2Z0Z_4 ;
    wire \u1.PIO_control.PIO_access_control.T1Z0Z_7 ;
    wire \u1.PIO_control.PIO_access_control.it2_1_iv_0_0_0_cascade_ ;
    wire \u1.PIO_control.PIO_access_control.T2Z0Z_0 ;
    wire \u1.PIO_control.PIO_access_control.it2_1_iv_i_i_0_1_cascade_ ;
    wire \u1.PIO_control.PIO_access_control.T2Z0Z_1 ;
    wire \u1.PIO_control.PIO_access_control.it2_1_iv_0_0_2_cascade_ ;
    wire \u1.PIO_control.PIO_access_control.T2Z0Z_2 ;
    wire \u1.PIO_control.PIO_access_control.it2_1_iv_i_i_0_3_cascade_ ;
    wire PIO_dport0_T2_3;
    wire \u1.PIO_control.PIO_access_control.T2Z0Z_3 ;
    wire \u1.PIO_control.PIO_access_control.it2_1_iv_0_0_4 ;
    wire \u1.PIO_control.PIO_access_control.it1_1_iv_i_i_0_7 ;
    wire \u1.PIO_control.PIO_access_control.it2_1_iv_0_0_5_cascade_ ;
    wire \u1.PIO_control.PIO_access_control.T2Z0Z_5 ;
    wire \u1.PIO_control.PIO_access_control.it2_1_iv_i_i_0_6_cascade_ ;
    wire \u1.PIO_control.PIO_access_control.T2Z0Z_6 ;
    wire \u1.PIO_control.PIO_access_control.it2_1_iv_i_i_0_7_cascade_ ;
    wire \u1.PIO_control.PIO_access_control.T2Z0Z_7 ;
    wire \u1.PIO_control.PIO_access_control.it4_1_iv_0_0_0_cascade_ ;
    wire \u1.PIO_control.PIO_access_control.T4Z0Z_0 ;
    wire \u1.PIO_control.PIO_access_control.TeocZ0Z_2 ;
    wire \u1.PIO_control.PIO_access_control.it4_1_iv_i_i_0_7_cascade_ ;
    wire \u1.PIO_control.PIO_access_control.T4Z0Z_7 ;
    wire \u1.PIO_control.PIO_access_control.iteoc_1_iv_i_i_0_5_cascade_ ;
    wire \u1.PIO_control.PIO_access_control.TeocZ0Z_5 ;
    wire \u1.PIO_control.PIO_access_control.iteoc_1_iv_i_i_0_2 ;
    wire \u1.DMA_control.Teoc_3 ;
    wire PIO_cmdport_T1_2;
    wire PIO_dport0_IORDYen;
    wire PIO_cmdport_T1_3;
    wire PIO_dport1_IORDYen;
    wire PIO_cmdport_T1_4;
    wire IDEctrl_ppen;
    wire IDEctrl_FATR0;
    wire PIO_cmdport_T1_1;
    wire \u0.CtrlRegZ0Z_20 ;
    wire \u0.dat_o_0_a2_i_2_20_cascade_ ;
    wire N_211_i;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIQI0RZ0Z_20_cascade_ ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.N_1386_i ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI2RHTZ0Z_20 ;
    wire iQ_RNIA4HM1_2;
    wire mem_mem_ram6__RNIULD71_20_cascade_;
    wire \u0.N_1559 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIEDOD1Z0Z_2_cascade_ ;
    wire DMAq_2_cascade_;
    wire \u0.dat_o_0_0_0_2 ;
    wire \u0.dat_o_0_0_1Z0Z_2_cascade_ ;
    wire \u0.dat_o_0_0_2_2 ;
    wire wb_dat_o_c_2;
    wire PIOq_2;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIQ0CMZ0Z_2 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIASNK1Z0Z_2 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI2PUQZ0Z_15 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_15 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_31 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_31 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIUO2RZ0Z_31 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_24 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_24 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_8 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_20 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_15 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_8 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_2 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_19 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_20 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_15 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_31 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_awe3 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_4 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_0 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_30 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_30 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_30 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI4VJTZ0Z_30_cascade_ ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_30 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_30 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNISM2RZ0Z_30 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI0BBKZ0Z_30_cascade_ ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_30 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_awe5 ;
    wire PIO_dport0_T2_4;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.QiZ0Z_0 ;
    wire bfn_12_18_0_;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.QiZ0Z_1 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_s_1 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_cry_0 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.QiZ0Z_2 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_s_2 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_cry_1 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.QiZ0Z_3 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_s_3 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_cry_2 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.QiZ0Z_4 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_s_4 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_cry_3 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.QiZ0Z_5 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_s_5 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_cry_4 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.QiZ0Z_6 ;
    wire CONSTANT_ONE_NET;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_s_6 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_cry_5 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.QiZ0Z_7 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_cry_6 ;
    wire \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_s_7 ;
    wire \u1.PIO_control.PIO_access_control.iteoc_1_iv_i_i_0_1 ;
    wire \u1.PIO_control.PIO_access_control.TeocZ0Z_1 ;
    wire \u1.PIO_control.PIO_access_control.it4_1_iv_0_0_1_cascade_ ;
    wire \u1.PIO_control.PIO_access_control.T4Z0Z_1 ;
    wire \u1.PIO_control.PIO_access_control.iteoc_1_iv_i_i_0_3 ;
    wire \u1.PIO_control.PIO_access_control.TeocZ0Z_3 ;
    wire \u1.PIO_control.PIO_access_control.N_1319 ;
    wire \u1.PIO_control.PIO_access_control.N_2112 ;
    wire \u1.PIO_control.PIO_access_control.iteoc_1_iv_i_i_0_4_cascade_ ;
    wire \u1.PIO_control.PIO_access_control.TeocZ0Z_4 ;
    wire \u1.PIO_control.PIO_access_control.it4_1_iv_i_i_0_6 ;
    wire \u1.PIO_control.PIO_access_control.T4Z0Z_6 ;
    wire \u1.PIO_control.PIO_access_control.N_2110 ;
    wire \u1.PIO_control.PIO_access_control.iteoc_1_iv_i_i_0_0 ;
    wire \u1.PIO_control.PIO_access_control.TeocZ0Z_0 ;
    wire PIO_cmdport_T2_5;
    wire PIO_cmdport_T2_7;
    wire PIO_cmdport_T4_3;
    wire PIO_cmdport_T4_4;
    wire \u0.dat_o_0_0_3_12 ;
    wire \u0.dat_o_0_0_2_12_cascade_ ;
    wire wb_dat_o_c_12;
    wire \u0.CtrlRegZ0Z_12 ;
    wire DMA_dev0_Td_4;
    wire \u0.dat_o_0_0_0_12 ;
    wire DMAq_12_cascade_;
    wire PIOq_12;
    wire \u0.dat_o_0_0_1Z0Z_12 ;
    wire \u0.dat_o_0_0_1Z0Z_4_cascade_ ;
    wire \u0.dat_o_0_0_2_4 ;
    wire wb_dat_o_c_4;
    wire PIO_dport1_T1_4;
    wire \u0.dat_o_0_0_0_4 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI2L4NZ0Z_4 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNII4OK1Z0Z_2_cascade_ ;
    wire DMAq_4;
    wire dd_pad_i_c_4;
    wire PIOq_4;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_4 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIKJOD1Z0Z_4 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_4 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIU4CMZ0Z_4 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_4 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_12 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_12 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI4RFTZ0Z_12_cascade_ ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI1MA71Z0Z_12 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_20 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_12 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_12 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI077KZ0Z_12_cascade_ ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNISIUQZ0Z_12 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIE4DM1Z0Z_2 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_14 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI8VFTZ0Z_14 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_2 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIUG4NZ0Z_2 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_2 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_1 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_1 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_2 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_2 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNI21TNZ0Z_2 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_3 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_3 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_4 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_4 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNI65TNZ0Z_4 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_5 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_5 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_7 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_7 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_17 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_17 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_1 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_1 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_18 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_18 ;
    wire \u1.DMA_control.readDlw_2 ;
    wire \u1.DMA_control.readDfw_2 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_14 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI4B7KZ0Z_14_cascade_ ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_14 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_30 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_26 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_26 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIE7ITZ0Z_26_cascade_ ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIG8E71Z0Z_26_cascade_ ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_23 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_23 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_9 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_9 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_11 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_11 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_20 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIU69KZ0Z_20 ;
    wire \u1.DMA_control.readDlw_4 ;
    wire \u1.DMA_control.readDfw_4 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_20 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_awe2 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_7 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_7 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_26 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_26 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_26 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIAJ9KZ0Z_26 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI6V0RZ0Z_26_cascade_ ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI2THM1Z0Z_2 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_28 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIA31RZ0Z_28_cascade_ ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_28 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_28 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_N_1197_cascade_ ;
    wire u1_DMA_control_gen_DMAbuf_Rxbuf_mem_N_1229_cascade_;
    wire u1_DMA_control_gen_DMAbuf_Rxbuf_mem_N_1165;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_28 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_28 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIEN9KZ0Z_28 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_28 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_12 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_6 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_6 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI6P4NZ0Z_6_cascade_ ;
    wire iQ_RNIQCOK1_2;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_6 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI29CMZ0Z_6 ;
    wire DMA_dev0_Tm_2;
    wire PIO_cmdport_T1_5;
    wire \u0.dat_o_0_0_0_8 ;
    wire \u0.dat_o_0_0_3_8 ;
    wire DMATxFull;
    wire PIO_dport1_T2_1;
    wire DMA_dev1_Td_7;
    wire \u0.dat_o_0_0_0_15 ;
    wire DMA_dev1_Td_0;
    wire DMA_dev1_Td_1;
    wire DMA_dev1_Td_3;
    wire DMA_dev1_Td_4;
    wire DMA_dev1_Td_5;
    wire PIO_dport1_T2_5;
    wire PIO_dport1_T2_7;
    wire DMA_dev1_Tm_1;
    wire PIO_dport0_T1_1;
    wire PIO_dport0_T1_2;
    wire DMA_dev1_Tm_2;
    wire \u0.dat_o_0_0_3_2 ;
    wire PIO_dport0_T1_3;
    wire \u1.DMA_control.Td_6 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNI87TNZ0Z_5 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_5 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI4N4NZ0Z_5 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNINMOD1Z0Z_5 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIM8OK1Z0Z_2_cascade_ ;
    wire DMAq_5_cascade_;
    wire \u0.dat_o_0_2_5 ;
    wire \u0.dat_o_0_1Z0Z_5_cascade_ ;
    wire \u0.dat_o_0_3_5 ;
    wire wb_dat_o_c_5;
    wire PIO_dport1_T1_5;
    wire \u0.dat_o_0_0_5 ;
    wire dd_pad_i_c_5;
    wire PIOq_5;
    wire \u1.DMA_control.Tm_3 ;
    wire \u1.DMA_control.Tm_4 ;
    wire \u1.DMA_control.Tm_5 ;
    wire \u1.DMA_control.Tm_6 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_5 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI07CMZ0Z_5 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_14 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_14 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI0NUQZ0Z_14 ;
    wire \u1.DMA_control.readDlw_12 ;
    wire \u1.DMA_control.readDfw_12 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_28 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_5 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_6 ;
    wire \u1.DMA_control.readDlw_14 ;
    wire \u1.DMA_control.readDfw_14 ;
    wire dd_pad_i_c_14;
    wire \u1.DMA_control.readDlw_6 ;
    wire \u1.DMA_control.readDfw_6 ;
    wire \u1.DMA_control.readDlw_15 ;
    wire \u1.DMA_control.readDfw_15 ;
    wire dd_pad_i_c_15;
    wire dd_pad_i_c_2;
    wire dd_pad_i_c_10;
    wire dd_pad_i_c_11;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_26 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_awe1 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_29 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_29 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_29 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_29 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIKDITZ0Z_29_cascade_ ;
    wire mem_mem_ram6__RNIPHE71_29_cascade_;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_29 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_29 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIGP9KZ0Z_29 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIC51RZ0Z_29_cascade_ ;
    wire iQ_RNIE9IM1_2;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_29 ;
    wire \u1.DMA_control.readDlw_13 ;
    wire \u1.DMA_control.readDfw_13 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_25 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_25 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_25 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI4T0RZ0Z_25 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI8H9KZ0Z_25_cascade_ ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_10 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_10 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_10 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_10 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIOEUQZ0Z_10 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIS27KZ0Z_10_cascade_ ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_10 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_10 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI0NFTZ0Z_10_cascade_ ;
    wire iQ_RNI6SCM1_2;
    wire mem_mem_ram6__RNIRFA71_10_cascade_;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_10 ;
    wire \u1.DMA_control.readDlw_10 ;
    wire \u1.DMA_control.readDfw_10 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_26 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_13 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_13 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI6TFTZ0Z_13_cascade_ ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_13 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI4PA71Z0Z_13_cascade_ ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_13 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_13 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI297KZ0Z_13_cascade_ ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNII8DM1Z0Z_2 ;
    wire DMAq_13;
    wire \u0.dat_o_0_0_1Z0Z_13 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_13 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_13 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIUKUQZ0Z_13 ;
    wire dd_pad_i_c_13;
    wire PIOq_13;
    wire PIO_cmdport_T2_1;
    wire PIO_cmdport_T2_0;
    wire PIO_dport1_T2_0;
    wire wb_dat_i_c_2;
    wire PIO_dport1_T1_2;
    wire wb_dat_i_c_13;
    wire PIO_dport0_T2_5;
    wire wb_dat_i_c_15;
    wire PIO_dport1_T4_3;
    wire \u0.dat_o_i_0_0_19 ;
    wire \u0.dat_o_0_0_3_4 ;
    wire PIO_dport0_T2_7;
    wire \u0.N_2033 ;
    wire wb_dat_i_c_19;
    wire PIO_dport0_T4_3;
    wire wb_dat_i_c_20;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIS2CMZ0Z_3 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI0J4NZ0Z_3 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIE0OK1Z0Z_2_cascade_ ;
    wire DMAq_3_cascade_;
    wire PIO_dport1_T1_3;
    wire \u0.dat_o_0_0_2_3 ;
    wire \u0.dat_o_0_0_3_3 ;
    wire \u0.dat_o_0_0_0_3_cascade_ ;
    wire \u0.dat_o_0_0_1Z0Z_3 ;
    wire wb_dat_o_c_3;
    wire dd_pad_i_c_3;
    wire PIOq_3;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_3 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNI43TNZ0Z_3 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIHGOD1Z0Z_3 ;
    wire DMA_dev0_Tm_3;
    wire DMA_dev0_Tm_4;
    wire DMA_dev0_Tm_5;
    wire PIO_cmdport_T4_2;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIG7GTZ0Z_18 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_18 ;
    wire mem_mem_ram6__RNIJ8B71_18_cascade_;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_18 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_18 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNICJ7KZ0Z_18 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI8VUQZ0Z_18_cascade_ ;
    wire iQ_RNI6TDM1_2;
    wire wb_dat_i_c_18;
    wire \u0.CtrlRegZ0Z_18 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI2R0RZ0Z_24 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI6F9KZ0Z_24 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_24 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIA3ITZ0Z_24_cascade_ ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_24 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIQKHM1Z0Z_2 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIA2E71Z0Z_24_cascade_ ;
    wire \u1.DMA_control.readDlw_5 ;
    wire \u1.DMA_control.readDfw_5 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_9 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_9 ;
    wire \u1.DMA_control.readDlw_9 ;
    wire \u1.DMA_control.readDfw_9 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_25 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_0 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_0 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_1 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_1 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_27 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_27 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_27 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI811RZ0Z_27 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNICL9KZ0Z_27_cascade_ ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI61IM1Z0Z_2_cascade_ ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_27 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_awe0 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_11 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_11 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIQGUQZ0Z_11_cascade_ ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIU47KZ0Z_11 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_16 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_16 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_11 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_11 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_27 ;
    wire \u1.DMA_control.readDlw_3 ;
    wire \u1.DMA_control.readDfw_3 ;
    wire \u1.DMA_control.rd_dstrb_g ;
    wire \u1.SelDev ;
    wire \u1.DMA_control.Tm_7 ;
    wire PIO_dport1_T1_7;
    wire PIO_dport0_T1_4;
    wire PIO_dport0_T2_0;
    wire wb_dat_i_c_9;
    wire wb_dat_i_c_12;
    wire PIO_cmdport_T2_4;
    wire DMA_dev1_Teoc_4;
    wire PIO_cmdport_Teoc_4;
    wire PIO_cmdport_T1_7;
    wire PIOtip;
    wire PIO_dport0_T1_7;
    wire \u0.dat_o_0_0_0_7 ;
    wire \u0.dat_o_0_0_3_7_cascade_ ;
    wire PIO_cmdport_T1_0;
    wire \u0.dat_o_0_0_0_0 ;
    wire \u0.dat_o_0_0_3_0_cascade_ ;
    wire wb_inta_o_c;
    wire PIO_dport0_T4_0;
    wire PIO_dport1_T4_0;
    wire PIO_dport1_T4_2;
    wire PIO_dport0_T4_2;
    wire PIO_dport1_T4_4;
    wire PIO_dport0_T4_4;
    wire \u0.dat_o_0_a2_i_0_20 ;
    wire PIO_dport1_T4_5;
    wire PIO_dport0_T4_5;
    wire PIO_dport1_T4_6;
    wire PIO_dport0_T4_6;
    wire wb_dat_i_c_3;
    wire DMA_dev1_Tm_3;
    wire wb_dat_i_c_4;
    wire DMA_dev1_Tm_4;
    wire DMA_dev1_Tm_5;
    wire PIO_cmdport_Teoc_3;
    wire \u0.dat_o_i_i_1_27_cascade_ ;
    wire PIO_dport0_Teoc_3;
    wire \u0.dat_o_i_i_4_27_cascade_ ;
    wire DMA_dev1_Teoc_3;
    wire N_269;
    wire wb_dat_i_c_27;
    wire \u0.CtrlRegZ0Z_27 ;
    wire PIO_dport1_Teoc_3;
    wire \u0.N_1682 ;
    wire DMA_dev0_Teoc_3;
    wire DMAq_27;
    wire \u0.dat_o_i_i_0_27 ;
    wire \u0.N_1636_cascade_ ;
    wire \u0.dat_o_i_0_21 ;
    wire N_259_i;
    wire wb_dat_i_c_21;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_21 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_21 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNISK0RZ0Z_21_cascade_ ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI099KZ0Z_21 ;
    wire iQ_RNIE8HM1_2;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI4THTZ0Z_21 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_21 ;
    wire mem_mem_ram6__RNI1PD71_21;
    wire \u0.CtrlRegZ0Z_21 ;
    wire PIO_cmdport_T4_5;
    wire \u0.dat_o_i_2_21 ;
    wire \u0.dat_o_0_0_6_7 ;
    wire \u0.N_1979_cascade_ ;
    wire wb_dat_o_c_7;
    wire dd_pad_i_c_7;
    wire PIOq_7;
    wire IDEctrl_IDEen;
    wire \u0.dat_o_0_0_2_7 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI8R4NZ0Z_7 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI4BCMZ0Z_7 ;
    wire iQ_RNIUGOK1_2;
    wire \u0.N_1980 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_7 ;
    wire mem_mem_ram6__RNITSOD1_7;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI6VHTZ0Z_22 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_22 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_22 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_22 ;
    wire wb_dat_i_c_22;
    wire \u0.CtrlRegZ0Z_22 ;
    wire PIO_cmdport_T4_6;
    wire \u0.dat_o_i_0_2_22_cascade_ ;
    wire \u0.dat_o_i_0_0_22 ;
    wire N_330_i;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_7 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNICBTNZ0Z_7 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_7 ;
    wire \u1.DMA_control.readDlw_7 ;
    wire \u1.DMA_control.readDfw_7 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_8 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_8 ;
    wire \u1.DMA_control.readDfw_8 ;
    wire \u1.DMA_control.readDlw_8 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_24 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_23 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_23 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_23 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI81ITZ0Z_23 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_9 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_9 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNIGFTNZ0Z_9_cascade_ ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_9 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_0 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_0 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIUOHM1Z0Z_2 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI4D9KZ0Z_23 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_23 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_23 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI0P0RZ0Z_23 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_25 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_25 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIC5ITZ0Z_25_cascade_ ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_25 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNID5E71Z0Z_25 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI2PFTZ0Z_11 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIUIA71Z0Z_11_cascade_ ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIA0DM1Z0Z_2 ;
    wire DMA_dev0_Tm_7;
    wire \u0.N_444 ;
    wire wb_dat_i_c_7;
    wire DMA_dev1_Tm_7;
    wire \u0.N_442 ;
    wire wb_dat_i_c_6;
    wire wb_dat_i_c_1;
    wire PIO_cmdport_IORDYen;
    wire \u0.N_446 ;
    wire PIO_cmdport_T2_2;
    wire \u0.dat_o_i_i_3_10_cascade_ ;
    wire PIO_dport0_T2_2;
    wire wb_dat_i_c_10;
    wire \u0.CtrlRegZ0Z_10 ;
    wire DMA_dev0_Td_2;
    wire \u0.N_1989 ;
    wire \u0.dat_o_i_i_2Z0Z_10 ;
    wire \u0.N_1990_cascade_ ;
    wire \u0.dat_o_i_i_6_10 ;
    wire N_1097;
    wire PIO_dport1_Teoc_0;
    wire \u0.N_1661_cascade_ ;
    wire PIO_dport0_Teoc_0;
    wire PIO_cmdport_Teoc_0;
    wire \u0.dat_o_i_i_1_24 ;
    wire wb_dat_i_c_24;
    wire \u0.CtrlRegZ0Z_24 ;
    wire wb_dat_i_c_31;
    wire DMAq_31;
    wire DMA_dev0_Teoc_7;
    wire \u0.dat_o_i_i_0_31_cascade_ ;
    wire DMA_dev1_Teoc_7;
    wire N_277;
    wire PIO_dport1_Teoc_7;
    wire \u0.CtrlRegZ0Z_31 ;
    wire PIO_cmdport_Teoc_7;
    wire \u0.N_1710 ;
    wire \u0.dat_o_i_i_1_31_cascade_ ;
    wire PIO_dport0_Teoc_7;
    wire \u0.dat_o_i_i_4_31 ;
    wire PIO_cmdport_Teoc_1;
    wire \u0.dat_o_i_i_1_25_cascade_ ;
    wire PIO_dport0_Teoc_1;
    wire PIO_dport1_Teoc_1;
    wire \u0.N_1668 ;
    wire wb_dat_i_c_25;
    wire \u0.CtrlRegZ0Z_25 ;
    wire DMAq_25;
    wire DMA_dev0_Teoc_1;
    wire DMA_dev0_Tm_6;
    wire PIO_dport1_T1_6;
    wire \u0.dat_o_0_0_0_6_cascade_ ;
    wire DMA_dev1_Tm_6;
    wire dd_pad_i_c_6;
    wire PIOq_6;
    wire \u0.N_1969 ;
    wire IDEctrl_FATR1;
    wire PIO_cmdport_T1_6;
    wire PIO_dport0_T1_6;
    wire \u0.dat_o_0_0_3_6 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNIEDTNZ0Z_8 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_8 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNI0VSNZ0Z_1 ;
    wire \u0.N_1971 ;
    wire \u0.N_1970 ;
    wire \u0.dat_o_0_0_6_6 ;
    wire \u0.dat_o_0_0_2_6 ;
    wire wb_dat_o_c_6;
    wire PIO_cmdport_T4_0;
    wire wb_dat_i_c_16;
    wire \u0.CtrlRegZ0Z_16 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_16 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_16 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIUM0RZ0Z_22 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI2B9KZ0Z_22 ;
    wire mem_mem_ram6__RNI4SD71_22;
    wire iQ_RNIICHM1_2_cascade_;
    wire \u0.N_1719 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI8F7KZ0Z_16 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI4RUQZ0Z_16 ;
    wire \u1.DMA_control.readDlw_0 ;
    wire \u1.DMA_control.readDfw_0 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_1 ;
    wire \u1.DMA_control.readDlw_1 ;
    wire \u1.DMA_control.readDfw_1 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_11 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_awe6 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIG9ITZ0Z_27 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_27 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIJBE71Z0Z_27 ;
    wire DMA_dev0_Tm_0;
    wire \u0.dat_o_0_0_6_0 ;
    wire \u0.N_1938_cascade_ ;
    wire wb_dat_o_c_0;
    wire dd_pad_i_c_0;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIMSBMZ0Z_0 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIQC4NZ0Z_0 ;
    wire iQ_RNI2KNK1_2_cascade_;
    wire \u0.N_1937 ;
    wire PIOq_0;
    wire IDEctrl_rst;
    wire \u0.dat_o_0_0_2_0 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_0 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNIUSSNZ0Z_0 ;
    wire mem_mem_ram6__RNI87OD1_0;
    wire \u1.DMA_control.readDfw_11 ;
    wire \u1.DMA_control.readDlw_11 ;
    wire \u1.DMA_control.N_1313 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_27 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_awe4 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI1SG71Z0Z_30 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIECLM1Z0Z_2 ;
    wire N_448;
    wire PIO_dport1_T2_3;
    wire DMA_dev0_Td_3;
    wire \u0.dat_o_0_0_0_11_cascade_ ;
    wire \u0.dat_o_0_0_3_11 ;
    wire wb_dat_o_c_11;
    wire wb_dat_i_c_11;
    wire \u0.CtrlRegZ0Z_11 ;
    wire PIO_cmdport_T2_3;
    wire \u0.dat_o_0_0_2_11 ;
    wire DMA_dev1_Td_2;
    wire PIO_dport1_T2_2;
    wire \u0.dat_o_i_i_0_10 ;
    wire PIO_dport0_T2_6;
    wire DMA_dev1_Td_6;
    wire \u0.dat_o_0_0_3_14_cascade_ ;
    wire wb_dat_o_c_14;
    wire PIOq_14;
    wire \u0.dat_o_0_0_1Z0Z_14 ;
    wire DMA_dev0_Td_6;
    wire PIO_dport1_T2_6;
    wire \u0.dat_o_0_0_0_14 ;
    wire wb_dat_i_c_14;
    wire \u0.CtrlRegZ0Z_14 ;
    wire PIO_cmdport_T2_6;
    wire \u0.dat_o_0_0_2_14 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI7SA71Z0Z_14 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIMCDM1Z0Z_2 ;
    wire DMAq_14;
    wire DMA_dev1_Teoc_5;
    wire DMA_dev0_Teoc_5;
    wire \u0.dat_o_i_i_0_29 ;
    wire PIO_dport0_Teoc_5;
    wire \u0.dat_o_i_i_a2_0_0_29_cascade_ ;
    wire PIO_dport1_Teoc_5;
    wire \u0.N_1696 ;
    wire \u0.dat_o_i_i_4_29 ;
    wire \u0.dat_o_i_i_2_29_cascade_ ;
    wire N_273;
    wire DMA_dev1_Teoc_2;
    wire \u0.N_1675_cascade_ ;
    wire PIO_dport0_Teoc_2;
    wire \u0.dat_o_i_i_4_26_cascade_ ;
    wire PIO_dport1_Teoc_2;
    wire N_267;
    wire wb_dat_i_c_26;
    wire DMAq_26;
    wire DMA_dev0_Teoc_2;
    wire \u0.dat_o_i_i_0_26 ;
    wire DMA_dev0_Tm_1;
    wire PIO_dport1_T1_1;
    wire \u0.dat_o_0_0_2_1 ;
    wire \u0.dat_o_0_0_3_1 ;
    wire \u0.dat_o_0_0_0_1_cascade_ ;
    wire wb_dat_o_c_1;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNISE4NZ0Z_1 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIOUBMZ0Z_1 ;
    wire dd_pad_i_c_1;
    wire \u0.N_1736 ;
    wire \u0.dat_o_0_0_6_8 ;
    wire \u0.dat_o_0_0_2_8_cascade_ ;
    wire wb_dat_o_c_8;
    wire dd_pad_i_c_8;
    wire PIOq_8;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI6DCMZ0Z_8 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIAT4NZ0Z_8 ;
    wire mem_mem_ram6__RNI00PD1_8;
    wire iQ_RNI2LOK1_2_cascade_;
    wire \u0.N_1735 ;
    wire dd_pad_i_c_9;
    wire \u1.PIO_control.PIO_access_control.dstrb ;
    wire PIO_cmdport_T4_1;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_17 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_17 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_0 ;
    wire wb_dat_i_c_17;
    wire \u0.CtrlRegZ0Z_17 ;
    wire \u0.N_2101 ;
    wire PIO_cmdport_T4_7;
    wire \u0.N_2142 ;
    wire wb_dat_i_c_23;
    wire \u0.CtrlRegZ0Z_23 ;
    wire u1_DMA_control_gen_DMAbuf_Rxbuf_mem_N_1224;
    wire u1_DMA_control_gen_DMAbuf_Rxbuf_mem_N_1160;
    wire DMActrl_BeLeC1;
    wire PIOq_9;
    wire DMAq_11;
    wire PIOq_11;
    wire \u0.dat_o_0_0_1Z0Z_11 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNICV4NZ0Z_9 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI8FCMZ0Z_9 ;
    wire mem_mem_ram6__RNI33PD1_9;
    wire iQ_RNI6POK1_2_cascade_;
    wire wb_dat_i_c_5;
    wire PIO_dport0_T1_5;
    wire wb_dat_i_c_28;
    wire \u0.N_1695 ;
    wire \u0.dat_o_0_0_0_9 ;
    wire \u0.dat_o_0_0_3_9 ;
    wire PIO_dport0_T2_1;
    wire \u0.CtrlRegZ0Z_28 ;
    wire PIO_dport0_Teoc_4;
    wire \u0.N_1688_cascade_ ;
    wire \u0.N_2137 ;
    wire PIO_dport1_Teoc_4;
    wire \u0.dat_o_i_i_1_28 ;
    wire \u0.N_2137_cascade_ ;
    wire \u0.dat_o_i_i_2_28 ;
    wire \u0.dat_o_i_i_4_28_cascade_ ;
    wire \u0.N_1689 ;
    wire N_271;
    wire \u0.N_1699 ;
    wire \u0.N_2095 ;
    wire \u0.N_2095_cascade_ ;
    wire PIO_cmdport_Teoc_2;
    wire \u0.N_2130_cascade_ ;
    wire \u0.CtrlRegZ0Z_26 ;
    wire \u0.dat_o_i_i_1_26 ;
    wire \u0.N_2122 ;
    wire PIO_dport1_Teoc_6;
    wire PIO_dport0_Teoc_6;
    wire \u0.N_1703_cascade_ ;
    wire \u0.N_2104 ;
    wire DMA_dev0_Teoc_4;
    wire \u0.N_1686 ;
    wire N_1321;
    wire DMAq_24;
    wire N_2119_cascade_;
    wire DMA_dev0_Teoc_0;
    wire \u0.N_2130 ;
    wire \u0.N_2123 ;
    wire PIO_cmdport_Teoc_6;
    wire \u0.dat_o_i_i_1_30 ;
    wire DMA_dev0_Teoc_6;
    wire DMAq_30;
    wire \u0.dat_o_i_i_4_30 ;
    wire \u0.dat_o_i_i_0_30_cascade_ ;
    wire DMA_dev1_Teoc_6;
    wire N_275;
    wire wb_dat_i_c_30;
    wire \u0.CtrlRegZ0Z_30 ;
    wire \u0.dat_o_0_a2_i_o2_0Z0Z_16 ;
    wire wb_adr_i_c_3;
    wire \u0.N_1714 ;
    wire \u0.dat_o_i_0_0_23 ;
    wire \u0.N_1374_cascade_ ;
    wire N_332_i;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI6ONK1Z0Z_2 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIBAOD1Z0Z_1 ;
    wire wb_adr_i_c_6;
    wire N_2119;
    wire DMAq_1_cascade_;
    wire PIOq_1;
    wire \u0.dat_o_0_0_1Z0Z_1 ;
    wire \u0.N_1729 ;
    wire \u0.dat_o_i_0_0_18 ;
    wire \u0.dat_o_i_0_2_18 ;
    wire N_325_i;
    wire iQ_RNIUKDM1_2;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIAH7KZ0Z_17 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI6TUQZ0Z_17 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIE5GTZ0Z_17 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_17 ;
    wire iQ_RNI2PDM1_2;
    wire mem_mem_ram6__RNIG5B71_17_cascade_;
    wire u1_DMA_control_gen_DMAbuf_Rxbuf_rd_ptr_2;
    wire \u0.N_1549 ;
    wire \u0.dat_o_0_a2_i_0_16 ;
    wire \u0.dat_o_0_a2_i_2_16 ;
    wire N_207_i;
    wire \u0.N_2128 ;
    wire DMA_dev0_Td_1;
    wire \u0.dat_o_0_0_2_9 ;
    wire \u0.dat_o_0_0_6_9 ;
    wire \u0.N_1651_cascade_ ;
    wire \u0.N_1650 ;
    wire wb_dat_o_c_9;
    wire \u1.DMA_control.rd_ptr_1 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_16 ;
    wire \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIC3GTZ0Z_16 ;
    wire mem_mem_ram6__RNID2B71_16;
    wire PIO_cmdport_Teoc_5;
    wire N_448_g;
    wire \u0.dat_o_0_a2_i_2_17 ;
    wire \u0.N_1374 ;
    wire \u0.N_1554 ;
    wire N_209_i;
    wire wb_dat_i_c_0;
    wire PIO_dport0_T1_0;
    wire N_77_g;
    wire wb_dat_i_c_29;
    wire \u0.CtrlRegZ0Z_29 ;
    wire PIO_dport0_T4_7;
    wire PIO_dport1_T4_7;
    wire \u0.dat_o_i_0_1_23 ;
    wire \u0.dat_o_i_i_0_25 ;
    wire \u0.dat_o_i_i_4_25 ;
    wire DMA_dev1_Teoc_1;
    wire N_265;
    wire \u0.dat_o_i_i_4_24 ;
    wire \u0.N_2124 ;
    wire \u0.dat_o_i_i_0_24 ;
    wire DMA_dev1_Teoc_0;
    wire N_263;
    wire wb_dat_i_c_8;
    wire DMActrl_BeLeC0;
    wire wb_clk_i_c_g;
    wire \u0.N_286 ;
    wire arst_i_c_i_g;
    wire wb_adr_i_c_4;
    wire \u0.N_2139 ;
    wire PIO_dport0_T4_1;
    wire PIO_dport1_T4_1;
    wire \u0.dat_o_0_a2_i_0_17 ;
    wire wb_rst_i_c;
    wire N_2140;
    wire \u0.N_2129 ;
    wire N_77;
    wire wb_adr_i_c_2;
    wire wb_adr_i_c_5;
    wire \u0.N_2143 ;
    wire _gnd_net_;

    PRE_IO_GBUF wb_clk_i_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__55910),
            .GLOBALBUFFEROUTPUT(wb_clk_i_c_g));
    IO_PAD wb_clk_i_ibuf_gb_io_iopad (
            .OE(N__55912),
            .DIN(N__55911),
            .DOUT(N__55910),
            .PACKAGEPIN(wb_clk_i));
    defparam wb_clk_i_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam wb_clk_i_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_clk_i_ibuf_gb_io_preio (
            .PADOEN(N__55912),
            .PADOUT(N__55911),
            .PADIN(N__55910),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD DMA_Ack_ibuf_iopad (
            .OE(N__55901),
            .DIN(N__55900),
            .DOUT(N__55899),
            .PACKAGEPIN(DMA_Ack));
    defparam DMA_Ack_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam DMA_Ack_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO DMA_Ack_ibuf_preio (
            .PADOEN(N__55901),
            .PADOUT(N__55900),
            .PADIN(N__55899),
            .CLOCKENABLE(),
            .DIN0(DMA_Ack_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD DMA_req_obuf_iopad (
            .OE(N__55892),
            .DIN(N__55891),
            .DOUT(N__55890),
            .PACKAGEPIN(DMA_req));
    defparam DMA_req_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DMA_req_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DMA_req_obuf_preio (
            .PADOEN(N__55892),
            .PADOUT(N__55891),
            .PADIN(N__55890),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__20209),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD arst_i_ibuf_iopad (
            .OE(N__55883),
            .DIN(N__55882),
            .DOUT(N__55881),
            .PACKAGEPIN(arst_i));
    defparam arst_i_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam arst_i_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO arst_i_ibuf_preio (
            .PADOEN(N__55883),
            .PADOUT(N__55882),
            .PADIN(N__55881),
            .CLOCKENABLE(),
            .DIN0(arst_i_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD cs0n_pad_o_obuf_iopad (
            .OE(N__55874),
            .DIN(N__55873),
            .DOUT(N__55872),
            .PACKAGEPIN(cs0n_pad_o));
    defparam cs0n_pad_o_obuf_preio.NEG_TRIGGER=1'b0;
    defparam cs0n_pad_o_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO cs0n_pad_o_obuf_preio (
            .PADOEN(N__55874),
            .PADOUT(N__55873),
            .PADIN(N__55872),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__26974),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD cs1n_pad_o_obuf_iopad (
            .OE(N__55865),
            .DIN(N__55864),
            .DOUT(N__55863),
            .PACKAGEPIN(cs1n_pad_o));
    defparam cs1n_pad_o_obuf_preio.NEG_TRIGGER=1'b0;
    defparam cs1n_pad_o_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO cs1n_pad_o_obuf_preio (
            .PADOEN(N__55865),
            .PADOUT(N__55864),
            .PADIN(N__55863),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__26695),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD da_pad_o_obuf_0_iopad (
            .OE(N__55856),
            .DIN(N__55855),
            .DOUT(N__55854),
            .PACKAGEPIN(da_pad_o[0]));
    defparam da_pad_o_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam da_pad_o_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO da_pad_o_obuf_0_preio (
            .PADOEN(N__55856),
            .PADOUT(N__55855),
            .PADIN(N__55854),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__26386),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD da_pad_o_obuf_1_iopad (
            .OE(N__55847),
            .DIN(N__55846),
            .DOUT(N__55845),
            .PACKAGEPIN(da_pad_o[1]));
    defparam da_pad_o_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam da_pad_o_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO da_pad_o_obuf_1_preio (
            .PADOEN(N__55847),
            .PADOUT(N__55846),
            .PADIN(N__55845),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__23566),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD da_pad_o_obuf_2_iopad (
            .OE(N__55838),
            .DIN(N__55837),
            .DOUT(N__55836),
            .PACKAGEPIN(da_pad_o[2]));
    defparam da_pad_o_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam da_pad_o_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO da_pad_o_obuf_2_preio (
            .PADOEN(N__55838),
            .PADOUT(N__55837),
            .PADIN(N__55836),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__20725),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD dd_pad_i_ibuf_0_iopad (
            .OE(N__55829),
            .DIN(N__55828),
            .DOUT(N__55827),
            .PACKAGEPIN(dd_pad_i[0]));
    defparam dd_pad_i_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam dd_pad_i_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO dd_pad_i_ibuf_0_preio (
            .PADOEN(N__55829),
            .PADOUT(N__55828),
            .PADIN(N__55827),
            .CLOCKENABLE(),
            .DIN0(dd_pad_i_c_0),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD dd_pad_i_ibuf_1_iopad (
            .OE(N__55820),
            .DIN(N__55819),
            .DOUT(N__55818),
            .PACKAGEPIN(dd_pad_i[1]));
    defparam dd_pad_i_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam dd_pad_i_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO dd_pad_i_ibuf_1_preio (
            .PADOEN(N__55820),
            .PADOUT(N__55819),
            .PADIN(N__55818),
            .CLOCKENABLE(),
            .DIN0(dd_pad_i_c_1),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD dd_pad_i_ibuf_10_iopad (
            .OE(N__55811),
            .DIN(N__55810),
            .DOUT(N__55809),
            .PACKAGEPIN(dd_pad_i[10]));
    defparam dd_pad_i_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam dd_pad_i_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO dd_pad_i_ibuf_10_preio (
            .PADOEN(N__55811),
            .PADOUT(N__55810),
            .PADIN(N__55809),
            .CLOCKENABLE(),
            .DIN0(dd_pad_i_c_10),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD dd_pad_i_ibuf_11_iopad (
            .OE(N__55802),
            .DIN(N__55801),
            .DOUT(N__55800),
            .PACKAGEPIN(dd_pad_i[11]));
    defparam dd_pad_i_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam dd_pad_i_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO dd_pad_i_ibuf_11_preio (
            .PADOEN(N__55802),
            .PADOUT(N__55801),
            .PADIN(N__55800),
            .CLOCKENABLE(),
            .DIN0(dd_pad_i_c_11),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD dd_pad_i_ibuf_12_iopad (
            .OE(N__55793),
            .DIN(N__55792),
            .DOUT(N__55791),
            .PACKAGEPIN(dd_pad_i[12]));
    defparam dd_pad_i_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam dd_pad_i_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO dd_pad_i_ibuf_12_preio (
            .PADOEN(N__55793),
            .PADOUT(N__55792),
            .PADIN(N__55791),
            .CLOCKENABLE(),
            .DIN0(dd_pad_i_c_12),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD dd_pad_i_ibuf_13_iopad (
            .OE(N__55784),
            .DIN(N__55783),
            .DOUT(N__55782),
            .PACKAGEPIN(dd_pad_i[13]));
    defparam dd_pad_i_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam dd_pad_i_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO dd_pad_i_ibuf_13_preio (
            .PADOEN(N__55784),
            .PADOUT(N__55783),
            .PADIN(N__55782),
            .CLOCKENABLE(),
            .DIN0(dd_pad_i_c_13),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD dd_pad_i_ibuf_14_iopad (
            .OE(N__55775),
            .DIN(N__55774),
            .DOUT(N__55773),
            .PACKAGEPIN(dd_pad_i[14]));
    defparam dd_pad_i_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam dd_pad_i_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO dd_pad_i_ibuf_14_preio (
            .PADOEN(N__55775),
            .PADOUT(N__55774),
            .PADIN(N__55773),
            .CLOCKENABLE(),
            .DIN0(dd_pad_i_c_14),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD dd_pad_i_ibuf_15_iopad (
            .OE(N__55766),
            .DIN(N__55765),
            .DOUT(N__55764),
            .PACKAGEPIN(dd_pad_i[15]));
    defparam dd_pad_i_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam dd_pad_i_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO dd_pad_i_ibuf_15_preio (
            .PADOEN(N__55766),
            .PADOUT(N__55765),
            .PADIN(N__55764),
            .CLOCKENABLE(),
            .DIN0(dd_pad_i_c_15),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD dd_pad_i_ibuf_2_iopad (
            .OE(N__55757),
            .DIN(N__55756),
            .DOUT(N__55755),
            .PACKAGEPIN(dd_pad_i[2]));
    defparam dd_pad_i_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam dd_pad_i_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO dd_pad_i_ibuf_2_preio (
            .PADOEN(N__55757),
            .PADOUT(N__55756),
            .PADIN(N__55755),
            .CLOCKENABLE(),
            .DIN0(dd_pad_i_c_2),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD dd_pad_i_ibuf_3_iopad (
            .OE(N__55748),
            .DIN(N__55747),
            .DOUT(N__55746),
            .PACKAGEPIN(dd_pad_i[3]));
    defparam dd_pad_i_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam dd_pad_i_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO dd_pad_i_ibuf_3_preio (
            .PADOEN(N__55748),
            .PADOUT(N__55747),
            .PADIN(N__55746),
            .CLOCKENABLE(),
            .DIN0(dd_pad_i_c_3),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD dd_pad_i_ibuf_4_iopad (
            .OE(N__55739),
            .DIN(N__55738),
            .DOUT(N__55737),
            .PACKAGEPIN(dd_pad_i[4]));
    defparam dd_pad_i_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam dd_pad_i_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO dd_pad_i_ibuf_4_preio (
            .PADOEN(N__55739),
            .PADOUT(N__55738),
            .PADIN(N__55737),
            .CLOCKENABLE(),
            .DIN0(dd_pad_i_c_4),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD dd_pad_i_ibuf_5_iopad (
            .OE(N__55730),
            .DIN(N__55729),
            .DOUT(N__55728),
            .PACKAGEPIN(dd_pad_i[5]));
    defparam dd_pad_i_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam dd_pad_i_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO dd_pad_i_ibuf_5_preio (
            .PADOEN(N__55730),
            .PADOUT(N__55729),
            .PADIN(N__55728),
            .CLOCKENABLE(),
            .DIN0(dd_pad_i_c_5),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD dd_pad_i_ibuf_6_iopad (
            .OE(N__55721),
            .DIN(N__55720),
            .DOUT(N__55719),
            .PACKAGEPIN(dd_pad_i[6]));
    defparam dd_pad_i_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam dd_pad_i_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO dd_pad_i_ibuf_6_preio (
            .PADOEN(N__55721),
            .PADOUT(N__55720),
            .PADIN(N__55719),
            .CLOCKENABLE(),
            .DIN0(dd_pad_i_c_6),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD dd_pad_i_ibuf_7_iopad (
            .OE(N__55712),
            .DIN(N__55711),
            .DOUT(N__55710),
            .PACKAGEPIN(dd_pad_i[7]));
    defparam dd_pad_i_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam dd_pad_i_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO dd_pad_i_ibuf_7_preio (
            .PADOEN(N__55712),
            .PADOUT(N__55711),
            .PADIN(N__55710),
            .CLOCKENABLE(),
            .DIN0(dd_pad_i_c_7),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD dd_pad_i_ibuf_8_iopad (
            .OE(N__55703),
            .DIN(N__55702),
            .DOUT(N__55701),
            .PACKAGEPIN(dd_pad_i[8]));
    defparam dd_pad_i_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam dd_pad_i_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO dd_pad_i_ibuf_8_preio (
            .PADOEN(N__55703),
            .PADOUT(N__55702),
            .PADIN(N__55701),
            .CLOCKENABLE(),
            .DIN0(dd_pad_i_c_8),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD dd_pad_i_ibuf_9_iopad (
            .OE(N__55694),
            .DIN(N__55693),
            .DOUT(N__55692),
            .PACKAGEPIN(dd_pad_i[9]));
    defparam dd_pad_i_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam dd_pad_i_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO dd_pad_i_ibuf_9_preio (
            .PADOEN(N__55694),
            .PADOUT(N__55693),
            .PADIN(N__55692),
            .CLOCKENABLE(),
            .DIN0(dd_pad_i_c_9),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD dd_pad_o_obuf_0_iopad (
            .OE(N__55685),
            .DIN(N__55684),
            .DOUT(N__55683),
            .PACKAGEPIN(dd_pad_o[0]));
    defparam dd_pad_o_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam dd_pad_o_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO dd_pad_o_obuf_0_preio (
            .PADOEN(N__55685),
            .PADOUT(N__55684),
            .PADIN(N__55683),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__27031),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD dd_pad_o_obuf_1_iopad (
            .OE(N__55676),
            .DIN(N__55675),
            .DOUT(N__55674),
            .PACKAGEPIN(dd_pad_o[1]));
    defparam dd_pad_o_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam dd_pad_o_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO dd_pad_o_obuf_1_preio (
            .PADOEN(N__55676),
            .PADOUT(N__55675),
            .PADIN(N__55674),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__26713),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD dd_pad_o_obuf_10_iopad (
            .OE(N__55667),
            .DIN(N__55666),
            .DOUT(N__55665),
            .PACKAGEPIN(dd_pad_o[10]));
    defparam dd_pad_o_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam dd_pad_o_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO dd_pad_o_obuf_10_preio (
            .PADOEN(N__55667),
            .PADOUT(N__55666),
            .PADIN(N__55665),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__21763),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD dd_pad_o_obuf_11_iopad (
            .OE(N__55658),
            .DIN(N__55657),
            .DOUT(N__55656),
            .PACKAGEPIN(dd_pad_o[11]));
    defparam dd_pad_o_obuf_11_preio.NEG_TRIGGER=1'b0;
    defparam dd_pad_o_obuf_11_preio.PIN_TYPE=6'b011001;
    PRE_IO dd_pad_o_obuf_11_preio (
            .PADOEN(N__55658),
            .PADOUT(N__55657),
            .PADIN(N__55656),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__22519),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD dd_pad_o_obuf_12_iopad (
            .OE(N__55649),
            .DIN(N__55648),
            .DOUT(N__55647),
            .PACKAGEPIN(dd_pad_o[12]));
    defparam dd_pad_o_obuf_12_preio.NEG_TRIGGER=1'b0;
    defparam dd_pad_o_obuf_12_preio.PIN_TYPE=6'b011001;
    PRE_IO dd_pad_o_obuf_12_preio (
            .PADOEN(N__55649),
            .PADOUT(N__55648),
            .PADIN(N__55647),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__22927),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD dd_pad_o_obuf_13_iopad (
            .OE(N__55640),
            .DIN(N__55639),
            .DOUT(N__55638),
            .PACKAGEPIN(dd_pad_o[13]));
    defparam dd_pad_o_obuf_13_preio.NEG_TRIGGER=1'b0;
    defparam dd_pad_o_obuf_13_preio.PIN_TYPE=6'b011001;
    PRE_IO dd_pad_o_obuf_13_preio (
            .PADOEN(N__55640),
            .PADOUT(N__55639),
            .PADIN(N__55638),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__21244),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD dd_pad_o_obuf_14_iopad (
            .OE(N__55631),
            .DIN(N__55630),
            .DOUT(N__55629),
            .PACKAGEPIN(dd_pad_o[14]));
    defparam dd_pad_o_obuf_14_preio.NEG_TRIGGER=1'b0;
    defparam dd_pad_o_obuf_14_preio.PIN_TYPE=6'b011001;
    PRE_IO dd_pad_o_obuf_14_preio (
            .PADOEN(N__55631),
            .PADOUT(N__55630),
            .PADIN(N__55629),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__22900),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD dd_pad_o_obuf_15_iopad (
            .OE(N__55622),
            .DIN(N__55621),
            .DOUT(N__55620),
            .PACKAGEPIN(dd_pad_o[15]));
    defparam dd_pad_o_obuf_15_preio.NEG_TRIGGER=1'b0;
    defparam dd_pad_o_obuf_15_preio.PIN_TYPE=6'b011001;
    PRE_IO dd_pad_o_obuf_15_preio (
            .PADOEN(N__55622),
            .PADOUT(N__55621),
            .PADIN(N__55620),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__20578),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD dd_pad_o_obuf_2_iopad (
            .OE(N__55613),
            .DIN(N__55612),
            .DOUT(N__55611),
            .PACKAGEPIN(dd_pad_o[2]));
    defparam dd_pad_o_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam dd_pad_o_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO dd_pad_o_obuf_2_preio (
            .PADOEN(N__55613),
            .PADOUT(N__55612),
            .PADIN(N__55611),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__20311),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD dd_pad_o_obuf_3_iopad (
            .OE(N__55604),
            .DIN(N__55603),
            .DOUT(N__55602),
            .PACKAGEPIN(dd_pad_o[3]));
    defparam dd_pad_o_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam dd_pad_o_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO dd_pad_o_obuf_3_preio (
            .PADOEN(N__55604),
            .PADOUT(N__55603),
            .PADIN(N__55602),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__20284),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD dd_pad_o_obuf_4_iopad (
            .OE(N__55595),
            .DIN(N__55594),
            .DOUT(N__55593),
            .PACKAGEPIN(dd_pad_o[4]));
    defparam dd_pad_o_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam dd_pad_o_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO dd_pad_o_obuf_4_preio (
            .PADOEN(N__55595),
            .PADOUT(N__55594),
            .PADIN(N__55593),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__21217),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD dd_pad_o_obuf_5_iopad (
            .OE(N__55586),
            .DIN(N__55585),
            .DOUT(N__55584),
            .PACKAGEPIN(dd_pad_o[5]));
    defparam dd_pad_o_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam dd_pad_o_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO dd_pad_o_obuf_5_preio (
            .PADOEN(N__55586),
            .PADOUT(N__55585),
            .PADIN(N__55584),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__21328),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD dd_pad_o_obuf_6_iopad (
            .OE(N__55577),
            .DIN(N__55576),
            .DOUT(N__55575),
            .PACKAGEPIN(dd_pad_o[6]));
    defparam dd_pad_o_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam dd_pad_o_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO dd_pad_o_obuf_6_preio (
            .PADOEN(N__55577),
            .PADOUT(N__55576),
            .PADIN(N__55575),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__21226),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD dd_pad_o_obuf_7_iopad (
            .OE(N__55568),
            .DIN(N__55567),
            .DOUT(N__55566),
            .PACKAGEPIN(dd_pad_o[7]));
    defparam dd_pad_o_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam dd_pad_o_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO dd_pad_o_obuf_7_preio (
            .PADOEN(N__55568),
            .PADOUT(N__55567),
            .PADIN(N__55566),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__22846),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD dd_pad_o_obuf_8_iopad (
            .OE(N__55559),
            .DIN(N__55558),
            .DOUT(N__55557),
            .PACKAGEPIN(dd_pad_o[8]));
    defparam dd_pad_o_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam dd_pad_o_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO dd_pad_o_obuf_8_preio (
            .PADOEN(N__55559),
            .PADOUT(N__55558),
            .PADIN(N__55557),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__22873),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD dd_pad_o_obuf_9_iopad (
            .OE(N__55550),
            .DIN(N__55549),
            .DOUT(N__55548),
            .PACKAGEPIN(dd_pad_o[9]));
    defparam dd_pad_o_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam dd_pad_o_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO dd_pad_o_obuf_9_preio (
            .PADOEN(N__55550),
            .PADOUT(N__55549),
            .PADIN(N__55548),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__19501),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD dd_padoe_o_obuf_iopad (
            .OE(N__55541),
            .DIN(N__55540),
            .DOUT(N__55539),
            .PACKAGEPIN(dd_padoe_o));
    defparam dd_padoe_o_obuf_preio.NEG_TRIGGER=1'b0;
    defparam dd_padoe_o_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO dd_padoe_o_obuf_preio (
            .PADOEN(N__55541),
            .PADOUT(N__55540),
            .PADIN(N__55539),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__19378),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD diorn_pad_o_obuf_iopad (
            .OE(N__55532),
            .DIN(N__55531),
            .DOUT(N__55530),
            .PACKAGEPIN(diorn_pad_o));
    defparam diorn_pad_o_obuf_preio.NEG_TRIGGER=1'b0;
    defparam diorn_pad_o_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO diorn_pad_o_obuf_preio (
            .PADOEN(N__55532),
            .PADOUT(N__55531),
            .PADIN(N__55530),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__19645),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD diown_pad_o_obuf_iopad (
            .OE(N__55523),
            .DIN(N__55522),
            .DOUT(N__55521),
            .PACKAGEPIN(diown_pad_o));
    defparam diown_pad_o_obuf_preio.NEG_TRIGGER=1'b0;
    defparam diown_pad_o_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO diown_pad_o_obuf_preio (
            .PADOEN(N__55523),
            .PADOUT(N__55522),
            .PADIN(N__55521),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__19336),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD dmackn_pad_o_obuf_iopad (
            .OE(N__55514),
            .DIN(N__55513),
            .DOUT(N__55512),
            .PACKAGEPIN(dmackn_pad_o));
    defparam dmackn_pad_o_obuf_preio.NEG_TRIGGER=1'b0;
    defparam dmackn_pad_o_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO dmackn_pad_o_obuf_preio (
            .PADOEN(N__55514),
            .PADOUT(N__55513),
            .PADIN(N__55512),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__21598),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD dmarq_pad_i_ibuf_iopad (
            .OE(N__55505),
            .DIN(N__55504),
            .DOUT(N__55503),
            .PACKAGEPIN(dmarq_pad_i));
    defparam dmarq_pad_i_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam dmarq_pad_i_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO dmarq_pad_i_ibuf_preio (
            .PADOEN(N__55505),
            .PADOUT(N__55504),
            .PADIN(N__55503),
            .CLOCKENABLE(),
            .DIN0(dmarq_pad_i_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD intrq_pad_i_ibuf_iopad (
            .OE(N__55496),
            .DIN(N__55495),
            .DOUT(N__55494),
            .PACKAGEPIN(intrq_pad_i));
    defparam intrq_pad_i_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam intrq_pad_i_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO intrq_pad_i_ibuf_preio (
            .PADOEN(N__55496),
            .PADOUT(N__55495),
            .PADIN(N__55494),
            .CLOCKENABLE(),
            .DIN0(intrq_pad_i_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD iordy_pad_i_ibuf_iopad (
            .OE(N__55487),
            .DIN(N__55486),
            .DOUT(N__55485),
            .PACKAGEPIN(iordy_pad_i));
    defparam iordy_pad_i_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam iordy_pad_i_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO iordy_pad_i_ibuf_preio (
            .PADOEN(N__55487),
            .PADOUT(N__55486),
            .PADIN(N__55485),
            .CLOCKENABLE(),
            .DIN0(iordy_pad_i_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD resetn_pad_o_obuf_iopad (
            .OE(N__55478),
            .DIN(N__55477),
            .DOUT(N__55476),
            .PACKAGEPIN(resetn_pad_o));
    defparam resetn_pad_o_obuf_preio.NEG_TRIGGER=1'b0;
    defparam resetn_pad_o_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO resetn_pad_o_obuf_preio (
            .PADOEN(N__55478),
            .PADOUT(N__55477),
            .PADIN(N__55476),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__23545),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_ack_o_obuf_iopad (
            .OE(N__55469),
            .DIN(N__55468),
            .DOUT(N__55467),
            .PACKAGEPIN(wb_ack_o));
    defparam wb_ack_o_obuf_preio.NEG_TRIGGER=1'b0;
    defparam wb_ack_o_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO wb_ack_o_obuf_preio (
            .PADOEN(N__55469),
            .PADOUT(N__55468),
            .PADIN(N__55467),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__21661),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_adr_i_ibuf_2_iopad (
            .OE(N__55460),
            .DIN(N__55459),
            .DOUT(N__55458),
            .PACKAGEPIN(wb_adr_i[2]));
    defparam wb_adr_i_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam wb_adr_i_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_adr_i_ibuf_2_preio (
            .PADOEN(N__55460),
            .PADOUT(N__55459),
            .PADIN(N__55458),
            .CLOCKENABLE(),
            .DIN0(wb_adr_i_c_2),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_adr_i_ibuf_3_iopad (
            .OE(N__55451),
            .DIN(N__55450),
            .DOUT(N__55449),
            .PACKAGEPIN(wb_adr_i[3]));
    defparam wb_adr_i_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam wb_adr_i_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_adr_i_ibuf_3_preio (
            .PADOEN(N__55451),
            .PADOUT(N__55450),
            .PADIN(N__55449),
            .CLOCKENABLE(),
            .DIN0(wb_adr_i_c_3),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_adr_i_ibuf_4_iopad (
            .OE(N__55442),
            .DIN(N__55441),
            .DOUT(N__55440),
            .PACKAGEPIN(wb_adr_i[4]));
    defparam wb_adr_i_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam wb_adr_i_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_adr_i_ibuf_4_preio (
            .PADOEN(N__55442),
            .PADOUT(N__55441),
            .PADIN(N__55440),
            .CLOCKENABLE(),
            .DIN0(wb_adr_i_c_4),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_adr_i_ibuf_5_iopad (
            .OE(N__55433),
            .DIN(N__55432),
            .DOUT(N__55431),
            .PACKAGEPIN(wb_adr_i[5]));
    defparam wb_adr_i_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam wb_adr_i_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_adr_i_ibuf_5_preio (
            .PADOEN(N__55433),
            .PADOUT(N__55432),
            .PADIN(N__55431),
            .CLOCKENABLE(),
            .DIN0(wb_adr_i_c_5),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_adr_i_ibuf_6_iopad (
            .OE(N__55424),
            .DIN(N__55423),
            .DOUT(N__55422),
            .PACKAGEPIN(wb_adr_i[6]));
    defparam wb_adr_i_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam wb_adr_i_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_adr_i_ibuf_6_preio (
            .PADOEN(N__55424),
            .PADOUT(N__55423),
            .PADIN(N__55422),
            .CLOCKENABLE(),
            .DIN0(wb_adr_i_c_6),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_cyc_i_ibuf_iopad (
            .OE(N__55415),
            .DIN(N__55414),
            .DOUT(N__55413),
            .PACKAGEPIN(wb_cyc_i));
    defparam wb_cyc_i_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam wb_cyc_i_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_cyc_i_ibuf_preio (
            .PADOEN(N__55415),
            .PADOUT(N__55414),
            .PADIN(N__55413),
            .CLOCKENABLE(),
            .DIN0(wb_cyc_i_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_i_ibuf_0_iopad (
            .OE(N__55406),
            .DIN(N__55405),
            .DOUT(N__55404),
            .PACKAGEPIN(wb_dat_i[0]));
    defparam wb_dat_i_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_i_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_dat_i_ibuf_0_preio (
            .PADOEN(N__55406),
            .PADOUT(N__55405),
            .PADIN(N__55404),
            .CLOCKENABLE(),
            .DIN0(wb_dat_i_c_0),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_i_ibuf_1_iopad (
            .OE(N__55397),
            .DIN(N__55396),
            .DOUT(N__55395),
            .PACKAGEPIN(wb_dat_i[1]));
    defparam wb_dat_i_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_i_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_dat_i_ibuf_1_preio (
            .PADOEN(N__55397),
            .PADOUT(N__55396),
            .PADIN(N__55395),
            .CLOCKENABLE(),
            .DIN0(wb_dat_i_c_1),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_i_ibuf_10_iopad (
            .OE(N__55388),
            .DIN(N__55387),
            .DOUT(N__55386),
            .PACKAGEPIN(wb_dat_i[10]));
    defparam wb_dat_i_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_i_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_dat_i_ibuf_10_preio (
            .PADOEN(N__55388),
            .PADOUT(N__55387),
            .PADIN(N__55386),
            .CLOCKENABLE(),
            .DIN0(wb_dat_i_c_10),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_i_ibuf_11_iopad (
            .OE(N__55379),
            .DIN(N__55378),
            .DOUT(N__55377),
            .PACKAGEPIN(wb_dat_i[11]));
    defparam wb_dat_i_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_i_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_dat_i_ibuf_11_preio (
            .PADOEN(N__55379),
            .PADOUT(N__55378),
            .PADIN(N__55377),
            .CLOCKENABLE(),
            .DIN0(wb_dat_i_c_11),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_i_ibuf_12_iopad (
            .OE(N__55370),
            .DIN(N__55369),
            .DOUT(N__55368),
            .PACKAGEPIN(wb_dat_i[12]));
    defparam wb_dat_i_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_i_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_dat_i_ibuf_12_preio (
            .PADOEN(N__55370),
            .PADOUT(N__55369),
            .PADIN(N__55368),
            .CLOCKENABLE(),
            .DIN0(wb_dat_i_c_12),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_i_ibuf_13_iopad (
            .OE(N__55361),
            .DIN(N__55360),
            .DOUT(N__55359),
            .PACKAGEPIN(wb_dat_i[13]));
    defparam wb_dat_i_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_i_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_dat_i_ibuf_13_preio (
            .PADOEN(N__55361),
            .PADOUT(N__55360),
            .PADIN(N__55359),
            .CLOCKENABLE(),
            .DIN0(wb_dat_i_c_13),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_i_ibuf_14_iopad (
            .OE(N__55352),
            .DIN(N__55351),
            .DOUT(N__55350),
            .PACKAGEPIN(wb_dat_i[14]));
    defparam wb_dat_i_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_i_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_dat_i_ibuf_14_preio (
            .PADOEN(N__55352),
            .PADOUT(N__55351),
            .PADIN(N__55350),
            .CLOCKENABLE(),
            .DIN0(wb_dat_i_c_14),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_i_ibuf_15_iopad (
            .OE(N__55343),
            .DIN(N__55342),
            .DOUT(N__55341),
            .PACKAGEPIN(wb_dat_i[15]));
    defparam wb_dat_i_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_i_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_dat_i_ibuf_15_preio (
            .PADOEN(N__55343),
            .PADOUT(N__55342),
            .PADIN(N__55341),
            .CLOCKENABLE(),
            .DIN0(wb_dat_i_c_15),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_i_ibuf_16_iopad (
            .OE(N__55334),
            .DIN(N__55333),
            .DOUT(N__55332),
            .PACKAGEPIN(wb_dat_i[16]));
    defparam wb_dat_i_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_i_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_dat_i_ibuf_16_preio (
            .PADOEN(N__55334),
            .PADOUT(N__55333),
            .PADIN(N__55332),
            .CLOCKENABLE(),
            .DIN0(wb_dat_i_c_16),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_i_ibuf_17_iopad (
            .OE(N__55325),
            .DIN(N__55324),
            .DOUT(N__55323),
            .PACKAGEPIN(wb_dat_i[17]));
    defparam wb_dat_i_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_i_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_dat_i_ibuf_17_preio (
            .PADOEN(N__55325),
            .PADOUT(N__55324),
            .PADIN(N__55323),
            .CLOCKENABLE(),
            .DIN0(wb_dat_i_c_17),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_i_ibuf_18_iopad (
            .OE(N__55316),
            .DIN(N__55315),
            .DOUT(N__55314),
            .PACKAGEPIN(wb_dat_i[18]));
    defparam wb_dat_i_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_i_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_dat_i_ibuf_18_preio (
            .PADOEN(N__55316),
            .PADOUT(N__55315),
            .PADIN(N__55314),
            .CLOCKENABLE(),
            .DIN0(wb_dat_i_c_18),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_i_ibuf_19_iopad (
            .OE(N__55307),
            .DIN(N__55306),
            .DOUT(N__55305),
            .PACKAGEPIN(wb_dat_i[19]));
    defparam wb_dat_i_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_i_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_dat_i_ibuf_19_preio (
            .PADOEN(N__55307),
            .PADOUT(N__55306),
            .PADIN(N__55305),
            .CLOCKENABLE(),
            .DIN0(wb_dat_i_c_19),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_i_ibuf_2_iopad (
            .OE(N__55298),
            .DIN(N__55297),
            .DOUT(N__55296),
            .PACKAGEPIN(wb_dat_i[2]));
    defparam wb_dat_i_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_i_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_dat_i_ibuf_2_preio (
            .PADOEN(N__55298),
            .PADOUT(N__55297),
            .PADIN(N__55296),
            .CLOCKENABLE(),
            .DIN0(wb_dat_i_c_2),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_i_ibuf_20_iopad (
            .OE(N__55289),
            .DIN(N__55288),
            .DOUT(N__55287),
            .PACKAGEPIN(wb_dat_i[20]));
    defparam wb_dat_i_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_i_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_dat_i_ibuf_20_preio (
            .PADOEN(N__55289),
            .PADOUT(N__55288),
            .PADIN(N__55287),
            .CLOCKENABLE(),
            .DIN0(wb_dat_i_c_20),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_i_ibuf_21_iopad (
            .OE(N__55280),
            .DIN(N__55279),
            .DOUT(N__55278),
            .PACKAGEPIN(wb_dat_i[21]));
    defparam wb_dat_i_ibuf_21_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_i_ibuf_21_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_dat_i_ibuf_21_preio (
            .PADOEN(N__55280),
            .PADOUT(N__55279),
            .PADIN(N__55278),
            .CLOCKENABLE(),
            .DIN0(wb_dat_i_c_21),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_i_ibuf_22_iopad (
            .OE(N__55271),
            .DIN(N__55270),
            .DOUT(N__55269),
            .PACKAGEPIN(wb_dat_i[22]));
    defparam wb_dat_i_ibuf_22_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_i_ibuf_22_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_dat_i_ibuf_22_preio (
            .PADOEN(N__55271),
            .PADOUT(N__55270),
            .PADIN(N__55269),
            .CLOCKENABLE(),
            .DIN0(wb_dat_i_c_22),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_i_ibuf_23_iopad (
            .OE(N__55262),
            .DIN(N__55261),
            .DOUT(N__55260),
            .PACKAGEPIN(wb_dat_i[23]));
    defparam wb_dat_i_ibuf_23_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_i_ibuf_23_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_dat_i_ibuf_23_preio (
            .PADOEN(N__55262),
            .PADOUT(N__55261),
            .PADIN(N__55260),
            .CLOCKENABLE(),
            .DIN0(wb_dat_i_c_23),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_i_ibuf_24_iopad (
            .OE(N__55253),
            .DIN(N__55252),
            .DOUT(N__55251),
            .PACKAGEPIN(wb_dat_i[24]));
    defparam wb_dat_i_ibuf_24_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_i_ibuf_24_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_dat_i_ibuf_24_preio (
            .PADOEN(N__55253),
            .PADOUT(N__55252),
            .PADIN(N__55251),
            .CLOCKENABLE(),
            .DIN0(wb_dat_i_c_24),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_i_ibuf_25_iopad (
            .OE(N__55244),
            .DIN(N__55243),
            .DOUT(N__55242),
            .PACKAGEPIN(wb_dat_i[25]));
    defparam wb_dat_i_ibuf_25_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_i_ibuf_25_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_dat_i_ibuf_25_preio (
            .PADOEN(N__55244),
            .PADOUT(N__55243),
            .PADIN(N__55242),
            .CLOCKENABLE(),
            .DIN0(wb_dat_i_c_25),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_i_ibuf_26_iopad (
            .OE(N__55235),
            .DIN(N__55234),
            .DOUT(N__55233),
            .PACKAGEPIN(wb_dat_i[26]));
    defparam wb_dat_i_ibuf_26_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_i_ibuf_26_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_dat_i_ibuf_26_preio (
            .PADOEN(N__55235),
            .PADOUT(N__55234),
            .PADIN(N__55233),
            .CLOCKENABLE(),
            .DIN0(wb_dat_i_c_26),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_i_ibuf_27_iopad (
            .OE(N__55226),
            .DIN(N__55225),
            .DOUT(N__55224),
            .PACKAGEPIN(wb_dat_i[27]));
    defparam wb_dat_i_ibuf_27_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_i_ibuf_27_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_dat_i_ibuf_27_preio (
            .PADOEN(N__55226),
            .PADOUT(N__55225),
            .PADIN(N__55224),
            .CLOCKENABLE(),
            .DIN0(wb_dat_i_c_27),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_i_ibuf_28_iopad (
            .OE(N__55217),
            .DIN(N__55216),
            .DOUT(N__55215),
            .PACKAGEPIN(wb_dat_i[28]));
    defparam wb_dat_i_ibuf_28_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_i_ibuf_28_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_dat_i_ibuf_28_preio (
            .PADOEN(N__55217),
            .PADOUT(N__55216),
            .PADIN(N__55215),
            .CLOCKENABLE(),
            .DIN0(wb_dat_i_c_28),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_i_ibuf_29_iopad (
            .OE(N__55208),
            .DIN(N__55207),
            .DOUT(N__55206),
            .PACKAGEPIN(wb_dat_i[29]));
    defparam wb_dat_i_ibuf_29_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_i_ibuf_29_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_dat_i_ibuf_29_preio (
            .PADOEN(N__55208),
            .PADOUT(N__55207),
            .PADIN(N__55206),
            .CLOCKENABLE(),
            .DIN0(wb_dat_i_c_29),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_i_ibuf_3_iopad (
            .OE(N__55199),
            .DIN(N__55198),
            .DOUT(N__55197),
            .PACKAGEPIN(wb_dat_i[3]));
    defparam wb_dat_i_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_i_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_dat_i_ibuf_3_preio (
            .PADOEN(N__55199),
            .PADOUT(N__55198),
            .PADIN(N__55197),
            .CLOCKENABLE(),
            .DIN0(wb_dat_i_c_3),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_i_ibuf_30_iopad (
            .OE(N__55190),
            .DIN(N__55189),
            .DOUT(N__55188),
            .PACKAGEPIN(wb_dat_i[30]));
    defparam wb_dat_i_ibuf_30_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_i_ibuf_30_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_dat_i_ibuf_30_preio (
            .PADOEN(N__55190),
            .PADOUT(N__55189),
            .PADIN(N__55188),
            .CLOCKENABLE(),
            .DIN0(wb_dat_i_c_30),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_i_ibuf_31_iopad (
            .OE(N__55181),
            .DIN(N__55180),
            .DOUT(N__55179),
            .PACKAGEPIN(wb_dat_i[31]));
    defparam wb_dat_i_ibuf_31_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_i_ibuf_31_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_dat_i_ibuf_31_preio (
            .PADOEN(N__55181),
            .PADOUT(N__55180),
            .PADIN(N__55179),
            .CLOCKENABLE(),
            .DIN0(wb_dat_i_c_31),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_i_ibuf_4_iopad (
            .OE(N__55172),
            .DIN(N__55171),
            .DOUT(N__55170),
            .PACKAGEPIN(wb_dat_i[4]));
    defparam wb_dat_i_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_i_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_dat_i_ibuf_4_preio (
            .PADOEN(N__55172),
            .PADOUT(N__55171),
            .PADIN(N__55170),
            .CLOCKENABLE(),
            .DIN0(wb_dat_i_c_4),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_i_ibuf_5_iopad (
            .OE(N__55163),
            .DIN(N__55162),
            .DOUT(N__55161),
            .PACKAGEPIN(wb_dat_i[5]));
    defparam wb_dat_i_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_i_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_dat_i_ibuf_5_preio (
            .PADOEN(N__55163),
            .PADOUT(N__55162),
            .PADIN(N__55161),
            .CLOCKENABLE(),
            .DIN0(wb_dat_i_c_5),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_i_ibuf_6_iopad (
            .OE(N__55154),
            .DIN(N__55153),
            .DOUT(N__55152),
            .PACKAGEPIN(wb_dat_i[6]));
    defparam wb_dat_i_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_i_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_dat_i_ibuf_6_preio (
            .PADOEN(N__55154),
            .PADOUT(N__55153),
            .PADIN(N__55152),
            .CLOCKENABLE(),
            .DIN0(wb_dat_i_c_6),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_i_ibuf_7_iopad (
            .OE(N__55145),
            .DIN(N__55144),
            .DOUT(N__55143),
            .PACKAGEPIN(wb_dat_i[7]));
    defparam wb_dat_i_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_i_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_dat_i_ibuf_7_preio (
            .PADOEN(N__55145),
            .PADOUT(N__55144),
            .PADIN(N__55143),
            .CLOCKENABLE(),
            .DIN0(wb_dat_i_c_7),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_i_ibuf_8_iopad (
            .OE(N__55136),
            .DIN(N__55135),
            .DOUT(N__55134),
            .PACKAGEPIN(wb_dat_i[8]));
    defparam wb_dat_i_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_i_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_dat_i_ibuf_8_preio (
            .PADOEN(N__55136),
            .PADOUT(N__55135),
            .PADIN(N__55134),
            .CLOCKENABLE(),
            .DIN0(wb_dat_i_c_8),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_i_ibuf_9_iopad (
            .OE(N__55127),
            .DIN(N__55126),
            .DOUT(N__55125),
            .PACKAGEPIN(wb_dat_i[9]));
    defparam wb_dat_i_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_i_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_dat_i_ibuf_9_preio (
            .PADOEN(N__55127),
            .PADOUT(N__55126),
            .PADIN(N__55125),
            .CLOCKENABLE(),
            .DIN0(wb_dat_i_c_9),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_o_obuf_0_iopad (
            .OE(N__55118),
            .DIN(N__55117),
            .DOUT(N__55116),
            .PACKAGEPIN(wb_dat_o[0]));
    defparam wb_dat_o_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_o_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO wb_dat_o_obuf_0_preio (
            .PADOEN(N__55118),
            .PADOUT(N__55117),
            .PADIN(N__55116),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__43405),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_o_obuf_1_iopad (
            .OE(N__55109),
            .DIN(N__55108),
            .DOUT(N__55107),
            .PACKAGEPIN(wb_dat_o[1]));
    defparam wb_dat_o_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_o_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO wb_dat_o_obuf_1_preio (
            .PADOEN(N__55109),
            .PADOUT(N__55108),
            .PADIN(N__55107),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__44617),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_o_obuf_10_iopad (
            .OE(N__55100),
            .DIN(N__55099),
            .DOUT(N__55098),
            .PACKAGEPIN(wb_dat_o[10]));
    defparam wb_dat_o_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_o_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO wb_dat_o_obuf_10_preio (
            .PADOEN(N__55100),
            .PADOUT(N__55099),
            .PADIN(N__55098),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__40012),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_o_obuf_11_iopad (
            .OE(N__55091),
            .DIN(N__55090),
            .DOUT(N__55089),
            .PACKAGEPIN(wb_dat_o[11]));
    defparam wb_dat_o_obuf_11_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_o_obuf_11_preio.PIN_TYPE=6'b011001;
    PRE_IO wb_dat_o_obuf_11_preio (
            .PADOEN(N__55091),
            .PADOUT(N__55090),
            .PADIN(N__55089),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__43723),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_o_obuf_12_iopad (
            .OE(N__55082),
            .DIN(N__55081),
            .DOUT(N__55080),
            .PACKAGEPIN(wb_dat_o[12]));
    defparam wb_dat_o_obuf_12_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_o_obuf_12_preio.PIN_TYPE=6'b011001;
    PRE_IO wb_dat_o_obuf_12_preio (
            .PADOEN(N__55082),
            .PADOUT(N__55081),
            .PADIN(N__55080),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__29725),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_o_obuf_13_iopad (
            .OE(N__55073),
            .DIN(N__55072),
            .DOUT(N__55071),
            .PACKAGEPIN(wb_dat_o[13]));
    defparam wb_dat_o_obuf_13_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_o_obuf_13_preio.PIN_TYPE=6'b011001;
    PRE_IO wb_dat_o_obuf_13_preio (
            .PADOEN(N__55073),
            .PADOUT(N__55072),
            .PADIN(N__55071),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__26095),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_o_obuf_14_iopad (
            .OE(N__55064),
            .DIN(N__55063),
            .DOUT(N__55062),
            .PACKAGEPIN(wb_dat_o[14]));
    defparam wb_dat_o_obuf_14_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_o_obuf_14_preio.PIN_TYPE=6'b011001;
    PRE_IO wb_dat_o_obuf_14_preio (
            .PADOEN(N__55064),
            .PADOUT(N__55063),
            .PADIN(N__55062),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__43465),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_o_obuf_15_iopad (
            .OE(N__55055),
            .DIN(N__55054),
            .DOUT(N__55053),
            .PACKAGEPIN(wb_dat_o[15]));
    defparam wb_dat_o_obuf_15_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_o_obuf_15_preio.PIN_TYPE=6'b011001;
    PRE_IO wb_dat_o_obuf_15_preio (
            .PADOEN(N__55055),
            .PADOUT(N__55054),
            .PADIN(N__55053),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__25183),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_o_obuf_16_iopad (
            .OE(N__55046),
            .DIN(N__55045),
            .DOUT(N__55044),
            .PACKAGEPIN(wb_dat_o[16]));
    defparam wb_dat_o_obuf_16_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_o_obuf_16_preio.PIN_TYPE=6'b011001;
    PRE_IO wb_dat_o_obuf_16_preio (
            .PADOEN(N__55046),
            .PADOUT(N__55045),
            .PADIN(N__55044),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__48619),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_o_obuf_17_iopad (
            .OE(N__55037),
            .DIN(N__55036),
            .DOUT(N__55035),
            .PACKAGEPIN(wb_dat_o[17]));
    defparam wb_dat_o_obuf_17_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_o_obuf_17_preio.PIN_TYPE=6'b011001;
    PRE_IO wb_dat_o_obuf_17_preio (
            .PADOEN(N__55037),
            .PADOUT(N__55036),
            .PADIN(N__55035),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__49567),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_o_obuf_18_iopad (
            .OE(N__55028),
            .DIN(N__55027),
            .DOUT(N__55026),
            .PACKAGEPIN(wb_dat_o[18]));
    defparam wb_dat_o_obuf_18_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_o_obuf_18_preio.PIN_TYPE=6'b011001;
    PRE_IO wb_dat_o_obuf_18_preio (
            .PADOEN(N__55028),
            .PADOUT(N__55027),
            .PADIN(N__55026),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__49075),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_o_obuf_19_iopad (
            .OE(N__55019),
            .DIN(N__55018),
            .DOUT(N__55017),
            .PACKAGEPIN(wb_dat_o[19]));
    defparam wb_dat_o_obuf_19_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_o_obuf_19_preio.PIN_TYPE=6'b011001;
    PRE_IO wb_dat_o_obuf_19_preio (
            .PADOEN(N__55019),
            .PADOUT(N__55018),
            .PADIN(N__55017),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__25255),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_o_obuf_2_iopad (
            .OE(N__55010),
            .DIN(N__55009),
            .DOUT(N__55008),
            .PACKAGEPIN(wb_dat_o[2]));
    defparam wb_dat_o_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_o_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO wb_dat_o_obuf_2_preio (
            .PADOEN(N__55010),
            .PADOUT(N__55009),
            .PADIN(N__55008),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__27895),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_o_obuf_20_iopad (
            .OE(N__55001),
            .DIN(N__55000),
            .DOUT(N__54999),
            .PACKAGEPIN(wb_dat_o[20]));
    defparam wb_dat_o_obuf_20_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_o_obuf_20_preio.PIN_TYPE=6'b011001;
    PRE_IO wb_dat_o_obuf_20_preio (
            .PADOEN(N__55001),
            .PADOUT(N__55000),
            .PADIN(N__54999),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__27616),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_o_obuf_21_iopad (
            .OE(N__54992),
            .DIN(N__54991),
            .DOUT(N__54990),
            .PACKAGEPIN(wb_dat_o[21]));
    defparam wb_dat_o_obuf_21_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_o_obuf_21_preio.PIN_TYPE=6'b011001;
    PRE_IO wb_dat_o_obuf_21_preio (
            .PADOEN(N__54992),
            .PADOUT(N__54991),
            .PADIN(N__54990),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__38101),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_o_obuf_22_iopad (
            .OE(N__54983),
            .DIN(N__54982),
            .DOUT(N__54981),
            .PACKAGEPIN(wb_dat_o[22]));
    defparam wb_dat_o_obuf_22_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_o_obuf_22_preio.PIN_TYPE=6'b011001;
    PRE_IO wb_dat_o_obuf_22_preio (
            .PADOEN(N__54983),
            .PADOUT(N__54982),
            .PADIN(N__54981),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__38905),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_o_obuf_23_iopad (
            .OE(N__54974),
            .DIN(N__54973),
            .DOUT(N__54972),
            .PACKAGEPIN(wb_dat_o[23]));
    defparam wb_dat_o_obuf_23_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_o_obuf_23_preio.PIN_TYPE=6'b011001;
    PRE_IO wb_dat_o_obuf_23_preio (
            .PADOEN(N__54974),
            .PADOUT(N__54973),
            .PADIN(N__54972),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__47554),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_o_obuf_24_iopad (
            .OE(N__54965),
            .DIN(N__54964),
            .DOUT(N__54963),
            .PACKAGEPIN(wb_dat_o[24]));
    defparam wb_dat_o_obuf_24_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_o_obuf_24_preio.PIN_TYPE=6'b011001;
    PRE_IO wb_dat_o_obuf_24_preio (
            .PADOEN(N__54965),
            .PADOUT(N__54964),
            .PADIN(N__54963),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__54493),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_o_obuf_25_iopad (
            .OE(N__54956),
            .DIN(N__54955),
            .DOUT(N__54954),
            .PACKAGEPIN(wb_dat_o[25]));
    defparam wb_dat_o_obuf_25_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_o_obuf_25_preio.PIN_TYPE=6'b011001;
    PRE_IO wb_dat_o_obuf_25_preio (
            .PADOEN(N__54956),
            .PADOUT(N__54955),
            .PADIN(N__54954),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__49129),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_o_obuf_26_iopad (
            .OE(N__54947),
            .DIN(N__54946),
            .DOUT(N__54945),
            .PACKAGEPIN(wb_dat_o[26]));
    defparam wb_dat_o_obuf_26_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_o_obuf_26_preio.PIN_TYPE=6'b011001;
    PRE_IO wb_dat_o_obuf_26_preio (
            .PADOEN(N__54947),
            .PADOUT(N__54946),
            .PADIN(N__54945),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__44260),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_o_obuf_27_iopad (
            .OE(N__54938),
            .DIN(N__54937),
            .DOUT(N__54936),
            .PACKAGEPIN(wb_dat_o[27]));
    defparam wb_dat_o_obuf_27_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_o_obuf_27_preio.PIN_TYPE=6'b011001;
    PRE_IO wb_dat_o_obuf_27_preio (
            .PADOEN(N__54938),
            .PADOUT(N__54937),
            .PADIN(N__54936),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__37735),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_o_obuf_28_iopad (
            .OE(N__54929),
            .DIN(N__54928),
            .DOUT(N__54927),
            .PACKAGEPIN(wb_dat_o[28]));
    defparam wb_dat_o_obuf_28_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_o_obuf_28_preio.PIN_TYPE=6'b011001;
    PRE_IO wb_dat_o_obuf_28_preio (
            .PADOEN(N__54929),
            .PADOUT(N__54928),
            .PADIN(N__54927),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__46450),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_o_obuf_29_iopad (
            .OE(N__54920),
            .DIN(N__54919),
            .DOUT(N__54918),
            .PACKAGEPIN(wb_dat_o[29]));
    defparam wb_dat_o_obuf_29_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_o_obuf_29_preio.PIN_TYPE=6'b011001;
    PRE_IO wb_dat_o_obuf_29_preio (
            .PADOEN(N__54920),
            .PADOUT(N__54919),
            .PADIN(N__54918),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__44362),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_o_obuf_3_iopad (
            .OE(N__54911),
            .DIN(N__54910),
            .DOUT(N__54909),
            .PACKAGEPIN(wb_dat_o[3]));
    defparam wb_dat_o_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_o_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO wb_dat_o_obuf_3_preio (
            .PADOEN(N__54911),
            .PADOUT(N__54910),
            .PADIN(N__54909),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__34924),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_o_obuf_30_iopad (
            .OE(N__54902),
            .DIN(N__54901),
            .DOUT(N__54900),
            .PACKAGEPIN(wb_dat_o[30]));
    defparam wb_dat_o_obuf_30_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_o_obuf_30_preio.PIN_TYPE=6'b011001;
    PRE_IO wb_dat_o_obuf_30_preio (
            .PADOEN(N__54902),
            .PADOUT(N__54901),
            .PADIN(N__54900),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__47857),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_o_obuf_31_iopad (
            .OE(N__54893),
            .DIN(N__54892),
            .DOUT(N__54891),
            .PACKAGEPIN(wb_dat_o[31]));
    defparam wb_dat_o_obuf_31_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_o_obuf_31_preio.PIN_TYPE=6'b011001;
    PRE_IO wb_dat_o_obuf_31_preio (
            .PADOEN(N__54893),
            .PADOUT(N__54892),
            .PADIN(N__54891),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__40384),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_o_obuf_4_iopad (
            .OE(N__54884),
            .DIN(N__54883),
            .DOUT(N__54882),
            .PACKAGEPIN(wb_dat_o[4]));
    defparam wb_dat_o_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_o_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO wb_dat_o_obuf_4_preio (
            .PADOEN(N__54884),
            .PADOUT(N__54883),
            .PADIN(N__54882),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__29893),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_o_obuf_5_iopad (
            .OE(N__54875),
            .DIN(N__54874),
            .DOUT(N__54873),
            .PACKAGEPIN(wb_dat_o[5]));
    defparam wb_dat_o_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_o_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO wb_dat_o_obuf_5_preio (
            .PADOEN(N__54875),
            .PADOUT(N__54874),
            .PADIN(N__54873),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__31930),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_o_obuf_6_iopad (
            .OE(N__54866),
            .DIN(N__54865),
            .DOUT(N__54864),
            .PACKAGEPIN(wb_dat_o[6]));
    defparam wb_dat_o_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_o_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO wb_dat_o_obuf_6_preio (
            .PADOEN(N__54866),
            .PADOUT(N__54865),
            .PADIN(N__54864),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__41062),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_o_obuf_7_iopad (
            .OE(N__54857),
            .DIN(N__54856),
            .DOUT(N__54855),
            .PACKAGEPIN(wb_dat_o[7]));
    defparam wb_dat_o_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_o_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO wb_dat_o_obuf_7_preio (
            .PADOEN(N__54857),
            .PADOUT(N__54856),
            .PADIN(N__54855),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__37876),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_o_obuf_8_iopad (
            .OE(N__54848),
            .DIN(N__54847),
            .DOUT(N__54846),
            .PACKAGEPIN(wb_dat_o[8]));
    defparam wb_dat_o_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_o_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO wb_dat_o_obuf_8_preio (
            .PADOEN(N__54848),
            .PADOUT(N__54847),
            .PADIN(N__54846),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__44503),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_dat_o_obuf_9_iopad (
            .OE(N__54839),
            .DIN(N__54838),
            .DOUT(N__54837),
            .PACKAGEPIN(wb_dat_o[9]));
    defparam wb_dat_o_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam wb_dat_o_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO wb_dat_o_obuf_9_preio (
            .PADOEN(N__54839),
            .PADOUT(N__54838),
            .PADIN(N__54837),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__50227),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_err_o_obuf_iopad (
            .OE(N__54830),
            .DIN(N__54829),
            .DOUT(N__54828),
            .PACKAGEPIN(wb_err_o));
    defparam wb_err_o_obuf_preio.NEG_TRIGGER=1'b0;
    defparam wb_err_o_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO wb_err_o_obuf_preio (
            .PADOEN(N__54830),
            .PADOUT(N__54829),
            .PADIN(N__54828),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__22753),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_inta_o_obuf_iopad (
            .OE(N__54821),
            .DIN(N__54820),
            .DOUT(N__54819),
            .PACKAGEPIN(wb_inta_o));
    defparam wb_inta_o_obuf_preio.NEG_TRIGGER=1'b0;
    defparam wb_inta_o_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO wb_inta_o_obuf_preio (
            .PADOEN(N__54821),
            .PADOUT(N__54820),
            .PADIN(N__54819),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__37095),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_rst_i_ibuf_iopad (
            .OE(N__54812),
            .DIN(N__54811),
            .DOUT(N__54810),
            .PACKAGEPIN(wb_rst_i));
    defparam wb_rst_i_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam wb_rst_i_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_rst_i_ibuf_preio (
            .PADOEN(N__54812),
            .PADOUT(N__54811),
            .PADIN(N__54810),
            .CLOCKENABLE(),
            .DIN0(wb_rst_i_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_rty_o_obuf_iopad (
            .OE(N__54803),
            .DIN(N__54802),
            .DOUT(N__54801),
            .PACKAGEPIN(wb_rty_o));
    defparam wb_rty_o_obuf_preio.NEG_TRIGGER=1'b0;
    defparam wb_rty_o_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO wb_rty_o_obuf_preio (
            .PADOEN(N__54803),
            .PADOUT(N__54802),
            .PADIN(N__54801),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__21625),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_sel_i_ibuf_0_iopad (
            .OE(N__54794),
            .DIN(N__54793),
            .DOUT(N__54792),
            .PACKAGEPIN(wb_sel_i[0]));
    defparam wb_sel_i_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam wb_sel_i_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_sel_i_ibuf_0_preio (
            .PADOEN(N__54794),
            .PADOUT(N__54793),
            .PADIN(N__54792),
            .CLOCKENABLE(),
            .DIN0(wb_sel_i_c_0),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_sel_i_ibuf_1_iopad (
            .OE(N__54785),
            .DIN(N__54784),
            .DOUT(N__54783),
            .PACKAGEPIN(wb_sel_i[1]));
    defparam wb_sel_i_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam wb_sel_i_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_sel_i_ibuf_1_preio (
            .PADOEN(N__54785),
            .PADOUT(N__54784),
            .PADIN(N__54783),
            .CLOCKENABLE(),
            .DIN0(wb_sel_i_c_1),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_sel_i_ibuf_2_iopad (
            .OE(N__54776),
            .DIN(N__54775),
            .DOUT(N__54774),
            .PACKAGEPIN(wb_sel_i[2]));
    defparam wb_sel_i_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam wb_sel_i_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_sel_i_ibuf_2_preio (
            .PADOEN(N__54776),
            .PADOUT(N__54775),
            .PADIN(N__54774),
            .CLOCKENABLE(),
            .DIN0(wb_sel_i_c_2),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_sel_i_ibuf_3_iopad (
            .OE(N__54767),
            .DIN(N__54766),
            .DOUT(N__54765),
            .PACKAGEPIN(wb_sel_i[3]));
    defparam wb_sel_i_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam wb_sel_i_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_sel_i_ibuf_3_preio (
            .PADOEN(N__54767),
            .PADOUT(N__54766),
            .PADIN(N__54765),
            .CLOCKENABLE(),
            .DIN0(wb_sel_i_c_3),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_stb_i_ibuf_iopad (
            .OE(N__54758),
            .DIN(N__54757),
            .DOUT(N__54756),
            .PACKAGEPIN(wb_stb_i));
    defparam wb_stb_i_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam wb_stb_i_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_stb_i_ibuf_preio (
            .PADOEN(N__54758),
            .PADOUT(N__54757),
            .PADIN(N__54756),
            .CLOCKENABLE(),
            .DIN0(wb_stb_i_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD wb_we_i_ibuf_iopad (
            .OE(N__54749),
            .DIN(N__54748),
            .DOUT(N__54747),
            .PACKAGEPIN(wb_we_i));
    defparam wb_we_i_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam wb_we_i_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO wb_we_i_ibuf_preio (
            .PADOEN(N__54749),
            .PADOUT(N__54748),
            .PADIN(N__54747),
            .CLOCKENABLE(),
            .DIN0(wb_we_i_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    InMux I__13692 (
            .O(N__54730),
            .I(N__54727));
    LocalMux I__13691 (
            .O(N__54727),
            .I(N__54724));
    Span4Mux_v I__13690 (
            .O(N__54724),
            .I(N__54721));
    Odrv4 I__13689 (
            .O(N__54721),
            .I(\u0.dat_o_i_i_4_24 ));
    CascadeMux I__13688 (
            .O(N__54718),
            .I(N__54709));
    InMux I__13687 (
            .O(N__54717),
            .I(N__54701));
    CascadeMux I__13686 (
            .O(N__54716),
            .I(N__54698));
    InMux I__13685 (
            .O(N__54715),
            .I(N__54693));
    InMux I__13684 (
            .O(N__54714),
            .I(N__54693));
    InMux I__13683 (
            .O(N__54713),
            .I(N__54690));
    InMux I__13682 (
            .O(N__54712),
            .I(N__54679));
    InMux I__13681 (
            .O(N__54709),
            .I(N__54679));
    InMux I__13680 (
            .O(N__54708),
            .I(N__54679));
    InMux I__13679 (
            .O(N__54707),
            .I(N__54676));
    InMux I__13678 (
            .O(N__54706),
            .I(N__54670));
    InMux I__13677 (
            .O(N__54705),
            .I(N__54667));
    InMux I__13676 (
            .O(N__54704),
            .I(N__54664));
    LocalMux I__13675 (
            .O(N__54701),
            .I(N__54661));
    InMux I__13674 (
            .O(N__54698),
            .I(N__54658));
    LocalMux I__13673 (
            .O(N__54693),
            .I(N__54655));
    LocalMux I__13672 (
            .O(N__54690),
            .I(N__54652));
    InMux I__13671 (
            .O(N__54689),
            .I(N__54643));
    InMux I__13670 (
            .O(N__54688),
            .I(N__54643));
    InMux I__13669 (
            .O(N__54687),
            .I(N__54643));
    InMux I__13668 (
            .O(N__54686),
            .I(N__54643));
    LocalMux I__13667 (
            .O(N__54679),
            .I(N__54638));
    LocalMux I__13666 (
            .O(N__54676),
            .I(N__54638));
    InMux I__13665 (
            .O(N__54675),
            .I(N__54635));
    InMux I__13664 (
            .O(N__54674),
            .I(N__54631));
    InMux I__13663 (
            .O(N__54673),
            .I(N__54626));
    LocalMux I__13662 (
            .O(N__54670),
            .I(N__54621));
    LocalMux I__13661 (
            .O(N__54667),
            .I(N__54621));
    LocalMux I__13660 (
            .O(N__54664),
            .I(N__54618));
    Span4Mux_v I__13659 (
            .O(N__54661),
            .I(N__54613));
    LocalMux I__13658 (
            .O(N__54658),
            .I(N__54613));
    Span4Mux_h I__13657 (
            .O(N__54655),
            .I(N__54606));
    Span4Mux_v I__13656 (
            .O(N__54652),
            .I(N__54606));
    LocalMux I__13655 (
            .O(N__54643),
            .I(N__54606));
    Span4Mux_v I__13654 (
            .O(N__54638),
            .I(N__54601));
    LocalMux I__13653 (
            .O(N__54635),
            .I(N__54601));
    InMux I__13652 (
            .O(N__54634),
            .I(N__54598));
    LocalMux I__13651 (
            .O(N__54631),
            .I(N__54595));
    InMux I__13650 (
            .O(N__54630),
            .I(N__54590));
    InMux I__13649 (
            .O(N__54629),
            .I(N__54590));
    LocalMux I__13648 (
            .O(N__54626),
            .I(N__54584));
    Span4Mux_v I__13647 (
            .O(N__54621),
            .I(N__54575));
    Span4Mux_v I__13646 (
            .O(N__54618),
            .I(N__54575));
    Span4Mux_v I__13645 (
            .O(N__54613),
            .I(N__54575));
    Span4Mux_h I__13644 (
            .O(N__54606),
            .I(N__54575));
    Span4Mux_h I__13643 (
            .O(N__54601),
            .I(N__54570));
    LocalMux I__13642 (
            .O(N__54598),
            .I(N__54570));
    Span4Mux_v I__13641 (
            .O(N__54595),
            .I(N__54565));
    LocalMux I__13640 (
            .O(N__54590),
            .I(N__54565));
    InMux I__13639 (
            .O(N__54589),
            .I(N__54562));
    InMux I__13638 (
            .O(N__54588),
            .I(N__54559));
    InMux I__13637 (
            .O(N__54587),
            .I(N__54556));
    Odrv12 I__13636 (
            .O(N__54584),
            .I(\u0.N_2124 ));
    Odrv4 I__13635 (
            .O(N__54575),
            .I(\u0.N_2124 ));
    Odrv4 I__13634 (
            .O(N__54570),
            .I(\u0.N_2124 ));
    Odrv4 I__13633 (
            .O(N__54565),
            .I(\u0.N_2124 ));
    LocalMux I__13632 (
            .O(N__54562),
            .I(\u0.N_2124 ));
    LocalMux I__13631 (
            .O(N__54559),
            .I(\u0.N_2124 ));
    LocalMux I__13630 (
            .O(N__54556),
            .I(\u0.N_2124 ));
    CascadeMux I__13629 (
            .O(N__54541),
            .I(N__54538));
    InMux I__13628 (
            .O(N__54538),
            .I(N__54535));
    LocalMux I__13627 (
            .O(N__54535),
            .I(N__54532));
    Span4Mux_v I__13626 (
            .O(N__54532),
            .I(N__54529));
    Odrv4 I__13625 (
            .O(N__54529),
            .I(\u0.dat_o_i_i_0_24 ));
    InMux I__13624 (
            .O(N__54526),
            .I(N__54523));
    LocalMux I__13623 (
            .O(N__54523),
            .I(N__54519));
    InMux I__13622 (
            .O(N__54522),
            .I(N__54516));
    Span4Mux_v I__13621 (
            .O(N__54519),
            .I(N__54513));
    LocalMux I__13620 (
            .O(N__54516),
            .I(N__54510));
    Sp12to4 I__13619 (
            .O(N__54513),
            .I(N__54507));
    Span4Mux_s3_h I__13618 (
            .O(N__54510),
            .I(N__54504));
    Span12Mux_h I__13617 (
            .O(N__54507),
            .I(N__54501));
    Span4Mux_h I__13616 (
            .O(N__54504),
            .I(N__54498));
    Odrv12 I__13615 (
            .O(N__54501),
            .I(DMA_dev1_Teoc_0));
    Odrv4 I__13614 (
            .O(N__54498),
            .I(DMA_dev1_Teoc_0));
    IoInMux I__13613 (
            .O(N__54493),
            .I(N__54490));
    LocalMux I__13612 (
            .O(N__54490),
            .I(N__54487));
    Span4Mux_s2_v I__13611 (
            .O(N__54487),
            .I(N__54484));
    Span4Mux_h I__13610 (
            .O(N__54484),
            .I(N__54481));
    Span4Mux_v I__13609 (
            .O(N__54481),
            .I(N__54478));
    Odrv4 I__13608 (
            .O(N__54478),
            .I(N_263));
    InMux I__13607 (
            .O(N__54475),
            .I(N__54472));
    LocalMux I__13606 (
            .O(N__54472),
            .I(N__54469));
    Span4Mux_h I__13605 (
            .O(N__54469),
            .I(N__54462));
    InMux I__13604 (
            .O(N__54468),
            .I(N__54456));
    InMux I__13603 (
            .O(N__54467),
            .I(N__54452));
    InMux I__13602 (
            .O(N__54466),
            .I(N__54449));
    InMux I__13601 (
            .O(N__54465),
            .I(N__54446));
    Span4Mux_h I__13600 (
            .O(N__54462),
            .I(N__54443));
    InMux I__13599 (
            .O(N__54461),
            .I(N__54440));
    InMux I__13598 (
            .O(N__54460),
            .I(N__54437));
    InMux I__13597 (
            .O(N__54459),
            .I(N__54434));
    LocalMux I__13596 (
            .O(N__54456),
            .I(N__54431));
    InMux I__13595 (
            .O(N__54455),
            .I(N__54428));
    LocalMux I__13594 (
            .O(N__54452),
            .I(N__54423));
    LocalMux I__13593 (
            .O(N__54449),
            .I(N__54423));
    LocalMux I__13592 (
            .O(N__54446),
            .I(N__54420));
    Span4Mux_h I__13591 (
            .O(N__54443),
            .I(N__54411));
    LocalMux I__13590 (
            .O(N__54440),
            .I(N__54411));
    LocalMux I__13589 (
            .O(N__54437),
            .I(N__54411));
    LocalMux I__13588 (
            .O(N__54434),
            .I(N__54411));
    Sp12to4 I__13587 (
            .O(N__54431),
            .I(N__54408));
    LocalMux I__13586 (
            .O(N__54428),
            .I(N__54405));
    Span12Mux_s11_v I__13585 (
            .O(N__54423),
            .I(N__54402));
    Span4Mux_h I__13584 (
            .O(N__54420),
            .I(N__54399));
    Span4Mux_v I__13583 (
            .O(N__54411),
            .I(N__54396));
    Span12Mux_v I__13582 (
            .O(N__54408),
            .I(N__54393));
    Span12Mux_s11_v I__13581 (
            .O(N__54405),
            .I(N__54390));
    Span12Mux_v I__13580 (
            .O(N__54402),
            .I(N__54387));
    Sp12to4 I__13579 (
            .O(N__54399),
            .I(N__54384));
    Span4Mux_v I__13578 (
            .O(N__54396),
            .I(N__54381));
    Span12Mux_h I__13577 (
            .O(N__54393),
            .I(N__54376));
    Span12Mux_v I__13576 (
            .O(N__54390),
            .I(N__54376));
    Span12Mux_h I__13575 (
            .O(N__54387),
            .I(N__54369));
    Span12Mux_v I__13574 (
            .O(N__54384),
            .I(N__54369));
    Sp12to4 I__13573 (
            .O(N__54381),
            .I(N__54369));
    Span12Mux_h I__13572 (
            .O(N__54376),
            .I(N__54366));
    Span12Mux_h I__13571 (
            .O(N__54369),
            .I(N__54363));
    Odrv12 I__13570 (
            .O(N__54366),
            .I(wb_dat_i_c_8));
    Odrv12 I__13569 (
            .O(N__54363),
            .I(wb_dat_i_c_8));
    InMux I__13568 (
            .O(N__54358),
            .I(N__54354));
    InMux I__13567 (
            .O(N__54357),
            .I(N__54351));
    LocalMux I__13566 (
            .O(N__54354),
            .I(N__54348));
    LocalMux I__13565 (
            .O(N__54351),
            .I(N__54345));
    Span4Mux_v I__13564 (
            .O(N__54348),
            .I(N__54342));
    Span12Mux_h I__13563 (
            .O(N__54345),
            .I(N__54339));
    Odrv4 I__13562 (
            .O(N__54342),
            .I(DMActrl_BeLeC0));
    Odrv12 I__13561 (
            .O(N__54339),
            .I(DMActrl_BeLeC0));
    ClkMux I__13560 (
            .O(N__54334),
            .I(N__53659));
    ClkMux I__13559 (
            .O(N__54333),
            .I(N__53659));
    ClkMux I__13558 (
            .O(N__54332),
            .I(N__53659));
    ClkMux I__13557 (
            .O(N__54331),
            .I(N__53659));
    ClkMux I__13556 (
            .O(N__54330),
            .I(N__53659));
    ClkMux I__13555 (
            .O(N__54329),
            .I(N__53659));
    ClkMux I__13554 (
            .O(N__54328),
            .I(N__53659));
    ClkMux I__13553 (
            .O(N__54327),
            .I(N__53659));
    ClkMux I__13552 (
            .O(N__54326),
            .I(N__53659));
    ClkMux I__13551 (
            .O(N__54325),
            .I(N__53659));
    ClkMux I__13550 (
            .O(N__54324),
            .I(N__53659));
    ClkMux I__13549 (
            .O(N__54323),
            .I(N__53659));
    ClkMux I__13548 (
            .O(N__54322),
            .I(N__53659));
    ClkMux I__13547 (
            .O(N__54321),
            .I(N__53659));
    ClkMux I__13546 (
            .O(N__54320),
            .I(N__53659));
    ClkMux I__13545 (
            .O(N__54319),
            .I(N__53659));
    ClkMux I__13544 (
            .O(N__54318),
            .I(N__53659));
    ClkMux I__13543 (
            .O(N__54317),
            .I(N__53659));
    ClkMux I__13542 (
            .O(N__54316),
            .I(N__53659));
    ClkMux I__13541 (
            .O(N__54315),
            .I(N__53659));
    ClkMux I__13540 (
            .O(N__54314),
            .I(N__53659));
    ClkMux I__13539 (
            .O(N__54313),
            .I(N__53659));
    ClkMux I__13538 (
            .O(N__54312),
            .I(N__53659));
    ClkMux I__13537 (
            .O(N__54311),
            .I(N__53659));
    ClkMux I__13536 (
            .O(N__54310),
            .I(N__53659));
    ClkMux I__13535 (
            .O(N__54309),
            .I(N__53659));
    ClkMux I__13534 (
            .O(N__54308),
            .I(N__53659));
    ClkMux I__13533 (
            .O(N__54307),
            .I(N__53659));
    ClkMux I__13532 (
            .O(N__54306),
            .I(N__53659));
    ClkMux I__13531 (
            .O(N__54305),
            .I(N__53659));
    ClkMux I__13530 (
            .O(N__54304),
            .I(N__53659));
    ClkMux I__13529 (
            .O(N__54303),
            .I(N__53659));
    ClkMux I__13528 (
            .O(N__54302),
            .I(N__53659));
    ClkMux I__13527 (
            .O(N__54301),
            .I(N__53659));
    ClkMux I__13526 (
            .O(N__54300),
            .I(N__53659));
    ClkMux I__13525 (
            .O(N__54299),
            .I(N__53659));
    ClkMux I__13524 (
            .O(N__54298),
            .I(N__53659));
    ClkMux I__13523 (
            .O(N__54297),
            .I(N__53659));
    ClkMux I__13522 (
            .O(N__54296),
            .I(N__53659));
    ClkMux I__13521 (
            .O(N__54295),
            .I(N__53659));
    ClkMux I__13520 (
            .O(N__54294),
            .I(N__53659));
    ClkMux I__13519 (
            .O(N__54293),
            .I(N__53659));
    ClkMux I__13518 (
            .O(N__54292),
            .I(N__53659));
    ClkMux I__13517 (
            .O(N__54291),
            .I(N__53659));
    ClkMux I__13516 (
            .O(N__54290),
            .I(N__53659));
    ClkMux I__13515 (
            .O(N__54289),
            .I(N__53659));
    ClkMux I__13514 (
            .O(N__54288),
            .I(N__53659));
    ClkMux I__13513 (
            .O(N__54287),
            .I(N__53659));
    ClkMux I__13512 (
            .O(N__54286),
            .I(N__53659));
    ClkMux I__13511 (
            .O(N__54285),
            .I(N__53659));
    ClkMux I__13510 (
            .O(N__54284),
            .I(N__53659));
    ClkMux I__13509 (
            .O(N__54283),
            .I(N__53659));
    ClkMux I__13508 (
            .O(N__54282),
            .I(N__53659));
    ClkMux I__13507 (
            .O(N__54281),
            .I(N__53659));
    ClkMux I__13506 (
            .O(N__54280),
            .I(N__53659));
    ClkMux I__13505 (
            .O(N__54279),
            .I(N__53659));
    ClkMux I__13504 (
            .O(N__54278),
            .I(N__53659));
    ClkMux I__13503 (
            .O(N__54277),
            .I(N__53659));
    ClkMux I__13502 (
            .O(N__54276),
            .I(N__53659));
    ClkMux I__13501 (
            .O(N__54275),
            .I(N__53659));
    ClkMux I__13500 (
            .O(N__54274),
            .I(N__53659));
    ClkMux I__13499 (
            .O(N__54273),
            .I(N__53659));
    ClkMux I__13498 (
            .O(N__54272),
            .I(N__53659));
    ClkMux I__13497 (
            .O(N__54271),
            .I(N__53659));
    ClkMux I__13496 (
            .O(N__54270),
            .I(N__53659));
    ClkMux I__13495 (
            .O(N__54269),
            .I(N__53659));
    ClkMux I__13494 (
            .O(N__54268),
            .I(N__53659));
    ClkMux I__13493 (
            .O(N__54267),
            .I(N__53659));
    ClkMux I__13492 (
            .O(N__54266),
            .I(N__53659));
    ClkMux I__13491 (
            .O(N__54265),
            .I(N__53659));
    ClkMux I__13490 (
            .O(N__54264),
            .I(N__53659));
    ClkMux I__13489 (
            .O(N__54263),
            .I(N__53659));
    ClkMux I__13488 (
            .O(N__54262),
            .I(N__53659));
    ClkMux I__13487 (
            .O(N__54261),
            .I(N__53659));
    ClkMux I__13486 (
            .O(N__54260),
            .I(N__53659));
    ClkMux I__13485 (
            .O(N__54259),
            .I(N__53659));
    ClkMux I__13484 (
            .O(N__54258),
            .I(N__53659));
    ClkMux I__13483 (
            .O(N__54257),
            .I(N__53659));
    ClkMux I__13482 (
            .O(N__54256),
            .I(N__53659));
    ClkMux I__13481 (
            .O(N__54255),
            .I(N__53659));
    ClkMux I__13480 (
            .O(N__54254),
            .I(N__53659));
    ClkMux I__13479 (
            .O(N__54253),
            .I(N__53659));
    ClkMux I__13478 (
            .O(N__54252),
            .I(N__53659));
    ClkMux I__13477 (
            .O(N__54251),
            .I(N__53659));
    ClkMux I__13476 (
            .O(N__54250),
            .I(N__53659));
    ClkMux I__13475 (
            .O(N__54249),
            .I(N__53659));
    ClkMux I__13474 (
            .O(N__54248),
            .I(N__53659));
    ClkMux I__13473 (
            .O(N__54247),
            .I(N__53659));
    ClkMux I__13472 (
            .O(N__54246),
            .I(N__53659));
    ClkMux I__13471 (
            .O(N__54245),
            .I(N__53659));
    ClkMux I__13470 (
            .O(N__54244),
            .I(N__53659));
    ClkMux I__13469 (
            .O(N__54243),
            .I(N__53659));
    ClkMux I__13468 (
            .O(N__54242),
            .I(N__53659));
    ClkMux I__13467 (
            .O(N__54241),
            .I(N__53659));
    ClkMux I__13466 (
            .O(N__54240),
            .I(N__53659));
    ClkMux I__13465 (
            .O(N__54239),
            .I(N__53659));
    ClkMux I__13464 (
            .O(N__54238),
            .I(N__53659));
    ClkMux I__13463 (
            .O(N__54237),
            .I(N__53659));
    ClkMux I__13462 (
            .O(N__54236),
            .I(N__53659));
    ClkMux I__13461 (
            .O(N__54235),
            .I(N__53659));
    ClkMux I__13460 (
            .O(N__54234),
            .I(N__53659));
    ClkMux I__13459 (
            .O(N__54233),
            .I(N__53659));
    ClkMux I__13458 (
            .O(N__54232),
            .I(N__53659));
    ClkMux I__13457 (
            .O(N__54231),
            .I(N__53659));
    ClkMux I__13456 (
            .O(N__54230),
            .I(N__53659));
    ClkMux I__13455 (
            .O(N__54229),
            .I(N__53659));
    ClkMux I__13454 (
            .O(N__54228),
            .I(N__53659));
    ClkMux I__13453 (
            .O(N__54227),
            .I(N__53659));
    ClkMux I__13452 (
            .O(N__54226),
            .I(N__53659));
    ClkMux I__13451 (
            .O(N__54225),
            .I(N__53659));
    ClkMux I__13450 (
            .O(N__54224),
            .I(N__53659));
    ClkMux I__13449 (
            .O(N__54223),
            .I(N__53659));
    ClkMux I__13448 (
            .O(N__54222),
            .I(N__53659));
    ClkMux I__13447 (
            .O(N__54221),
            .I(N__53659));
    ClkMux I__13446 (
            .O(N__54220),
            .I(N__53659));
    ClkMux I__13445 (
            .O(N__54219),
            .I(N__53659));
    ClkMux I__13444 (
            .O(N__54218),
            .I(N__53659));
    ClkMux I__13443 (
            .O(N__54217),
            .I(N__53659));
    ClkMux I__13442 (
            .O(N__54216),
            .I(N__53659));
    ClkMux I__13441 (
            .O(N__54215),
            .I(N__53659));
    ClkMux I__13440 (
            .O(N__54214),
            .I(N__53659));
    ClkMux I__13439 (
            .O(N__54213),
            .I(N__53659));
    ClkMux I__13438 (
            .O(N__54212),
            .I(N__53659));
    ClkMux I__13437 (
            .O(N__54211),
            .I(N__53659));
    ClkMux I__13436 (
            .O(N__54210),
            .I(N__53659));
    ClkMux I__13435 (
            .O(N__54209),
            .I(N__53659));
    ClkMux I__13434 (
            .O(N__54208),
            .I(N__53659));
    ClkMux I__13433 (
            .O(N__54207),
            .I(N__53659));
    ClkMux I__13432 (
            .O(N__54206),
            .I(N__53659));
    ClkMux I__13431 (
            .O(N__54205),
            .I(N__53659));
    ClkMux I__13430 (
            .O(N__54204),
            .I(N__53659));
    ClkMux I__13429 (
            .O(N__54203),
            .I(N__53659));
    ClkMux I__13428 (
            .O(N__54202),
            .I(N__53659));
    ClkMux I__13427 (
            .O(N__54201),
            .I(N__53659));
    ClkMux I__13426 (
            .O(N__54200),
            .I(N__53659));
    ClkMux I__13425 (
            .O(N__54199),
            .I(N__53659));
    ClkMux I__13424 (
            .O(N__54198),
            .I(N__53659));
    ClkMux I__13423 (
            .O(N__54197),
            .I(N__53659));
    ClkMux I__13422 (
            .O(N__54196),
            .I(N__53659));
    ClkMux I__13421 (
            .O(N__54195),
            .I(N__53659));
    ClkMux I__13420 (
            .O(N__54194),
            .I(N__53659));
    ClkMux I__13419 (
            .O(N__54193),
            .I(N__53659));
    ClkMux I__13418 (
            .O(N__54192),
            .I(N__53659));
    ClkMux I__13417 (
            .O(N__54191),
            .I(N__53659));
    ClkMux I__13416 (
            .O(N__54190),
            .I(N__53659));
    ClkMux I__13415 (
            .O(N__54189),
            .I(N__53659));
    ClkMux I__13414 (
            .O(N__54188),
            .I(N__53659));
    ClkMux I__13413 (
            .O(N__54187),
            .I(N__53659));
    ClkMux I__13412 (
            .O(N__54186),
            .I(N__53659));
    ClkMux I__13411 (
            .O(N__54185),
            .I(N__53659));
    ClkMux I__13410 (
            .O(N__54184),
            .I(N__53659));
    ClkMux I__13409 (
            .O(N__54183),
            .I(N__53659));
    ClkMux I__13408 (
            .O(N__54182),
            .I(N__53659));
    ClkMux I__13407 (
            .O(N__54181),
            .I(N__53659));
    ClkMux I__13406 (
            .O(N__54180),
            .I(N__53659));
    ClkMux I__13405 (
            .O(N__54179),
            .I(N__53659));
    ClkMux I__13404 (
            .O(N__54178),
            .I(N__53659));
    ClkMux I__13403 (
            .O(N__54177),
            .I(N__53659));
    ClkMux I__13402 (
            .O(N__54176),
            .I(N__53659));
    ClkMux I__13401 (
            .O(N__54175),
            .I(N__53659));
    ClkMux I__13400 (
            .O(N__54174),
            .I(N__53659));
    ClkMux I__13399 (
            .O(N__54173),
            .I(N__53659));
    ClkMux I__13398 (
            .O(N__54172),
            .I(N__53659));
    ClkMux I__13397 (
            .O(N__54171),
            .I(N__53659));
    ClkMux I__13396 (
            .O(N__54170),
            .I(N__53659));
    ClkMux I__13395 (
            .O(N__54169),
            .I(N__53659));
    ClkMux I__13394 (
            .O(N__54168),
            .I(N__53659));
    ClkMux I__13393 (
            .O(N__54167),
            .I(N__53659));
    ClkMux I__13392 (
            .O(N__54166),
            .I(N__53659));
    ClkMux I__13391 (
            .O(N__54165),
            .I(N__53659));
    ClkMux I__13390 (
            .O(N__54164),
            .I(N__53659));
    ClkMux I__13389 (
            .O(N__54163),
            .I(N__53659));
    ClkMux I__13388 (
            .O(N__54162),
            .I(N__53659));
    ClkMux I__13387 (
            .O(N__54161),
            .I(N__53659));
    ClkMux I__13386 (
            .O(N__54160),
            .I(N__53659));
    ClkMux I__13385 (
            .O(N__54159),
            .I(N__53659));
    ClkMux I__13384 (
            .O(N__54158),
            .I(N__53659));
    ClkMux I__13383 (
            .O(N__54157),
            .I(N__53659));
    ClkMux I__13382 (
            .O(N__54156),
            .I(N__53659));
    ClkMux I__13381 (
            .O(N__54155),
            .I(N__53659));
    ClkMux I__13380 (
            .O(N__54154),
            .I(N__53659));
    ClkMux I__13379 (
            .O(N__54153),
            .I(N__53659));
    ClkMux I__13378 (
            .O(N__54152),
            .I(N__53659));
    ClkMux I__13377 (
            .O(N__54151),
            .I(N__53659));
    ClkMux I__13376 (
            .O(N__54150),
            .I(N__53659));
    ClkMux I__13375 (
            .O(N__54149),
            .I(N__53659));
    ClkMux I__13374 (
            .O(N__54148),
            .I(N__53659));
    ClkMux I__13373 (
            .O(N__54147),
            .I(N__53659));
    ClkMux I__13372 (
            .O(N__54146),
            .I(N__53659));
    ClkMux I__13371 (
            .O(N__54145),
            .I(N__53659));
    ClkMux I__13370 (
            .O(N__54144),
            .I(N__53659));
    ClkMux I__13369 (
            .O(N__54143),
            .I(N__53659));
    ClkMux I__13368 (
            .O(N__54142),
            .I(N__53659));
    ClkMux I__13367 (
            .O(N__54141),
            .I(N__53659));
    ClkMux I__13366 (
            .O(N__54140),
            .I(N__53659));
    ClkMux I__13365 (
            .O(N__54139),
            .I(N__53659));
    ClkMux I__13364 (
            .O(N__54138),
            .I(N__53659));
    ClkMux I__13363 (
            .O(N__54137),
            .I(N__53659));
    ClkMux I__13362 (
            .O(N__54136),
            .I(N__53659));
    ClkMux I__13361 (
            .O(N__54135),
            .I(N__53659));
    ClkMux I__13360 (
            .O(N__54134),
            .I(N__53659));
    ClkMux I__13359 (
            .O(N__54133),
            .I(N__53659));
    ClkMux I__13358 (
            .O(N__54132),
            .I(N__53659));
    ClkMux I__13357 (
            .O(N__54131),
            .I(N__53659));
    ClkMux I__13356 (
            .O(N__54130),
            .I(N__53659));
    ClkMux I__13355 (
            .O(N__54129),
            .I(N__53659));
    ClkMux I__13354 (
            .O(N__54128),
            .I(N__53659));
    ClkMux I__13353 (
            .O(N__54127),
            .I(N__53659));
    ClkMux I__13352 (
            .O(N__54126),
            .I(N__53659));
    ClkMux I__13351 (
            .O(N__54125),
            .I(N__53659));
    ClkMux I__13350 (
            .O(N__54124),
            .I(N__53659));
    ClkMux I__13349 (
            .O(N__54123),
            .I(N__53659));
    ClkMux I__13348 (
            .O(N__54122),
            .I(N__53659));
    ClkMux I__13347 (
            .O(N__54121),
            .I(N__53659));
    ClkMux I__13346 (
            .O(N__54120),
            .I(N__53659));
    ClkMux I__13345 (
            .O(N__54119),
            .I(N__53659));
    ClkMux I__13344 (
            .O(N__54118),
            .I(N__53659));
    ClkMux I__13343 (
            .O(N__54117),
            .I(N__53659));
    ClkMux I__13342 (
            .O(N__54116),
            .I(N__53659));
    ClkMux I__13341 (
            .O(N__54115),
            .I(N__53659));
    ClkMux I__13340 (
            .O(N__54114),
            .I(N__53659));
    ClkMux I__13339 (
            .O(N__54113),
            .I(N__53659));
    ClkMux I__13338 (
            .O(N__54112),
            .I(N__53659));
    ClkMux I__13337 (
            .O(N__54111),
            .I(N__53659));
    ClkMux I__13336 (
            .O(N__54110),
            .I(N__53659));
    GlobalMux I__13335 (
            .O(N__53659),
            .I(N__53656));
    gio2CtrlBuf I__13334 (
            .O(N__53656),
            .I(wb_clk_i_c_g));
    CEMux I__13333 (
            .O(N__53653),
            .I(N__53648));
    CEMux I__13332 (
            .O(N__53652),
            .I(N__53638));
    CEMux I__13331 (
            .O(N__53651),
            .I(N__53635));
    LocalMux I__13330 (
            .O(N__53648),
            .I(N__53631));
    CEMux I__13329 (
            .O(N__53647),
            .I(N__53628));
    CEMux I__13328 (
            .O(N__53646),
            .I(N__53625));
    CEMux I__13327 (
            .O(N__53645),
            .I(N__53622));
    CEMux I__13326 (
            .O(N__53644),
            .I(N__53619));
    CEMux I__13325 (
            .O(N__53643),
            .I(N__53616));
    CEMux I__13324 (
            .O(N__53642),
            .I(N__53611));
    CEMux I__13323 (
            .O(N__53641),
            .I(N__53607));
    LocalMux I__13322 (
            .O(N__53638),
            .I(N__53601));
    LocalMux I__13321 (
            .O(N__53635),
            .I(N__53601));
    CEMux I__13320 (
            .O(N__53634),
            .I(N__53598));
    Span4Mux_v I__13319 (
            .O(N__53631),
            .I(N__53591));
    LocalMux I__13318 (
            .O(N__53628),
            .I(N__53591));
    LocalMux I__13317 (
            .O(N__53625),
            .I(N__53591));
    LocalMux I__13316 (
            .O(N__53622),
            .I(N__53588));
    LocalMux I__13315 (
            .O(N__53619),
            .I(N__53582));
    LocalMux I__13314 (
            .O(N__53616),
            .I(N__53582));
    CEMux I__13313 (
            .O(N__53615),
            .I(N__53579));
    CEMux I__13312 (
            .O(N__53614),
            .I(N__53576));
    LocalMux I__13311 (
            .O(N__53611),
            .I(N__53572));
    CEMux I__13310 (
            .O(N__53610),
            .I(N__53569));
    LocalMux I__13309 (
            .O(N__53607),
            .I(N__53566));
    CEMux I__13308 (
            .O(N__53606),
            .I(N__53562));
    Span4Mux_v I__13307 (
            .O(N__53601),
            .I(N__53555));
    LocalMux I__13306 (
            .O(N__53598),
            .I(N__53555));
    Span4Mux_v I__13305 (
            .O(N__53591),
            .I(N__53550));
    Span4Mux_v I__13304 (
            .O(N__53588),
            .I(N__53550));
    CEMux I__13303 (
            .O(N__53587),
            .I(N__53546));
    Span4Mux_v I__13302 (
            .O(N__53582),
            .I(N__53539));
    LocalMux I__13301 (
            .O(N__53579),
            .I(N__53539));
    LocalMux I__13300 (
            .O(N__53576),
            .I(N__53539));
    CEMux I__13299 (
            .O(N__53575),
            .I(N__53536));
    Span4Mux_h I__13298 (
            .O(N__53572),
            .I(N__53531));
    LocalMux I__13297 (
            .O(N__53569),
            .I(N__53531));
    Span4Mux_v I__13296 (
            .O(N__53566),
            .I(N__53527));
    CEMux I__13295 (
            .O(N__53565),
            .I(N__53524));
    LocalMux I__13294 (
            .O(N__53562),
            .I(N__53521));
    CEMux I__13293 (
            .O(N__53561),
            .I(N__53518));
    CEMux I__13292 (
            .O(N__53560),
            .I(N__53515));
    Span4Mux_v I__13291 (
            .O(N__53555),
            .I(N__53510));
    Span4Mux_h I__13290 (
            .O(N__53550),
            .I(N__53507));
    CEMux I__13289 (
            .O(N__53549),
            .I(N__53504));
    LocalMux I__13288 (
            .O(N__53546),
            .I(N__53501));
    Span4Mux_v I__13287 (
            .O(N__53539),
            .I(N__53496));
    LocalMux I__13286 (
            .O(N__53536),
            .I(N__53496));
    Span4Mux_h I__13285 (
            .O(N__53531),
            .I(N__53493));
    CEMux I__13284 (
            .O(N__53530),
            .I(N__53490));
    Span4Mux_h I__13283 (
            .O(N__53527),
            .I(N__53487));
    LocalMux I__13282 (
            .O(N__53524),
            .I(N__53484));
    Span4Mux_h I__13281 (
            .O(N__53521),
            .I(N__53477));
    LocalMux I__13280 (
            .O(N__53518),
            .I(N__53477));
    LocalMux I__13279 (
            .O(N__53515),
            .I(N__53477));
    CEMux I__13278 (
            .O(N__53514),
            .I(N__53474));
    CEMux I__13277 (
            .O(N__53513),
            .I(N__53471));
    Span4Mux_h I__13276 (
            .O(N__53510),
            .I(N__53464));
    Span4Mux_v I__13275 (
            .O(N__53507),
            .I(N__53464));
    LocalMux I__13274 (
            .O(N__53504),
            .I(N__53464));
    Span4Mux_h I__13273 (
            .O(N__53501),
            .I(N__53459));
    Span4Mux_v I__13272 (
            .O(N__53496),
            .I(N__53459));
    Span4Mux_v I__13271 (
            .O(N__53493),
            .I(N__53454));
    LocalMux I__13270 (
            .O(N__53490),
            .I(N__53454));
    Span4Mux_h I__13269 (
            .O(N__53487),
            .I(N__53447));
    Span4Mux_h I__13268 (
            .O(N__53484),
            .I(N__53447));
    Span4Mux_v I__13267 (
            .O(N__53477),
            .I(N__53447));
    LocalMux I__13266 (
            .O(N__53474),
            .I(N__53444));
    LocalMux I__13265 (
            .O(N__53471),
            .I(N__53441));
    Span4Mux_h I__13264 (
            .O(N__53464),
            .I(N__53438));
    Span4Mux_h I__13263 (
            .O(N__53459),
            .I(N__53433));
    Span4Mux_v I__13262 (
            .O(N__53454),
            .I(N__53433));
    Sp12to4 I__13261 (
            .O(N__53447),
            .I(N__53430));
    Span4Mux_h I__13260 (
            .O(N__53444),
            .I(N__53425));
    Span4Mux_v I__13259 (
            .O(N__53441),
            .I(N__53425));
    Span4Mux_v I__13258 (
            .O(N__53438),
            .I(N__53422));
    Odrv4 I__13257 (
            .O(N__53433),
            .I(\u0.N_286 ));
    Odrv12 I__13256 (
            .O(N__53430),
            .I(\u0.N_286 ));
    Odrv4 I__13255 (
            .O(N__53425),
            .I(\u0.N_286 ));
    Odrv4 I__13254 (
            .O(N__53422),
            .I(\u0.N_286 ));
    SRMux I__13253 (
            .O(N__53413),
            .I(N__53086));
    SRMux I__13252 (
            .O(N__53412),
            .I(N__53086));
    SRMux I__13251 (
            .O(N__53411),
            .I(N__53086));
    SRMux I__13250 (
            .O(N__53410),
            .I(N__53086));
    SRMux I__13249 (
            .O(N__53409),
            .I(N__53086));
    SRMux I__13248 (
            .O(N__53408),
            .I(N__53086));
    SRMux I__13247 (
            .O(N__53407),
            .I(N__53086));
    SRMux I__13246 (
            .O(N__53406),
            .I(N__53086));
    SRMux I__13245 (
            .O(N__53405),
            .I(N__53086));
    SRMux I__13244 (
            .O(N__53404),
            .I(N__53086));
    SRMux I__13243 (
            .O(N__53403),
            .I(N__53086));
    SRMux I__13242 (
            .O(N__53402),
            .I(N__53086));
    SRMux I__13241 (
            .O(N__53401),
            .I(N__53086));
    SRMux I__13240 (
            .O(N__53400),
            .I(N__53086));
    SRMux I__13239 (
            .O(N__53399),
            .I(N__53086));
    SRMux I__13238 (
            .O(N__53398),
            .I(N__53086));
    SRMux I__13237 (
            .O(N__53397),
            .I(N__53086));
    SRMux I__13236 (
            .O(N__53396),
            .I(N__53086));
    SRMux I__13235 (
            .O(N__53395),
            .I(N__53086));
    SRMux I__13234 (
            .O(N__53394),
            .I(N__53086));
    SRMux I__13233 (
            .O(N__53393),
            .I(N__53086));
    SRMux I__13232 (
            .O(N__53392),
            .I(N__53086));
    SRMux I__13231 (
            .O(N__53391),
            .I(N__53086));
    SRMux I__13230 (
            .O(N__53390),
            .I(N__53086));
    SRMux I__13229 (
            .O(N__53389),
            .I(N__53086));
    SRMux I__13228 (
            .O(N__53388),
            .I(N__53086));
    SRMux I__13227 (
            .O(N__53387),
            .I(N__53086));
    SRMux I__13226 (
            .O(N__53386),
            .I(N__53086));
    SRMux I__13225 (
            .O(N__53385),
            .I(N__53086));
    SRMux I__13224 (
            .O(N__53384),
            .I(N__53086));
    SRMux I__13223 (
            .O(N__53383),
            .I(N__53086));
    SRMux I__13222 (
            .O(N__53382),
            .I(N__53086));
    SRMux I__13221 (
            .O(N__53381),
            .I(N__53086));
    SRMux I__13220 (
            .O(N__53380),
            .I(N__53086));
    SRMux I__13219 (
            .O(N__53379),
            .I(N__53086));
    SRMux I__13218 (
            .O(N__53378),
            .I(N__53086));
    SRMux I__13217 (
            .O(N__53377),
            .I(N__53086));
    SRMux I__13216 (
            .O(N__53376),
            .I(N__53086));
    SRMux I__13215 (
            .O(N__53375),
            .I(N__53086));
    SRMux I__13214 (
            .O(N__53374),
            .I(N__53086));
    SRMux I__13213 (
            .O(N__53373),
            .I(N__53086));
    SRMux I__13212 (
            .O(N__53372),
            .I(N__53086));
    SRMux I__13211 (
            .O(N__53371),
            .I(N__53086));
    SRMux I__13210 (
            .O(N__53370),
            .I(N__53086));
    SRMux I__13209 (
            .O(N__53369),
            .I(N__53086));
    SRMux I__13208 (
            .O(N__53368),
            .I(N__53086));
    SRMux I__13207 (
            .O(N__53367),
            .I(N__53086));
    SRMux I__13206 (
            .O(N__53366),
            .I(N__53086));
    SRMux I__13205 (
            .O(N__53365),
            .I(N__53086));
    SRMux I__13204 (
            .O(N__53364),
            .I(N__53086));
    SRMux I__13203 (
            .O(N__53363),
            .I(N__53086));
    SRMux I__13202 (
            .O(N__53362),
            .I(N__53086));
    SRMux I__13201 (
            .O(N__53361),
            .I(N__53086));
    SRMux I__13200 (
            .O(N__53360),
            .I(N__53086));
    SRMux I__13199 (
            .O(N__53359),
            .I(N__53086));
    SRMux I__13198 (
            .O(N__53358),
            .I(N__53086));
    SRMux I__13197 (
            .O(N__53357),
            .I(N__53086));
    SRMux I__13196 (
            .O(N__53356),
            .I(N__53086));
    SRMux I__13195 (
            .O(N__53355),
            .I(N__53086));
    SRMux I__13194 (
            .O(N__53354),
            .I(N__53086));
    SRMux I__13193 (
            .O(N__53353),
            .I(N__53086));
    SRMux I__13192 (
            .O(N__53352),
            .I(N__53086));
    SRMux I__13191 (
            .O(N__53351),
            .I(N__53086));
    SRMux I__13190 (
            .O(N__53350),
            .I(N__53086));
    SRMux I__13189 (
            .O(N__53349),
            .I(N__53086));
    SRMux I__13188 (
            .O(N__53348),
            .I(N__53086));
    SRMux I__13187 (
            .O(N__53347),
            .I(N__53086));
    SRMux I__13186 (
            .O(N__53346),
            .I(N__53086));
    SRMux I__13185 (
            .O(N__53345),
            .I(N__53086));
    SRMux I__13184 (
            .O(N__53344),
            .I(N__53086));
    SRMux I__13183 (
            .O(N__53343),
            .I(N__53086));
    SRMux I__13182 (
            .O(N__53342),
            .I(N__53086));
    SRMux I__13181 (
            .O(N__53341),
            .I(N__53086));
    SRMux I__13180 (
            .O(N__53340),
            .I(N__53086));
    SRMux I__13179 (
            .O(N__53339),
            .I(N__53086));
    SRMux I__13178 (
            .O(N__53338),
            .I(N__53086));
    SRMux I__13177 (
            .O(N__53337),
            .I(N__53086));
    SRMux I__13176 (
            .O(N__53336),
            .I(N__53086));
    SRMux I__13175 (
            .O(N__53335),
            .I(N__53086));
    SRMux I__13174 (
            .O(N__53334),
            .I(N__53086));
    SRMux I__13173 (
            .O(N__53333),
            .I(N__53086));
    SRMux I__13172 (
            .O(N__53332),
            .I(N__53086));
    SRMux I__13171 (
            .O(N__53331),
            .I(N__53086));
    SRMux I__13170 (
            .O(N__53330),
            .I(N__53086));
    SRMux I__13169 (
            .O(N__53329),
            .I(N__53086));
    SRMux I__13168 (
            .O(N__53328),
            .I(N__53086));
    SRMux I__13167 (
            .O(N__53327),
            .I(N__53086));
    SRMux I__13166 (
            .O(N__53326),
            .I(N__53086));
    SRMux I__13165 (
            .O(N__53325),
            .I(N__53086));
    SRMux I__13164 (
            .O(N__53324),
            .I(N__53086));
    SRMux I__13163 (
            .O(N__53323),
            .I(N__53086));
    SRMux I__13162 (
            .O(N__53322),
            .I(N__53086));
    SRMux I__13161 (
            .O(N__53321),
            .I(N__53086));
    SRMux I__13160 (
            .O(N__53320),
            .I(N__53086));
    SRMux I__13159 (
            .O(N__53319),
            .I(N__53086));
    SRMux I__13158 (
            .O(N__53318),
            .I(N__53086));
    SRMux I__13157 (
            .O(N__53317),
            .I(N__53086));
    SRMux I__13156 (
            .O(N__53316),
            .I(N__53086));
    SRMux I__13155 (
            .O(N__53315),
            .I(N__53086));
    SRMux I__13154 (
            .O(N__53314),
            .I(N__53086));
    SRMux I__13153 (
            .O(N__53313),
            .I(N__53086));
    SRMux I__13152 (
            .O(N__53312),
            .I(N__53086));
    SRMux I__13151 (
            .O(N__53311),
            .I(N__53086));
    SRMux I__13150 (
            .O(N__53310),
            .I(N__53086));
    SRMux I__13149 (
            .O(N__53309),
            .I(N__53086));
    SRMux I__13148 (
            .O(N__53308),
            .I(N__53086));
    SRMux I__13147 (
            .O(N__53307),
            .I(N__53086));
    SRMux I__13146 (
            .O(N__53306),
            .I(N__53086));
    SRMux I__13145 (
            .O(N__53305),
            .I(N__53086));
    GlobalMux I__13144 (
            .O(N__53086),
            .I(N__53083));
    gio2CtrlBuf I__13143 (
            .O(N__53083),
            .I(arst_i_c_i_g));
    CascadeMux I__13142 (
            .O(N__53080),
            .I(N__53074));
    CascadeMux I__13141 (
            .O(N__53079),
            .I(N__53071));
    CascadeMux I__13140 (
            .O(N__53078),
            .I(N__53062));
    CascadeMux I__13139 (
            .O(N__53077),
            .I(N__53059));
    InMux I__13138 (
            .O(N__53074),
            .I(N__53047));
    InMux I__13137 (
            .O(N__53071),
            .I(N__53047));
    InMux I__13136 (
            .O(N__53070),
            .I(N__53047));
    InMux I__13135 (
            .O(N__53069),
            .I(N__53047));
    InMux I__13134 (
            .O(N__53068),
            .I(N__53044));
    InMux I__13133 (
            .O(N__53067),
            .I(N__53041));
    InMux I__13132 (
            .O(N__53066),
            .I(N__53038));
    InMux I__13131 (
            .O(N__53065),
            .I(N__53031));
    InMux I__13130 (
            .O(N__53062),
            .I(N__53031));
    InMux I__13129 (
            .O(N__53059),
            .I(N__53031));
    InMux I__13128 (
            .O(N__53058),
            .I(N__53028));
    CascadeMux I__13127 (
            .O(N__53057),
            .I(N__53025));
    CascadeMux I__13126 (
            .O(N__53056),
            .I(N__53020));
    LocalMux I__13125 (
            .O(N__53047),
            .I(N__53016));
    LocalMux I__13124 (
            .O(N__53044),
            .I(N__53012));
    LocalMux I__13123 (
            .O(N__53041),
            .I(N__53007));
    LocalMux I__13122 (
            .O(N__53038),
            .I(N__53007));
    LocalMux I__13121 (
            .O(N__53031),
            .I(N__53003));
    LocalMux I__13120 (
            .O(N__53028),
            .I(N__53000));
    InMux I__13119 (
            .O(N__53025),
            .I(N__52991));
    InMux I__13118 (
            .O(N__53024),
            .I(N__52991));
    InMux I__13117 (
            .O(N__53023),
            .I(N__52991));
    InMux I__13116 (
            .O(N__53020),
            .I(N__52991));
    InMux I__13115 (
            .O(N__53019),
            .I(N__52988));
    Span4Mux_v I__13114 (
            .O(N__53016),
            .I(N__52985));
    InMux I__13113 (
            .O(N__53015),
            .I(N__52982));
    Span4Mux_v I__13112 (
            .O(N__53012),
            .I(N__52979));
    Span4Mux_v I__13111 (
            .O(N__53007),
            .I(N__52976));
    InMux I__13110 (
            .O(N__53006),
            .I(N__52973));
    Span4Mux_v I__13109 (
            .O(N__53003),
            .I(N__52964));
    Span4Mux_v I__13108 (
            .O(N__53000),
            .I(N__52964));
    LocalMux I__13107 (
            .O(N__52991),
            .I(N__52964));
    LocalMux I__13106 (
            .O(N__52988),
            .I(N__52964));
    Span4Mux_h I__13105 (
            .O(N__52985),
            .I(N__52959));
    LocalMux I__13104 (
            .O(N__52982),
            .I(N__52959));
    Sp12to4 I__13103 (
            .O(N__52979),
            .I(N__52956));
    Sp12to4 I__13102 (
            .O(N__52976),
            .I(N__52951));
    LocalMux I__13101 (
            .O(N__52973),
            .I(N__52951));
    Span4Mux_v I__13100 (
            .O(N__52964),
            .I(N__52948));
    Span4Mux_v I__13099 (
            .O(N__52959),
            .I(N__52945));
    Span12Mux_h I__13098 (
            .O(N__52956),
            .I(N__52942));
    Span12Mux_h I__13097 (
            .O(N__52951),
            .I(N__52939));
    Sp12to4 I__13096 (
            .O(N__52948),
            .I(N__52934));
    Sp12to4 I__13095 (
            .O(N__52945),
            .I(N__52934));
    Span12Mux_v I__13094 (
            .O(N__52942),
            .I(N__52931));
    Span12Mux_v I__13093 (
            .O(N__52939),
            .I(N__52928));
    Span12Mux_h I__13092 (
            .O(N__52934),
            .I(N__52925));
    Span12Mux_h I__13091 (
            .O(N__52931),
            .I(N__52922));
    Span12Mux_h I__13090 (
            .O(N__52928),
            .I(N__52917));
    Span12Mux_v I__13089 (
            .O(N__52925),
            .I(N__52917));
    Odrv12 I__13088 (
            .O(N__52922),
            .I(wb_adr_i_c_4));
    Odrv12 I__13087 (
            .O(N__52917),
            .I(wb_adr_i_c_4));
    InMux I__13086 (
            .O(N__52912),
            .I(N__52904));
    InMux I__13085 (
            .O(N__52911),
            .I(N__52893));
    InMux I__13084 (
            .O(N__52910),
            .I(N__52893));
    InMux I__13083 (
            .O(N__52909),
            .I(N__52893));
    InMux I__13082 (
            .O(N__52908),
            .I(N__52893));
    InMux I__13081 (
            .O(N__52907),
            .I(N__52893));
    LocalMux I__13080 (
            .O(N__52904),
            .I(N__52888));
    LocalMux I__13079 (
            .O(N__52893),
            .I(N__52888));
    Span4Mux_v I__13078 (
            .O(N__52888),
            .I(N__52883));
    InMux I__13077 (
            .O(N__52887),
            .I(N__52880));
    InMux I__13076 (
            .O(N__52886),
            .I(N__52877));
    Span4Mux_h I__13075 (
            .O(N__52883),
            .I(N__52874));
    LocalMux I__13074 (
            .O(N__52880),
            .I(N__52869));
    LocalMux I__13073 (
            .O(N__52877),
            .I(N__52869));
    Odrv4 I__13072 (
            .O(N__52874),
            .I(\u0.N_2139 ));
    Odrv4 I__13071 (
            .O(N__52869),
            .I(\u0.N_2139 ));
    CascadeMux I__13070 (
            .O(N__52864),
            .I(N__52861));
    InMux I__13069 (
            .O(N__52861),
            .I(N__52857));
    CascadeMux I__13068 (
            .O(N__52860),
            .I(N__52854));
    LocalMux I__13067 (
            .O(N__52857),
            .I(N__52851));
    InMux I__13066 (
            .O(N__52854),
            .I(N__52848));
    Sp12to4 I__13065 (
            .O(N__52851),
            .I(N__52845));
    LocalMux I__13064 (
            .O(N__52848),
            .I(N__52842));
    Span12Mux_v I__13063 (
            .O(N__52845),
            .I(N__52839));
    Span4Mux_h I__13062 (
            .O(N__52842),
            .I(N__52836));
    Odrv12 I__13061 (
            .O(N__52839),
            .I(PIO_dport0_T4_1));
    Odrv4 I__13060 (
            .O(N__52836),
            .I(PIO_dport0_T4_1));
    InMux I__13059 (
            .O(N__52831),
            .I(N__52828));
    LocalMux I__13058 (
            .O(N__52828),
            .I(N__52824));
    InMux I__13057 (
            .O(N__52827),
            .I(N__52821));
    Span4Mux_v I__13056 (
            .O(N__52824),
            .I(N__52818));
    LocalMux I__13055 (
            .O(N__52821),
            .I(N__52815));
    Sp12to4 I__13054 (
            .O(N__52818),
            .I(N__52812));
    Span4Mux_v I__13053 (
            .O(N__52815),
            .I(N__52809));
    Odrv12 I__13052 (
            .O(N__52812),
            .I(PIO_dport1_T4_1));
    Odrv4 I__13051 (
            .O(N__52809),
            .I(PIO_dport1_T4_1));
    CascadeMux I__13050 (
            .O(N__52804),
            .I(N__52801));
    InMux I__13049 (
            .O(N__52801),
            .I(N__52798));
    LocalMux I__13048 (
            .O(N__52798),
            .I(N__52795));
    Span4Mux_v I__13047 (
            .O(N__52795),
            .I(N__52792));
    Odrv4 I__13046 (
            .O(N__52792),
            .I(\u0.dat_o_0_a2_i_0_17 ));
    InMux I__13045 (
            .O(N__52789),
            .I(N__52784));
    CascadeMux I__13044 (
            .O(N__52788),
            .I(N__52775));
    CascadeMux I__13043 (
            .O(N__52787),
            .I(N__52764));
    LocalMux I__13042 (
            .O(N__52784),
            .I(N__52758));
    InMux I__13041 (
            .O(N__52783),
            .I(N__52751));
    InMux I__13040 (
            .O(N__52782),
            .I(N__52751));
    InMux I__13039 (
            .O(N__52781),
            .I(N__52751));
    InMux I__13038 (
            .O(N__52780),
            .I(N__52742));
    InMux I__13037 (
            .O(N__52779),
            .I(N__52742));
    InMux I__13036 (
            .O(N__52778),
            .I(N__52742));
    InMux I__13035 (
            .O(N__52775),
            .I(N__52742));
    CascadeMux I__13034 (
            .O(N__52774),
            .I(N__52739));
    CascadeMux I__13033 (
            .O(N__52773),
            .I(N__52736));
    CascadeMux I__13032 (
            .O(N__52772),
            .I(N__52733));
    CascadeMux I__13031 (
            .O(N__52771),
            .I(N__52729));
    CascadeMux I__13030 (
            .O(N__52770),
            .I(N__52726));
    CascadeMux I__13029 (
            .O(N__52769),
            .I(N__52723));
    CascadeMux I__13028 (
            .O(N__52768),
            .I(N__52720));
    CascadeMux I__13027 (
            .O(N__52767),
            .I(N__52717));
    InMux I__13026 (
            .O(N__52764),
            .I(N__52714));
    InMux I__13025 (
            .O(N__52763),
            .I(N__52711));
    CascadeMux I__13024 (
            .O(N__52762),
            .I(N__52704));
    CascadeMux I__13023 (
            .O(N__52761),
            .I(N__52701));
    Span4Mux_v I__13022 (
            .O(N__52758),
            .I(N__52685));
    LocalMux I__13021 (
            .O(N__52751),
            .I(N__52685));
    LocalMux I__13020 (
            .O(N__52742),
            .I(N__52685));
    InMux I__13019 (
            .O(N__52739),
            .I(N__52680));
    InMux I__13018 (
            .O(N__52736),
            .I(N__52680));
    InMux I__13017 (
            .O(N__52733),
            .I(N__52677));
    InMux I__13016 (
            .O(N__52732),
            .I(N__52670));
    InMux I__13015 (
            .O(N__52729),
            .I(N__52670));
    InMux I__13014 (
            .O(N__52726),
            .I(N__52670));
    InMux I__13013 (
            .O(N__52723),
            .I(N__52667));
    InMux I__13012 (
            .O(N__52720),
            .I(N__52664));
    InMux I__13011 (
            .O(N__52717),
            .I(N__52661));
    LocalMux I__13010 (
            .O(N__52714),
            .I(N__52656));
    LocalMux I__13009 (
            .O(N__52711),
            .I(N__52656));
    InMux I__13008 (
            .O(N__52710),
            .I(N__52653));
    CascadeMux I__13007 (
            .O(N__52709),
            .I(N__52648));
    CascadeMux I__13006 (
            .O(N__52708),
            .I(N__52632));
    CascadeMux I__13005 (
            .O(N__52707),
            .I(N__52624));
    InMux I__13004 (
            .O(N__52704),
            .I(N__52618));
    InMux I__13003 (
            .O(N__52701),
            .I(N__52618));
    CascadeMux I__13002 (
            .O(N__52700),
            .I(N__52615));
    CascadeMux I__13001 (
            .O(N__52699),
            .I(N__52612));
    CascadeMux I__13000 (
            .O(N__52698),
            .I(N__52603));
    CascadeMux I__12999 (
            .O(N__52697),
            .I(N__52598));
    CascadeMux I__12998 (
            .O(N__52696),
            .I(N__52595));
    CascadeMux I__12997 (
            .O(N__52695),
            .I(N__52592));
    CascadeMux I__12996 (
            .O(N__52694),
            .I(N__52589));
    CascadeMux I__12995 (
            .O(N__52693),
            .I(N__52585));
    CascadeMux I__12994 (
            .O(N__52692),
            .I(N__52582));
    Span4Mux_v I__12993 (
            .O(N__52685),
            .I(N__52560));
    LocalMux I__12992 (
            .O(N__52680),
            .I(N__52560));
    LocalMux I__12991 (
            .O(N__52677),
            .I(N__52560));
    LocalMux I__12990 (
            .O(N__52670),
            .I(N__52560));
    LocalMux I__12989 (
            .O(N__52667),
            .I(N__52560));
    LocalMux I__12988 (
            .O(N__52664),
            .I(N__52560));
    LocalMux I__12987 (
            .O(N__52661),
            .I(N__52553));
    Span4Mux_s3_v I__12986 (
            .O(N__52656),
            .I(N__52553));
    LocalMux I__12985 (
            .O(N__52653),
            .I(N__52553));
    InMux I__12984 (
            .O(N__52652),
            .I(N__52550));
    InMux I__12983 (
            .O(N__52651),
            .I(N__52547));
    InMux I__12982 (
            .O(N__52648),
            .I(N__52544));
    InMux I__12981 (
            .O(N__52647),
            .I(N__52537));
    InMux I__12980 (
            .O(N__52646),
            .I(N__52537));
    InMux I__12979 (
            .O(N__52645),
            .I(N__52537));
    InMux I__12978 (
            .O(N__52644),
            .I(N__52526));
    InMux I__12977 (
            .O(N__52643),
            .I(N__52526));
    InMux I__12976 (
            .O(N__52642),
            .I(N__52526));
    InMux I__12975 (
            .O(N__52641),
            .I(N__52526));
    InMux I__12974 (
            .O(N__52640),
            .I(N__52526));
    InMux I__12973 (
            .O(N__52639),
            .I(N__52519));
    InMux I__12972 (
            .O(N__52638),
            .I(N__52519));
    InMux I__12971 (
            .O(N__52637),
            .I(N__52519));
    CascadeMux I__12970 (
            .O(N__52636),
            .I(N__52498));
    CascadeMux I__12969 (
            .O(N__52635),
            .I(N__52495));
    InMux I__12968 (
            .O(N__52632),
            .I(N__52490));
    InMux I__12967 (
            .O(N__52631),
            .I(N__52485));
    InMux I__12966 (
            .O(N__52630),
            .I(N__52485));
    CascadeMux I__12965 (
            .O(N__52629),
            .I(N__52482));
    CascadeMux I__12964 (
            .O(N__52628),
            .I(N__52479));
    InMux I__12963 (
            .O(N__52627),
            .I(N__52476));
    InMux I__12962 (
            .O(N__52624),
            .I(N__52473));
    CascadeMux I__12961 (
            .O(N__52623),
            .I(N__52464));
    LocalMux I__12960 (
            .O(N__52618),
            .I(N__52456));
    InMux I__12959 (
            .O(N__52615),
            .I(N__52451));
    InMux I__12958 (
            .O(N__52612),
            .I(N__52451));
    CascadeMux I__12957 (
            .O(N__52611),
            .I(N__52446));
    CascadeMux I__12956 (
            .O(N__52610),
            .I(N__52441));
    CascadeMux I__12955 (
            .O(N__52609),
            .I(N__52437));
    CascadeMux I__12954 (
            .O(N__52608),
            .I(N__52433));
    CascadeMux I__12953 (
            .O(N__52607),
            .I(N__52430));
    CascadeMux I__12952 (
            .O(N__52606),
            .I(N__52427));
    InMux I__12951 (
            .O(N__52603),
            .I(N__52417));
    InMux I__12950 (
            .O(N__52602),
            .I(N__52417));
    InMux I__12949 (
            .O(N__52601),
            .I(N__52414));
    InMux I__12948 (
            .O(N__52598),
            .I(N__52405));
    InMux I__12947 (
            .O(N__52595),
            .I(N__52405));
    InMux I__12946 (
            .O(N__52592),
            .I(N__52405));
    InMux I__12945 (
            .O(N__52589),
            .I(N__52405));
    InMux I__12944 (
            .O(N__52588),
            .I(N__52396));
    InMux I__12943 (
            .O(N__52585),
            .I(N__52396));
    InMux I__12942 (
            .O(N__52582),
            .I(N__52396));
    InMux I__12941 (
            .O(N__52581),
            .I(N__52396));
    CascadeMux I__12940 (
            .O(N__52580),
            .I(N__52393));
    CascadeMux I__12939 (
            .O(N__52579),
            .I(N__52390));
    CascadeMux I__12938 (
            .O(N__52578),
            .I(N__52387));
    CascadeMux I__12937 (
            .O(N__52577),
            .I(N__52384));
    CascadeMux I__12936 (
            .O(N__52576),
            .I(N__52381));
    CascadeMux I__12935 (
            .O(N__52575),
            .I(N__52378));
    CascadeMux I__12934 (
            .O(N__52574),
            .I(N__52375));
    CascadeMux I__12933 (
            .O(N__52573),
            .I(N__52372));
    Span4Mux_v I__12932 (
            .O(N__52560),
            .I(N__52369));
    Span4Mux_v I__12931 (
            .O(N__52553),
            .I(N__52354));
    LocalMux I__12930 (
            .O(N__52550),
            .I(N__52354));
    LocalMux I__12929 (
            .O(N__52547),
            .I(N__52354));
    LocalMux I__12928 (
            .O(N__52544),
            .I(N__52354));
    LocalMux I__12927 (
            .O(N__52537),
            .I(N__52354));
    LocalMux I__12926 (
            .O(N__52526),
            .I(N__52354));
    LocalMux I__12925 (
            .O(N__52519),
            .I(N__52354));
    InMux I__12924 (
            .O(N__52518),
            .I(N__52337));
    InMux I__12923 (
            .O(N__52517),
            .I(N__52337));
    InMux I__12922 (
            .O(N__52516),
            .I(N__52337));
    InMux I__12921 (
            .O(N__52515),
            .I(N__52337));
    InMux I__12920 (
            .O(N__52514),
            .I(N__52337));
    InMux I__12919 (
            .O(N__52513),
            .I(N__52337));
    InMux I__12918 (
            .O(N__52512),
            .I(N__52337));
    InMux I__12917 (
            .O(N__52511),
            .I(N__52337));
    InMux I__12916 (
            .O(N__52510),
            .I(N__52322));
    InMux I__12915 (
            .O(N__52509),
            .I(N__52322));
    InMux I__12914 (
            .O(N__52508),
            .I(N__52322));
    InMux I__12913 (
            .O(N__52507),
            .I(N__52322));
    InMux I__12912 (
            .O(N__52506),
            .I(N__52322));
    InMux I__12911 (
            .O(N__52505),
            .I(N__52322));
    InMux I__12910 (
            .O(N__52504),
            .I(N__52322));
    InMux I__12909 (
            .O(N__52503),
            .I(N__52319));
    InMux I__12908 (
            .O(N__52502),
            .I(N__52312));
    InMux I__12907 (
            .O(N__52501),
            .I(N__52312));
    InMux I__12906 (
            .O(N__52498),
            .I(N__52312));
    InMux I__12905 (
            .O(N__52495),
            .I(N__52309));
    CascadeMux I__12904 (
            .O(N__52494),
            .I(N__52302));
    CascadeMux I__12903 (
            .O(N__52493),
            .I(N__52298));
    LocalMux I__12902 (
            .O(N__52490),
            .I(N__52292));
    LocalMux I__12901 (
            .O(N__52485),
            .I(N__52292));
    InMux I__12900 (
            .O(N__52482),
            .I(N__52287));
    InMux I__12899 (
            .O(N__52479),
            .I(N__52287));
    LocalMux I__12898 (
            .O(N__52476),
            .I(N__52282));
    LocalMux I__12897 (
            .O(N__52473),
            .I(N__52282));
    InMux I__12896 (
            .O(N__52472),
            .I(N__52275));
    InMux I__12895 (
            .O(N__52471),
            .I(N__52275));
    InMux I__12894 (
            .O(N__52470),
            .I(N__52275));
    InMux I__12893 (
            .O(N__52469),
            .I(N__52264));
    InMux I__12892 (
            .O(N__52468),
            .I(N__52264));
    InMux I__12891 (
            .O(N__52467),
            .I(N__52264));
    InMux I__12890 (
            .O(N__52464),
            .I(N__52264));
    InMux I__12889 (
            .O(N__52463),
            .I(N__52264));
    CascadeMux I__12888 (
            .O(N__52462),
            .I(N__52259));
    CascadeMux I__12887 (
            .O(N__52461),
            .I(N__52256));
    CascadeMux I__12886 (
            .O(N__52460),
            .I(N__52249));
    CascadeMux I__12885 (
            .O(N__52459),
            .I(N__52246));
    Span4Mux_s3_v I__12884 (
            .O(N__52456),
            .I(N__52236));
    LocalMux I__12883 (
            .O(N__52451),
            .I(N__52236));
    InMux I__12882 (
            .O(N__52450),
            .I(N__52233));
    InMux I__12881 (
            .O(N__52449),
            .I(N__52230));
    InMux I__12880 (
            .O(N__52446),
            .I(N__52227));
    InMux I__12879 (
            .O(N__52445),
            .I(N__52218));
    InMux I__12878 (
            .O(N__52444),
            .I(N__52218));
    InMux I__12877 (
            .O(N__52441),
            .I(N__52218));
    InMux I__12876 (
            .O(N__52440),
            .I(N__52218));
    InMux I__12875 (
            .O(N__52437),
            .I(N__52213));
    InMux I__12874 (
            .O(N__52436),
            .I(N__52213));
    InMux I__12873 (
            .O(N__52433),
            .I(N__52206));
    InMux I__12872 (
            .O(N__52430),
            .I(N__52206));
    InMux I__12871 (
            .O(N__52427),
            .I(N__52206));
    CascadeMux I__12870 (
            .O(N__52426),
            .I(N__52201));
    InMux I__12869 (
            .O(N__52425),
            .I(N__52187));
    InMux I__12868 (
            .O(N__52424),
            .I(N__52187));
    InMux I__12867 (
            .O(N__52423),
            .I(N__52187));
    CascadeMux I__12866 (
            .O(N__52422),
            .I(N__52183));
    LocalMux I__12865 (
            .O(N__52417),
            .I(N__52169));
    LocalMux I__12864 (
            .O(N__52414),
            .I(N__52169));
    LocalMux I__12863 (
            .O(N__52405),
            .I(N__52169));
    LocalMux I__12862 (
            .O(N__52396),
            .I(N__52169));
    InMux I__12861 (
            .O(N__52393),
            .I(N__52160));
    InMux I__12860 (
            .O(N__52390),
            .I(N__52160));
    InMux I__12859 (
            .O(N__52387),
            .I(N__52160));
    InMux I__12858 (
            .O(N__52384),
            .I(N__52160));
    InMux I__12857 (
            .O(N__52381),
            .I(N__52151));
    InMux I__12856 (
            .O(N__52378),
            .I(N__52151));
    InMux I__12855 (
            .O(N__52375),
            .I(N__52151));
    InMux I__12854 (
            .O(N__52372),
            .I(N__52151));
    Span4Mux_h I__12853 (
            .O(N__52369),
            .I(N__52136));
    Span4Mux_v I__12852 (
            .O(N__52354),
            .I(N__52136));
    LocalMux I__12851 (
            .O(N__52337),
            .I(N__52136));
    LocalMux I__12850 (
            .O(N__52322),
            .I(N__52136));
    LocalMux I__12849 (
            .O(N__52319),
            .I(N__52136));
    LocalMux I__12848 (
            .O(N__52312),
            .I(N__52136));
    LocalMux I__12847 (
            .O(N__52309),
            .I(N__52136));
    CascadeMux I__12846 (
            .O(N__52308),
            .I(N__52133));
    CascadeMux I__12845 (
            .O(N__52307),
            .I(N__52130));
    CascadeMux I__12844 (
            .O(N__52306),
            .I(N__52127));
    CascadeMux I__12843 (
            .O(N__52305),
            .I(N__52124));
    InMux I__12842 (
            .O(N__52302),
            .I(N__52119));
    InMux I__12841 (
            .O(N__52301),
            .I(N__52119));
    InMux I__12840 (
            .O(N__52298),
            .I(N__52116));
    CascadeMux I__12839 (
            .O(N__52297),
            .I(N__52107));
    Span4Mux_v I__12838 (
            .O(N__52292),
            .I(N__52100));
    LocalMux I__12837 (
            .O(N__52287),
            .I(N__52100));
    Span4Mux_v I__12836 (
            .O(N__52282),
            .I(N__52093));
    LocalMux I__12835 (
            .O(N__52275),
            .I(N__52093));
    LocalMux I__12834 (
            .O(N__52264),
            .I(N__52093));
    InMux I__12833 (
            .O(N__52263),
            .I(N__52088));
    InMux I__12832 (
            .O(N__52262),
            .I(N__52088));
    InMux I__12831 (
            .O(N__52259),
            .I(N__52081));
    InMux I__12830 (
            .O(N__52256),
            .I(N__52081));
    InMux I__12829 (
            .O(N__52255),
            .I(N__52081));
    InMux I__12828 (
            .O(N__52254),
            .I(N__52078));
    InMux I__12827 (
            .O(N__52253),
            .I(N__52069));
    InMux I__12826 (
            .O(N__52252),
            .I(N__52069));
    InMux I__12825 (
            .O(N__52249),
            .I(N__52069));
    InMux I__12824 (
            .O(N__52246),
            .I(N__52069));
    InMux I__12823 (
            .O(N__52245),
            .I(N__52066));
    InMux I__12822 (
            .O(N__52244),
            .I(N__52063));
    CascadeMux I__12821 (
            .O(N__52243),
            .I(N__52060));
    CascadeMux I__12820 (
            .O(N__52242),
            .I(N__52055));
    CascadeMux I__12819 (
            .O(N__52241),
            .I(N__52052));
    Span4Mux_v I__12818 (
            .O(N__52236),
            .I(N__52046));
    LocalMux I__12817 (
            .O(N__52233),
            .I(N__52046));
    LocalMux I__12816 (
            .O(N__52230),
            .I(N__52039));
    LocalMux I__12815 (
            .O(N__52227),
            .I(N__52039));
    LocalMux I__12814 (
            .O(N__52218),
            .I(N__52039));
    LocalMux I__12813 (
            .O(N__52213),
            .I(N__52034));
    LocalMux I__12812 (
            .O(N__52206),
            .I(N__52034));
    InMux I__12811 (
            .O(N__52205),
            .I(N__52031));
    InMux I__12810 (
            .O(N__52204),
            .I(N__52026));
    InMux I__12809 (
            .O(N__52201),
            .I(N__52026));
    InMux I__12808 (
            .O(N__52200),
            .I(N__52021));
    InMux I__12807 (
            .O(N__52199),
            .I(N__52021));
    CascadeMux I__12806 (
            .O(N__52198),
            .I(N__52018));
    CascadeMux I__12805 (
            .O(N__52197),
            .I(N__52015));
    CascadeMux I__12804 (
            .O(N__52196),
            .I(N__52012));
    CascadeMux I__12803 (
            .O(N__52195),
            .I(N__52008));
    CascadeMux I__12802 (
            .O(N__52194),
            .I(N__52004));
    LocalMux I__12801 (
            .O(N__52187),
            .I(N__52000));
    InMux I__12800 (
            .O(N__52186),
            .I(N__51991));
    InMux I__12799 (
            .O(N__52183),
            .I(N__51991));
    InMux I__12798 (
            .O(N__52182),
            .I(N__51991));
    InMux I__12797 (
            .O(N__52181),
            .I(N__51991));
    CascadeMux I__12796 (
            .O(N__52180),
            .I(N__51988));
    CascadeMux I__12795 (
            .O(N__52179),
            .I(N__51983));
    CascadeMux I__12794 (
            .O(N__52178),
            .I(N__51979));
    Span4Mux_v I__12793 (
            .O(N__52169),
            .I(N__51974));
    LocalMux I__12792 (
            .O(N__52160),
            .I(N__51974));
    LocalMux I__12791 (
            .O(N__52151),
            .I(N__51969));
    Span4Mux_v I__12790 (
            .O(N__52136),
            .I(N__51969));
    InMux I__12789 (
            .O(N__52133),
            .I(N__51962));
    InMux I__12788 (
            .O(N__52130),
            .I(N__51962));
    InMux I__12787 (
            .O(N__52127),
            .I(N__51962));
    InMux I__12786 (
            .O(N__52124),
            .I(N__51959));
    LocalMux I__12785 (
            .O(N__52119),
            .I(N__51954));
    LocalMux I__12784 (
            .O(N__52116),
            .I(N__51954));
    InMux I__12783 (
            .O(N__52115),
            .I(N__51951));
    InMux I__12782 (
            .O(N__52114),
            .I(N__51943));
    CascadeMux I__12781 (
            .O(N__52113),
            .I(N__51935));
    CascadeMux I__12780 (
            .O(N__52112),
            .I(N__51929));
    CascadeMux I__12779 (
            .O(N__52111),
            .I(N__51925));
    CascadeMux I__12778 (
            .O(N__52110),
            .I(N__51919));
    InMux I__12777 (
            .O(N__52107),
            .I(N__51914));
    InMux I__12776 (
            .O(N__52106),
            .I(N__51911));
    InMux I__12775 (
            .O(N__52105),
            .I(N__51908));
    Span4Mux_v I__12774 (
            .O(N__52100),
            .I(N__51900));
    Span4Mux_v I__12773 (
            .O(N__52093),
            .I(N__51900));
    LocalMux I__12772 (
            .O(N__52088),
            .I(N__51900));
    LocalMux I__12771 (
            .O(N__52081),
            .I(N__51893));
    LocalMux I__12770 (
            .O(N__52078),
            .I(N__51893));
    LocalMux I__12769 (
            .O(N__52069),
            .I(N__51893));
    LocalMux I__12768 (
            .O(N__52066),
            .I(N__51890));
    LocalMux I__12767 (
            .O(N__52063),
            .I(N__51887));
    InMux I__12766 (
            .O(N__52060),
            .I(N__51884));
    InMux I__12765 (
            .O(N__52059),
            .I(N__51881));
    InMux I__12764 (
            .O(N__52058),
            .I(N__51864));
    InMux I__12763 (
            .O(N__52055),
            .I(N__51859));
    InMux I__12762 (
            .O(N__52052),
            .I(N__51856));
    CascadeMux I__12761 (
            .O(N__52051),
            .I(N__51845));
    Span4Mux_v I__12760 (
            .O(N__52046),
            .I(N__51826));
    Span4Mux_v I__12759 (
            .O(N__52039),
            .I(N__51826));
    Span4Mux_h I__12758 (
            .O(N__52034),
            .I(N__51826));
    LocalMux I__12757 (
            .O(N__52031),
            .I(N__51826));
    LocalMux I__12756 (
            .O(N__52026),
            .I(N__51826));
    LocalMux I__12755 (
            .O(N__52021),
            .I(N__51826));
    InMux I__12754 (
            .O(N__52018),
            .I(N__51819));
    InMux I__12753 (
            .O(N__52015),
            .I(N__51819));
    InMux I__12752 (
            .O(N__52012),
            .I(N__51819));
    InMux I__12751 (
            .O(N__52011),
            .I(N__51810));
    InMux I__12750 (
            .O(N__52008),
            .I(N__51810));
    InMux I__12749 (
            .O(N__52007),
            .I(N__51810));
    InMux I__12748 (
            .O(N__52004),
            .I(N__51810));
    InMux I__12747 (
            .O(N__52003),
            .I(N__51803));
    Span4Mux_v I__12746 (
            .O(N__52000),
            .I(N__51797));
    LocalMux I__12745 (
            .O(N__51991),
            .I(N__51797));
    InMux I__12744 (
            .O(N__51988),
            .I(N__51784));
    InMux I__12743 (
            .O(N__51987),
            .I(N__51784));
    InMux I__12742 (
            .O(N__51986),
            .I(N__51784));
    InMux I__12741 (
            .O(N__51983),
            .I(N__51784));
    InMux I__12740 (
            .O(N__51982),
            .I(N__51784));
    InMux I__12739 (
            .O(N__51979),
            .I(N__51784));
    Span4Mux_h I__12738 (
            .O(N__51974),
            .I(N__51773));
    Span4Mux_h I__12737 (
            .O(N__51969),
            .I(N__51773));
    LocalMux I__12736 (
            .O(N__51962),
            .I(N__51773));
    LocalMux I__12735 (
            .O(N__51959),
            .I(N__51773));
    Span4Mux_v I__12734 (
            .O(N__51954),
            .I(N__51768));
    LocalMux I__12733 (
            .O(N__51951),
            .I(N__51768));
    InMux I__12732 (
            .O(N__51950),
            .I(N__51761));
    InMux I__12731 (
            .O(N__51949),
            .I(N__51761));
    InMux I__12730 (
            .O(N__51948),
            .I(N__51761));
    InMux I__12729 (
            .O(N__51947),
            .I(N__51758));
    InMux I__12728 (
            .O(N__51946),
            .I(N__51755));
    LocalMux I__12727 (
            .O(N__51943),
            .I(N__51751));
    InMux I__12726 (
            .O(N__51942),
            .I(N__51748));
    InMux I__12725 (
            .O(N__51941),
            .I(N__51745));
    InMux I__12724 (
            .O(N__51940),
            .I(N__51742));
    InMux I__12723 (
            .O(N__51939),
            .I(N__51725));
    InMux I__12722 (
            .O(N__51938),
            .I(N__51725));
    InMux I__12721 (
            .O(N__51935),
            .I(N__51725));
    InMux I__12720 (
            .O(N__51934),
            .I(N__51725));
    InMux I__12719 (
            .O(N__51933),
            .I(N__51725));
    InMux I__12718 (
            .O(N__51932),
            .I(N__51725));
    InMux I__12717 (
            .O(N__51929),
            .I(N__51725));
    InMux I__12716 (
            .O(N__51928),
            .I(N__51725));
    InMux I__12715 (
            .O(N__51925),
            .I(N__51697));
    InMux I__12714 (
            .O(N__51924),
            .I(N__51697));
    InMux I__12713 (
            .O(N__51923),
            .I(N__51697));
    InMux I__12712 (
            .O(N__51922),
            .I(N__51697));
    InMux I__12711 (
            .O(N__51919),
            .I(N__51697));
    InMux I__12710 (
            .O(N__51918),
            .I(N__51697));
    InMux I__12709 (
            .O(N__51917),
            .I(N__51697));
    LocalMux I__12708 (
            .O(N__51914),
            .I(N__51689));
    LocalMux I__12707 (
            .O(N__51911),
            .I(N__51689));
    LocalMux I__12706 (
            .O(N__51908),
            .I(N__51689));
    InMux I__12705 (
            .O(N__51907),
            .I(N__51686));
    Span4Mux_v I__12704 (
            .O(N__51900),
            .I(N__51678));
    Span4Mux_v I__12703 (
            .O(N__51893),
            .I(N__51678));
    Span4Mux_v I__12702 (
            .O(N__51890),
            .I(N__51675));
    Span4Mux_v I__12701 (
            .O(N__51887),
            .I(N__51670));
    LocalMux I__12700 (
            .O(N__51884),
            .I(N__51670));
    LocalMux I__12699 (
            .O(N__51881),
            .I(N__51667));
    InMux I__12698 (
            .O(N__51880),
            .I(N__51654));
    InMux I__12697 (
            .O(N__51879),
            .I(N__51654));
    InMux I__12696 (
            .O(N__51878),
            .I(N__51654));
    InMux I__12695 (
            .O(N__51877),
            .I(N__51654));
    InMux I__12694 (
            .O(N__51876),
            .I(N__51654));
    InMux I__12693 (
            .O(N__51875),
            .I(N__51654));
    InMux I__12692 (
            .O(N__51874),
            .I(N__51639));
    InMux I__12691 (
            .O(N__51873),
            .I(N__51639));
    InMux I__12690 (
            .O(N__51872),
            .I(N__51639));
    InMux I__12689 (
            .O(N__51871),
            .I(N__51639));
    InMux I__12688 (
            .O(N__51870),
            .I(N__51639));
    InMux I__12687 (
            .O(N__51869),
            .I(N__51639));
    InMux I__12686 (
            .O(N__51868),
            .I(N__51639));
    CascadeMux I__12685 (
            .O(N__51867),
            .I(N__51628));
    LocalMux I__12684 (
            .O(N__51864),
            .I(N__51623));
    InMux I__12683 (
            .O(N__51863),
            .I(N__51618));
    InMux I__12682 (
            .O(N__51862),
            .I(N__51615));
    LocalMux I__12681 (
            .O(N__51859),
            .I(N__51607));
    LocalMux I__12680 (
            .O(N__51856),
            .I(N__51604));
    CascadeMux I__12679 (
            .O(N__51855),
            .I(N__51601));
    CascadeMux I__12678 (
            .O(N__51854),
            .I(N__51598));
    CascadeMux I__12677 (
            .O(N__51853),
            .I(N__51595));
    CascadeMux I__12676 (
            .O(N__51852),
            .I(N__51591));
    CascadeMux I__12675 (
            .O(N__51851),
            .I(N__51588));
    CascadeMux I__12674 (
            .O(N__51850),
            .I(N__51585));
    InMux I__12673 (
            .O(N__51849),
            .I(N__51569));
    InMux I__12672 (
            .O(N__51848),
            .I(N__51569));
    InMux I__12671 (
            .O(N__51845),
            .I(N__51569));
    InMux I__12670 (
            .O(N__51844),
            .I(N__51569));
    InMux I__12669 (
            .O(N__51843),
            .I(N__51569));
    InMux I__12668 (
            .O(N__51842),
            .I(N__51569));
    InMux I__12667 (
            .O(N__51841),
            .I(N__51569));
    CascadeMux I__12666 (
            .O(N__51840),
            .I(N__51566));
    CascadeMux I__12665 (
            .O(N__51839),
            .I(N__51561));
    Span4Mux_v I__12664 (
            .O(N__51826),
            .I(N__51553));
    LocalMux I__12663 (
            .O(N__51819),
            .I(N__51553));
    LocalMux I__12662 (
            .O(N__51810),
            .I(N__51553));
    InMux I__12661 (
            .O(N__51809),
            .I(N__51532));
    InMux I__12660 (
            .O(N__51808),
            .I(N__51532));
    InMux I__12659 (
            .O(N__51807),
            .I(N__51532));
    InMux I__12658 (
            .O(N__51806),
            .I(N__51532));
    LocalMux I__12657 (
            .O(N__51803),
            .I(N__51529));
    InMux I__12656 (
            .O(N__51802),
            .I(N__51526));
    Span4Mux_v I__12655 (
            .O(N__51797),
            .I(N__51521));
    LocalMux I__12654 (
            .O(N__51784),
            .I(N__51521));
    InMux I__12653 (
            .O(N__51783),
            .I(N__51516));
    InMux I__12652 (
            .O(N__51782),
            .I(N__51516));
    Span4Mux_v I__12651 (
            .O(N__51773),
            .I(N__51511));
    Span4Mux_v I__12650 (
            .O(N__51768),
            .I(N__51511));
    LocalMux I__12649 (
            .O(N__51761),
            .I(N__51504));
    LocalMux I__12648 (
            .O(N__51758),
            .I(N__51504));
    LocalMux I__12647 (
            .O(N__51755),
            .I(N__51504));
    InMux I__12646 (
            .O(N__51754),
            .I(N__51501));
    Span4Mux_v I__12645 (
            .O(N__51751),
            .I(N__51489));
    LocalMux I__12644 (
            .O(N__51748),
            .I(N__51489));
    LocalMux I__12643 (
            .O(N__51745),
            .I(N__51489));
    LocalMux I__12642 (
            .O(N__51742),
            .I(N__51489));
    LocalMux I__12641 (
            .O(N__51725),
            .I(N__51489));
    InMux I__12640 (
            .O(N__51724),
            .I(N__51474));
    InMux I__12639 (
            .O(N__51723),
            .I(N__51474));
    InMux I__12638 (
            .O(N__51722),
            .I(N__51474));
    InMux I__12637 (
            .O(N__51721),
            .I(N__51474));
    InMux I__12636 (
            .O(N__51720),
            .I(N__51474));
    InMux I__12635 (
            .O(N__51719),
            .I(N__51474));
    InMux I__12634 (
            .O(N__51718),
            .I(N__51474));
    InMux I__12633 (
            .O(N__51717),
            .I(N__51471));
    InMux I__12632 (
            .O(N__51716),
            .I(N__51460));
    InMux I__12631 (
            .O(N__51715),
            .I(N__51460));
    InMux I__12630 (
            .O(N__51714),
            .I(N__51460));
    InMux I__12629 (
            .O(N__51713),
            .I(N__51460));
    InMux I__12628 (
            .O(N__51712),
            .I(N__51460));
    LocalMux I__12627 (
            .O(N__51697),
            .I(N__51454));
    InMux I__12626 (
            .O(N__51696),
            .I(N__51451));
    Span4Mux_v I__12625 (
            .O(N__51689),
            .I(N__51446));
    LocalMux I__12624 (
            .O(N__51686),
            .I(N__51446));
    InMux I__12623 (
            .O(N__51685),
            .I(N__51443));
    InMux I__12622 (
            .O(N__51684),
            .I(N__51440));
    InMux I__12621 (
            .O(N__51683),
            .I(N__51437));
    Span4Mux_h I__12620 (
            .O(N__51678),
            .I(N__51433));
    Span4Mux_h I__12619 (
            .O(N__51675),
            .I(N__51428));
    Span4Mux_v I__12618 (
            .O(N__51670),
            .I(N__51428));
    Span4Mux_v I__12617 (
            .O(N__51667),
            .I(N__51421));
    LocalMux I__12616 (
            .O(N__51654),
            .I(N__51421));
    LocalMux I__12615 (
            .O(N__51639),
            .I(N__51421));
    InMux I__12614 (
            .O(N__51638),
            .I(N__51408));
    InMux I__12613 (
            .O(N__51637),
            .I(N__51408));
    InMux I__12612 (
            .O(N__51636),
            .I(N__51408));
    InMux I__12611 (
            .O(N__51635),
            .I(N__51408));
    InMux I__12610 (
            .O(N__51634),
            .I(N__51408));
    InMux I__12609 (
            .O(N__51633),
            .I(N__51408));
    InMux I__12608 (
            .O(N__51632),
            .I(N__51397));
    InMux I__12607 (
            .O(N__51631),
            .I(N__51397));
    InMux I__12606 (
            .O(N__51628),
            .I(N__51397));
    InMux I__12605 (
            .O(N__51627),
            .I(N__51397));
    InMux I__12604 (
            .O(N__51626),
            .I(N__51397));
    Span4Mux_v I__12603 (
            .O(N__51623),
            .I(N__51394));
    InMux I__12602 (
            .O(N__51622),
            .I(N__51391));
    InMux I__12601 (
            .O(N__51621),
            .I(N__51388));
    LocalMux I__12600 (
            .O(N__51618),
            .I(N__51383));
    LocalMux I__12599 (
            .O(N__51615),
            .I(N__51383));
    InMux I__12598 (
            .O(N__51614),
            .I(N__51380));
    InMux I__12597 (
            .O(N__51613),
            .I(N__51377));
    InMux I__12596 (
            .O(N__51612),
            .I(N__51374));
    InMux I__12595 (
            .O(N__51611),
            .I(N__51370));
    InMux I__12594 (
            .O(N__51610),
            .I(N__51367));
    Span4Mux_v I__12593 (
            .O(N__51607),
            .I(N__51358));
    Span4Mux_v I__12592 (
            .O(N__51604),
            .I(N__51358));
    InMux I__12591 (
            .O(N__51601),
            .I(N__51349));
    InMux I__12590 (
            .O(N__51598),
            .I(N__51349));
    InMux I__12589 (
            .O(N__51595),
            .I(N__51349));
    InMux I__12588 (
            .O(N__51594),
            .I(N__51349));
    InMux I__12587 (
            .O(N__51591),
            .I(N__51340));
    InMux I__12586 (
            .O(N__51588),
            .I(N__51340));
    InMux I__12585 (
            .O(N__51585),
            .I(N__51340));
    InMux I__12584 (
            .O(N__51584),
            .I(N__51340));
    LocalMux I__12583 (
            .O(N__51569),
            .I(N__51337));
    InMux I__12582 (
            .O(N__51566),
            .I(N__51334));
    InMux I__12581 (
            .O(N__51565),
            .I(N__51325));
    InMux I__12580 (
            .O(N__51564),
            .I(N__51325));
    InMux I__12579 (
            .O(N__51561),
            .I(N__51325));
    InMux I__12578 (
            .O(N__51560),
            .I(N__51325));
    Span4Mux_v I__12577 (
            .O(N__51553),
            .I(N__51322));
    InMux I__12576 (
            .O(N__51552),
            .I(N__51315));
    InMux I__12575 (
            .O(N__51551),
            .I(N__51315));
    InMux I__12574 (
            .O(N__51550),
            .I(N__51315));
    InMux I__12573 (
            .O(N__51549),
            .I(N__51312));
    InMux I__12572 (
            .O(N__51548),
            .I(N__51283));
    InMux I__12571 (
            .O(N__51547),
            .I(N__51283));
    InMux I__12570 (
            .O(N__51546),
            .I(N__51283));
    InMux I__12569 (
            .O(N__51545),
            .I(N__51283));
    InMux I__12568 (
            .O(N__51544),
            .I(N__51283));
    InMux I__12567 (
            .O(N__51543),
            .I(N__51283));
    InMux I__12566 (
            .O(N__51542),
            .I(N__51283));
    InMux I__12565 (
            .O(N__51541),
            .I(N__51280));
    LocalMux I__12564 (
            .O(N__51532),
            .I(N__51261));
    Span4Mux_h I__12563 (
            .O(N__51529),
            .I(N__51256));
    LocalMux I__12562 (
            .O(N__51526),
            .I(N__51256));
    Span4Mux_v I__12561 (
            .O(N__51521),
            .I(N__51251));
    LocalMux I__12560 (
            .O(N__51516),
            .I(N__51251));
    Span4Mux_h I__12559 (
            .O(N__51511),
            .I(N__51244));
    Span4Mux_v I__12558 (
            .O(N__51504),
            .I(N__51244));
    LocalMux I__12557 (
            .O(N__51501),
            .I(N__51244));
    InMux I__12556 (
            .O(N__51500),
            .I(N__51241));
    Span4Mux_v I__12555 (
            .O(N__51489),
            .I(N__51232));
    LocalMux I__12554 (
            .O(N__51474),
            .I(N__51232));
    LocalMux I__12553 (
            .O(N__51471),
            .I(N__51232));
    LocalMux I__12552 (
            .O(N__51460),
            .I(N__51232));
    InMux I__12551 (
            .O(N__51459),
            .I(N__51229));
    InMux I__12550 (
            .O(N__51458),
            .I(N__51226));
    InMux I__12549 (
            .O(N__51457),
            .I(N__51223));
    Span4Mux_v I__12548 (
            .O(N__51454),
            .I(N__51218));
    LocalMux I__12547 (
            .O(N__51451),
            .I(N__51218));
    Span4Mux_v I__12546 (
            .O(N__51446),
            .I(N__51213));
    LocalMux I__12545 (
            .O(N__51443),
            .I(N__51213));
    LocalMux I__12544 (
            .O(N__51440),
            .I(N__51207));
    LocalMux I__12543 (
            .O(N__51437),
            .I(N__51207));
    InMux I__12542 (
            .O(N__51436),
            .I(N__51204));
    Span4Mux_h I__12541 (
            .O(N__51433),
            .I(N__51191));
    Span4Mux_h I__12540 (
            .O(N__51428),
            .I(N__51191));
    Span4Mux_v I__12539 (
            .O(N__51421),
            .I(N__51191));
    LocalMux I__12538 (
            .O(N__51408),
            .I(N__51191));
    LocalMux I__12537 (
            .O(N__51397),
            .I(N__51191));
    Span4Mux_v I__12536 (
            .O(N__51394),
            .I(N__51184));
    LocalMux I__12535 (
            .O(N__51391),
            .I(N__51184));
    LocalMux I__12534 (
            .O(N__51388),
            .I(N__51184));
    Span4Mux_v I__12533 (
            .O(N__51383),
            .I(N__51175));
    LocalMux I__12532 (
            .O(N__51380),
            .I(N__51175));
    LocalMux I__12531 (
            .O(N__51377),
            .I(N__51175));
    LocalMux I__12530 (
            .O(N__51374),
            .I(N__51175));
    InMux I__12529 (
            .O(N__51373),
            .I(N__51172));
    LocalMux I__12528 (
            .O(N__51370),
            .I(N__51167));
    LocalMux I__12527 (
            .O(N__51367),
            .I(N__51167));
    InMux I__12526 (
            .O(N__51366),
            .I(N__51164));
    InMux I__12525 (
            .O(N__51365),
            .I(N__51161));
    InMux I__12524 (
            .O(N__51364),
            .I(N__51158));
    InMux I__12523 (
            .O(N__51363),
            .I(N__51155));
    Span4Mux_v I__12522 (
            .O(N__51358),
            .I(N__51152));
    LocalMux I__12521 (
            .O(N__51349),
            .I(N__51141));
    LocalMux I__12520 (
            .O(N__51340),
            .I(N__51141));
    Sp12to4 I__12519 (
            .O(N__51337),
            .I(N__51141));
    LocalMux I__12518 (
            .O(N__51334),
            .I(N__51141));
    LocalMux I__12517 (
            .O(N__51325),
            .I(N__51141));
    Span4Mux_h I__12516 (
            .O(N__51322),
            .I(N__51138));
    LocalMux I__12515 (
            .O(N__51315),
            .I(N__51133));
    LocalMux I__12514 (
            .O(N__51312),
            .I(N__51133));
    InMux I__12513 (
            .O(N__51311),
            .I(N__51130));
    InMux I__12512 (
            .O(N__51310),
            .I(N__51117));
    InMux I__12511 (
            .O(N__51309),
            .I(N__51117));
    InMux I__12510 (
            .O(N__51308),
            .I(N__51117));
    InMux I__12509 (
            .O(N__51307),
            .I(N__51117));
    InMux I__12508 (
            .O(N__51306),
            .I(N__51117));
    InMux I__12507 (
            .O(N__51305),
            .I(N__51117));
    InMux I__12506 (
            .O(N__51304),
            .I(N__51114));
    InMux I__12505 (
            .O(N__51303),
            .I(N__51101));
    InMux I__12504 (
            .O(N__51302),
            .I(N__51101));
    InMux I__12503 (
            .O(N__51301),
            .I(N__51101));
    InMux I__12502 (
            .O(N__51300),
            .I(N__51101));
    InMux I__12501 (
            .O(N__51299),
            .I(N__51101));
    InMux I__12500 (
            .O(N__51298),
            .I(N__51101));
    LocalMux I__12499 (
            .O(N__51283),
            .I(N__51096));
    LocalMux I__12498 (
            .O(N__51280),
            .I(N__51096));
    InMux I__12497 (
            .O(N__51279),
            .I(N__51081));
    InMux I__12496 (
            .O(N__51278),
            .I(N__51081));
    InMux I__12495 (
            .O(N__51277),
            .I(N__51081));
    InMux I__12494 (
            .O(N__51276),
            .I(N__51081));
    InMux I__12493 (
            .O(N__51275),
            .I(N__51081));
    InMux I__12492 (
            .O(N__51274),
            .I(N__51081));
    InMux I__12491 (
            .O(N__51273),
            .I(N__51081));
    InMux I__12490 (
            .O(N__51272),
            .I(N__51074));
    InMux I__12489 (
            .O(N__51271),
            .I(N__51074));
    InMux I__12488 (
            .O(N__51270),
            .I(N__51074));
    InMux I__12487 (
            .O(N__51269),
            .I(N__51063));
    InMux I__12486 (
            .O(N__51268),
            .I(N__51063));
    InMux I__12485 (
            .O(N__51267),
            .I(N__51063));
    InMux I__12484 (
            .O(N__51266),
            .I(N__51063));
    InMux I__12483 (
            .O(N__51265),
            .I(N__51063));
    InMux I__12482 (
            .O(N__51264),
            .I(N__51060));
    Span4Mux_h I__12481 (
            .O(N__51261),
            .I(N__51055));
    Span4Mux_v I__12480 (
            .O(N__51256),
            .I(N__51055));
    Span4Mux_v I__12479 (
            .O(N__51251),
            .I(N__51050));
    Span4Mux_v I__12478 (
            .O(N__51244),
            .I(N__51050));
    LocalMux I__12477 (
            .O(N__51241),
            .I(N__51039));
    Span4Mux_v I__12476 (
            .O(N__51232),
            .I(N__51039));
    LocalMux I__12475 (
            .O(N__51229),
            .I(N__51039));
    LocalMux I__12474 (
            .O(N__51226),
            .I(N__51039));
    LocalMux I__12473 (
            .O(N__51223),
            .I(N__51039));
    Span4Mux_v I__12472 (
            .O(N__51218),
            .I(N__51034));
    Span4Mux_h I__12471 (
            .O(N__51213),
            .I(N__51034));
    InMux I__12470 (
            .O(N__51212),
            .I(N__51031));
    Span4Mux_v I__12469 (
            .O(N__51207),
            .I(N__51026));
    LocalMux I__12468 (
            .O(N__51204),
            .I(N__51026));
    InMux I__12467 (
            .O(N__51203),
            .I(N__51023));
    InMux I__12466 (
            .O(N__51202),
            .I(N__51020));
    Span4Mux_v I__12465 (
            .O(N__51191),
            .I(N__51017));
    Span4Mux_v I__12464 (
            .O(N__51184),
            .I(N__51014));
    Span4Mux_v I__12463 (
            .O(N__51175),
            .I(N__50999));
    LocalMux I__12462 (
            .O(N__51172),
            .I(N__50999));
    Span4Mux_v I__12461 (
            .O(N__51167),
            .I(N__50999));
    LocalMux I__12460 (
            .O(N__51164),
            .I(N__50999));
    LocalMux I__12459 (
            .O(N__51161),
            .I(N__50999));
    LocalMux I__12458 (
            .O(N__51158),
            .I(N__50999));
    LocalMux I__12457 (
            .O(N__51155),
            .I(N__50999));
    Sp12to4 I__12456 (
            .O(N__51152),
            .I(N__50992));
    Span12Mux_v I__12455 (
            .O(N__51141),
            .I(N__50992));
    Span4Mux_h I__12454 (
            .O(N__51138),
            .I(N__50987));
    Span4Mux_v I__12453 (
            .O(N__51133),
            .I(N__50987));
    LocalMux I__12452 (
            .O(N__51130),
            .I(N__50968));
    LocalMux I__12451 (
            .O(N__51117),
            .I(N__50968));
    LocalMux I__12450 (
            .O(N__51114),
            .I(N__50968));
    LocalMux I__12449 (
            .O(N__51101),
            .I(N__50968));
    Sp12to4 I__12448 (
            .O(N__51096),
            .I(N__50968));
    LocalMux I__12447 (
            .O(N__51081),
            .I(N__50968));
    LocalMux I__12446 (
            .O(N__51074),
            .I(N__50968));
    LocalMux I__12445 (
            .O(N__51063),
            .I(N__50968));
    LocalMux I__12444 (
            .O(N__51060),
            .I(N__50968));
    Span4Mux_v I__12443 (
            .O(N__51055),
            .I(N__50961));
    Span4Mux_h I__12442 (
            .O(N__51050),
            .I(N__50961));
    Span4Mux_v I__12441 (
            .O(N__51039),
            .I(N__50961));
    Span4Mux_h I__12440 (
            .O(N__51034),
            .I(N__50958));
    LocalMux I__12439 (
            .O(N__51031),
            .I(N__50949));
    Sp12to4 I__12438 (
            .O(N__51026),
            .I(N__50949));
    LocalMux I__12437 (
            .O(N__51023),
            .I(N__50949));
    LocalMux I__12436 (
            .O(N__51020),
            .I(N__50949));
    Span4Mux_h I__12435 (
            .O(N__51017),
            .I(N__50942));
    Span4Mux_v I__12434 (
            .O(N__51014),
            .I(N__50942));
    Span4Mux_v I__12433 (
            .O(N__50999),
            .I(N__50942));
    InMux I__12432 (
            .O(N__50998),
            .I(N__50939));
    InMux I__12431 (
            .O(N__50997),
            .I(N__50936));
    Span12Mux_v I__12430 (
            .O(N__50992),
            .I(N__50933));
    Sp12to4 I__12429 (
            .O(N__50987),
            .I(N__50928));
    Span12Mux_v I__12428 (
            .O(N__50968),
            .I(N__50928));
    Sp12to4 I__12427 (
            .O(N__50961),
            .I(N__50925));
    Sp12to4 I__12426 (
            .O(N__50958),
            .I(N__50920));
    Span12Mux_v I__12425 (
            .O(N__50949),
            .I(N__50920));
    Sp12to4 I__12424 (
            .O(N__50942),
            .I(N__50917));
    LocalMux I__12423 (
            .O(N__50939),
            .I(N__50914));
    LocalMux I__12422 (
            .O(N__50936),
            .I(N__50911));
    Span12Mux_h I__12421 (
            .O(N__50933),
            .I(N__50906));
    Span12Mux_v I__12420 (
            .O(N__50928),
            .I(N__50906));
    Span12Mux_h I__12419 (
            .O(N__50925),
            .I(N__50903));
    Span12Mux_v I__12418 (
            .O(N__50920),
            .I(N__50900));
    Span12Mux_h I__12417 (
            .O(N__50917),
            .I(N__50897));
    Span12Mux_h I__12416 (
            .O(N__50914),
            .I(N__50892));
    Span12Mux_v I__12415 (
            .O(N__50911),
            .I(N__50892));
    Span12Mux_h I__12414 (
            .O(N__50906),
            .I(N__50887));
    Span12Mux_v I__12413 (
            .O(N__50903),
            .I(N__50887));
    Span12Mux_h I__12412 (
            .O(N__50900),
            .I(N__50882));
    Span12Mux_v I__12411 (
            .O(N__50897),
            .I(N__50882));
    Span12Mux_v I__12410 (
            .O(N__50892),
            .I(N__50879));
    Odrv12 I__12409 (
            .O(N__50887),
            .I(wb_rst_i_c));
    Odrv12 I__12408 (
            .O(N__50882),
            .I(wb_rst_i_c));
    Odrv12 I__12407 (
            .O(N__50879),
            .I(wb_rst_i_c));
    InMux I__12406 (
            .O(N__50872),
            .I(N__50869));
    LocalMux I__12405 (
            .O(N__50869),
            .I(N__50865));
    InMux I__12404 (
            .O(N__50868),
            .I(N__50860));
    Span4Mux_h I__12403 (
            .O(N__50865),
            .I(N__50857));
    InMux I__12402 (
            .O(N__50864),
            .I(N__50854));
    CascadeMux I__12401 (
            .O(N__50863),
            .I(N__50851));
    LocalMux I__12400 (
            .O(N__50860),
            .I(N__50847));
    Span4Mux_h I__12399 (
            .O(N__50857),
            .I(N__50842));
    LocalMux I__12398 (
            .O(N__50854),
            .I(N__50842));
    InMux I__12397 (
            .O(N__50851),
            .I(N__50839));
    InMux I__12396 (
            .O(N__50850),
            .I(N__50835));
    Span4Mux_v I__12395 (
            .O(N__50847),
            .I(N__50832));
    Span4Mux_h I__12394 (
            .O(N__50842),
            .I(N__50826));
    LocalMux I__12393 (
            .O(N__50839),
            .I(N__50826));
    InMux I__12392 (
            .O(N__50838),
            .I(N__50823));
    LocalMux I__12391 (
            .O(N__50835),
            .I(N__50819));
    Span4Mux_h I__12390 (
            .O(N__50832),
            .I(N__50816));
    InMux I__12389 (
            .O(N__50831),
            .I(N__50813));
    Span4Mux_h I__12388 (
            .O(N__50826),
            .I(N__50810));
    LocalMux I__12387 (
            .O(N__50823),
            .I(N__50807));
    InMux I__12386 (
            .O(N__50822),
            .I(N__50804));
    Span4Mux_v I__12385 (
            .O(N__50819),
            .I(N__50801));
    Span4Mux_v I__12384 (
            .O(N__50816),
            .I(N__50796));
    LocalMux I__12383 (
            .O(N__50813),
            .I(N__50796));
    Span4Mux_h I__12382 (
            .O(N__50810),
            .I(N__50793));
    Span4Mux_v I__12381 (
            .O(N__50807),
            .I(N__50790));
    LocalMux I__12380 (
            .O(N__50804),
            .I(N__50787));
    Span4Mux_h I__12379 (
            .O(N__50801),
            .I(N__50784));
    Span4Mux_v I__12378 (
            .O(N__50796),
            .I(N__50781));
    Span4Mux_v I__12377 (
            .O(N__50793),
            .I(N__50774));
    Span4Mux_h I__12376 (
            .O(N__50790),
            .I(N__50774));
    Span4Mux_h I__12375 (
            .O(N__50787),
            .I(N__50774));
    Odrv4 I__12374 (
            .O(N__50784),
            .I(N_2140));
    Odrv4 I__12373 (
            .O(N__50781),
            .I(N_2140));
    Odrv4 I__12372 (
            .O(N__50774),
            .I(N_2140));
    CascadeMux I__12371 (
            .O(N__50767),
            .I(N__50762));
    InMux I__12370 (
            .O(N__50766),
            .I(N__50758));
    InMux I__12369 (
            .O(N__50765),
            .I(N__50752));
    InMux I__12368 (
            .O(N__50762),
            .I(N__50752));
    InMux I__12367 (
            .O(N__50761),
            .I(N__50744));
    LocalMux I__12366 (
            .O(N__50758),
            .I(N__50741));
    InMux I__12365 (
            .O(N__50757),
            .I(N__50738));
    LocalMux I__12364 (
            .O(N__50752),
            .I(N__50735));
    InMux I__12363 (
            .O(N__50751),
            .I(N__50726));
    InMux I__12362 (
            .O(N__50750),
            .I(N__50726));
    InMux I__12361 (
            .O(N__50749),
            .I(N__50726));
    InMux I__12360 (
            .O(N__50748),
            .I(N__50726));
    CascadeMux I__12359 (
            .O(N__50747),
            .I(N__50721));
    LocalMux I__12358 (
            .O(N__50744),
            .I(N__50713));
    Span4Mux_h I__12357 (
            .O(N__50741),
            .I(N__50708));
    LocalMux I__12356 (
            .O(N__50738),
            .I(N__50708));
    Span4Mux_h I__12355 (
            .O(N__50735),
            .I(N__50703));
    LocalMux I__12354 (
            .O(N__50726),
            .I(N__50703));
    InMux I__12353 (
            .O(N__50725),
            .I(N__50699));
    InMux I__12352 (
            .O(N__50724),
            .I(N__50696));
    InMux I__12351 (
            .O(N__50721),
            .I(N__50693));
    InMux I__12350 (
            .O(N__50720),
            .I(N__50690));
    InMux I__12349 (
            .O(N__50719),
            .I(N__50687));
    InMux I__12348 (
            .O(N__50718),
            .I(N__50682));
    InMux I__12347 (
            .O(N__50717),
            .I(N__50682));
    InMux I__12346 (
            .O(N__50716),
            .I(N__50679));
    Span4Mux_h I__12345 (
            .O(N__50713),
            .I(N__50673));
    Span4Mux_v I__12344 (
            .O(N__50708),
            .I(N__50670));
    Span4Mux_h I__12343 (
            .O(N__50703),
            .I(N__50667));
    InMux I__12342 (
            .O(N__50702),
            .I(N__50664));
    LocalMux I__12341 (
            .O(N__50699),
            .I(N__50660));
    LocalMux I__12340 (
            .O(N__50696),
            .I(N__50651));
    LocalMux I__12339 (
            .O(N__50693),
            .I(N__50651));
    LocalMux I__12338 (
            .O(N__50690),
            .I(N__50651));
    LocalMux I__12337 (
            .O(N__50687),
            .I(N__50651));
    LocalMux I__12336 (
            .O(N__50682),
            .I(N__50646));
    LocalMux I__12335 (
            .O(N__50679),
            .I(N__50646));
    InMux I__12334 (
            .O(N__50678),
            .I(N__50643));
    InMux I__12333 (
            .O(N__50677),
            .I(N__50640));
    CascadeMux I__12332 (
            .O(N__50676),
            .I(N__50637));
    Span4Mux_v I__12331 (
            .O(N__50673),
            .I(N__50632));
    Span4Mux_h I__12330 (
            .O(N__50670),
            .I(N__50632));
    Span4Mux_h I__12329 (
            .O(N__50667),
            .I(N__50629));
    LocalMux I__12328 (
            .O(N__50664),
            .I(N__50626));
    InMux I__12327 (
            .O(N__50663),
            .I(N__50623));
    Span4Mux_h I__12326 (
            .O(N__50660),
            .I(N__50614));
    Span4Mux_v I__12325 (
            .O(N__50651),
            .I(N__50614));
    Span4Mux_v I__12324 (
            .O(N__50646),
            .I(N__50614));
    LocalMux I__12323 (
            .O(N__50643),
            .I(N__50614));
    LocalMux I__12322 (
            .O(N__50640),
            .I(N__50611));
    InMux I__12321 (
            .O(N__50637),
            .I(N__50608));
    Odrv4 I__12320 (
            .O(N__50632),
            .I(\u0.N_2129 ));
    Odrv4 I__12319 (
            .O(N__50629),
            .I(\u0.N_2129 ));
    Odrv4 I__12318 (
            .O(N__50626),
            .I(\u0.N_2129 ));
    LocalMux I__12317 (
            .O(N__50623),
            .I(\u0.N_2129 ));
    Odrv4 I__12316 (
            .O(N__50614),
            .I(\u0.N_2129 ));
    Odrv12 I__12315 (
            .O(N__50611),
            .I(\u0.N_2129 ));
    LocalMux I__12314 (
            .O(N__50608),
            .I(\u0.N_2129 ));
    IoInMux I__12313 (
            .O(N__50593),
            .I(N__50590));
    LocalMux I__12312 (
            .O(N__50590),
            .I(N__50587));
    Span12Mux_s4_h I__12311 (
            .O(N__50587),
            .I(N__50584));
    Odrv12 I__12310 (
            .O(N__50584),
            .I(N_77));
    InMux I__12309 (
            .O(N__50581),
            .I(N__50578));
    LocalMux I__12308 (
            .O(N__50578),
            .I(N__50570));
    InMux I__12307 (
            .O(N__50577),
            .I(N__50563));
    InMux I__12306 (
            .O(N__50576),
            .I(N__50563));
    InMux I__12305 (
            .O(N__50575),
            .I(N__50563));
    InMux I__12304 (
            .O(N__50574),
            .I(N__50554));
    InMux I__12303 (
            .O(N__50573),
            .I(N__50551));
    Span4Mux_v I__12302 (
            .O(N__50570),
            .I(N__50548));
    LocalMux I__12301 (
            .O(N__50563),
            .I(N__50545));
    InMux I__12300 (
            .O(N__50562),
            .I(N__50542));
    InMux I__12299 (
            .O(N__50561),
            .I(N__50531));
    InMux I__12298 (
            .O(N__50560),
            .I(N__50531));
    InMux I__12297 (
            .O(N__50559),
            .I(N__50531));
    InMux I__12296 (
            .O(N__50558),
            .I(N__50531));
    InMux I__12295 (
            .O(N__50557),
            .I(N__50531));
    LocalMux I__12294 (
            .O(N__50554),
            .I(N__50526));
    LocalMux I__12293 (
            .O(N__50551),
            .I(N__50526));
    Span4Mux_h I__12292 (
            .O(N__50548),
            .I(N__50522));
    Span4Mux_v I__12291 (
            .O(N__50545),
            .I(N__50519));
    LocalMux I__12290 (
            .O(N__50542),
            .I(N__50514));
    LocalMux I__12289 (
            .O(N__50531),
            .I(N__50514));
    Span4Mux_v I__12288 (
            .O(N__50526),
            .I(N__50511));
    InMux I__12287 (
            .O(N__50525),
            .I(N__50508));
    Sp12to4 I__12286 (
            .O(N__50522),
            .I(N__50505));
    Sp12to4 I__12285 (
            .O(N__50519),
            .I(N__50500));
    Span12Mux_v I__12284 (
            .O(N__50514),
            .I(N__50500));
    Sp12to4 I__12283 (
            .O(N__50511),
            .I(N__50497));
    LocalMux I__12282 (
            .O(N__50508),
            .I(N__50494));
    Span12Mux_h I__12281 (
            .O(N__50505),
            .I(N__50491));
    Span12Mux_v I__12280 (
            .O(N__50500),
            .I(N__50488));
    Span12Mux_v I__12279 (
            .O(N__50497),
            .I(N__50485));
    Span12Mux_v I__12278 (
            .O(N__50494),
            .I(N__50482));
    Span12Mux_v I__12277 (
            .O(N__50491),
            .I(N__50477));
    Span12Mux_h I__12276 (
            .O(N__50488),
            .I(N__50477));
    Span12Mux_h I__12275 (
            .O(N__50485),
            .I(N__50472));
    Span12Mux_v I__12274 (
            .O(N__50482),
            .I(N__50472));
    Odrv12 I__12273 (
            .O(N__50477),
            .I(wb_adr_i_c_2));
    Odrv12 I__12272 (
            .O(N__50472),
            .I(wb_adr_i_c_2));
    InMux I__12271 (
            .O(N__50467),
            .I(N__50460));
    InMux I__12270 (
            .O(N__50466),
            .I(N__50454));
    InMux I__12269 (
            .O(N__50465),
            .I(N__50451));
    InMux I__12268 (
            .O(N__50464),
            .I(N__50448));
    InMux I__12267 (
            .O(N__50463),
            .I(N__50445));
    LocalMux I__12266 (
            .O(N__50460),
            .I(N__50439));
    InMux I__12265 (
            .O(N__50459),
            .I(N__50436));
    InMux I__12264 (
            .O(N__50458),
            .I(N__50433));
    InMux I__12263 (
            .O(N__50457),
            .I(N__50430));
    LocalMux I__12262 (
            .O(N__50454),
            .I(N__50427));
    LocalMux I__12261 (
            .O(N__50451),
            .I(N__50422));
    LocalMux I__12260 (
            .O(N__50448),
            .I(N__50422));
    LocalMux I__12259 (
            .O(N__50445),
            .I(N__50419));
    InMux I__12258 (
            .O(N__50444),
            .I(N__50416));
    CascadeMux I__12257 (
            .O(N__50443),
            .I(N__50413));
    CascadeMux I__12256 (
            .O(N__50442),
            .I(N__50410));
    Span4Mux_v I__12255 (
            .O(N__50439),
            .I(N__50401));
    LocalMux I__12254 (
            .O(N__50436),
            .I(N__50401));
    LocalMux I__12253 (
            .O(N__50433),
            .I(N__50401));
    LocalMux I__12252 (
            .O(N__50430),
            .I(N__50398));
    Span4Mux_h I__12251 (
            .O(N__50427),
            .I(N__50393));
    Span4Mux_v I__12250 (
            .O(N__50422),
            .I(N__50393));
    Span4Mux_v I__12249 (
            .O(N__50419),
            .I(N__50388));
    LocalMux I__12248 (
            .O(N__50416),
            .I(N__50388));
    InMux I__12247 (
            .O(N__50413),
            .I(N__50385));
    InMux I__12246 (
            .O(N__50410),
            .I(N__50378));
    InMux I__12245 (
            .O(N__50409),
            .I(N__50378));
    InMux I__12244 (
            .O(N__50408),
            .I(N__50378));
    Span4Mux_v I__12243 (
            .O(N__50401),
            .I(N__50374));
    Span4Mux_v I__12242 (
            .O(N__50398),
            .I(N__50371));
    Span4Mux_h I__12241 (
            .O(N__50393),
            .I(N__50360));
    Span4Mux_v I__12240 (
            .O(N__50388),
            .I(N__50360));
    LocalMux I__12239 (
            .O(N__50385),
            .I(N__50360));
    LocalMux I__12238 (
            .O(N__50378),
            .I(N__50360));
    InMux I__12237 (
            .O(N__50377),
            .I(N__50357));
    Span4Mux_h I__12236 (
            .O(N__50374),
            .I(N__50354));
    Span4Mux_h I__12235 (
            .O(N__50371),
            .I(N__50351));
    InMux I__12234 (
            .O(N__50370),
            .I(N__50348));
    InMux I__12233 (
            .O(N__50369),
            .I(N__50345));
    Span4Mux_v I__12232 (
            .O(N__50360),
            .I(N__50342));
    LocalMux I__12231 (
            .O(N__50357),
            .I(N__50339));
    Span4Mux_h I__12230 (
            .O(N__50354),
            .I(N__50336));
    Span4Mux_v I__12229 (
            .O(N__50351),
            .I(N__50331));
    LocalMux I__12228 (
            .O(N__50348),
            .I(N__50331));
    LocalMux I__12227 (
            .O(N__50345),
            .I(N__50328));
    Span4Mux_h I__12226 (
            .O(N__50342),
            .I(N__50323));
    Span4Mux_v I__12225 (
            .O(N__50339),
            .I(N__50323));
    Span4Mux_h I__12224 (
            .O(N__50336),
            .I(N__50318));
    Span4Mux_v I__12223 (
            .O(N__50331),
            .I(N__50318));
    Span12Mux_v I__12222 (
            .O(N__50328),
            .I(N__50315));
    Sp12to4 I__12221 (
            .O(N__50323),
            .I(N__50310));
    Sp12to4 I__12220 (
            .O(N__50318),
            .I(N__50310));
    Span12Mux_v I__12219 (
            .O(N__50315),
            .I(N__50307));
    Span12Mux_h I__12218 (
            .O(N__50310),
            .I(N__50304));
    Span12Mux_h I__12217 (
            .O(N__50307),
            .I(N__50301));
    Span12Mux_v I__12216 (
            .O(N__50304),
            .I(N__50298));
    Odrv12 I__12215 (
            .O(N__50301),
            .I(wb_adr_i_c_5));
    Odrv12 I__12214 (
            .O(N__50298),
            .I(wb_adr_i_c_5));
    CascadeMux I__12213 (
            .O(N__50293),
            .I(N__50285));
    InMux I__12212 (
            .O(N__50292),
            .I(N__50273));
    InMux I__12211 (
            .O(N__50291),
            .I(N__50273));
    InMux I__12210 (
            .O(N__50290),
            .I(N__50273));
    InMux I__12209 (
            .O(N__50289),
            .I(N__50273));
    InMux I__12208 (
            .O(N__50288),
            .I(N__50273));
    InMux I__12207 (
            .O(N__50285),
            .I(N__50270));
    CascadeMux I__12206 (
            .O(N__50284),
            .I(N__50267));
    LocalMux I__12205 (
            .O(N__50273),
            .I(N__50264));
    LocalMux I__12204 (
            .O(N__50270),
            .I(N__50261));
    InMux I__12203 (
            .O(N__50267),
            .I(N__50258));
    Span4Mux_v I__12202 (
            .O(N__50264),
            .I(N__50254));
    Span4Mux_h I__12201 (
            .O(N__50261),
            .I(N__50251));
    LocalMux I__12200 (
            .O(N__50258),
            .I(N__50248));
    InMux I__12199 (
            .O(N__50257),
            .I(N__50245));
    Span4Mux_h I__12198 (
            .O(N__50254),
            .I(N__50242));
    Span4Mux_h I__12197 (
            .O(N__50251),
            .I(N__50237));
    Span4Mux_v I__12196 (
            .O(N__50248),
            .I(N__50237));
    LocalMux I__12195 (
            .O(N__50245),
            .I(N__50234));
    Odrv4 I__12194 (
            .O(N__50242),
            .I(\u0.N_2143 ));
    Odrv4 I__12193 (
            .O(N__50237),
            .I(\u0.N_2143 ));
    Odrv4 I__12192 (
            .O(N__50234),
            .I(\u0.N_2143 ));
    IoInMux I__12191 (
            .O(N__50227),
            .I(N__50224));
    LocalMux I__12190 (
            .O(N__50224),
            .I(N__50221));
    Span12Mux_s4_v I__12189 (
            .O(N__50221),
            .I(N__50218));
    Span12Mux_h I__12188 (
            .O(N__50218),
            .I(N__50215));
    Odrv12 I__12187 (
            .O(N__50215),
            .I(wb_dat_o_c_9));
    InMux I__12186 (
            .O(N__50212),
            .I(N__50209));
    LocalMux I__12185 (
            .O(N__50209),
            .I(N__50202));
    InMux I__12184 (
            .O(N__50208),
            .I(N__50199));
    InMux I__12183 (
            .O(N__50207),
            .I(N__50195));
    InMux I__12182 (
            .O(N__50206),
            .I(N__50190));
    InMux I__12181 (
            .O(N__50205),
            .I(N__50185));
    Span4Mux_h I__12180 (
            .O(N__50202),
            .I(N__50180));
    LocalMux I__12179 (
            .O(N__50199),
            .I(N__50180));
    InMux I__12178 (
            .O(N__50198),
            .I(N__50176));
    LocalMux I__12177 (
            .O(N__50195),
            .I(N__50162));
    InMux I__12176 (
            .O(N__50194),
            .I(N__50157));
    InMux I__12175 (
            .O(N__50193),
            .I(N__50157));
    LocalMux I__12174 (
            .O(N__50190),
            .I(N__50154));
    InMux I__12173 (
            .O(N__50189),
            .I(N__50147));
    InMux I__12172 (
            .O(N__50188),
            .I(N__50147));
    LocalMux I__12171 (
            .O(N__50185),
            .I(N__50142));
    Span4Mux_h I__12170 (
            .O(N__50180),
            .I(N__50142));
    InMux I__12169 (
            .O(N__50179),
            .I(N__50131));
    LocalMux I__12168 (
            .O(N__50176),
            .I(N__50128));
    InMux I__12167 (
            .O(N__50175),
            .I(N__50125));
    InMux I__12166 (
            .O(N__50174),
            .I(N__50120));
    InMux I__12165 (
            .O(N__50173),
            .I(N__50120));
    InMux I__12164 (
            .O(N__50172),
            .I(N__50115));
    InMux I__12163 (
            .O(N__50171),
            .I(N__50115));
    InMux I__12162 (
            .O(N__50170),
            .I(N__50106));
    InMux I__12161 (
            .O(N__50169),
            .I(N__50106));
    InMux I__12160 (
            .O(N__50168),
            .I(N__50101));
    InMux I__12159 (
            .O(N__50167),
            .I(N__50101));
    InMux I__12158 (
            .O(N__50166),
            .I(N__50096));
    InMux I__12157 (
            .O(N__50165),
            .I(N__50096));
    Span4Mux_h I__12156 (
            .O(N__50162),
            .I(N__50089));
    LocalMux I__12155 (
            .O(N__50157),
            .I(N__50089));
    Span4Mux_h I__12154 (
            .O(N__50154),
            .I(N__50089));
    InMux I__12153 (
            .O(N__50153),
            .I(N__50084));
    InMux I__12152 (
            .O(N__50152),
            .I(N__50084));
    LocalMux I__12151 (
            .O(N__50147),
            .I(N__50081));
    IoSpan4Mux I__12150 (
            .O(N__50142),
            .I(N__50078));
    InMux I__12149 (
            .O(N__50141),
            .I(N__50075));
    InMux I__12148 (
            .O(N__50140),
            .I(N__50070));
    InMux I__12147 (
            .O(N__50139),
            .I(N__50070));
    InMux I__12146 (
            .O(N__50138),
            .I(N__50065));
    InMux I__12145 (
            .O(N__50137),
            .I(N__50065));
    CascadeMux I__12144 (
            .O(N__50136),
            .I(N__50061));
    InMux I__12143 (
            .O(N__50135),
            .I(N__50053));
    InMux I__12142 (
            .O(N__50134),
            .I(N__50053));
    LocalMux I__12141 (
            .O(N__50131),
            .I(N__50049));
    Span4Mux_h I__12140 (
            .O(N__50128),
            .I(N__50040));
    LocalMux I__12139 (
            .O(N__50125),
            .I(N__50040));
    LocalMux I__12138 (
            .O(N__50120),
            .I(N__50040));
    LocalMux I__12137 (
            .O(N__50115),
            .I(N__50040));
    InMux I__12136 (
            .O(N__50114),
            .I(N__50033));
    InMux I__12135 (
            .O(N__50113),
            .I(N__50030));
    InMux I__12134 (
            .O(N__50112),
            .I(N__50027));
    InMux I__12133 (
            .O(N__50111),
            .I(N__50024));
    LocalMux I__12132 (
            .O(N__50106),
            .I(N__50021));
    LocalMux I__12131 (
            .O(N__50101),
            .I(N__50003));
    LocalMux I__12130 (
            .O(N__50096),
            .I(N__50003));
    Span4Mux_v I__12129 (
            .O(N__50089),
            .I(N__50003));
    LocalMux I__12128 (
            .O(N__50084),
            .I(N__50003));
    Span4Mux_h I__12127 (
            .O(N__50081),
            .I(N__49996));
    Span4Mux_s1_v I__12126 (
            .O(N__50078),
            .I(N__49996));
    LocalMux I__12125 (
            .O(N__50075),
            .I(N__49996));
    LocalMux I__12124 (
            .O(N__50070),
            .I(N__49991));
    LocalMux I__12123 (
            .O(N__50065),
            .I(N__49991));
    InMux I__12122 (
            .O(N__50064),
            .I(N__49984));
    InMux I__12121 (
            .O(N__50061),
            .I(N__49984));
    InMux I__12120 (
            .O(N__50060),
            .I(N__49984));
    InMux I__12119 (
            .O(N__50059),
            .I(N__49979));
    InMux I__12118 (
            .O(N__50058),
            .I(N__49979));
    LocalMux I__12117 (
            .O(N__50053),
            .I(N__49974));
    InMux I__12116 (
            .O(N__50052),
            .I(N__49971));
    Span4Mux_h I__12115 (
            .O(N__50049),
            .I(N__49966));
    Span4Mux_v I__12114 (
            .O(N__50040),
            .I(N__49966));
    InMux I__12113 (
            .O(N__50039),
            .I(N__49961));
    InMux I__12112 (
            .O(N__50038),
            .I(N__49961));
    InMux I__12111 (
            .O(N__50037),
            .I(N__49956));
    InMux I__12110 (
            .O(N__50036),
            .I(N__49956));
    LocalMux I__12109 (
            .O(N__50033),
            .I(N__49953));
    LocalMux I__12108 (
            .O(N__50030),
            .I(N__49944));
    LocalMux I__12107 (
            .O(N__50027),
            .I(N__49944));
    LocalMux I__12106 (
            .O(N__50024),
            .I(N__49944));
    Span4Mux_h I__12105 (
            .O(N__50021),
            .I(N__49944));
    InMux I__12104 (
            .O(N__50020),
            .I(N__49939));
    InMux I__12103 (
            .O(N__50019),
            .I(N__49939));
    InMux I__12102 (
            .O(N__50018),
            .I(N__49934));
    InMux I__12101 (
            .O(N__50017),
            .I(N__49929));
    InMux I__12100 (
            .O(N__50016),
            .I(N__49929));
    InMux I__12099 (
            .O(N__50015),
            .I(N__49924));
    InMux I__12098 (
            .O(N__50014),
            .I(N__49924));
    InMux I__12097 (
            .O(N__50013),
            .I(N__49919));
    InMux I__12096 (
            .O(N__50012),
            .I(N__49919));
    Span4Mux_h I__12095 (
            .O(N__50003),
            .I(N__49912));
    Span4Mux_v I__12094 (
            .O(N__49996),
            .I(N__49905));
    Span4Mux_v I__12093 (
            .O(N__49991),
            .I(N__49905));
    LocalMux I__12092 (
            .O(N__49984),
            .I(N__49905));
    LocalMux I__12091 (
            .O(N__49979),
            .I(N__49902));
    InMux I__12090 (
            .O(N__49978),
            .I(N__49897));
    InMux I__12089 (
            .O(N__49977),
            .I(N__49897));
    Span4Mux_h I__12088 (
            .O(N__49974),
            .I(N__49892));
    LocalMux I__12087 (
            .O(N__49971),
            .I(N__49892));
    Span4Mux_h I__12086 (
            .O(N__49966),
            .I(N__49885));
    LocalMux I__12085 (
            .O(N__49961),
            .I(N__49885));
    LocalMux I__12084 (
            .O(N__49956),
            .I(N__49885));
    Span4Mux_h I__12083 (
            .O(N__49953),
            .I(N__49878));
    Span4Mux_v I__12082 (
            .O(N__49944),
            .I(N__49878));
    LocalMux I__12081 (
            .O(N__49939),
            .I(N__49878));
    InMux I__12080 (
            .O(N__49938),
            .I(N__49873));
    InMux I__12079 (
            .O(N__49937),
            .I(N__49873));
    LocalMux I__12078 (
            .O(N__49934),
            .I(N__49864));
    LocalMux I__12077 (
            .O(N__49929),
            .I(N__49864));
    LocalMux I__12076 (
            .O(N__49924),
            .I(N__49864));
    LocalMux I__12075 (
            .O(N__49919),
            .I(N__49864));
    InMux I__12074 (
            .O(N__49918),
            .I(N__49859));
    InMux I__12073 (
            .O(N__49917),
            .I(N__49859));
    InMux I__12072 (
            .O(N__49916),
            .I(N__49854));
    InMux I__12071 (
            .O(N__49915),
            .I(N__49854));
    Span4Mux_h I__12070 (
            .O(N__49912),
            .I(N__49848));
    Span4Mux_v I__12069 (
            .O(N__49905),
            .I(N__49841));
    Span4Mux_h I__12068 (
            .O(N__49902),
            .I(N__49841));
    LocalMux I__12067 (
            .O(N__49897),
            .I(N__49841));
    Span4Mux_v I__12066 (
            .O(N__49892),
            .I(N__49836));
    Span4Mux_h I__12065 (
            .O(N__49885),
            .I(N__49836));
    Span4Mux_v I__12064 (
            .O(N__49878),
            .I(N__49829));
    LocalMux I__12063 (
            .O(N__49873),
            .I(N__49829));
    Span4Mux_v I__12062 (
            .O(N__49864),
            .I(N__49824));
    LocalMux I__12061 (
            .O(N__49859),
            .I(N__49824));
    LocalMux I__12060 (
            .O(N__49854),
            .I(N__49821));
    InMux I__12059 (
            .O(N__49853),
            .I(N__49814));
    InMux I__12058 (
            .O(N__49852),
            .I(N__49814));
    InMux I__12057 (
            .O(N__49851),
            .I(N__49814));
    Span4Mux_v I__12056 (
            .O(N__49848),
            .I(N__49811));
    Span4Mux_h I__12055 (
            .O(N__49841),
            .I(N__49806));
    Span4Mux_v I__12054 (
            .O(N__49836),
            .I(N__49806));
    CascadeMux I__12053 (
            .O(N__49835),
            .I(N__49803));
    CascadeMux I__12052 (
            .O(N__49834),
            .I(N__49798));
    Span4Mux_h I__12051 (
            .O(N__49829),
            .I(N__49794));
    Span4Mux_h I__12050 (
            .O(N__49824),
            .I(N__49787));
    Span4Mux_h I__12049 (
            .O(N__49821),
            .I(N__49787));
    LocalMux I__12048 (
            .O(N__49814),
            .I(N__49787));
    Span4Mux_v I__12047 (
            .O(N__49811),
            .I(N__49784));
    Span4Mux_v I__12046 (
            .O(N__49806),
            .I(N__49781));
    InMux I__12045 (
            .O(N__49803),
            .I(N__49778));
    InMux I__12044 (
            .O(N__49802),
            .I(N__49775));
    InMux I__12043 (
            .O(N__49801),
            .I(N__49768));
    InMux I__12042 (
            .O(N__49798),
            .I(N__49768));
    InMux I__12041 (
            .O(N__49797),
            .I(N__49768));
    Span4Mux_v I__12040 (
            .O(N__49794),
            .I(N__49763));
    Span4Mux_v I__12039 (
            .O(N__49787),
            .I(N__49763));
    Odrv4 I__12038 (
            .O(N__49784),
            .I(\u1.DMA_control.rd_ptr_1 ));
    Odrv4 I__12037 (
            .O(N__49781),
            .I(\u1.DMA_control.rd_ptr_1 ));
    LocalMux I__12036 (
            .O(N__49778),
            .I(\u1.DMA_control.rd_ptr_1 ));
    LocalMux I__12035 (
            .O(N__49775),
            .I(\u1.DMA_control.rd_ptr_1 ));
    LocalMux I__12034 (
            .O(N__49768),
            .I(\u1.DMA_control.rd_ptr_1 ));
    Odrv4 I__12033 (
            .O(N__49763),
            .I(\u1.DMA_control.rd_ptr_1 ));
    InMux I__12032 (
            .O(N__49750),
            .I(N__49747));
    LocalMux I__12031 (
            .O(N__49747),
            .I(N__49744));
    Span4Mux_v I__12030 (
            .O(N__49744),
            .I(N__49741));
    Odrv4 I__12029 (
            .O(N__49741),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_16 ));
    InMux I__12028 (
            .O(N__49738),
            .I(N__49735));
    LocalMux I__12027 (
            .O(N__49735),
            .I(N__49732));
    Odrv12 I__12026 (
            .O(N__49732),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIC3GTZ0Z_16 ));
    InMux I__12025 (
            .O(N__49729),
            .I(N__49726));
    LocalMux I__12024 (
            .O(N__49726),
            .I(N__49723));
    Odrv12 I__12023 (
            .O(N__49723),
            .I(mem_mem_ram6__RNID2B71_16));
    InMux I__12022 (
            .O(N__49720),
            .I(N__49717));
    LocalMux I__12021 (
            .O(N__49717),
            .I(N__49713));
    InMux I__12020 (
            .O(N__49716),
            .I(N__49710));
    Span12Mux_h I__12019 (
            .O(N__49713),
            .I(N__49707));
    LocalMux I__12018 (
            .O(N__49710),
            .I(PIO_cmdport_Teoc_5));
    Odrv12 I__12017 (
            .O(N__49707),
            .I(PIO_cmdport_Teoc_5));
    CEMux I__12016 (
            .O(N__49702),
            .I(N__49663));
    CEMux I__12015 (
            .O(N__49701),
            .I(N__49663));
    CEMux I__12014 (
            .O(N__49700),
            .I(N__49663));
    CEMux I__12013 (
            .O(N__49699),
            .I(N__49663));
    CEMux I__12012 (
            .O(N__49698),
            .I(N__49663));
    CEMux I__12011 (
            .O(N__49697),
            .I(N__49663));
    CEMux I__12010 (
            .O(N__49696),
            .I(N__49663));
    CEMux I__12009 (
            .O(N__49695),
            .I(N__49663));
    CEMux I__12008 (
            .O(N__49694),
            .I(N__49663));
    CEMux I__12007 (
            .O(N__49693),
            .I(N__49663));
    CEMux I__12006 (
            .O(N__49692),
            .I(N__49663));
    CEMux I__12005 (
            .O(N__49691),
            .I(N__49663));
    CEMux I__12004 (
            .O(N__49690),
            .I(N__49663));
    GlobalMux I__12003 (
            .O(N__49663),
            .I(N__49660));
    gio2CtrlBuf I__12002 (
            .O(N__49660),
            .I(N_448_g));
    InMux I__12001 (
            .O(N__49657),
            .I(N__49654));
    LocalMux I__12000 (
            .O(N__49654),
            .I(N__49651));
    Span4Mux_v I__11999 (
            .O(N__49651),
            .I(N__49648));
    Odrv4 I__11998 (
            .O(N__49648),
            .I(\u0.dat_o_0_a2_i_2_17 ));
    InMux I__11997 (
            .O(N__49645),
            .I(N__49641));
    InMux I__11996 (
            .O(N__49644),
            .I(N__49638));
    LocalMux I__11995 (
            .O(N__49641),
            .I(N__49634));
    LocalMux I__11994 (
            .O(N__49638),
            .I(N__49631));
    InMux I__11993 (
            .O(N__49637),
            .I(N__49628));
    Span4Mux_v I__11992 (
            .O(N__49634),
            .I(N__49625));
    Span4Mux_v I__11991 (
            .O(N__49631),
            .I(N__49620));
    LocalMux I__11990 (
            .O(N__49628),
            .I(N__49617));
    Span4Mux_h I__11989 (
            .O(N__49625),
            .I(N__49614));
    InMux I__11988 (
            .O(N__49624),
            .I(N__49611));
    InMux I__11987 (
            .O(N__49623),
            .I(N__49608));
    Span4Mux_h I__11986 (
            .O(N__49620),
            .I(N__49601));
    Span4Mux_v I__11985 (
            .O(N__49617),
            .I(N__49601));
    Sp12to4 I__11984 (
            .O(N__49614),
            .I(N__49596));
    LocalMux I__11983 (
            .O(N__49611),
            .I(N__49596));
    LocalMux I__11982 (
            .O(N__49608),
            .I(N__49593));
    InMux I__11981 (
            .O(N__49607),
            .I(N__49590));
    InMux I__11980 (
            .O(N__49606),
            .I(N__49587));
    Odrv4 I__11979 (
            .O(N__49601),
            .I(\u0.N_1374 ));
    Odrv12 I__11978 (
            .O(N__49596),
            .I(\u0.N_1374 ));
    Odrv12 I__11977 (
            .O(N__49593),
            .I(\u0.N_1374 ));
    LocalMux I__11976 (
            .O(N__49590),
            .I(\u0.N_1374 ));
    LocalMux I__11975 (
            .O(N__49587),
            .I(\u0.N_1374 ));
    InMux I__11974 (
            .O(N__49576),
            .I(N__49573));
    LocalMux I__11973 (
            .O(N__49573),
            .I(N__49570));
    Odrv4 I__11972 (
            .O(N__49570),
            .I(\u0.N_1554 ));
    IoInMux I__11971 (
            .O(N__49567),
            .I(N__49564));
    LocalMux I__11970 (
            .O(N__49564),
            .I(N__49561));
    IoSpan4Mux I__11969 (
            .O(N__49561),
            .I(N__49558));
    Span4Mux_s2_h I__11968 (
            .O(N__49558),
            .I(N__49555));
    Sp12to4 I__11967 (
            .O(N__49555),
            .I(N__49552));
    Odrv12 I__11966 (
            .O(N__49552),
            .I(N_209_i));
    InMux I__11965 (
            .O(N__49549),
            .I(N__49546));
    LocalMux I__11964 (
            .O(N__49546),
            .I(N__49541));
    InMux I__11963 (
            .O(N__49545),
            .I(N__49538));
    InMux I__11962 (
            .O(N__49544),
            .I(N__49535));
    Span4Mux_v I__11961 (
            .O(N__49541),
            .I(N__49530));
    LocalMux I__11960 (
            .O(N__49538),
            .I(N__49527));
    LocalMux I__11959 (
            .O(N__49535),
            .I(N__49523));
    InMux I__11958 (
            .O(N__49534),
            .I(N__49520));
    InMux I__11957 (
            .O(N__49533),
            .I(N__49517));
    Span4Mux_h I__11956 (
            .O(N__49530),
            .I(N__49512));
    Span4Mux_v I__11955 (
            .O(N__49527),
            .I(N__49512));
    InMux I__11954 (
            .O(N__49526),
            .I(N__49509));
    Span4Mux_v I__11953 (
            .O(N__49523),
            .I(N__49502));
    LocalMux I__11952 (
            .O(N__49520),
            .I(N__49502));
    LocalMux I__11951 (
            .O(N__49517),
            .I(N__49502));
    Span4Mux_h I__11950 (
            .O(N__49512),
            .I(N__49497));
    LocalMux I__11949 (
            .O(N__49509),
            .I(N__49494));
    Span4Mux_v I__11948 (
            .O(N__49502),
            .I(N__49490));
    InMux I__11947 (
            .O(N__49501),
            .I(N__49485));
    InMux I__11946 (
            .O(N__49500),
            .I(N__49485));
    Span4Mux_v I__11945 (
            .O(N__49497),
            .I(N__49480));
    Span4Mux_v I__11944 (
            .O(N__49494),
            .I(N__49480));
    InMux I__11943 (
            .O(N__49493),
            .I(N__49477));
    Span4Mux_h I__11942 (
            .O(N__49490),
            .I(N__49472));
    LocalMux I__11941 (
            .O(N__49485),
            .I(N__49472));
    Span4Mux_h I__11940 (
            .O(N__49480),
            .I(N__49469));
    LocalMux I__11939 (
            .O(N__49477),
            .I(N__49466));
    Span4Mux_v I__11938 (
            .O(N__49472),
            .I(N__49462));
    Span4Mux_v I__11937 (
            .O(N__49469),
            .I(N__49457));
    Span4Mux_v I__11936 (
            .O(N__49466),
            .I(N__49457));
    InMux I__11935 (
            .O(N__49465),
            .I(N__49454));
    Span4Mux_v I__11934 (
            .O(N__49462),
            .I(N__49451));
    Span4Mux_v I__11933 (
            .O(N__49457),
            .I(N__49448));
    LocalMux I__11932 (
            .O(N__49454),
            .I(N__49445));
    Span4Mux_v I__11931 (
            .O(N__49451),
            .I(N__49442));
    Span4Mux_v I__11930 (
            .O(N__49448),
            .I(N__49439));
    Span12Mux_v I__11929 (
            .O(N__49445),
            .I(N__49436));
    Sp12to4 I__11928 (
            .O(N__49442),
            .I(N__49431));
    Sp12to4 I__11927 (
            .O(N__49439),
            .I(N__49431));
    Span12Mux_v I__11926 (
            .O(N__49436),
            .I(N__49428));
    Span12Mux_h I__11925 (
            .O(N__49431),
            .I(N__49425));
    Span12Mux_h I__11924 (
            .O(N__49428),
            .I(N__49422));
    Odrv12 I__11923 (
            .O(N__49425),
            .I(wb_dat_i_c_0));
    Odrv12 I__11922 (
            .O(N__49422),
            .I(wb_dat_i_c_0));
    InMux I__11921 (
            .O(N__49417),
            .I(N__49413));
    InMux I__11920 (
            .O(N__49416),
            .I(N__49410));
    LocalMux I__11919 (
            .O(N__49413),
            .I(N__49407));
    LocalMux I__11918 (
            .O(N__49410),
            .I(N__49404));
    Span4Mux_v I__11917 (
            .O(N__49407),
            .I(N__49401));
    Span4Mux_v I__11916 (
            .O(N__49404),
            .I(N__49398));
    Span4Mux_h I__11915 (
            .O(N__49401),
            .I(N__49395));
    Span4Mux_h I__11914 (
            .O(N__49398),
            .I(N__49392));
    Span4Mux_h I__11913 (
            .O(N__49395),
            .I(N__49389));
    Odrv4 I__11912 (
            .O(N__49392),
            .I(PIO_dport0_T1_0));
    Odrv4 I__11911 (
            .O(N__49389),
            .I(PIO_dport0_T1_0));
    CEMux I__11910 (
            .O(N__49384),
            .I(N__49354));
    CEMux I__11909 (
            .O(N__49383),
            .I(N__49354));
    CEMux I__11908 (
            .O(N__49382),
            .I(N__49354));
    CEMux I__11907 (
            .O(N__49381),
            .I(N__49354));
    CEMux I__11906 (
            .O(N__49380),
            .I(N__49354));
    CEMux I__11905 (
            .O(N__49379),
            .I(N__49354));
    CEMux I__11904 (
            .O(N__49378),
            .I(N__49354));
    CEMux I__11903 (
            .O(N__49377),
            .I(N__49354));
    CEMux I__11902 (
            .O(N__49376),
            .I(N__49354));
    CEMux I__11901 (
            .O(N__49375),
            .I(N__49354));
    GlobalMux I__11900 (
            .O(N__49354),
            .I(N__49351));
    gio2CtrlBuf I__11899 (
            .O(N__49351),
            .I(N_77_g));
    InMux I__11898 (
            .O(N__49348),
            .I(N__49345));
    LocalMux I__11897 (
            .O(N__49345),
            .I(N__49339));
    InMux I__11896 (
            .O(N__49344),
            .I(N__49336));
    InMux I__11895 (
            .O(N__49343),
            .I(N__49332));
    InMux I__11894 (
            .O(N__49342),
            .I(N__49329));
    Span4Mux_v I__11893 (
            .O(N__49339),
            .I(N__49326));
    LocalMux I__11892 (
            .O(N__49336),
            .I(N__49323));
    InMux I__11891 (
            .O(N__49335),
            .I(N__49320));
    LocalMux I__11890 (
            .O(N__49332),
            .I(N__49315));
    LocalMux I__11889 (
            .O(N__49329),
            .I(N__49315));
    Span4Mux_v I__11888 (
            .O(N__49326),
            .I(N__49311));
    Span4Mux_h I__11887 (
            .O(N__49323),
            .I(N__49306));
    LocalMux I__11886 (
            .O(N__49320),
            .I(N__49306));
    Span4Mux_v I__11885 (
            .O(N__49315),
            .I(N__49303));
    InMux I__11884 (
            .O(N__49314),
            .I(N__49300));
    Sp12to4 I__11883 (
            .O(N__49311),
            .I(N__49297));
    Span4Mux_v I__11882 (
            .O(N__49306),
            .I(N__49294));
    Span4Mux_h I__11881 (
            .O(N__49303),
            .I(N__49289));
    LocalMux I__11880 (
            .O(N__49300),
            .I(N__49289));
    Span12Mux_h I__11879 (
            .O(N__49297),
            .I(N__49285));
    Span4Mux_h I__11878 (
            .O(N__49294),
            .I(N__49282));
    Sp12to4 I__11877 (
            .O(N__49289),
            .I(N__49279));
    InMux I__11876 (
            .O(N__49288),
            .I(N__49276));
    Span12Mux_h I__11875 (
            .O(N__49285),
            .I(N__49273));
    Sp12to4 I__11874 (
            .O(N__49282),
            .I(N__49266));
    Span12Mux_v I__11873 (
            .O(N__49279),
            .I(N__49266));
    LocalMux I__11872 (
            .O(N__49276),
            .I(N__49266));
    Span12Mux_v I__11871 (
            .O(N__49273),
            .I(N__49263));
    Span12Mux_h I__11870 (
            .O(N__49266),
            .I(N__49260));
    Odrv12 I__11869 (
            .O(N__49263),
            .I(wb_dat_i_c_29));
    Odrv12 I__11868 (
            .O(N__49260),
            .I(wb_dat_i_c_29));
    InMux I__11867 (
            .O(N__49255),
            .I(N__49252));
    LocalMux I__11866 (
            .O(N__49252),
            .I(N__49249));
    Odrv4 I__11865 (
            .O(N__49249),
            .I(\u0.CtrlRegZ0Z_29 ));
    InMux I__11864 (
            .O(N__49246),
            .I(N__49243));
    LocalMux I__11863 (
            .O(N__49243),
            .I(N__49239));
    InMux I__11862 (
            .O(N__49242),
            .I(N__49236));
    Span4Mux_v I__11861 (
            .O(N__49239),
            .I(N__49233));
    LocalMux I__11860 (
            .O(N__49236),
            .I(N__49230));
    Span4Mux_h I__11859 (
            .O(N__49233),
            .I(N__49227));
    Span4Mux_h I__11858 (
            .O(N__49230),
            .I(N__49224));
    Odrv4 I__11857 (
            .O(N__49227),
            .I(PIO_dport0_T4_7));
    Odrv4 I__11856 (
            .O(N__49224),
            .I(PIO_dport0_T4_7));
    InMux I__11855 (
            .O(N__49219),
            .I(N__49215));
    CascadeMux I__11854 (
            .O(N__49218),
            .I(N__49212));
    LocalMux I__11853 (
            .O(N__49215),
            .I(N__49209));
    InMux I__11852 (
            .O(N__49212),
            .I(N__49206));
    Span12Mux_h I__11851 (
            .O(N__49209),
            .I(N__49203));
    LocalMux I__11850 (
            .O(N__49206),
            .I(N__49200));
    Odrv12 I__11849 (
            .O(N__49203),
            .I(PIO_dport1_T4_7));
    Odrv12 I__11848 (
            .O(N__49200),
            .I(PIO_dport1_T4_7));
    InMux I__11847 (
            .O(N__49195),
            .I(N__49192));
    LocalMux I__11846 (
            .O(N__49192),
            .I(N__49189));
    Span4Mux_v I__11845 (
            .O(N__49189),
            .I(N__49186));
    Odrv4 I__11844 (
            .O(N__49186),
            .I(\u0.dat_o_i_0_1_23 ));
    InMux I__11843 (
            .O(N__49183),
            .I(N__49180));
    LocalMux I__11842 (
            .O(N__49180),
            .I(N__49177));
    Odrv12 I__11841 (
            .O(N__49177),
            .I(\u0.dat_o_i_i_0_25 ));
    InMux I__11840 (
            .O(N__49174),
            .I(N__49171));
    LocalMux I__11839 (
            .O(N__49171),
            .I(N__49168));
    Odrv12 I__11838 (
            .O(N__49168),
            .I(\u0.dat_o_i_i_4_25 ));
    CascadeMux I__11837 (
            .O(N__49165),
            .I(N__49162));
    InMux I__11836 (
            .O(N__49162),
            .I(N__49159));
    LocalMux I__11835 (
            .O(N__49159),
            .I(N__49155));
    InMux I__11834 (
            .O(N__49158),
            .I(N__49152));
    Span4Mux_v I__11833 (
            .O(N__49155),
            .I(N__49149));
    LocalMux I__11832 (
            .O(N__49152),
            .I(N__49146));
    Sp12to4 I__11831 (
            .O(N__49149),
            .I(N__49143));
    Span4Mux_s3_h I__11830 (
            .O(N__49146),
            .I(N__49140));
    Span12Mux_h I__11829 (
            .O(N__49143),
            .I(N__49137));
    Span4Mux_h I__11828 (
            .O(N__49140),
            .I(N__49134));
    Odrv12 I__11827 (
            .O(N__49137),
            .I(DMA_dev1_Teoc_1));
    Odrv4 I__11826 (
            .O(N__49134),
            .I(DMA_dev1_Teoc_1));
    IoInMux I__11825 (
            .O(N__49129),
            .I(N__49126));
    LocalMux I__11824 (
            .O(N__49126),
            .I(N__49123));
    Span4Mux_s3_v I__11823 (
            .O(N__49123),
            .I(N__49120));
    Span4Mux_h I__11822 (
            .O(N__49120),
            .I(N__49117));
    Span4Mux_v I__11821 (
            .O(N__49117),
            .I(N__49114));
    Odrv4 I__11820 (
            .O(N__49114),
            .I(N_265));
    InMux I__11819 (
            .O(N__49111),
            .I(N__49108));
    LocalMux I__11818 (
            .O(N__49108),
            .I(N__49105));
    Odrv12 I__11817 (
            .O(N__49105),
            .I(\u0.N_1729 ));
    InMux I__11816 (
            .O(N__49102),
            .I(N__49099));
    LocalMux I__11815 (
            .O(N__49099),
            .I(N__49096));
    Span4Mux_v I__11814 (
            .O(N__49096),
            .I(N__49093));
    Span4Mux_h I__11813 (
            .O(N__49093),
            .I(N__49090));
    Odrv4 I__11812 (
            .O(N__49090),
            .I(\u0.dat_o_i_0_0_18 ));
    CascadeMux I__11811 (
            .O(N__49087),
            .I(N__49084));
    InMux I__11810 (
            .O(N__49084),
            .I(N__49081));
    LocalMux I__11809 (
            .O(N__49081),
            .I(N__49078));
    Odrv12 I__11808 (
            .O(N__49078),
            .I(\u0.dat_o_i_0_2_18 ));
    IoInMux I__11807 (
            .O(N__49075),
            .I(N__49072));
    LocalMux I__11806 (
            .O(N__49072),
            .I(N__49069));
    IoSpan4Mux I__11805 (
            .O(N__49069),
            .I(N__49066));
    Span4Mux_s3_h I__11804 (
            .O(N__49066),
            .I(N__49063));
    Span4Mux_h I__11803 (
            .O(N__49063),
            .I(N__49060));
    Span4Mux_h I__11802 (
            .O(N__49060),
            .I(N__49057));
    Odrv4 I__11801 (
            .O(N__49057),
            .I(N_325_i));
    CascadeMux I__11800 (
            .O(N__49054),
            .I(N__49051));
    InMux I__11799 (
            .O(N__49051),
            .I(N__49048));
    LocalMux I__11798 (
            .O(N__49048),
            .I(N__49045));
    Odrv4 I__11797 (
            .O(N__49045),
            .I(iQ_RNIUKDM1_2));
    InMux I__11796 (
            .O(N__49042),
            .I(N__49039));
    LocalMux I__11795 (
            .O(N__49039),
            .I(N__49036));
    Span12Mux_h I__11794 (
            .O(N__49036),
            .I(N__49033));
    Odrv12 I__11793 (
            .O(N__49033),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIAH7KZ0Z_17 ));
    InMux I__11792 (
            .O(N__49030),
            .I(N__49027));
    LocalMux I__11791 (
            .O(N__49027),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI6TUQZ0Z_17 ));
    InMux I__11790 (
            .O(N__49024),
            .I(N__49021));
    LocalMux I__11789 (
            .O(N__49021),
            .I(N__49018));
    Span4Mux_v I__11788 (
            .O(N__49018),
            .I(N__49015));
    Span4Mux_h I__11787 (
            .O(N__49015),
            .I(N__49012));
    Span4Mux_h I__11786 (
            .O(N__49012),
            .I(N__49009));
    Odrv4 I__11785 (
            .O(N__49009),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIE5GTZ0Z_17 ));
    InMux I__11784 (
            .O(N__49006),
            .I(N__49003));
    LocalMux I__11783 (
            .O(N__49003),
            .I(N__49000));
    Odrv4 I__11782 (
            .O(N__49000),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_17 ));
    InMux I__11781 (
            .O(N__48997),
            .I(N__48994));
    LocalMux I__11780 (
            .O(N__48994),
            .I(iQ_RNI2PDM1_2));
    CascadeMux I__11779 (
            .O(N__48991),
            .I(mem_mem_ram6__RNIG5B71_17_cascade_));
    InMux I__11778 (
            .O(N__48988),
            .I(N__48982));
    InMux I__11777 (
            .O(N__48987),
            .I(N__48979));
    InMux I__11776 (
            .O(N__48986),
            .I(N__48976));
    InMux I__11775 (
            .O(N__48985),
            .I(N__48972));
    LocalMux I__11774 (
            .O(N__48982),
            .I(N__48964));
    LocalMux I__11773 (
            .O(N__48979),
            .I(N__48959));
    LocalMux I__11772 (
            .O(N__48976),
            .I(N__48959));
    InMux I__11771 (
            .O(N__48975),
            .I(N__48955));
    LocalMux I__11770 (
            .O(N__48972),
            .I(N__48952));
    InMux I__11769 (
            .O(N__48971),
            .I(N__48949));
    InMux I__11768 (
            .O(N__48970),
            .I(N__48946));
    InMux I__11767 (
            .O(N__48969),
            .I(N__48941));
    InMux I__11766 (
            .O(N__48968),
            .I(N__48934));
    InMux I__11765 (
            .O(N__48967),
            .I(N__48931));
    Span4Mux_v I__11764 (
            .O(N__48964),
            .I(N__48924));
    Span4Mux_h I__11763 (
            .O(N__48959),
            .I(N__48924));
    InMux I__11762 (
            .O(N__48958),
            .I(N__48921));
    LocalMux I__11761 (
            .O(N__48955),
            .I(N__48918));
    Span4Mux_h I__11760 (
            .O(N__48952),
            .I(N__48911));
    LocalMux I__11759 (
            .O(N__48949),
            .I(N__48911));
    LocalMux I__11758 (
            .O(N__48946),
            .I(N__48911));
    InMux I__11757 (
            .O(N__48945),
            .I(N__48907));
    InMux I__11756 (
            .O(N__48944),
            .I(N__48904));
    LocalMux I__11755 (
            .O(N__48941),
            .I(N__48901));
    InMux I__11754 (
            .O(N__48940),
            .I(N__48898));
    InMux I__11753 (
            .O(N__48939),
            .I(N__48895));
    CascadeMux I__11752 (
            .O(N__48938),
            .I(N__48892));
    InMux I__11751 (
            .O(N__48937),
            .I(N__48886));
    LocalMux I__11750 (
            .O(N__48934),
            .I(N__48883));
    LocalMux I__11749 (
            .O(N__48931),
            .I(N__48880));
    InMux I__11748 (
            .O(N__48930),
            .I(N__48877));
    InMux I__11747 (
            .O(N__48929),
            .I(N__48874));
    Span4Mux_v I__11746 (
            .O(N__48924),
            .I(N__48869));
    LocalMux I__11745 (
            .O(N__48921),
            .I(N__48869));
    Span4Mux_h I__11744 (
            .O(N__48918),
            .I(N__48865));
    Span4Mux_h I__11743 (
            .O(N__48911),
            .I(N__48862));
    InMux I__11742 (
            .O(N__48910),
            .I(N__48859));
    LocalMux I__11741 (
            .O(N__48907),
            .I(N__48851));
    LocalMux I__11740 (
            .O(N__48904),
            .I(N__48851));
    Span4Mux_h I__11739 (
            .O(N__48901),
            .I(N__48851));
    LocalMux I__11738 (
            .O(N__48898),
            .I(N__48846));
    LocalMux I__11737 (
            .O(N__48895),
            .I(N__48846));
    InMux I__11736 (
            .O(N__48892),
            .I(N__48843));
    InMux I__11735 (
            .O(N__48891),
            .I(N__48840));
    InMux I__11734 (
            .O(N__48890),
            .I(N__48837));
    InMux I__11733 (
            .O(N__48889),
            .I(N__48834));
    LocalMux I__11732 (
            .O(N__48886),
            .I(N__48826));
    Span4Mux_h I__11731 (
            .O(N__48883),
            .I(N__48817));
    Span4Mux_h I__11730 (
            .O(N__48880),
            .I(N__48817));
    LocalMux I__11729 (
            .O(N__48877),
            .I(N__48817));
    LocalMux I__11728 (
            .O(N__48874),
            .I(N__48817));
    Span4Mux_h I__11727 (
            .O(N__48869),
            .I(N__48814));
    InMux I__11726 (
            .O(N__48868),
            .I(N__48810));
    Span4Mux_v I__11725 (
            .O(N__48865),
            .I(N__48807));
    Span4Mux_v I__11724 (
            .O(N__48862),
            .I(N__48804));
    LocalMux I__11723 (
            .O(N__48859),
            .I(N__48801));
    InMux I__11722 (
            .O(N__48858),
            .I(N__48798));
    Span4Mux_v I__11721 (
            .O(N__48851),
            .I(N__48785));
    Span4Mux_h I__11720 (
            .O(N__48846),
            .I(N__48785));
    LocalMux I__11719 (
            .O(N__48843),
            .I(N__48785));
    LocalMux I__11718 (
            .O(N__48840),
            .I(N__48785));
    LocalMux I__11717 (
            .O(N__48837),
            .I(N__48785));
    LocalMux I__11716 (
            .O(N__48834),
            .I(N__48785));
    InMux I__11715 (
            .O(N__48833),
            .I(N__48782));
    InMux I__11714 (
            .O(N__48832),
            .I(N__48779));
    InMux I__11713 (
            .O(N__48831),
            .I(N__48776));
    InMux I__11712 (
            .O(N__48830),
            .I(N__48773));
    InMux I__11711 (
            .O(N__48829),
            .I(N__48770));
    Span4Mux_h I__11710 (
            .O(N__48826),
            .I(N__48763));
    Span4Mux_h I__11709 (
            .O(N__48817),
            .I(N__48763));
    Span4Mux_h I__11708 (
            .O(N__48814),
            .I(N__48760));
    InMux I__11707 (
            .O(N__48813),
            .I(N__48757));
    LocalMux I__11706 (
            .O(N__48810),
            .I(N__48754));
    Span4Mux_h I__11705 (
            .O(N__48807),
            .I(N__48745));
    Span4Mux_v I__11704 (
            .O(N__48804),
            .I(N__48745));
    Span4Mux_h I__11703 (
            .O(N__48801),
            .I(N__48745));
    LocalMux I__11702 (
            .O(N__48798),
            .I(N__48745));
    Span4Mux_v I__11701 (
            .O(N__48785),
            .I(N__48736));
    LocalMux I__11700 (
            .O(N__48782),
            .I(N__48736));
    LocalMux I__11699 (
            .O(N__48779),
            .I(N__48736));
    LocalMux I__11698 (
            .O(N__48776),
            .I(N__48736));
    LocalMux I__11697 (
            .O(N__48773),
            .I(N__48733));
    LocalMux I__11696 (
            .O(N__48770),
            .I(N__48730));
    InMux I__11695 (
            .O(N__48769),
            .I(N__48725));
    InMux I__11694 (
            .O(N__48768),
            .I(N__48725));
    Span4Mux_h I__11693 (
            .O(N__48763),
            .I(N__48722));
    Span4Mux_h I__11692 (
            .O(N__48760),
            .I(N__48719));
    LocalMux I__11691 (
            .O(N__48757),
            .I(N__48716));
    Span4Mux_h I__11690 (
            .O(N__48754),
            .I(N__48713));
    Span4Mux_h I__11689 (
            .O(N__48745),
            .I(N__48710));
    Span4Mux_h I__11688 (
            .O(N__48736),
            .I(N__48702));
    Span4Mux_v I__11687 (
            .O(N__48733),
            .I(N__48695));
    Span4Mux_h I__11686 (
            .O(N__48730),
            .I(N__48695));
    LocalMux I__11685 (
            .O(N__48725),
            .I(N__48695));
    Sp12to4 I__11684 (
            .O(N__48722),
            .I(N__48688));
    Sp12to4 I__11683 (
            .O(N__48719),
            .I(N__48688));
    Span12Mux_s4_v I__11682 (
            .O(N__48716),
            .I(N__48688));
    Span4Mux_v I__11681 (
            .O(N__48713),
            .I(N__48683));
    Span4Mux_v I__11680 (
            .O(N__48710),
            .I(N__48683));
    InMux I__11679 (
            .O(N__48709),
            .I(N__48678));
    InMux I__11678 (
            .O(N__48708),
            .I(N__48678));
    InMux I__11677 (
            .O(N__48707),
            .I(N__48671));
    InMux I__11676 (
            .O(N__48706),
            .I(N__48671));
    InMux I__11675 (
            .O(N__48705),
            .I(N__48671));
    Span4Mux_v I__11674 (
            .O(N__48702),
            .I(N__48666));
    Span4Mux_v I__11673 (
            .O(N__48695),
            .I(N__48666));
    Odrv12 I__11672 (
            .O(N__48688),
            .I(u1_DMA_control_gen_DMAbuf_Rxbuf_rd_ptr_2));
    Odrv4 I__11671 (
            .O(N__48683),
            .I(u1_DMA_control_gen_DMAbuf_Rxbuf_rd_ptr_2));
    LocalMux I__11670 (
            .O(N__48678),
            .I(u1_DMA_control_gen_DMAbuf_Rxbuf_rd_ptr_2));
    LocalMux I__11669 (
            .O(N__48671),
            .I(u1_DMA_control_gen_DMAbuf_Rxbuf_rd_ptr_2));
    Odrv4 I__11668 (
            .O(N__48666),
            .I(u1_DMA_control_gen_DMAbuf_Rxbuf_rd_ptr_2));
    InMux I__11667 (
            .O(N__48655),
            .I(N__48652));
    LocalMux I__11666 (
            .O(N__48652),
            .I(\u0.N_1549 ));
    InMux I__11665 (
            .O(N__48649),
            .I(N__48646));
    LocalMux I__11664 (
            .O(N__48646),
            .I(N__48643));
    Span4Mux_v I__11663 (
            .O(N__48643),
            .I(N__48640));
    Span4Mux_v I__11662 (
            .O(N__48640),
            .I(N__48637));
    Odrv4 I__11661 (
            .O(N__48637),
            .I(\u0.dat_o_0_a2_i_0_16 ));
    CascadeMux I__11660 (
            .O(N__48634),
            .I(N__48631));
    InMux I__11659 (
            .O(N__48631),
            .I(N__48628));
    LocalMux I__11658 (
            .O(N__48628),
            .I(N__48625));
    Span4Mux_v I__11657 (
            .O(N__48625),
            .I(N__48622));
    Odrv4 I__11656 (
            .O(N__48622),
            .I(\u0.dat_o_0_a2_i_2_16 ));
    IoInMux I__11655 (
            .O(N__48619),
            .I(N__48616));
    LocalMux I__11654 (
            .O(N__48616),
            .I(N__48613));
    Span12Mux_s5_v I__11653 (
            .O(N__48613),
            .I(N__48610));
    Span12Mux_h I__11652 (
            .O(N__48610),
            .I(N__48607));
    Odrv12 I__11651 (
            .O(N__48607),
            .I(N_207_i));
    InMux I__11650 (
            .O(N__48604),
            .I(N__48601));
    LocalMux I__11649 (
            .O(N__48601),
            .I(N__48594));
    InMux I__11648 (
            .O(N__48600),
            .I(N__48591));
    InMux I__11647 (
            .O(N__48599),
            .I(N__48588));
    InMux I__11646 (
            .O(N__48598),
            .I(N__48584));
    CascadeMux I__11645 (
            .O(N__48597),
            .I(N__48579));
    Span4Mux_v I__11644 (
            .O(N__48594),
            .I(N__48574));
    LocalMux I__11643 (
            .O(N__48591),
            .I(N__48571));
    LocalMux I__11642 (
            .O(N__48588),
            .I(N__48567));
    CascadeMux I__11641 (
            .O(N__48587),
            .I(N__48562));
    LocalMux I__11640 (
            .O(N__48584),
            .I(N__48559));
    InMux I__11639 (
            .O(N__48583),
            .I(N__48556));
    InMux I__11638 (
            .O(N__48582),
            .I(N__48553));
    InMux I__11637 (
            .O(N__48579),
            .I(N__48550));
    InMux I__11636 (
            .O(N__48578),
            .I(N__48545));
    CascadeMux I__11635 (
            .O(N__48577),
            .I(N__48541));
    Span4Mux_h I__11634 (
            .O(N__48574),
            .I(N__48535));
    Span4Mux_v I__11633 (
            .O(N__48571),
            .I(N__48535));
    InMux I__11632 (
            .O(N__48570),
            .I(N__48532));
    Span4Mux_v I__11631 (
            .O(N__48567),
            .I(N__48528));
    InMux I__11630 (
            .O(N__48566),
            .I(N__48525));
    InMux I__11629 (
            .O(N__48565),
            .I(N__48522));
    InMux I__11628 (
            .O(N__48562),
            .I(N__48518));
    Span4Mux_v I__11627 (
            .O(N__48559),
            .I(N__48515));
    LocalMux I__11626 (
            .O(N__48556),
            .I(N__48512));
    LocalMux I__11625 (
            .O(N__48553),
            .I(N__48507));
    LocalMux I__11624 (
            .O(N__48550),
            .I(N__48507));
    InMux I__11623 (
            .O(N__48549),
            .I(N__48504));
    CascadeMux I__11622 (
            .O(N__48548),
            .I(N__48501));
    LocalMux I__11621 (
            .O(N__48545),
            .I(N__48498));
    InMux I__11620 (
            .O(N__48544),
            .I(N__48495));
    InMux I__11619 (
            .O(N__48541),
            .I(N__48492));
    InMux I__11618 (
            .O(N__48540),
            .I(N__48489));
    Span4Mux_h I__11617 (
            .O(N__48535),
            .I(N__48484));
    LocalMux I__11616 (
            .O(N__48532),
            .I(N__48484));
    InMux I__11615 (
            .O(N__48531),
            .I(N__48481));
    Sp12to4 I__11614 (
            .O(N__48528),
            .I(N__48473));
    LocalMux I__11613 (
            .O(N__48525),
            .I(N__48473));
    LocalMux I__11612 (
            .O(N__48522),
            .I(N__48473));
    InMux I__11611 (
            .O(N__48521),
            .I(N__48470));
    LocalMux I__11610 (
            .O(N__48518),
            .I(N__48465));
    Span4Mux_h I__11609 (
            .O(N__48515),
            .I(N__48456));
    Span4Mux_h I__11608 (
            .O(N__48512),
            .I(N__48456));
    Span4Mux_v I__11607 (
            .O(N__48507),
            .I(N__48456));
    LocalMux I__11606 (
            .O(N__48504),
            .I(N__48456));
    InMux I__11605 (
            .O(N__48501),
            .I(N__48453));
    Span4Mux_v I__11604 (
            .O(N__48498),
            .I(N__48440));
    LocalMux I__11603 (
            .O(N__48495),
            .I(N__48440));
    LocalMux I__11602 (
            .O(N__48492),
            .I(N__48440));
    LocalMux I__11601 (
            .O(N__48489),
            .I(N__48440));
    Span4Mux_v I__11600 (
            .O(N__48484),
            .I(N__48440));
    LocalMux I__11599 (
            .O(N__48481),
            .I(N__48440));
    InMux I__11598 (
            .O(N__48480),
            .I(N__48437));
    Span12Mux_h I__11597 (
            .O(N__48473),
            .I(N__48433));
    LocalMux I__11596 (
            .O(N__48470),
            .I(N__48430));
    InMux I__11595 (
            .O(N__48469),
            .I(N__48427));
    InMux I__11594 (
            .O(N__48468),
            .I(N__48424));
    Span4Mux_v I__11593 (
            .O(N__48465),
            .I(N__48417));
    Span4Mux_h I__11592 (
            .O(N__48456),
            .I(N__48417));
    LocalMux I__11591 (
            .O(N__48453),
            .I(N__48417));
    Span4Mux_v I__11590 (
            .O(N__48440),
            .I(N__48412));
    LocalMux I__11589 (
            .O(N__48437),
            .I(N__48412));
    InMux I__11588 (
            .O(N__48436),
            .I(N__48409));
    Odrv12 I__11587 (
            .O(N__48433),
            .I(\u0.N_2128 ));
    Odrv12 I__11586 (
            .O(N__48430),
            .I(\u0.N_2128 ));
    LocalMux I__11585 (
            .O(N__48427),
            .I(\u0.N_2128 ));
    LocalMux I__11584 (
            .O(N__48424),
            .I(\u0.N_2128 ));
    Odrv4 I__11583 (
            .O(N__48417),
            .I(\u0.N_2128 ));
    Odrv4 I__11582 (
            .O(N__48412),
            .I(\u0.N_2128 ));
    LocalMux I__11581 (
            .O(N__48409),
            .I(\u0.N_2128 ));
    InMux I__11580 (
            .O(N__48394),
            .I(N__48391));
    LocalMux I__11579 (
            .O(N__48391),
            .I(N__48388));
    Sp12to4 I__11578 (
            .O(N__48388),
            .I(N__48385));
    Span12Mux_v I__11577 (
            .O(N__48385),
            .I(N__48381));
    InMux I__11576 (
            .O(N__48384),
            .I(N__48378));
    Span12Mux_h I__11575 (
            .O(N__48381),
            .I(N__48375));
    LocalMux I__11574 (
            .O(N__48378),
            .I(N__48372));
    Odrv12 I__11573 (
            .O(N__48375),
            .I(DMA_dev0_Td_1));
    Odrv4 I__11572 (
            .O(N__48372),
            .I(DMA_dev0_Td_1));
    InMux I__11571 (
            .O(N__48367),
            .I(N__48364));
    LocalMux I__11570 (
            .O(N__48364),
            .I(\u0.dat_o_0_0_2_9 ));
    InMux I__11569 (
            .O(N__48361),
            .I(N__48358));
    LocalMux I__11568 (
            .O(N__48358),
            .I(N__48355));
    Span4Mux_v I__11567 (
            .O(N__48355),
            .I(N__48352));
    Span4Mux_v I__11566 (
            .O(N__48352),
            .I(N__48349));
    Odrv4 I__11565 (
            .O(N__48349),
            .I(\u0.dat_o_0_0_6_9 ));
    CascadeMux I__11564 (
            .O(N__48346),
            .I(\u0.N_1651_cascade_ ));
    InMux I__11563 (
            .O(N__48343),
            .I(N__48340));
    LocalMux I__11562 (
            .O(N__48340),
            .I(\u0.N_1650 ));
    InMux I__11561 (
            .O(N__48337),
            .I(N__48334));
    LocalMux I__11560 (
            .O(N__48334),
            .I(N__48321));
    InMux I__11559 (
            .O(N__48333),
            .I(N__48318));
    CascadeMux I__11558 (
            .O(N__48332),
            .I(N__48315));
    InMux I__11557 (
            .O(N__48331),
            .I(N__48312));
    CascadeMux I__11556 (
            .O(N__48330),
            .I(N__48308));
    InMux I__11555 (
            .O(N__48329),
            .I(N__48305));
    InMux I__11554 (
            .O(N__48328),
            .I(N__48302));
    InMux I__11553 (
            .O(N__48327),
            .I(N__48299));
    CascadeMux I__11552 (
            .O(N__48326),
            .I(N__48296));
    InMux I__11551 (
            .O(N__48325),
            .I(N__48293));
    CascadeMux I__11550 (
            .O(N__48324),
            .I(N__48290));
    Span4Mux_v I__11549 (
            .O(N__48321),
            .I(N__48284));
    LocalMux I__11548 (
            .O(N__48318),
            .I(N__48284));
    InMux I__11547 (
            .O(N__48315),
            .I(N__48280));
    LocalMux I__11546 (
            .O(N__48312),
            .I(N__48272));
    InMux I__11545 (
            .O(N__48311),
            .I(N__48269));
    InMux I__11544 (
            .O(N__48308),
            .I(N__48266));
    LocalMux I__11543 (
            .O(N__48305),
            .I(N__48263));
    LocalMux I__11542 (
            .O(N__48302),
            .I(N__48258));
    LocalMux I__11541 (
            .O(N__48299),
            .I(N__48258));
    InMux I__11540 (
            .O(N__48296),
            .I(N__48255));
    LocalMux I__11539 (
            .O(N__48293),
            .I(N__48250));
    InMux I__11538 (
            .O(N__48290),
            .I(N__48247));
    InMux I__11537 (
            .O(N__48289),
            .I(N__48244));
    Span4Mux_v I__11536 (
            .O(N__48284),
            .I(N__48241));
    InMux I__11535 (
            .O(N__48283),
            .I(N__48238));
    LocalMux I__11534 (
            .O(N__48280),
            .I(N__48234));
    InMux I__11533 (
            .O(N__48279),
            .I(N__48223));
    InMux I__11532 (
            .O(N__48278),
            .I(N__48223));
    InMux I__11531 (
            .O(N__48277),
            .I(N__48223));
    InMux I__11530 (
            .O(N__48276),
            .I(N__48223));
    InMux I__11529 (
            .O(N__48275),
            .I(N__48223));
    Span4Mux_v I__11528 (
            .O(N__48272),
            .I(N__48218));
    LocalMux I__11527 (
            .O(N__48269),
            .I(N__48218));
    LocalMux I__11526 (
            .O(N__48266),
            .I(N__48215));
    Span4Mux_h I__11525 (
            .O(N__48263),
            .I(N__48208));
    Span4Mux_v I__11524 (
            .O(N__48258),
            .I(N__48208));
    LocalMux I__11523 (
            .O(N__48255),
            .I(N__48208));
    CascadeMux I__11522 (
            .O(N__48254),
            .I(N__48205));
    InMux I__11521 (
            .O(N__48253),
            .I(N__48202));
    Span4Mux_h I__11520 (
            .O(N__48250),
            .I(N__48197));
    LocalMux I__11519 (
            .O(N__48247),
            .I(N__48197));
    LocalMux I__11518 (
            .O(N__48244),
            .I(N__48194));
    Span4Mux_h I__11517 (
            .O(N__48241),
            .I(N__48189));
    LocalMux I__11516 (
            .O(N__48238),
            .I(N__48189));
    InMux I__11515 (
            .O(N__48237),
            .I(N__48186));
    Span12Mux_s10_h I__11514 (
            .O(N__48234),
            .I(N__48181));
    LocalMux I__11513 (
            .O(N__48223),
            .I(N__48181));
    Span4Mux_v I__11512 (
            .O(N__48218),
            .I(N__48176));
    Span4Mux_v I__11511 (
            .O(N__48215),
            .I(N__48176));
    Span4Mux_h I__11510 (
            .O(N__48208),
            .I(N__48173));
    InMux I__11509 (
            .O(N__48205),
            .I(N__48170));
    LocalMux I__11508 (
            .O(N__48202),
            .I(N__48167));
    Span4Mux_v I__11507 (
            .O(N__48197),
            .I(N__48158));
    Span4Mux_h I__11506 (
            .O(N__48194),
            .I(N__48158));
    Span4Mux_h I__11505 (
            .O(N__48189),
            .I(N__48158));
    LocalMux I__11504 (
            .O(N__48186),
            .I(N__48158));
    Odrv12 I__11503 (
            .O(N__48181),
            .I(\u0.N_2130 ));
    Odrv4 I__11502 (
            .O(N__48176),
            .I(\u0.N_2130 ));
    Odrv4 I__11501 (
            .O(N__48173),
            .I(\u0.N_2130 ));
    LocalMux I__11500 (
            .O(N__48170),
            .I(\u0.N_2130 ));
    Odrv4 I__11499 (
            .O(N__48167),
            .I(\u0.N_2130 ));
    Odrv4 I__11498 (
            .O(N__48158),
            .I(\u0.N_2130 ));
    InMux I__11497 (
            .O(N__48145),
            .I(N__48141));
    InMux I__11496 (
            .O(N__48144),
            .I(N__48138));
    LocalMux I__11495 (
            .O(N__48141),
            .I(N__48135));
    LocalMux I__11494 (
            .O(N__48138),
            .I(N__48129));
    Span4Mux_v I__11493 (
            .O(N__48135),
            .I(N__48121));
    InMux I__11492 (
            .O(N__48134),
            .I(N__48115));
    InMux I__11491 (
            .O(N__48133),
            .I(N__48115));
    CascadeMux I__11490 (
            .O(N__48132),
            .I(N__48107));
    Span4Mux_h I__11489 (
            .O(N__48129),
            .I(N__48103));
    InMux I__11488 (
            .O(N__48128),
            .I(N__48092));
    InMux I__11487 (
            .O(N__48127),
            .I(N__48092));
    InMux I__11486 (
            .O(N__48126),
            .I(N__48092));
    InMux I__11485 (
            .O(N__48125),
            .I(N__48092));
    InMux I__11484 (
            .O(N__48124),
            .I(N__48092));
    Sp12to4 I__11483 (
            .O(N__48121),
            .I(N__48089));
    InMux I__11482 (
            .O(N__48120),
            .I(N__48086));
    LocalMux I__11481 (
            .O(N__48115),
            .I(N__48082));
    InMux I__11480 (
            .O(N__48114),
            .I(N__48075));
    InMux I__11479 (
            .O(N__48113),
            .I(N__48075));
    InMux I__11478 (
            .O(N__48112),
            .I(N__48075));
    InMux I__11477 (
            .O(N__48111),
            .I(N__48072));
    InMux I__11476 (
            .O(N__48110),
            .I(N__48069));
    InMux I__11475 (
            .O(N__48107),
            .I(N__48066));
    CascadeMux I__11474 (
            .O(N__48106),
            .I(N__48062));
    Span4Mux_h I__11473 (
            .O(N__48103),
            .I(N__48055));
    LocalMux I__11472 (
            .O(N__48092),
            .I(N__48055));
    Span12Mux_s4_h I__11471 (
            .O(N__48089),
            .I(N__48050));
    LocalMux I__11470 (
            .O(N__48086),
            .I(N__48050));
    InMux I__11469 (
            .O(N__48085),
            .I(N__48047));
    Span4Mux_v I__11468 (
            .O(N__48082),
            .I(N__48042));
    LocalMux I__11467 (
            .O(N__48075),
            .I(N__48042));
    LocalMux I__11466 (
            .O(N__48072),
            .I(N__48037));
    LocalMux I__11465 (
            .O(N__48069),
            .I(N__48037));
    LocalMux I__11464 (
            .O(N__48066),
            .I(N__48034));
    InMux I__11463 (
            .O(N__48065),
            .I(N__48031));
    InMux I__11462 (
            .O(N__48062),
            .I(N__48028));
    CascadeMux I__11461 (
            .O(N__48061),
            .I(N__48024));
    CascadeMux I__11460 (
            .O(N__48060),
            .I(N__48021));
    Span4Mux_h I__11459 (
            .O(N__48055),
            .I(N__48015));
    Span12Mux_h I__11458 (
            .O(N__48050),
            .I(N__48010));
    LocalMux I__11457 (
            .O(N__48047),
            .I(N__48010));
    Span4Mux_h I__11456 (
            .O(N__48042),
            .I(N__48003));
    Span4Mux_h I__11455 (
            .O(N__48037),
            .I(N__48003));
    Span4Mux_h I__11454 (
            .O(N__48034),
            .I(N__48003));
    LocalMux I__11453 (
            .O(N__48031),
            .I(N__47998));
    LocalMux I__11452 (
            .O(N__48028),
            .I(N__47998));
    InMux I__11451 (
            .O(N__48027),
            .I(N__47995));
    InMux I__11450 (
            .O(N__48024),
            .I(N__47992));
    InMux I__11449 (
            .O(N__48021),
            .I(N__47989));
    InMux I__11448 (
            .O(N__48020),
            .I(N__47984));
    InMux I__11447 (
            .O(N__48019),
            .I(N__47984));
    InMux I__11446 (
            .O(N__48018),
            .I(N__47981));
    Odrv4 I__11445 (
            .O(N__48015),
            .I(\u0.N_2123 ));
    Odrv12 I__11444 (
            .O(N__48010),
            .I(\u0.N_2123 ));
    Odrv4 I__11443 (
            .O(N__48003),
            .I(\u0.N_2123 ));
    Odrv4 I__11442 (
            .O(N__47998),
            .I(\u0.N_2123 ));
    LocalMux I__11441 (
            .O(N__47995),
            .I(\u0.N_2123 ));
    LocalMux I__11440 (
            .O(N__47992),
            .I(\u0.N_2123 ));
    LocalMux I__11439 (
            .O(N__47989),
            .I(\u0.N_2123 ));
    LocalMux I__11438 (
            .O(N__47984),
            .I(\u0.N_2123 ));
    LocalMux I__11437 (
            .O(N__47981),
            .I(\u0.N_2123 ));
    InMux I__11436 (
            .O(N__47962),
            .I(N__47959));
    LocalMux I__11435 (
            .O(N__47959),
            .I(N__47956));
    Span4Mux_v I__11434 (
            .O(N__47956),
            .I(N__47952));
    InMux I__11433 (
            .O(N__47955),
            .I(N__47949));
    Span4Mux_h I__11432 (
            .O(N__47952),
            .I(N__47946));
    LocalMux I__11431 (
            .O(N__47949),
            .I(N__47943));
    Odrv4 I__11430 (
            .O(N__47946),
            .I(PIO_cmdport_Teoc_6));
    Odrv12 I__11429 (
            .O(N__47943),
            .I(PIO_cmdport_Teoc_6));
    InMux I__11428 (
            .O(N__47938),
            .I(N__47935));
    LocalMux I__11427 (
            .O(N__47935),
            .I(\u0.dat_o_i_i_1_30 ));
    InMux I__11426 (
            .O(N__47932),
            .I(N__47929));
    LocalMux I__11425 (
            .O(N__47929),
            .I(N__47926));
    Span4Mux_v I__11424 (
            .O(N__47926),
            .I(N__47923));
    Sp12to4 I__11423 (
            .O(N__47923),
            .I(N__47920));
    Span12Mux_h I__11422 (
            .O(N__47920),
            .I(N__47916));
    InMux I__11421 (
            .O(N__47919),
            .I(N__47913));
    Odrv12 I__11420 (
            .O(N__47916),
            .I(DMA_dev0_Teoc_6));
    LocalMux I__11419 (
            .O(N__47913),
            .I(DMA_dev0_Teoc_6));
    InMux I__11418 (
            .O(N__47908),
            .I(N__47905));
    LocalMux I__11417 (
            .O(N__47905),
            .I(N__47902));
    Span12Mux_v I__11416 (
            .O(N__47902),
            .I(N__47899));
    Odrv12 I__11415 (
            .O(N__47899),
            .I(DMAq_30));
    InMux I__11414 (
            .O(N__47896),
            .I(N__47893));
    LocalMux I__11413 (
            .O(N__47893),
            .I(N__47890));
    Odrv4 I__11412 (
            .O(N__47890),
            .I(\u0.dat_o_i_i_4_30 ));
    CascadeMux I__11411 (
            .O(N__47887),
            .I(\u0.dat_o_i_i_0_30_cascade_ ));
    InMux I__11410 (
            .O(N__47884),
            .I(N__47880));
    InMux I__11409 (
            .O(N__47883),
            .I(N__47877));
    LocalMux I__11408 (
            .O(N__47880),
            .I(N__47874));
    LocalMux I__11407 (
            .O(N__47877),
            .I(N__47871));
    Sp12to4 I__11406 (
            .O(N__47874),
            .I(N__47868));
    Span4Mux_v I__11405 (
            .O(N__47871),
            .I(N__47865));
    Span12Mux_s7_h I__11404 (
            .O(N__47868),
            .I(N__47862));
    Odrv4 I__11403 (
            .O(N__47865),
            .I(DMA_dev1_Teoc_6));
    Odrv12 I__11402 (
            .O(N__47862),
            .I(DMA_dev1_Teoc_6));
    IoInMux I__11401 (
            .O(N__47857),
            .I(N__47854));
    LocalMux I__11400 (
            .O(N__47854),
            .I(N__47851));
    Span4Mux_s2_v I__11399 (
            .O(N__47851),
            .I(N__47848));
    Span4Mux_h I__11398 (
            .O(N__47848),
            .I(N__47845));
    Span4Mux_v I__11397 (
            .O(N__47845),
            .I(N__47842));
    Odrv4 I__11396 (
            .O(N__47842),
            .I(N_275));
    InMux I__11395 (
            .O(N__47839),
            .I(N__47835));
    InMux I__11394 (
            .O(N__47838),
            .I(N__47832));
    LocalMux I__11393 (
            .O(N__47835),
            .I(N__47826));
    LocalMux I__11392 (
            .O(N__47832),
            .I(N__47826));
    InMux I__11391 (
            .O(N__47831),
            .I(N__47823));
    Span4Mux_h I__11390 (
            .O(N__47826),
            .I(N__47816));
    LocalMux I__11389 (
            .O(N__47823),
            .I(N__47816));
    InMux I__11388 (
            .O(N__47822),
            .I(N__47813));
    InMux I__11387 (
            .O(N__47821),
            .I(N__47810));
    Span4Mux_v I__11386 (
            .O(N__47816),
            .I(N__47807));
    LocalMux I__11385 (
            .O(N__47813),
            .I(N__47804));
    LocalMux I__11384 (
            .O(N__47810),
            .I(N__47801));
    Span4Mux_v I__11383 (
            .O(N__47807),
            .I(N__47796));
    Span4Mux_v I__11382 (
            .O(N__47804),
            .I(N__47796));
    Span4Mux_v I__11381 (
            .O(N__47801),
            .I(N__47791));
    Span4Mux_h I__11380 (
            .O(N__47796),
            .I(N__47788));
    InMux I__11379 (
            .O(N__47795),
            .I(N__47785));
    InMux I__11378 (
            .O(N__47794),
            .I(N__47782));
    Sp12to4 I__11377 (
            .O(N__47791),
            .I(N__47779));
    Span4Mux_h I__11376 (
            .O(N__47788),
            .I(N__47776));
    LocalMux I__11375 (
            .O(N__47785),
            .I(N__47773));
    LocalMux I__11374 (
            .O(N__47782),
            .I(N__47770));
    Span12Mux_h I__11373 (
            .O(N__47779),
            .I(N__47767));
    Span4Mux_h I__11372 (
            .O(N__47776),
            .I(N__47762));
    Span4Mux_v I__11371 (
            .O(N__47773),
            .I(N__47762));
    Span4Mux_v I__11370 (
            .O(N__47770),
            .I(N__47759));
    Odrv12 I__11369 (
            .O(N__47767),
            .I(wb_dat_i_c_30));
    Odrv4 I__11368 (
            .O(N__47762),
            .I(wb_dat_i_c_30));
    Odrv4 I__11367 (
            .O(N__47759),
            .I(wb_dat_i_c_30));
    InMux I__11366 (
            .O(N__47752),
            .I(N__47749));
    LocalMux I__11365 (
            .O(N__47749),
            .I(\u0.CtrlRegZ0Z_30 ));
    InMux I__11364 (
            .O(N__47746),
            .I(N__47743));
    LocalMux I__11363 (
            .O(N__47743),
            .I(N__47740));
    Odrv4 I__11362 (
            .O(N__47740),
            .I(\u0.dat_o_0_a2_i_o2_0Z0Z_16 ));
    InMux I__11361 (
            .O(N__47737),
            .I(N__47732));
    CascadeMux I__11360 (
            .O(N__47736),
            .I(N__47728));
    InMux I__11359 (
            .O(N__47735),
            .I(N__47724));
    LocalMux I__11358 (
            .O(N__47732),
            .I(N__47721));
    CascadeMux I__11357 (
            .O(N__47731),
            .I(N__47716));
    InMux I__11356 (
            .O(N__47728),
            .I(N__47712));
    InMux I__11355 (
            .O(N__47727),
            .I(N__47709));
    LocalMux I__11354 (
            .O(N__47724),
            .I(N__47697));
    Span4Mux_v I__11353 (
            .O(N__47721),
            .I(N__47694));
    InMux I__11352 (
            .O(N__47720),
            .I(N__47685));
    InMux I__11351 (
            .O(N__47719),
            .I(N__47685));
    InMux I__11350 (
            .O(N__47716),
            .I(N__47685));
    InMux I__11349 (
            .O(N__47715),
            .I(N__47685));
    LocalMux I__11348 (
            .O(N__47712),
            .I(N__47682));
    LocalMux I__11347 (
            .O(N__47709),
            .I(N__47679));
    InMux I__11346 (
            .O(N__47708),
            .I(N__47674));
    InMux I__11345 (
            .O(N__47707),
            .I(N__47674));
    InMux I__11344 (
            .O(N__47706),
            .I(N__47667));
    InMux I__11343 (
            .O(N__47705),
            .I(N__47667));
    InMux I__11342 (
            .O(N__47704),
            .I(N__47667));
    InMux I__11341 (
            .O(N__47703),
            .I(N__47660));
    InMux I__11340 (
            .O(N__47702),
            .I(N__47660));
    InMux I__11339 (
            .O(N__47701),
            .I(N__47660));
    InMux I__11338 (
            .O(N__47700),
            .I(N__47657));
    Span4Mux_h I__11337 (
            .O(N__47697),
            .I(N__47654));
    Span4Mux_h I__11336 (
            .O(N__47694),
            .I(N__47650));
    LocalMux I__11335 (
            .O(N__47685),
            .I(N__47647));
    Span4Mux_v I__11334 (
            .O(N__47682),
            .I(N__47644));
    Span4Mux_v I__11333 (
            .O(N__47679),
            .I(N__47635));
    LocalMux I__11332 (
            .O(N__47674),
            .I(N__47635));
    LocalMux I__11331 (
            .O(N__47667),
            .I(N__47635));
    LocalMux I__11330 (
            .O(N__47660),
            .I(N__47635));
    LocalMux I__11329 (
            .O(N__47657),
            .I(N__47631));
    Span4Mux_v I__11328 (
            .O(N__47654),
            .I(N__47628));
    InMux I__11327 (
            .O(N__47653),
            .I(N__47625));
    Span4Mux_h I__11326 (
            .O(N__47650),
            .I(N__47620));
    Span4Mux_v I__11325 (
            .O(N__47647),
            .I(N__47620));
    Span4Mux_h I__11324 (
            .O(N__47644),
            .I(N__47615));
    Span4Mux_v I__11323 (
            .O(N__47635),
            .I(N__47615));
    InMux I__11322 (
            .O(N__47634),
            .I(N__47612));
    Span12Mux_s11_h I__11321 (
            .O(N__47631),
            .I(N__47605));
    Sp12to4 I__11320 (
            .O(N__47628),
            .I(N__47605));
    LocalMux I__11319 (
            .O(N__47625),
            .I(N__47605));
    Sp12to4 I__11318 (
            .O(N__47620),
            .I(N__47598));
    Sp12to4 I__11317 (
            .O(N__47615),
            .I(N__47598));
    LocalMux I__11316 (
            .O(N__47612),
            .I(N__47598));
    Span12Mux_v I__11315 (
            .O(N__47605),
            .I(N__47595));
    Span12Mux_h I__11314 (
            .O(N__47598),
            .I(N__47592));
    Span12Mux_h I__11313 (
            .O(N__47595),
            .I(N__47589));
    Span12Mux_v I__11312 (
            .O(N__47592),
            .I(N__47586));
    Odrv12 I__11311 (
            .O(N__47589),
            .I(wb_adr_i_c_3));
    Odrv12 I__11310 (
            .O(N__47586),
            .I(wb_adr_i_c_3));
    InMux I__11309 (
            .O(N__47581),
            .I(N__47578));
    LocalMux I__11308 (
            .O(N__47578),
            .I(N__47575));
    Span4Mux_v I__11307 (
            .O(N__47575),
            .I(N__47572));
    Odrv4 I__11306 (
            .O(N__47572),
            .I(\u0.N_1714 ));
    InMux I__11305 (
            .O(N__47569),
            .I(N__47566));
    LocalMux I__11304 (
            .O(N__47566),
            .I(N__47563));
    Span4Mux_h I__11303 (
            .O(N__47563),
            .I(N__47560));
    Odrv4 I__11302 (
            .O(N__47560),
            .I(\u0.dat_o_i_0_0_23 ));
    CascadeMux I__11301 (
            .O(N__47557),
            .I(\u0.N_1374_cascade_ ));
    IoInMux I__11300 (
            .O(N__47554),
            .I(N__47551));
    LocalMux I__11299 (
            .O(N__47551),
            .I(N__47548));
    IoSpan4Mux I__11298 (
            .O(N__47548),
            .I(N__47545));
    Span4Mux_s3_h I__11297 (
            .O(N__47545),
            .I(N__47542));
    Span4Mux_h I__11296 (
            .O(N__47542),
            .I(N__47539));
    Span4Mux_h I__11295 (
            .O(N__47539),
            .I(N__47536));
    Odrv4 I__11294 (
            .O(N__47536),
            .I(N_332_i));
    InMux I__11293 (
            .O(N__47533),
            .I(N__47530));
    LocalMux I__11292 (
            .O(N__47530),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI6ONK1Z0Z_2 ));
    InMux I__11291 (
            .O(N__47527),
            .I(N__47524));
    LocalMux I__11290 (
            .O(N__47524),
            .I(N__47521));
    Odrv12 I__11289 (
            .O(N__47521),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIBAOD1Z0Z_1 ));
    CascadeMux I__11288 (
            .O(N__47518),
            .I(N__47513));
    InMux I__11287 (
            .O(N__47517),
            .I(N__47505));
    InMux I__11286 (
            .O(N__47516),
            .I(N__47505));
    InMux I__11285 (
            .O(N__47513),
            .I(N__47498));
    InMux I__11284 (
            .O(N__47512),
            .I(N__47498));
    InMux I__11283 (
            .O(N__47511),
            .I(N__47498));
    CascadeMux I__11282 (
            .O(N__47510),
            .I(N__47494));
    LocalMux I__11281 (
            .O(N__47505),
            .I(N__47488));
    LocalMux I__11280 (
            .O(N__47498),
            .I(N__47488));
    CascadeMux I__11279 (
            .O(N__47497),
            .I(N__47484));
    InMux I__11278 (
            .O(N__47494),
            .I(N__47478));
    InMux I__11277 (
            .O(N__47493),
            .I(N__47475));
    Span4Mux_v I__11276 (
            .O(N__47488),
            .I(N__47472));
    InMux I__11275 (
            .O(N__47487),
            .I(N__47469));
    InMux I__11274 (
            .O(N__47484),
            .I(N__47464));
    InMux I__11273 (
            .O(N__47483),
            .I(N__47461));
    InMux I__11272 (
            .O(N__47482),
            .I(N__47458));
    InMux I__11271 (
            .O(N__47481),
            .I(N__47455));
    LocalMux I__11270 (
            .O(N__47478),
            .I(N__47450));
    LocalMux I__11269 (
            .O(N__47475),
            .I(N__47447));
    Span4Mux_h I__11268 (
            .O(N__47472),
            .I(N__47442));
    LocalMux I__11267 (
            .O(N__47469),
            .I(N__47442));
    InMux I__11266 (
            .O(N__47468),
            .I(N__47439));
    InMux I__11265 (
            .O(N__47467),
            .I(N__47436));
    LocalMux I__11264 (
            .O(N__47464),
            .I(N__47432));
    LocalMux I__11263 (
            .O(N__47461),
            .I(N__47429));
    LocalMux I__11262 (
            .O(N__47458),
            .I(N__47424));
    LocalMux I__11261 (
            .O(N__47455),
            .I(N__47424));
    InMux I__11260 (
            .O(N__47454),
            .I(N__47420));
    CascadeMux I__11259 (
            .O(N__47453),
            .I(N__47417));
    Span4Mux_v I__11258 (
            .O(N__47450),
            .I(N__47411));
    Span4Mux_h I__11257 (
            .O(N__47447),
            .I(N__47411));
    Span4Mux_h I__11256 (
            .O(N__47442),
            .I(N__47406));
    LocalMux I__11255 (
            .O(N__47439),
            .I(N__47406));
    LocalMux I__11254 (
            .O(N__47436),
            .I(N__47402));
    InMux I__11253 (
            .O(N__47435),
            .I(N__47399));
    Span4Mux_v I__11252 (
            .O(N__47432),
            .I(N__47395));
    Span4Mux_v I__11251 (
            .O(N__47429),
            .I(N__47392));
    Span4Mux_v I__11250 (
            .O(N__47424),
            .I(N__47389));
    InMux I__11249 (
            .O(N__47423),
            .I(N__47386));
    LocalMux I__11248 (
            .O(N__47420),
            .I(N__47383));
    InMux I__11247 (
            .O(N__47417),
            .I(N__47380));
    CascadeMux I__11246 (
            .O(N__47416),
            .I(N__47377));
    Span4Mux_h I__11245 (
            .O(N__47411),
            .I(N__47370));
    Span4Mux_h I__11244 (
            .O(N__47406),
            .I(N__47367));
    InMux I__11243 (
            .O(N__47405),
            .I(N__47364));
    Span4Mux_v I__11242 (
            .O(N__47402),
            .I(N__47361));
    LocalMux I__11241 (
            .O(N__47399),
            .I(N__47358));
    InMux I__11240 (
            .O(N__47398),
            .I(N__47355));
    Span4Mux_v I__11239 (
            .O(N__47395),
            .I(N__47348));
    Span4Mux_v I__11238 (
            .O(N__47392),
            .I(N__47348));
    Span4Mux_h I__11237 (
            .O(N__47389),
            .I(N__47348));
    LocalMux I__11236 (
            .O(N__47386),
            .I(N__47345));
    Span4Mux_h I__11235 (
            .O(N__47383),
            .I(N__47340));
    LocalMux I__11234 (
            .O(N__47380),
            .I(N__47340));
    InMux I__11233 (
            .O(N__47377),
            .I(N__47335));
    InMux I__11232 (
            .O(N__47376),
            .I(N__47335));
    InMux I__11231 (
            .O(N__47375),
            .I(N__47332));
    InMux I__11230 (
            .O(N__47374),
            .I(N__47327));
    InMux I__11229 (
            .O(N__47373),
            .I(N__47327));
    Span4Mux_h I__11228 (
            .O(N__47370),
            .I(N__47320));
    Span4Mux_v I__11227 (
            .O(N__47367),
            .I(N__47320));
    LocalMux I__11226 (
            .O(N__47364),
            .I(N__47320));
    Sp12to4 I__11225 (
            .O(N__47361),
            .I(N__47313));
    Sp12to4 I__11224 (
            .O(N__47358),
            .I(N__47313));
    LocalMux I__11223 (
            .O(N__47355),
            .I(N__47313));
    Span4Mux_v I__11222 (
            .O(N__47348),
            .I(N__47310));
    Sp12to4 I__11221 (
            .O(N__47345),
            .I(N__47299));
    Sp12to4 I__11220 (
            .O(N__47340),
            .I(N__47299));
    LocalMux I__11219 (
            .O(N__47335),
            .I(N__47299));
    LocalMux I__11218 (
            .O(N__47332),
            .I(N__47299));
    LocalMux I__11217 (
            .O(N__47327),
            .I(N__47299));
    Span4Mux_v I__11216 (
            .O(N__47320),
            .I(N__47296));
    Span12Mux_v I__11215 (
            .O(N__47313),
            .I(N__47293));
    Sp12to4 I__11214 (
            .O(N__47310),
            .I(N__47290));
    Span12Mux_v I__11213 (
            .O(N__47299),
            .I(N__47285));
    Sp12to4 I__11212 (
            .O(N__47296),
            .I(N__47285));
    Span12Mux_v I__11211 (
            .O(N__47293),
            .I(N__47282));
    Span12Mux_h I__11210 (
            .O(N__47290),
            .I(N__47279));
    Span12Mux_v I__11209 (
            .O(N__47285),
            .I(N__47276));
    Span12Mux_h I__11208 (
            .O(N__47282),
            .I(N__47273));
    Span12Mux_v I__11207 (
            .O(N__47279),
            .I(N__47268));
    Span12Mux_h I__11206 (
            .O(N__47276),
            .I(N__47268));
    Odrv12 I__11205 (
            .O(N__47273),
            .I(wb_adr_i_c_6));
    Odrv12 I__11204 (
            .O(N__47268),
            .I(wb_adr_i_c_6));
    CascadeMux I__11203 (
            .O(N__47263),
            .I(N__47259));
    InMux I__11202 (
            .O(N__47262),
            .I(N__47256));
    InMux I__11201 (
            .O(N__47259),
            .I(N__47250));
    LocalMux I__11200 (
            .O(N__47256),
            .I(N__47246));
    InMux I__11199 (
            .O(N__47255),
            .I(N__47242));
    InMux I__11198 (
            .O(N__47254),
            .I(N__47239));
    InMux I__11197 (
            .O(N__47253),
            .I(N__47235));
    LocalMux I__11196 (
            .O(N__47250),
            .I(N__47232));
    InMux I__11195 (
            .O(N__47249),
            .I(N__47229));
    Span4Mux_h I__11194 (
            .O(N__47246),
            .I(N__47225));
    InMux I__11193 (
            .O(N__47245),
            .I(N__47221));
    LocalMux I__11192 (
            .O(N__47242),
            .I(N__47217));
    LocalMux I__11191 (
            .O(N__47239),
            .I(N__47214));
    CascadeMux I__11190 (
            .O(N__47238),
            .I(N__47210));
    LocalMux I__11189 (
            .O(N__47235),
            .I(N__47206));
    Span4Mux_v I__11188 (
            .O(N__47232),
            .I(N__47201));
    LocalMux I__11187 (
            .O(N__47229),
            .I(N__47201));
    InMux I__11186 (
            .O(N__47228),
            .I(N__47198));
    Span4Mux_h I__11185 (
            .O(N__47225),
            .I(N__47193));
    CascadeMux I__11184 (
            .O(N__47224),
            .I(N__47190));
    LocalMux I__11183 (
            .O(N__47221),
            .I(N__47187));
    InMux I__11182 (
            .O(N__47220),
            .I(N__47184));
    Span4Mux_v I__11181 (
            .O(N__47217),
            .I(N__47178));
    Span4Mux_s2_v I__11180 (
            .O(N__47214),
            .I(N__47175));
    InMux I__11179 (
            .O(N__47213),
            .I(N__47172));
    InMux I__11178 (
            .O(N__47210),
            .I(N__47169));
    CascadeMux I__11177 (
            .O(N__47209),
            .I(N__47164));
    Span4Mux_v I__11176 (
            .O(N__47206),
            .I(N__47157));
    Span4Mux_h I__11175 (
            .O(N__47201),
            .I(N__47157));
    LocalMux I__11174 (
            .O(N__47198),
            .I(N__47157));
    InMux I__11173 (
            .O(N__47197),
            .I(N__47152));
    InMux I__11172 (
            .O(N__47196),
            .I(N__47152));
    Span4Mux_h I__11171 (
            .O(N__47193),
            .I(N__47149));
    InMux I__11170 (
            .O(N__47190),
            .I(N__47146));
    Span4Mux_v I__11169 (
            .O(N__47187),
            .I(N__47139));
    LocalMux I__11168 (
            .O(N__47184),
            .I(N__47139));
    InMux I__11167 (
            .O(N__47183),
            .I(N__47136));
    InMux I__11166 (
            .O(N__47182),
            .I(N__47133));
    InMux I__11165 (
            .O(N__47181),
            .I(N__47130));
    Span4Mux_h I__11164 (
            .O(N__47178),
            .I(N__47121));
    Span4Mux_v I__11163 (
            .O(N__47175),
            .I(N__47121));
    LocalMux I__11162 (
            .O(N__47172),
            .I(N__47121));
    LocalMux I__11161 (
            .O(N__47169),
            .I(N__47121));
    InMux I__11160 (
            .O(N__47168),
            .I(N__47118));
    InMux I__11159 (
            .O(N__47167),
            .I(N__47115));
    InMux I__11158 (
            .O(N__47164),
            .I(N__47112));
    Span4Mux_h I__11157 (
            .O(N__47157),
            .I(N__47106));
    LocalMux I__11156 (
            .O(N__47152),
            .I(N__47106));
    Span4Mux_h I__11155 (
            .O(N__47149),
            .I(N__47101));
    LocalMux I__11154 (
            .O(N__47146),
            .I(N__47101));
    InMux I__11153 (
            .O(N__47145),
            .I(N__47098));
    InMux I__11152 (
            .O(N__47144),
            .I(N__47095));
    Span4Mux_h I__11151 (
            .O(N__47139),
            .I(N__47090));
    LocalMux I__11150 (
            .O(N__47136),
            .I(N__47090));
    LocalMux I__11149 (
            .O(N__47133),
            .I(N__47085));
    LocalMux I__11148 (
            .O(N__47130),
            .I(N__47085));
    Span4Mux_v I__11147 (
            .O(N__47121),
            .I(N__47078));
    LocalMux I__11146 (
            .O(N__47118),
            .I(N__47078));
    LocalMux I__11145 (
            .O(N__47115),
            .I(N__47078));
    LocalMux I__11144 (
            .O(N__47112),
            .I(N__47075));
    InMux I__11143 (
            .O(N__47111),
            .I(N__47072));
    Span4Mux_v I__11142 (
            .O(N__47106),
            .I(N__47061));
    Span4Mux_v I__11141 (
            .O(N__47101),
            .I(N__47061));
    LocalMux I__11140 (
            .O(N__47098),
            .I(N__47061));
    LocalMux I__11139 (
            .O(N__47095),
            .I(N__47061));
    Span4Mux_h I__11138 (
            .O(N__47090),
            .I(N__47050));
    Span4Mux_v I__11137 (
            .O(N__47085),
            .I(N__47050));
    Span4Mux_h I__11136 (
            .O(N__47078),
            .I(N__47050));
    Span4Mux_v I__11135 (
            .O(N__47075),
            .I(N__47050));
    LocalMux I__11134 (
            .O(N__47072),
            .I(N__47050));
    InMux I__11133 (
            .O(N__47071),
            .I(N__47047));
    InMux I__11132 (
            .O(N__47070),
            .I(N__47044));
    Odrv4 I__11131 (
            .O(N__47061),
            .I(N_2119));
    Odrv4 I__11130 (
            .O(N__47050),
            .I(N_2119));
    LocalMux I__11129 (
            .O(N__47047),
            .I(N_2119));
    LocalMux I__11128 (
            .O(N__47044),
            .I(N_2119));
    CascadeMux I__11127 (
            .O(N__47035),
            .I(DMAq_1_cascade_));
    InMux I__11126 (
            .O(N__47032),
            .I(N__47029));
    LocalMux I__11125 (
            .O(N__47029),
            .I(PIOq_1));
    InMux I__11124 (
            .O(N__47026),
            .I(N__47023));
    LocalMux I__11123 (
            .O(N__47023),
            .I(\u0.dat_o_0_0_1Z0Z_1 ));
    InMux I__11122 (
            .O(N__47020),
            .I(N__47017));
    LocalMux I__11121 (
            .O(N__47017),
            .I(N__47014));
    Span4Mux_v I__11120 (
            .O(N__47014),
            .I(N__47011));
    Span4Mux_h I__11119 (
            .O(N__47011),
            .I(N__47007));
    InMux I__11118 (
            .O(N__47010),
            .I(N__47004));
    Odrv4 I__11117 (
            .O(N__47007),
            .I(PIO_cmdport_Teoc_2));
    LocalMux I__11116 (
            .O(N__47004),
            .I(PIO_cmdport_Teoc_2));
    CascadeMux I__11115 (
            .O(N__46999),
            .I(\u0.N_2130_cascade_ ));
    InMux I__11114 (
            .O(N__46996),
            .I(N__46993));
    LocalMux I__11113 (
            .O(N__46993),
            .I(\u0.CtrlRegZ0Z_26 ));
    InMux I__11112 (
            .O(N__46990),
            .I(N__46987));
    LocalMux I__11111 (
            .O(N__46987),
            .I(\u0.dat_o_i_i_1_26 ));
    InMux I__11110 (
            .O(N__46984),
            .I(N__46980));
    InMux I__11109 (
            .O(N__46983),
            .I(N__46975));
    LocalMux I__11108 (
            .O(N__46980),
            .I(N__46972));
    InMux I__11107 (
            .O(N__46979),
            .I(N__46969));
    InMux I__11106 (
            .O(N__46978),
            .I(N__46966));
    LocalMux I__11105 (
            .O(N__46975),
            .I(N__46963));
    Span4Mux_h I__11104 (
            .O(N__46972),
            .I(N__46955));
    LocalMux I__11103 (
            .O(N__46969),
            .I(N__46955));
    LocalMux I__11102 (
            .O(N__46966),
            .I(N__46952));
    Span4Mux_v I__11101 (
            .O(N__46963),
            .I(N__46948));
    InMux I__11100 (
            .O(N__46962),
            .I(N__46941));
    InMux I__11099 (
            .O(N__46961),
            .I(N__46941));
    InMux I__11098 (
            .O(N__46960),
            .I(N__46941));
    Span4Mux_h I__11097 (
            .O(N__46955),
            .I(N__46931));
    Span4Mux_v I__11096 (
            .O(N__46952),
            .I(N__46931));
    InMux I__11095 (
            .O(N__46951),
            .I(N__46928));
    Span4Mux_h I__11094 (
            .O(N__46948),
            .I(N__46923));
    LocalMux I__11093 (
            .O(N__46941),
            .I(N__46923));
    InMux I__11092 (
            .O(N__46940),
            .I(N__46920));
    InMux I__11091 (
            .O(N__46939),
            .I(N__46917));
    InMux I__11090 (
            .O(N__46938),
            .I(N__46912));
    InMux I__11089 (
            .O(N__46937),
            .I(N__46912));
    InMux I__11088 (
            .O(N__46936),
            .I(N__46909));
    Span4Mux_h I__11087 (
            .O(N__46931),
            .I(N__46899));
    LocalMux I__11086 (
            .O(N__46928),
            .I(N__46899));
    Span4Mux_v I__11085 (
            .O(N__46923),
            .I(N__46894));
    LocalMux I__11084 (
            .O(N__46920),
            .I(N__46894));
    LocalMux I__11083 (
            .O(N__46917),
            .I(N__46891));
    LocalMux I__11082 (
            .O(N__46912),
            .I(N__46883));
    LocalMux I__11081 (
            .O(N__46909),
            .I(N__46883));
    InMux I__11080 (
            .O(N__46908),
            .I(N__46880));
    InMux I__11079 (
            .O(N__46907),
            .I(N__46877));
    InMux I__11078 (
            .O(N__46906),
            .I(N__46874));
    InMux I__11077 (
            .O(N__46905),
            .I(N__46871));
    InMux I__11076 (
            .O(N__46904),
            .I(N__46868));
    Span4Mux_v I__11075 (
            .O(N__46899),
            .I(N__46861));
    Span4Mux_v I__11074 (
            .O(N__46894),
            .I(N__46856));
    Span4Mux_v I__11073 (
            .O(N__46891),
            .I(N__46856));
    InMux I__11072 (
            .O(N__46890),
            .I(N__46853));
    InMux I__11071 (
            .O(N__46889),
            .I(N__46850));
    InMux I__11070 (
            .O(N__46888),
            .I(N__46847));
    Span12Mux_h I__11069 (
            .O(N__46883),
            .I(N__46840));
    LocalMux I__11068 (
            .O(N__46880),
            .I(N__46840));
    LocalMux I__11067 (
            .O(N__46877),
            .I(N__46840));
    LocalMux I__11066 (
            .O(N__46874),
            .I(N__46833));
    LocalMux I__11065 (
            .O(N__46871),
            .I(N__46833));
    LocalMux I__11064 (
            .O(N__46868),
            .I(N__46833));
    InMux I__11063 (
            .O(N__46867),
            .I(N__46830));
    InMux I__11062 (
            .O(N__46866),
            .I(N__46827));
    InMux I__11061 (
            .O(N__46865),
            .I(N__46824));
    InMux I__11060 (
            .O(N__46864),
            .I(N__46821));
    Odrv4 I__11059 (
            .O(N__46861),
            .I(\u0.N_2122 ));
    Odrv4 I__11058 (
            .O(N__46856),
            .I(\u0.N_2122 ));
    LocalMux I__11057 (
            .O(N__46853),
            .I(\u0.N_2122 ));
    LocalMux I__11056 (
            .O(N__46850),
            .I(\u0.N_2122 ));
    LocalMux I__11055 (
            .O(N__46847),
            .I(\u0.N_2122 ));
    Odrv12 I__11054 (
            .O(N__46840),
            .I(\u0.N_2122 ));
    Odrv4 I__11053 (
            .O(N__46833),
            .I(\u0.N_2122 ));
    LocalMux I__11052 (
            .O(N__46830),
            .I(\u0.N_2122 ));
    LocalMux I__11051 (
            .O(N__46827),
            .I(\u0.N_2122 ));
    LocalMux I__11050 (
            .O(N__46824),
            .I(\u0.N_2122 ));
    LocalMux I__11049 (
            .O(N__46821),
            .I(\u0.N_2122 ));
    InMux I__11048 (
            .O(N__46798),
            .I(N__46794));
    InMux I__11047 (
            .O(N__46797),
            .I(N__46791));
    LocalMux I__11046 (
            .O(N__46794),
            .I(N__46788));
    LocalMux I__11045 (
            .O(N__46791),
            .I(N__46785));
    Span4Mux_h I__11044 (
            .O(N__46788),
            .I(N__46782));
    Span4Mux_v I__11043 (
            .O(N__46785),
            .I(N__46779));
    Span4Mux_h I__11042 (
            .O(N__46782),
            .I(N__46776));
    Odrv4 I__11041 (
            .O(N__46779),
            .I(PIO_dport1_Teoc_6));
    Odrv4 I__11040 (
            .O(N__46776),
            .I(PIO_dport1_Teoc_6));
    InMux I__11039 (
            .O(N__46771),
            .I(N__46768));
    LocalMux I__11038 (
            .O(N__46768),
            .I(N__46764));
    InMux I__11037 (
            .O(N__46767),
            .I(N__46761));
    Span4Mux_v I__11036 (
            .O(N__46764),
            .I(N__46758));
    LocalMux I__11035 (
            .O(N__46761),
            .I(N__46755));
    Span4Mux_v I__11034 (
            .O(N__46758),
            .I(N__46752));
    Span12Mux_s10_h I__11033 (
            .O(N__46755),
            .I(N__46749));
    Odrv4 I__11032 (
            .O(N__46752),
            .I(PIO_dport0_Teoc_6));
    Odrv12 I__11031 (
            .O(N__46749),
            .I(PIO_dport0_Teoc_6));
    CascadeMux I__11030 (
            .O(N__46744),
            .I(\u0.N_1703_cascade_ ));
    InMux I__11029 (
            .O(N__46741),
            .I(N__46738));
    LocalMux I__11028 (
            .O(N__46738),
            .I(N__46735));
    Span4Mux_h I__11027 (
            .O(N__46735),
            .I(N__46726));
    InMux I__11026 (
            .O(N__46734),
            .I(N__46719));
    InMux I__11025 (
            .O(N__46733),
            .I(N__46719));
    InMux I__11024 (
            .O(N__46732),
            .I(N__46719));
    InMux I__11023 (
            .O(N__46731),
            .I(N__46714));
    InMux I__11022 (
            .O(N__46730),
            .I(N__46714));
    InMux I__11021 (
            .O(N__46729),
            .I(N__46711));
    Odrv4 I__11020 (
            .O(N__46726),
            .I(\u0.N_2104 ));
    LocalMux I__11019 (
            .O(N__46719),
            .I(\u0.N_2104 ));
    LocalMux I__11018 (
            .O(N__46714),
            .I(\u0.N_2104 ));
    LocalMux I__11017 (
            .O(N__46711),
            .I(\u0.N_2104 ));
    InMux I__11016 (
            .O(N__46702),
            .I(N__46698));
    InMux I__11015 (
            .O(N__46701),
            .I(N__46695));
    LocalMux I__11014 (
            .O(N__46698),
            .I(N__46692));
    LocalMux I__11013 (
            .O(N__46695),
            .I(N__46689));
    Span12Mux_v I__11012 (
            .O(N__46692),
            .I(N__46686));
    Span4Mux_v I__11011 (
            .O(N__46689),
            .I(N__46683));
    Span12Mux_h I__11010 (
            .O(N__46686),
            .I(N__46680));
    Odrv4 I__11009 (
            .O(N__46683),
            .I(DMA_dev0_Teoc_4));
    Odrv12 I__11008 (
            .O(N__46680),
            .I(DMA_dev0_Teoc_4));
    InMux I__11007 (
            .O(N__46675),
            .I(N__46672));
    LocalMux I__11006 (
            .O(N__46672),
            .I(N__46669));
    Odrv4 I__11005 (
            .O(N__46669),
            .I(\u0.N_1686 ));
    InMux I__11004 (
            .O(N__46666),
            .I(N__46663));
    LocalMux I__11003 (
            .O(N__46663),
            .I(N_1321));
    InMux I__11002 (
            .O(N__46660),
            .I(N__46657));
    LocalMux I__11001 (
            .O(N__46657),
            .I(N__46654));
    Span4Mux_h I__11000 (
            .O(N__46654),
            .I(N__46651));
    Odrv4 I__10999 (
            .O(N__46651),
            .I(DMAq_24));
    CascadeMux I__10998 (
            .O(N__46648),
            .I(N_2119_cascade_));
    InMux I__10997 (
            .O(N__46645),
            .I(N__46642));
    LocalMux I__10996 (
            .O(N__46642),
            .I(N__46639));
    Span12Mux_h I__10995 (
            .O(N__46639),
            .I(N__46635));
    InMux I__10994 (
            .O(N__46638),
            .I(N__46632));
    Odrv12 I__10993 (
            .O(N__46635),
            .I(DMA_dev0_Teoc_0));
    LocalMux I__10992 (
            .O(N__46632),
            .I(DMA_dev0_Teoc_0));
    InMux I__10991 (
            .O(N__46627),
            .I(N__46624));
    LocalMux I__10990 (
            .O(N__46624),
            .I(N__46620));
    InMux I__10989 (
            .O(N__46623),
            .I(N__46617));
    Span4Mux_v I__10988 (
            .O(N__46620),
            .I(N__46614));
    LocalMux I__10987 (
            .O(N__46617),
            .I(N__46611));
    Odrv4 I__10986 (
            .O(N__46614),
            .I(PIO_dport0_Teoc_4));
    Odrv12 I__10985 (
            .O(N__46611),
            .I(PIO_dport0_Teoc_4));
    CascadeMux I__10984 (
            .O(N__46606),
            .I(\u0.N_1688_cascade_ ));
    InMux I__10983 (
            .O(N__46603),
            .I(N__46598));
    InMux I__10982 (
            .O(N__46602),
            .I(N__46595));
    InMux I__10981 (
            .O(N__46601),
            .I(N__46590));
    LocalMux I__10980 (
            .O(N__46598),
            .I(N__46586));
    LocalMux I__10979 (
            .O(N__46595),
            .I(N__46583));
    InMux I__10978 (
            .O(N__46594),
            .I(N__46580));
    InMux I__10977 (
            .O(N__46593),
            .I(N__46577));
    LocalMux I__10976 (
            .O(N__46590),
            .I(N__46574));
    InMux I__10975 (
            .O(N__46589),
            .I(N__46571));
    Span4Mux_v I__10974 (
            .O(N__46586),
            .I(N__46568));
    Span4Mux_v I__10973 (
            .O(N__46583),
            .I(N__46559));
    LocalMux I__10972 (
            .O(N__46580),
            .I(N__46559));
    LocalMux I__10971 (
            .O(N__46577),
            .I(N__46559));
    Span4Mux_h I__10970 (
            .O(N__46574),
            .I(N__46554));
    LocalMux I__10969 (
            .O(N__46571),
            .I(N__46554));
    Span4Mux_h I__10968 (
            .O(N__46568),
            .I(N__46551));
    InMux I__10967 (
            .O(N__46567),
            .I(N__46546));
    InMux I__10966 (
            .O(N__46566),
            .I(N__46546));
    Span4Mux_h I__10965 (
            .O(N__46559),
            .I(N__46541));
    Span4Mux_v I__10964 (
            .O(N__46554),
            .I(N__46541));
    Span4Mux_h I__10963 (
            .O(N__46551),
            .I(N__46536));
    LocalMux I__10962 (
            .O(N__46546),
            .I(N__46536));
    Sp12to4 I__10961 (
            .O(N__46541),
            .I(N__46532));
    Span4Mux_v I__10960 (
            .O(N__46536),
            .I(N__46529));
    InMux I__10959 (
            .O(N__46535),
            .I(N__46526));
    Odrv12 I__10958 (
            .O(N__46532),
            .I(\u0.N_2137 ));
    Odrv4 I__10957 (
            .O(N__46529),
            .I(\u0.N_2137 ));
    LocalMux I__10956 (
            .O(N__46526),
            .I(\u0.N_2137 ));
    InMux I__10955 (
            .O(N__46519),
            .I(N__46515));
    InMux I__10954 (
            .O(N__46518),
            .I(N__46512));
    LocalMux I__10953 (
            .O(N__46515),
            .I(N__46509));
    LocalMux I__10952 (
            .O(N__46512),
            .I(N__46506));
    Span4Mux_v I__10951 (
            .O(N__46509),
            .I(N__46503));
    Span4Mux_h I__10950 (
            .O(N__46506),
            .I(N__46500));
    Odrv4 I__10949 (
            .O(N__46503),
            .I(PIO_dport1_Teoc_4));
    Odrv4 I__10948 (
            .O(N__46500),
            .I(PIO_dport1_Teoc_4));
    InMux I__10947 (
            .O(N__46495),
            .I(N__46492));
    LocalMux I__10946 (
            .O(N__46492),
            .I(N__46489));
    Span4Mux_v I__10945 (
            .O(N__46489),
            .I(N__46486));
    Span4Mux_h I__10944 (
            .O(N__46486),
            .I(N__46483));
    Odrv4 I__10943 (
            .O(N__46483),
            .I(\u0.dat_o_i_i_1_28 ));
    CascadeMux I__10942 (
            .O(N__46480),
            .I(\u0.N_2137_cascade_ ));
    InMux I__10941 (
            .O(N__46477),
            .I(N__46474));
    LocalMux I__10940 (
            .O(N__46474),
            .I(\u0.dat_o_i_i_2_28 ));
    CascadeMux I__10939 (
            .O(N__46471),
            .I(\u0.dat_o_i_i_4_28_cascade_ ));
    InMux I__10938 (
            .O(N__46468),
            .I(N__46465));
    LocalMux I__10937 (
            .O(N__46465),
            .I(N__46462));
    Span4Mux_v I__10936 (
            .O(N__46462),
            .I(N__46459));
    Sp12to4 I__10935 (
            .O(N__46459),
            .I(N__46456));
    Span12Mux_h I__10934 (
            .O(N__46456),
            .I(N__46453));
    Odrv12 I__10933 (
            .O(N__46453),
            .I(\u0.N_1689 ));
    IoInMux I__10932 (
            .O(N__46450),
            .I(N__46447));
    LocalMux I__10931 (
            .O(N__46447),
            .I(N__46444));
    Span4Mux_s0_v I__10930 (
            .O(N__46444),
            .I(N__46441));
    Span4Mux_v I__10929 (
            .O(N__46441),
            .I(N__46438));
    Span4Mux_v I__10928 (
            .O(N__46438),
            .I(N__46435));
    Span4Mux_v I__10927 (
            .O(N__46435),
            .I(N__46432));
    Odrv4 I__10926 (
            .O(N__46432),
            .I(N_271));
    InMux I__10925 (
            .O(N__46429),
            .I(N__46426));
    LocalMux I__10924 (
            .O(N__46426),
            .I(\u0.N_1699 ));
    CascadeMux I__10923 (
            .O(N__46423),
            .I(N__46420));
    InMux I__10922 (
            .O(N__46420),
            .I(N__46417));
    LocalMux I__10921 (
            .O(N__46417),
            .I(N__46409));
    InMux I__10920 (
            .O(N__46416),
            .I(N__46402));
    InMux I__10919 (
            .O(N__46415),
            .I(N__46402));
    InMux I__10918 (
            .O(N__46414),
            .I(N__46402));
    InMux I__10917 (
            .O(N__46413),
            .I(N__46399));
    InMux I__10916 (
            .O(N__46412),
            .I(N__46396));
    Odrv4 I__10915 (
            .O(N__46409),
            .I(\u0.N_2095 ));
    LocalMux I__10914 (
            .O(N__46402),
            .I(\u0.N_2095 ));
    LocalMux I__10913 (
            .O(N__46399),
            .I(\u0.N_2095 ));
    LocalMux I__10912 (
            .O(N__46396),
            .I(\u0.N_2095 ));
    CascadeMux I__10911 (
            .O(N__46387),
            .I(\u0.N_2095_cascade_ ));
    CascadeMux I__10910 (
            .O(N__46384),
            .I(N__46381));
    InMux I__10909 (
            .O(N__46381),
            .I(N__46378));
    LocalMux I__10908 (
            .O(N__46378),
            .I(N__46375));
    Span4Mux_v I__10907 (
            .O(N__46375),
            .I(N__46372));
    Odrv4 I__10906 (
            .O(N__46372),
            .I(DMAq_11));
    InMux I__10905 (
            .O(N__46369),
            .I(N__46366));
    LocalMux I__10904 (
            .O(N__46366),
            .I(N__46363));
    Span12Mux_s11_v I__10903 (
            .O(N__46363),
            .I(N__46360));
    Span12Mux_h I__10902 (
            .O(N__46360),
            .I(N__46357));
    Odrv12 I__10901 (
            .O(N__46357),
            .I(PIOq_11));
    InMux I__10900 (
            .O(N__46354),
            .I(N__46351));
    LocalMux I__10899 (
            .O(N__46351),
            .I(N__46348));
    Span12Mux_h I__10898 (
            .O(N__46348),
            .I(N__46345));
    Odrv12 I__10897 (
            .O(N__46345),
            .I(\u0.dat_o_0_0_1Z0Z_11 ));
    InMux I__10896 (
            .O(N__46342),
            .I(N__46339));
    LocalMux I__10895 (
            .O(N__46339),
            .I(N__46336));
    Span4Mux_v I__10894 (
            .O(N__46336),
            .I(N__46333));
    Span4Mux_h I__10893 (
            .O(N__46333),
            .I(N__46330));
    Odrv4 I__10892 (
            .O(N__46330),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNICV4NZ0Z_9 ));
    InMux I__10891 (
            .O(N__46327),
            .I(N__46324));
    LocalMux I__10890 (
            .O(N__46324),
            .I(N__46321));
    Span4Mux_v I__10889 (
            .O(N__46321),
            .I(N__46318));
    Odrv4 I__10888 (
            .O(N__46318),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI8FCMZ0Z_9 ));
    InMux I__10887 (
            .O(N__46315),
            .I(N__46312));
    LocalMux I__10886 (
            .O(N__46312),
            .I(N__46309));
    Odrv4 I__10885 (
            .O(N__46309),
            .I(mem_mem_ram6__RNI33PD1_9));
    CascadeMux I__10884 (
            .O(N__46306),
            .I(iQ_RNI6POK1_2_cascade_));
    InMux I__10883 (
            .O(N__46303),
            .I(N__46299));
    InMux I__10882 (
            .O(N__46302),
            .I(N__46296));
    LocalMux I__10881 (
            .O(N__46299),
            .I(N__46291));
    LocalMux I__10880 (
            .O(N__46296),
            .I(N__46291));
    Span4Mux_v I__10879 (
            .O(N__46291),
            .I(N__46285));
    InMux I__10878 (
            .O(N__46290),
            .I(N__46282));
    InMux I__10877 (
            .O(N__46289),
            .I(N__46279));
    InMux I__10876 (
            .O(N__46288),
            .I(N__46276));
    Span4Mux_h I__10875 (
            .O(N__46285),
            .I(N__46273));
    LocalMux I__10874 (
            .O(N__46282),
            .I(N__46266));
    LocalMux I__10873 (
            .O(N__46279),
            .I(N__46266));
    LocalMux I__10872 (
            .O(N__46276),
            .I(N__46261));
    Span4Mux_h I__10871 (
            .O(N__46273),
            .I(N__46258));
    InMux I__10870 (
            .O(N__46272),
            .I(N__46255));
    InMux I__10869 (
            .O(N__46271),
            .I(N__46252));
    Span4Mux_v I__10868 (
            .O(N__46266),
            .I(N__46249));
    InMux I__10867 (
            .O(N__46265),
            .I(N__46246));
    InMux I__10866 (
            .O(N__46264),
            .I(N__46243));
    Span4Mux_v I__10865 (
            .O(N__46261),
            .I(N__46240));
    Span4Mux_v I__10864 (
            .O(N__46258),
            .I(N__46233));
    LocalMux I__10863 (
            .O(N__46255),
            .I(N__46233));
    LocalMux I__10862 (
            .O(N__46252),
            .I(N__46233));
    Span4Mux_h I__10861 (
            .O(N__46249),
            .I(N__46228));
    LocalMux I__10860 (
            .O(N__46246),
            .I(N__46228));
    LocalMux I__10859 (
            .O(N__46243),
            .I(N__46225));
    Sp12to4 I__10858 (
            .O(N__46240),
            .I(N__46222));
    Span4Mux_v I__10857 (
            .O(N__46233),
            .I(N__46219));
    Span4Mux_v I__10856 (
            .O(N__46228),
            .I(N__46216));
    Span12Mux_h I__10855 (
            .O(N__46225),
            .I(N__46213));
    Span12Mux_s11_h I__10854 (
            .O(N__46222),
            .I(N__46210));
    Span4Mux_v I__10853 (
            .O(N__46219),
            .I(N__46207));
    Span4Mux_v I__10852 (
            .O(N__46216),
            .I(N__46204));
    Span12Mux_v I__10851 (
            .O(N__46213),
            .I(N__46201));
    Span12Mux_v I__10850 (
            .O(N__46210),
            .I(N__46196));
    Sp12to4 I__10849 (
            .O(N__46207),
            .I(N__46196));
    Sp12to4 I__10848 (
            .O(N__46204),
            .I(N__46193));
    Span12Mux_h I__10847 (
            .O(N__46201),
            .I(N__46190));
    Span12Mux_h I__10846 (
            .O(N__46196),
            .I(N__46187));
    Span12Mux_h I__10845 (
            .O(N__46193),
            .I(N__46184));
    Odrv12 I__10844 (
            .O(N__46190),
            .I(wb_dat_i_c_5));
    Odrv12 I__10843 (
            .O(N__46187),
            .I(wb_dat_i_c_5));
    Odrv12 I__10842 (
            .O(N__46184),
            .I(wb_dat_i_c_5));
    CascadeMux I__10841 (
            .O(N__46177),
            .I(N__46174));
    InMux I__10840 (
            .O(N__46174),
            .I(N__46170));
    InMux I__10839 (
            .O(N__46173),
            .I(N__46167));
    LocalMux I__10838 (
            .O(N__46170),
            .I(N__46164));
    LocalMux I__10837 (
            .O(N__46167),
            .I(N__46161));
    Span4Mux_v I__10836 (
            .O(N__46164),
            .I(N__46156));
    Span4Mux_h I__10835 (
            .O(N__46161),
            .I(N__46156));
    Span4Mux_h I__10834 (
            .O(N__46156),
            .I(N__46153));
    Odrv4 I__10833 (
            .O(N__46153),
            .I(PIO_dport0_T1_5));
    InMux I__10832 (
            .O(N__46150),
            .I(N__46146));
    InMux I__10831 (
            .O(N__46149),
            .I(N__46143));
    LocalMux I__10830 (
            .O(N__46146),
            .I(N__46140));
    LocalMux I__10829 (
            .O(N__46143),
            .I(N__46137));
    Span4Mux_h I__10828 (
            .O(N__46140),
            .I(N__46132));
    Span4Mux_v I__10827 (
            .O(N__46137),
            .I(N__46132));
    Span4Mux_h I__10826 (
            .O(N__46132),
            .I(N__46128));
    InMux I__10825 (
            .O(N__46131),
            .I(N__46125));
    Span4Mux_h I__10824 (
            .O(N__46128),
            .I(N__46118));
    LocalMux I__10823 (
            .O(N__46125),
            .I(N__46118));
    InMux I__10822 (
            .O(N__46124),
            .I(N__46115));
    InMux I__10821 (
            .O(N__46123),
            .I(N__46112));
    Span4Mux_v I__10820 (
            .O(N__46118),
            .I(N__46106));
    LocalMux I__10819 (
            .O(N__46115),
            .I(N__46106));
    LocalMux I__10818 (
            .O(N__46112),
            .I(N__46102));
    InMux I__10817 (
            .O(N__46111),
            .I(N__46099));
    Span4Mux_v I__10816 (
            .O(N__46106),
            .I(N__46096));
    InMux I__10815 (
            .O(N__46105),
            .I(N__46093));
    Span4Mux_v I__10814 (
            .O(N__46102),
            .I(N__46090));
    LocalMux I__10813 (
            .O(N__46099),
            .I(N__46087));
    Sp12to4 I__10812 (
            .O(N__46096),
            .I(N__46084));
    LocalMux I__10811 (
            .O(N__46093),
            .I(N__46081));
    Sp12to4 I__10810 (
            .O(N__46090),
            .I(N__46076));
    Span12Mux_v I__10809 (
            .O(N__46087),
            .I(N__46076));
    Span12Mux_h I__10808 (
            .O(N__46084),
            .I(N__46073));
    Span12Mux_h I__10807 (
            .O(N__46081),
            .I(N__46070));
    Span12Mux_h I__10806 (
            .O(N__46076),
            .I(N__46067));
    Odrv12 I__10805 (
            .O(N__46073),
            .I(wb_dat_i_c_28));
    Odrv12 I__10804 (
            .O(N__46070),
            .I(wb_dat_i_c_28));
    Odrv12 I__10803 (
            .O(N__46067),
            .I(wb_dat_i_c_28));
    InMux I__10802 (
            .O(N__46060),
            .I(N__46057));
    LocalMux I__10801 (
            .O(N__46057),
            .I(N__46054));
    Odrv4 I__10800 (
            .O(N__46054),
            .I(\u0.N_1695 ));
    InMux I__10799 (
            .O(N__46051),
            .I(N__46048));
    LocalMux I__10798 (
            .O(N__46048),
            .I(N__46045));
    Span4Mux_v I__10797 (
            .O(N__46045),
            .I(N__46042));
    Sp12to4 I__10796 (
            .O(N__46042),
            .I(N__46039));
    Odrv12 I__10795 (
            .O(N__46039),
            .I(\u0.dat_o_0_0_0_9 ));
    InMux I__10794 (
            .O(N__46036),
            .I(N__46033));
    LocalMux I__10793 (
            .O(N__46033),
            .I(N__46030));
    Span4Mux_v I__10792 (
            .O(N__46030),
            .I(N__46027));
    Span4Mux_h I__10791 (
            .O(N__46027),
            .I(N__46024));
    Odrv4 I__10790 (
            .O(N__46024),
            .I(\u0.dat_o_0_0_3_9 ));
    InMux I__10789 (
            .O(N__46021),
            .I(N__46018));
    LocalMux I__10788 (
            .O(N__46018),
            .I(N__46014));
    InMux I__10787 (
            .O(N__46017),
            .I(N__46011));
    Span4Mux_v I__10786 (
            .O(N__46014),
            .I(N__46008));
    LocalMux I__10785 (
            .O(N__46011),
            .I(N__46005));
    Odrv4 I__10784 (
            .O(N__46008),
            .I(PIO_dport0_T2_1));
    Odrv12 I__10783 (
            .O(N__46005),
            .I(PIO_dport0_T2_1));
    InMux I__10782 (
            .O(N__46000),
            .I(N__45997));
    LocalMux I__10781 (
            .O(N__45997),
            .I(N__45994));
    Odrv4 I__10780 (
            .O(N__45994),
            .I(\u0.CtrlRegZ0Z_28 ));
    InMux I__10779 (
            .O(N__45991),
            .I(N__45988));
    LocalMux I__10778 (
            .O(N__45988),
            .I(mem_mem_ram6__RNI00PD1_8));
    CascadeMux I__10777 (
            .O(N__45985),
            .I(iQ_RNI2LOK1_2_cascade_));
    InMux I__10776 (
            .O(N__45982),
            .I(N__45979));
    LocalMux I__10775 (
            .O(N__45979),
            .I(\u0.N_1735 ));
    InMux I__10774 (
            .O(N__45976),
            .I(N__45971));
    InMux I__10773 (
            .O(N__45975),
            .I(N__45966));
    InMux I__10772 (
            .O(N__45974),
            .I(N__45966));
    LocalMux I__10771 (
            .O(N__45971),
            .I(N__45963));
    LocalMux I__10770 (
            .O(N__45966),
            .I(N__45960));
    Span4Mux_h I__10769 (
            .O(N__45963),
            .I(N__45955));
    Span4Mux_v I__10768 (
            .O(N__45960),
            .I(N__45955));
    Span4Mux_h I__10767 (
            .O(N__45955),
            .I(N__45952));
    Span4Mux_v I__10766 (
            .O(N__45952),
            .I(N__45949));
    Span4Mux_v I__10765 (
            .O(N__45949),
            .I(N__45946));
    Span4Mux_v I__10764 (
            .O(N__45946),
            .I(N__45943));
    Sp12to4 I__10763 (
            .O(N__45943),
            .I(N__45940));
    Odrv12 I__10762 (
            .O(N__45940),
            .I(dd_pad_i_c_9));
    CEMux I__10761 (
            .O(N__45937),
            .I(N__45933));
    CEMux I__10760 (
            .O(N__45936),
            .I(N__45928));
    LocalMux I__10759 (
            .O(N__45933),
            .I(N__45922));
    CEMux I__10758 (
            .O(N__45932),
            .I(N__45919));
    CEMux I__10757 (
            .O(N__45931),
            .I(N__45916));
    LocalMux I__10756 (
            .O(N__45928),
            .I(N__45913));
    CEMux I__10755 (
            .O(N__45927),
            .I(N__45910));
    CEMux I__10754 (
            .O(N__45926),
            .I(N__45904));
    CEMux I__10753 (
            .O(N__45925),
            .I(N__45900));
    Span4Mux_h I__10752 (
            .O(N__45922),
            .I(N__45896));
    LocalMux I__10751 (
            .O(N__45919),
            .I(N__45893));
    LocalMux I__10750 (
            .O(N__45916),
            .I(N__45890));
    Span4Mux_v I__10749 (
            .O(N__45913),
            .I(N__45885));
    LocalMux I__10748 (
            .O(N__45910),
            .I(N__45885));
    CEMux I__10747 (
            .O(N__45909),
            .I(N__45882));
    CEMux I__10746 (
            .O(N__45908),
            .I(N__45877));
    CEMux I__10745 (
            .O(N__45907),
            .I(N__45874));
    LocalMux I__10744 (
            .O(N__45904),
            .I(N__45870));
    CEMux I__10743 (
            .O(N__45903),
            .I(N__45867));
    LocalMux I__10742 (
            .O(N__45900),
            .I(N__45864));
    CEMux I__10741 (
            .O(N__45899),
            .I(N__45861));
    Span4Mux_v I__10740 (
            .O(N__45896),
            .I(N__45856));
    Span4Mux_v I__10739 (
            .O(N__45893),
            .I(N__45856));
    Span4Mux_v I__10738 (
            .O(N__45890),
            .I(N__45853));
    Span4Mux_v I__10737 (
            .O(N__45885),
            .I(N__45848));
    LocalMux I__10736 (
            .O(N__45882),
            .I(N__45848));
    CEMux I__10735 (
            .O(N__45881),
            .I(N__45845));
    CEMux I__10734 (
            .O(N__45880),
            .I(N__45842));
    LocalMux I__10733 (
            .O(N__45877),
            .I(N__45839));
    LocalMux I__10732 (
            .O(N__45874),
            .I(N__45836));
    CEMux I__10731 (
            .O(N__45873),
            .I(N__45833));
    Span4Mux_v I__10730 (
            .O(N__45870),
            .I(N__45830));
    LocalMux I__10729 (
            .O(N__45867),
            .I(N__45823));
    Span4Mux_h I__10728 (
            .O(N__45864),
            .I(N__45823));
    LocalMux I__10727 (
            .O(N__45861),
            .I(N__45823));
    Sp12to4 I__10726 (
            .O(N__45856),
            .I(N__45820));
    Span4Mux_v I__10725 (
            .O(N__45853),
            .I(N__45817));
    Span4Mux_h I__10724 (
            .O(N__45848),
            .I(N__45814));
    LocalMux I__10723 (
            .O(N__45845),
            .I(N__45811));
    LocalMux I__10722 (
            .O(N__45842),
            .I(N__45808));
    Span4Mux_h I__10721 (
            .O(N__45839),
            .I(N__45805));
    Span4Mux_h I__10720 (
            .O(N__45836),
            .I(N__45802));
    LocalMux I__10719 (
            .O(N__45833),
            .I(N__45797));
    Span4Mux_h I__10718 (
            .O(N__45830),
            .I(N__45797));
    Span4Mux_v I__10717 (
            .O(N__45823),
            .I(N__45794));
    Span12Mux_h I__10716 (
            .O(N__45820),
            .I(N__45791));
    Span4Mux_v I__10715 (
            .O(N__45817),
            .I(N__45788));
    Sp12to4 I__10714 (
            .O(N__45814),
            .I(N__45785));
    Span12Mux_v I__10713 (
            .O(N__45811),
            .I(N__45782));
    Span4Mux_v I__10712 (
            .O(N__45808),
            .I(N__45775));
    Span4Mux_h I__10711 (
            .O(N__45805),
            .I(N__45775));
    Span4Mux_v I__10710 (
            .O(N__45802),
            .I(N__45775));
    Span4Mux_h I__10709 (
            .O(N__45797),
            .I(N__45770));
    Span4Mux_h I__10708 (
            .O(N__45794),
            .I(N__45770));
    Span12Mux_v I__10707 (
            .O(N__45791),
            .I(N__45763));
    Sp12to4 I__10706 (
            .O(N__45788),
            .I(N__45763));
    Span12Mux_v I__10705 (
            .O(N__45785),
            .I(N__45763));
    Odrv12 I__10704 (
            .O(N__45782),
            .I(\u1.PIO_control.PIO_access_control.dstrb ));
    Odrv4 I__10703 (
            .O(N__45775),
            .I(\u1.PIO_control.PIO_access_control.dstrb ));
    Odrv4 I__10702 (
            .O(N__45770),
            .I(\u1.PIO_control.PIO_access_control.dstrb ));
    Odrv12 I__10701 (
            .O(N__45763),
            .I(\u1.PIO_control.PIO_access_control.dstrb ));
    InMux I__10700 (
            .O(N__45754),
            .I(N__45751));
    LocalMux I__10699 (
            .O(N__45751),
            .I(N__45747));
    InMux I__10698 (
            .O(N__45750),
            .I(N__45744));
    Span4Mux_v I__10697 (
            .O(N__45747),
            .I(N__45741));
    LocalMux I__10696 (
            .O(N__45744),
            .I(N__45738));
    Span4Mux_v I__10695 (
            .O(N__45741),
            .I(N__45735));
    Span4Mux_h I__10694 (
            .O(N__45738),
            .I(N__45732));
    Odrv4 I__10693 (
            .O(N__45735),
            .I(PIO_cmdport_T4_1));
    Odrv4 I__10692 (
            .O(N__45732),
            .I(PIO_cmdport_T4_1));
    InMux I__10691 (
            .O(N__45727),
            .I(N__45724));
    LocalMux I__10690 (
            .O(N__45724),
            .I(N__45721));
    Span4Mux_h I__10689 (
            .O(N__45721),
            .I(N__45718));
    Odrv4 I__10688 (
            .O(N__45718),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_17 ));
    InMux I__10687 (
            .O(N__45715),
            .I(N__45712));
    LocalMux I__10686 (
            .O(N__45712),
            .I(N__45709));
    Span4Mux_h I__10685 (
            .O(N__45709),
            .I(N__45706));
    Odrv4 I__10684 (
            .O(N__45706),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_17 ));
    CascadeMux I__10683 (
            .O(N__45703),
            .I(N__45677));
    InMux I__10682 (
            .O(N__45702),
            .I(N__45670));
    InMux I__10681 (
            .O(N__45701),
            .I(N__45664));
    InMux I__10680 (
            .O(N__45700),
            .I(N__45645));
    InMux I__10679 (
            .O(N__45699),
            .I(N__45645));
    InMux I__10678 (
            .O(N__45698),
            .I(N__45638));
    InMux I__10677 (
            .O(N__45697),
            .I(N__45638));
    InMux I__10676 (
            .O(N__45696),
            .I(N__45638));
    InMux I__10675 (
            .O(N__45695),
            .I(N__45625));
    InMux I__10674 (
            .O(N__45694),
            .I(N__45625));
    InMux I__10673 (
            .O(N__45693),
            .I(N__45625));
    InMux I__10672 (
            .O(N__45692),
            .I(N__45620));
    InMux I__10671 (
            .O(N__45691),
            .I(N__45620));
    InMux I__10670 (
            .O(N__45690),
            .I(N__45610));
    InMux I__10669 (
            .O(N__45689),
            .I(N__45610));
    InMux I__10668 (
            .O(N__45688),
            .I(N__45607));
    InMux I__10667 (
            .O(N__45687),
            .I(N__45604));
    InMux I__10666 (
            .O(N__45686),
            .I(N__45595));
    InMux I__10665 (
            .O(N__45685),
            .I(N__45595));
    InMux I__10664 (
            .O(N__45684),
            .I(N__45595));
    InMux I__10663 (
            .O(N__45683),
            .I(N__45595));
    InMux I__10662 (
            .O(N__45682),
            .I(N__45588));
    InMux I__10661 (
            .O(N__45681),
            .I(N__45588));
    InMux I__10660 (
            .O(N__45680),
            .I(N__45588));
    InMux I__10659 (
            .O(N__45677),
            .I(N__45583));
    InMux I__10658 (
            .O(N__45676),
            .I(N__45583));
    InMux I__10657 (
            .O(N__45675),
            .I(N__45576));
    InMux I__10656 (
            .O(N__45674),
            .I(N__45576));
    InMux I__10655 (
            .O(N__45673),
            .I(N__45576));
    LocalMux I__10654 (
            .O(N__45670),
            .I(N__45573));
    InMux I__10653 (
            .O(N__45669),
            .I(N__45566));
    InMux I__10652 (
            .O(N__45668),
            .I(N__45566));
    InMux I__10651 (
            .O(N__45667),
            .I(N__45566));
    LocalMux I__10650 (
            .O(N__45664),
            .I(N__45563));
    InMux I__10649 (
            .O(N__45663),
            .I(N__45560));
    InMux I__10648 (
            .O(N__45662),
            .I(N__45553));
    InMux I__10647 (
            .O(N__45661),
            .I(N__45553));
    InMux I__10646 (
            .O(N__45660),
            .I(N__45553));
    InMux I__10645 (
            .O(N__45659),
            .I(N__45546));
    InMux I__10644 (
            .O(N__45658),
            .I(N__45539));
    InMux I__10643 (
            .O(N__45657),
            .I(N__45539));
    InMux I__10642 (
            .O(N__45656),
            .I(N__45539));
    InMux I__10641 (
            .O(N__45655),
            .I(N__45532));
    InMux I__10640 (
            .O(N__45654),
            .I(N__45532));
    InMux I__10639 (
            .O(N__45653),
            .I(N__45532));
    InMux I__10638 (
            .O(N__45652),
            .I(N__45525));
    InMux I__10637 (
            .O(N__45651),
            .I(N__45525));
    InMux I__10636 (
            .O(N__45650),
            .I(N__45525));
    LocalMux I__10635 (
            .O(N__45645),
            .I(N__45520));
    LocalMux I__10634 (
            .O(N__45638),
            .I(N__45520));
    InMux I__10633 (
            .O(N__45637),
            .I(N__45515));
    InMux I__10632 (
            .O(N__45636),
            .I(N__45515));
    InMux I__10631 (
            .O(N__45635),
            .I(N__45496));
    InMux I__10630 (
            .O(N__45634),
            .I(N__45496));
    InMux I__10629 (
            .O(N__45633),
            .I(N__45496));
    InMux I__10628 (
            .O(N__45632),
            .I(N__45496));
    LocalMux I__10627 (
            .O(N__45625),
            .I(N__45489));
    LocalMux I__10626 (
            .O(N__45620),
            .I(N__45486));
    InMux I__10625 (
            .O(N__45619),
            .I(N__45481));
    InMux I__10624 (
            .O(N__45618),
            .I(N__45481));
    InMux I__10623 (
            .O(N__45617),
            .I(N__45474));
    InMux I__10622 (
            .O(N__45616),
            .I(N__45474));
    InMux I__10621 (
            .O(N__45615),
            .I(N__45474));
    LocalMux I__10620 (
            .O(N__45610),
            .I(N__45467));
    LocalMux I__10619 (
            .O(N__45607),
            .I(N__45467));
    LocalMux I__10618 (
            .O(N__45604),
            .I(N__45467));
    LocalMux I__10617 (
            .O(N__45595),
            .I(N__45458));
    LocalMux I__10616 (
            .O(N__45588),
            .I(N__45453));
    LocalMux I__10615 (
            .O(N__45583),
            .I(N__45453));
    LocalMux I__10614 (
            .O(N__45576),
            .I(N__45440));
    Span4Mux_h I__10613 (
            .O(N__45573),
            .I(N__45440));
    LocalMux I__10612 (
            .O(N__45566),
            .I(N__45440));
    Span4Mux_h I__10611 (
            .O(N__45563),
            .I(N__45440));
    LocalMux I__10610 (
            .O(N__45560),
            .I(N__45440));
    LocalMux I__10609 (
            .O(N__45553),
            .I(N__45440));
    InMux I__10608 (
            .O(N__45552),
            .I(N__45437));
    InMux I__10607 (
            .O(N__45551),
            .I(N__45434));
    CascadeMux I__10606 (
            .O(N__45550),
            .I(N__45431));
    CascadeMux I__10605 (
            .O(N__45549),
            .I(N__45427));
    LocalMux I__10604 (
            .O(N__45546),
            .I(N__45408));
    LocalMux I__10603 (
            .O(N__45539),
            .I(N__45408));
    LocalMux I__10602 (
            .O(N__45532),
            .I(N__45408));
    LocalMux I__10601 (
            .O(N__45525),
            .I(N__45408));
    Span4Mux_v I__10600 (
            .O(N__45520),
            .I(N__45403));
    LocalMux I__10599 (
            .O(N__45515),
            .I(N__45403));
    InMux I__10598 (
            .O(N__45514),
            .I(N__45394));
    InMux I__10597 (
            .O(N__45513),
            .I(N__45394));
    InMux I__10596 (
            .O(N__45512),
            .I(N__45394));
    InMux I__10595 (
            .O(N__45511),
            .I(N__45394));
    InMux I__10594 (
            .O(N__45510),
            .I(N__45381));
    InMux I__10593 (
            .O(N__45509),
            .I(N__45381));
    InMux I__10592 (
            .O(N__45508),
            .I(N__45381));
    InMux I__10591 (
            .O(N__45507),
            .I(N__45381));
    InMux I__10590 (
            .O(N__45506),
            .I(N__45381));
    InMux I__10589 (
            .O(N__45505),
            .I(N__45381));
    LocalMux I__10588 (
            .O(N__45496),
            .I(N__45378));
    InMux I__10587 (
            .O(N__45495),
            .I(N__45369));
    InMux I__10586 (
            .O(N__45494),
            .I(N__45369));
    InMux I__10585 (
            .O(N__45493),
            .I(N__45369));
    InMux I__10584 (
            .O(N__45492),
            .I(N__45369));
    Span4Mux_h I__10583 (
            .O(N__45489),
            .I(N__45360));
    Span4Mux_s1_v I__10582 (
            .O(N__45486),
            .I(N__45360));
    LocalMux I__10581 (
            .O(N__45481),
            .I(N__45360));
    LocalMux I__10580 (
            .O(N__45474),
            .I(N__45360));
    Span4Mux_v I__10579 (
            .O(N__45467),
            .I(N__45357));
    InMux I__10578 (
            .O(N__45466),
            .I(N__45350));
    InMux I__10577 (
            .O(N__45465),
            .I(N__45350));
    InMux I__10576 (
            .O(N__45464),
            .I(N__45350));
    InMux I__10575 (
            .O(N__45463),
            .I(N__45347));
    InMux I__10574 (
            .O(N__45462),
            .I(N__45344));
    CascadeMux I__10573 (
            .O(N__45461),
            .I(N__45341));
    Span4Mux_v I__10572 (
            .O(N__45458),
            .I(N__45334));
    Span4Mux_v I__10571 (
            .O(N__45453),
            .I(N__45325));
    Span4Mux_v I__10570 (
            .O(N__45440),
            .I(N__45325));
    LocalMux I__10569 (
            .O(N__45437),
            .I(N__45325));
    LocalMux I__10568 (
            .O(N__45434),
            .I(N__45325));
    InMux I__10567 (
            .O(N__45431),
            .I(N__45318));
    InMux I__10566 (
            .O(N__45430),
            .I(N__45318));
    InMux I__10565 (
            .O(N__45427),
            .I(N__45318));
    InMux I__10564 (
            .O(N__45426),
            .I(N__45311));
    InMux I__10563 (
            .O(N__45425),
            .I(N__45311));
    InMux I__10562 (
            .O(N__45424),
            .I(N__45311));
    InMux I__10561 (
            .O(N__45423),
            .I(N__45302));
    InMux I__10560 (
            .O(N__45422),
            .I(N__45302));
    InMux I__10559 (
            .O(N__45421),
            .I(N__45302));
    InMux I__10558 (
            .O(N__45420),
            .I(N__45302));
    InMux I__10557 (
            .O(N__45419),
            .I(N__45295));
    InMux I__10556 (
            .O(N__45418),
            .I(N__45295));
    InMux I__10555 (
            .O(N__45417),
            .I(N__45295));
    Span4Mux_v I__10554 (
            .O(N__45408),
            .I(N__45285));
    Span4Mux_h I__10553 (
            .O(N__45403),
            .I(N__45285));
    LocalMux I__10552 (
            .O(N__45394),
            .I(N__45285));
    LocalMux I__10551 (
            .O(N__45381),
            .I(N__45285));
    Span4Mux_h I__10550 (
            .O(N__45378),
            .I(N__45280));
    LocalMux I__10549 (
            .O(N__45369),
            .I(N__45280));
    Span4Mux_v I__10548 (
            .O(N__45360),
            .I(N__45273));
    Span4Mux_h I__10547 (
            .O(N__45357),
            .I(N__45273));
    LocalMux I__10546 (
            .O(N__45350),
            .I(N__45273));
    LocalMux I__10545 (
            .O(N__45347),
            .I(N__45268));
    LocalMux I__10544 (
            .O(N__45344),
            .I(N__45268));
    InMux I__10543 (
            .O(N__45341),
            .I(N__45265));
    InMux I__10542 (
            .O(N__45340),
            .I(N__45262));
    InMux I__10541 (
            .O(N__45339),
            .I(N__45259));
    InMux I__10540 (
            .O(N__45338),
            .I(N__45254));
    InMux I__10539 (
            .O(N__45337),
            .I(N__45254));
    Span4Mux_h I__10538 (
            .O(N__45334),
            .I(N__45250));
    Span4Mux_v I__10537 (
            .O(N__45325),
            .I(N__45247));
    LocalMux I__10536 (
            .O(N__45318),
            .I(N__45244));
    LocalMux I__10535 (
            .O(N__45311),
            .I(N__45237));
    LocalMux I__10534 (
            .O(N__45302),
            .I(N__45237));
    LocalMux I__10533 (
            .O(N__45295),
            .I(N__45237));
    InMux I__10532 (
            .O(N__45294),
            .I(N__45234));
    Span4Mux_v I__10531 (
            .O(N__45285),
            .I(N__45231));
    Span4Mux_v I__10530 (
            .O(N__45280),
            .I(N__45228));
    Span4Mux_v I__10529 (
            .O(N__45273),
            .I(N__45219));
    Span4Mux_h I__10528 (
            .O(N__45268),
            .I(N__45219));
    LocalMux I__10527 (
            .O(N__45265),
            .I(N__45219));
    LocalMux I__10526 (
            .O(N__45262),
            .I(N__45219));
    LocalMux I__10525 (
            .O(N__45259),
            .I(N__45214));
    LocalMux I__10524 (
            .O(N__45254),
            .I(N__45214));
    CascadeMux I__10523 (
            .O(N__45253),
            .I(N__45211));
    Span4Mux_v I__10522 (
            .O(N__45250),
            .I(N__45203));
    Span4Mux_h I__10521 (
            .O(N__45247),
            .I(N__45203));
    Span4Mux_v I__10520 (
            .O(N__45244),
            .I(N__45203));
    Span4Mux_v I__10519 (
            .O(N__45237),
            .I(N__45198));
    LocalMux I__10518 (
            .O(N__45234),
            .I(N__45198));
    Span4Mux_h I__10517 (
            .O(N__45231),
            .I(N__45191));
    Span4Mux_v I__10516 (
            .O(N__45228),
            .I(N__45191));
    Span4Mux_h I__10515 (
            .O(N__45219),
            .I(N__45191));
    Span4Mux_v I__10514 (
            .O(N__45214),
            .I(N__45188));
    InMux I__10513 (
            .O(N__45211),
            .I(N__45183));
    InMux I__10512 (
            .O(N__45210),
            .I(N__45183));
    Span4Mux_v I__10511 (
            .O(N__45203),
            .I(N__45178));
    Span4Mux_v I__10510 (
            .O(N__45198),
            .I(N__45175));
    Span4Mux_v I__10509 (
            .O(N__45191),
            .I(N__45172));
    Span4Mux_v I__10508 (
            .O(N__45188),
            .I(N__45169));
    LocalMux I__10507 (
            .O(N__45183),
            .I(N__45166));
    InMux I__10506 (
            .O(N__45182),
            .I(N__45163));
    InMux I__10505 (
            .O(N__45181),
            .I(N__45160));
    Odrv4 I__10504 (
            .O(N__45178),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_0 ));
    Odrv4 I__10503 (
            .O(N__45175),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_0 ));
    Odrv4 I__10502 (
            .O(N__45172),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_0 ));
    Odrv4 I__10501 (
            .O(N__45169),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_0 ));
    Odrv4 I__10500 (
            .O(N__45166),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_0 ));
    LocalMux I__10499 (
            .O(N__45163),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_0 ));
    LocalMux I__10498 (
            .O(N__45160),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_0 ));
    InMux I__10497 (
            .O(N__45145),
            .I(N__45142));
    LocalMux I__10496 (
            .O(N__45142),
            .I(N__45138));
    InMux I__10495 (
            .O(N__45141),
            .I(N__45135));
    Span4Mux_v I__10494 (
            .O(N__45138),
            .I(N__45130));
    LocalMux I__10493 (
            .O(N__45135),
            .I(N__45127));
    InMux I__10492 (
            .O(N__45134),
            .I(N__45124));
    InMux I__10491 (
            .O(N__45133),
            .I(N__45121));
    Span4Mux_v I__10490 (
            .O(N__45130),
            .I(N__45118));
    Span4Mux_v I__10489 (
            .O(N__45127),
            .I(N__45114));
    LocalMux I__10488 (
            .O(N__45124),
            .I(N__45111));
    LocalMux I__10487 (
            .O(N__45121),
            .I(N__45108));
    Span4Mux_h I__10486 (
            .O(N__45118),
            .I(N__45105));
    InMux I__10485 (
            .O(N__45117),
            .I(N__45102));
    Span4Mux_h I__10484 (
            .O(N__45114),
            .I(N__45099));
    Span4Mux_v I__10483 (
            .O(N__45111),
            .I(N__45096));
    Span4Mux_v I__10482 (
            .O(N__45108),
            .I(N__45093));
    Span4Mux_h I__10481 (
            .O(N__45105),
            .I(N__45088));
    LocalMux I__10480 (
            .O(N__45102),
            .I(N__45088));
    Span4Mux_h I__10479 (
            .O(N__45099),
            .I(N__45083));
    Span4Mux_h I__10478 (
            .O(N__45096),
            .I(N__45083));
    Span4Mux_v I__10477 (
            .O(N__45093),
            .I(N__45080));
    Span4Mux_v I__10476 (
            .O(N__45088),
            .I(N__45077));
    Sp12to4 I__10475 (
            .O(N__45083),
            .I(N__45074));
    Sp12to4 I__10474 (
            .O(N__45080),
            .I(N__45071));
    Span4Mux_v I__10473 (
            .O(N__45077),
            .I(N__45068));
    Span12Mux_v I__10472 (
            .O(N__45074),
            .I(N__45063));
    Span12Mux_h I__10471 (
            .O(N__45071),
            .I(N__45063));
    Span4Mux_h I__10470 (
            .O(N__45068),
            .I(N__45060));
    Odrv12 I__10469 (
            .O(N__45063),
            .I(wb_dat_i_c_17));
    Odrv4 I__10468 (
            .O(N__45060),
            .I(wb_dat_i_c_17));
    InMux I__10467 (
            .O(N__45055),
            .I(N__45052));
    LocalMux I__10466 (
            .O(N__45052),
            .I(\u0.CtrlRegZ0Z_17 ));
    InMux I__10465 (
            .O(N__45049),
            .I(N__45043));
    InMux I__10464 (
            .O(N__45048),
            .I(N__45040));
    InMux I__10463 (
            .O(N__45047),
            .I(N__45037));
    InMux I__10462 (
            .O(N__45046),
            .I(N__45034));
    LocalMux I__10461 (
            .O(N__45043),
            .I(N__45031));
    LocalMux I__10460 (
            .O(N__45040),
            .I(N__45026));
    LocalMux I__10459 (
            .O(N__45037),
            .I(N__45020));
    LocalMux I__10458 (
            .O(N__45034),
            .I(N__45020));
    Span4Mux_v I__10457 (
            .O(N__45031),
            .I(N__45017));
    InMux I__10456 (
            .O(N__45030),
            .I(N__45014));
    InMux I__10455 (
            .O(N__45029),
            .I(N__45011));
    Span4Mux_v I__10454 (
            .O(N__45026),
            .I(N__45008));
    InMux I__10453 (
            .O(N__45025),
            .I(N__45005));
    Span4Mux_v I__10452 (
            .O(N__45020),
            .I(N__44996));
    Span4Mux_h I__10451 (
            .O(N__45017),
            .I(N__44996));
    LocalMux I__10450 (
            .O(N__45014),
            .I(N__44996));
    LocalMux I__10449 (
            .O(N__45011),
            .I(N__44996));
    Span4Mux_h I__10448 (
            .O(N__45008),
            .I(N__44990));
    LocalMux I__10447 (
            .O(N__45005),
            .I(N__44990));
    Span4Mux_h I__10446 (
            .O(N__44996),
            .I(N__44987));
    InMux I__10445 (
            .O(N__44995),
            .I(N__44984));
    Span4Mux_v I__10444 (
            .O(N__44990),
            .I(N__44981));
    Span4Mux_h I__10443 (
            .O(N__44987),
            .I(N__44976));
    LocalMux I__10442 (
            .O(N__44984),
            .I(N__44976));
    Span4Mux_v I__10441 (
            .O(N__44981),
            .I(N__44973));
    Span4Mux_v I__10440 (
            .O(N__44976),
            .I(N__44970));
    Odrv4 I__10439 (
            .O(N__44973),
            .I(\u0.N_2101 ));
    Odrv4 I__10438 (
            .O(N__44970),
            .I(\u0.N_2101 ));
    CascadeMux I__10437 (
            .O(N__44965),
            .I(N__44962));
    InMux I__10436 (
            .O(N__44962),
            .I(N__44959));
    LocalMux I__10435 (
            .O(N__44959),
            .I(N__44956));
    Span4Mux_v I__10434 (
            .O(N__44956),
            .I(N__44953));
    Span4Mux_v I__10433 (
            .O(N__44953),
            .I(N__44950));
    Span4Mux_h I__10432 (
            .O(N__44950),
            .I(N__44946));
    InMux I__10431 (
            .O(N__44949),
            .I(N__44943));
    Odrv4 I__10430 (
            .O(N__44946),
            .I(PIO_cmdport_T4_7));
    LocalMux I__10429 (
            .O(N__44943),
            .I(PIO_cmdport_T4_7));
    CascadeMux I__10428 (
            .O(N__44938),
            .I(N__44932));
    CascadeMux I__10427 (
            .O(N__44937),
            .I(N__44929));
    CascadeMux I__10426 (
            .O(N__44936),
            .I(N__44924));
    CascadeMux I__10425 (
            .O(N__44935),
            .I(N__44921));
    InMux I__10424 (
            .O(N__44932),
            .I(N__44918));
    InMux I__10423 (
            .O(N__44929),
            .I(N__44915));
    InMux I__10422 (
            .O(N__44928),
            .I(N__44912));
    InMux I__10421 (
            .O(N__44927),
            .I(N__44908));
    InMux I__10420 (
            .O(N__44924),
            .I(N__44905));
    InMux I__10419 (
            .O(N__44921),
            .I(N__44901));
    LocalMux I__10418 (
            .O(N__44918),
            .I(N__44894));
    LocalMux I__10417 (
            .O(N__44915),
            .I(N__44894));
    LocalMux I__10416 (
            .O(N__44912),
            .I(N__44894));
    CascadeMux I__10415 (
            .O(N__44911),
            .I(N__44891));
    LocalMux I__10414 (
            .O(N__44908),
            .I(N__44886));
    LocalMux I__10413 (
            .O(N__44905),
            .I(N__44886));
    CascadeMux I__10412 (
            .O(N__44904),
            .I(N__44883));
    LocalMux I__10411 (
            .O(N__44901),
            .I(N__44880));
    Span4Mux_v I__10410 (
            .O(N__44894),
            .I(N__44877));
    InMux I__10409 (
            .O(N__44891),
            .I(N__44874));
    Span4Mux_v I__10408 (
            .O(N__44886),
            .I(N__44871));
    InMux I__10407 (
            .O(N__44883),
            .I(N__44868));
    Span4Mux_h I__10406 (
            .O(N__44880),
            .I(N__44861));
    Span4Mux_h I__10405 (
            .O(N__44877),
            .I(N__44861));
    LocalMux I__10404 (
            .O(N__44874),
            .I(N__44861));
    Sp12to4 I__10403 (
            .O(N__44871),
            .I(N__44856));
    LocalMux I__10402 (
            .O(N__44868),
            .I(N__44856));
    Span4Mux_v I__10401 (
            .O(N__44861),
            .I(N__44853));
    Span12Mux_h I__10400 (
            .O(N__44856),
            .I(N__44850));
    Span4Mux_v I__10399 (
            .O(N__44853),
            .I(N__44847));
    Odrv12 I__10398 (
            .O(N__44850),
            .I(\u0.N_2142 ));
    Odrv4 I__10397 (
            .O(N__44847),
            .I(\u0.N_2142 ));
    InMux I__10396 (
            .O(N__44842),
            .I(N__44839));
    LocalMux I__10395 (
            .O(N__44839),
            .I(N__44835));
    InMux I__10394 (
            .O(N__44838),
            .I(N__44832));
    Span4Mux_h I__10393 (
            .O(N__44835),
            .I(N__44826));
    LocalMux I__10392 (
            .O(N__44832),
            .I(N__44826));
    InMux I__10391 (
            .O(N__44831),
            .I(N__44823));
    Span4Mux_v I__10390 (
            .O(N__44826),
            .I(N__44820));
    LocalMux I__10389 (
            .O(N__44823),
            .I(N__44815));
    Span4Mux_h I__10388 (
            .O(N__44820),
            .I(N__44812));
    InMux I__10387 (
            .O(N__44819),
            .I(N__44809));
    InMux I__10386 (
            .O(N__44818),
            .I(N__44806));
    Span4Mux_v I__10385 (
            .O(N__44815),
            .I(N__44803));
    Span4Mux_h I__10384 (
            .O(N__44812),
            .I(N__44798));
    LocalMux I__10383 (
            .O(N__44809),
            .I(N__44798));
    LocalMux I__10382 (
            .O(N__44806),
            .I(N__44795));
    Sp12to4 I__10381 (
            .O(N__44803),
            .I(N__44792));
    Span4Mux_h I__10380 (
            .O(N__44798),
            .I(N__44789));
    Span12Mux_v I__10379 (
            .O(N__44795),
            .I(N__44786));
    Span12Mux_h I__10378 (
            .O(N__44792),
            .I(N__44783));
    Span4Mux_v I__10377 (
            .O(N__44789),
            .I(N__44780));
    Odrv12 I__10376 (
            .O(N__44786),
            .I(wb_dat_i_c_23));
    Odrv12 I__10375 (
            .O(N__44783),
            .I(wb_dat_i_c_23));
    Odrv4 I__10374 (
            .O(N__44780),
            .I(wb_dat_i_c_23));
    InMux I__10373 (
            .O(N__44773),
            .I(N__44770));
    LocalMux I__10372 (
            .O(N__44770),
            .I(\u0.CtrlRegZ0Z_23 ));
    InMux I__10371 (
            .O(N__44767),
            .I(N__44764));
    LocalMux I__10370 (
            .O(N__44764),
            .I(N__44761));
    Span4Mux_v I__10369 (
            .O(N__44761),
            .I(N__44758));
    Odrv4 I__10368 (
            .O(N__44758),
            .I(u1_DMA_control_gen_DMAbuf_Rxbuf_mem_N_1224));
    CascadeMux I__10367 (
            .O(N__44755),
            .I(N__44752));
    InMux I__10366 (
            .O(N__44752),
            .I(N__44749));
    LocalMux I__10365 (
            .O(N__44749),
            .I(N__44746));
    Span4Mux_h I__10364 (
            .O(N__44746),
            .I(N__44743));
    Odrv4 I__10363 (
            .O(N__44743),
            .I(u1_DMA_control_gen_DMAbuf_Rxbuf_mem_N_1160));
    InMux I__10362 (
            .O(N__44740),
            .I(N__44737));
    LocalMux I__10361 (
            .O(N__44737),
            .I(N__44734));
    Span4Mux_v I__10360 (
            .O(N__44734),
            .I(N__44731));
    Span4Mux_h I__10359 (
            .O(N__44731),
            .I(N__44727));
    InMux I__10358 (
            .O(N__44730),
            .I(N__44724));
    Span4Mux_h I__10357 (
            .O(N__44727),
            .I(N__44719));
    LocalMux I__10356 (
            .O(N__44724),
            .I(N__44719));
    Span4Mux_v I__10355 (
            .O(N__44719),
            .I(N__44716));
    Odrv4 I__10354 (
            .O(N__44716),
            .I(DMActrl_BeLeC1));
    InMux I__10353 (
            .O(N__44713),
            .I(N__44710));
    LocalMux I__10352 (
            .O(N__44710),
            .I(N__44707));
    Odrv12 I__10351 (
            .O(N__44707),
            .I(PIOq_9));
    CascadeMux I__10350 (
            .O(N__44704),
            .I(N__44701));
    InMux I__10349 (
            .O(N__44701),
            .I(N__44698));
    LocalMux I__10348 (
            .O(N__44698),
            .I(N__44695));
    Span4Mux_v I__10347 (
            .O(N__44695),
            .I(N__44692));
    Span4Mux_v I__10346 (
            .O(N__44692),
            .I(N__44688));
    InMux I__10345 (
            .O(N__44691),
            .I(N__44685));
    Span4Mux_h I__10344 (
            .O(N__44688),
            .I(N__44682));
    LocalMux I__10343 (
            .O(N__44685),
            .I(N__44679));
    Odrv4 I__10342 (
            .O(N__44682),
            .I(DMA_dev0_Tm_1));
    Odrv4 I__10341 (
            .O(N__44679),
            .I(DMA_dev0_Tm_1));
    InMux I__10340 (
            .O(N__44674),
            .I(N__44670));
    CascadeMux I__10339 (
            .O(N__44673),
            .I(N__44667));
    LocalMux I__10338 (
            .O(N__44670),
            .I(N__44664));
    InMux I__10337 (
            .O(N__44667),
            .I(N__44661));
    Span4Mux_v I__10336 (
            .O(N__44664),
            .I(N__44658));
    LocalMux I__10335 (
            .O(N__44661),
            .I(N__44655));
    Span4Mux_h I__10334 (
            .O(N__44658),
            .I(N__44650));
    Span4Mux_h I__10333 (
            .O(N__44655),
            .I(N__44650));
    Odrv4 I__10332 (
            .O(N__44650),
            .I(PIO_dport1_T1_1));
    InMux I__10331 (
            .O(N__44647),
            .I(N__44644));
    LocalMux I__10330 (
            .O(N__44644),
            .I(N__44641));
    Span4Mux_v I__10329 (
            .O(N__44641),
            .I(N__44638));
    Span4Mux_h I__10328 (
            .O(N__44638),
            .I(N__44635));
    Odrv4 I__10327 (
            .O(N__44635),
            .I(\u0.dat_o_0_0_2_1 ));
    InMux I__10326 (
            .O(N__44632),
            .I(N__44629));
    LocalMux I__10325 (
            .O(N__44629),
            .I(N__44626));
    Span4Mux_v I__10324 (
            .O(N__44626),
            .I(N__44623));
    Odrv4 I__10323 (
            .O(N__44623),
            .I(\u0.dat_o_0_0_3_1 ));
    CascadeMux I__10322 (
            .O(N__44620),
            .I(\u0.dat_o_0_0_0_1_cascade_ ));
    IoInMux I__10321 (
            .O(N__44617),
            .I(N__44614));
    LocalMux I__10320 (
            .O(N__44614),
            .I(N__44611));
    Span12Mux_s3_h I__10319 (
            .O(N__44611),
            .I(N__44608));
    Span12Mux_h I__10318 (
            .O(N__44608),
            .I(N__44605));
    Odrv12 I__10317 (
            .O(N__44605),
            .I(wb_dat_o_c_1));
    InMux I__10316 (
            .O(N__44602),
            .I(N__44599));
    LocalMux I__10315 (
            .O(N__44599),
            .I(N__44596));
    Span4Mux_v I__10314 (
            .O(N__44596),
            .I(N__44593));
    Span4Mux_h I__10313 (
            .O(N__44593),
            .I(N__44590));
    Odrv4 I__10312 (
            .O(N__44590),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNISE4NZ0Z_1 ));
    InMux I__10311 (
            .O(N__44587),
            .I(N__44584));
    LocalMux I__10310 (
            .O(N__44584),
            .I(N__44581));
    Span4Mux_h I__10309 (
            .O(N__44581),
            .I(N__44578));
    Span4Mux_v I__10308 (
            .O(N__44578),
            .I(N__44575));
    Odrv4 I__10307 (
            .O(N__44575),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIOUBMZ0Z_1 ));
    InMux I__10306 (
            .O(N__44572),
            .I(N__44567));
    InMux I__10305 (
            .O(N__44571),
            .I(N__44562));
    InMux I__10304 (
            .O(N__44570),
            .I(N__44562));
    LocalMux I__10303 (
            .O(N__44567),
            .I(N__44559));
    LocalMux I__10302 (
            .O(N__44562),
            .I(N__44556));
    Span4Mux_v I__10301 (
            .O(N__44559),
            .I(N__44553));
    Span4Mux_v I__10300 (
            .O(N__44556),
            .I(N__44550));
    Sp12to4 I__10299 (
            .O(N__44553),
            .I(N__44545));
    Sp12to4 I__10298 (
            .O(N__44550),
            .I(N__44545));
    Span12Mux_h I__10297 (
            .O(N__44545),
            .I(N__44542));
    Span12Mux_v I__10296 (
            .O(N__44542),
            .I(N__44539));
    Span12Mux_h I__10295 (
            .O(N__44539),
            .I(N__44536));
    Odrv12 I__10294 (
            .O(N__44536),
            .I(dd_pad_i_c_1));
    InMux I__10293 (
            .O(N__44533),
            .I(N__44530));
    LocalMux I__10292 (
            .O(N__44530),
            .I(N__44527));
    Span12Mux_v I__10291 (
            .O(N__44527),
            .I(N__44524));
    Odrv12 I__10290 (
            .O(N__44524),
            .I(\u0.N_1736 ));
    InMux I__10289 (
            .O(N__44521),
            .I(N__44518));
    LocalMux I__10288 (
            .O(N__44518),
            .I(N__44515));
    Span12Mux_s9_v I__10287 (
            .O(N__44515),
            .I(N__44512));
    Span12Mux_h I__10286 (
            .O(N__44512),
            .I(N__44509));
    Odrv12 I__10285 (
            .O(N__44509),
            .I(\u0.dat_o_0_0_6_8 ));
    CascadeMux I__10284 (
            .O(N__44506),
            .I(\u0.dat_o_0_0_2_8_cascade_ ));
    IoInMux I__10283 (
            .O(N__44503),
            .I(N__44500));
    LocalMux I__10282 (
            .O(N__44500),
            .I(N__44497));
    IoSpan4Mux I__10281 (
            .O(N__44497),
            .I(N__44494));
    Span4Mux_s1_h I__10280 (
            .O(N__44494),
            .I(N__44491));
    Sp12to4 I__10279 (
            .O(N__44491),
            .I(N__44488));
    Span12Mux_h I__10278 (
            .O(N__44488),
            .I(N__44485));
    Odrv12 I__10277 (
            .O(N__44485),
            .I(wb_dat_o_c_8));
    InMux I__10276 (
            .O(N__44482),
            .I(N__44477));
    InMux I__10275 (
            .O(N__44481),
            .I(N__44472));
    InMux I__10274 (
            .O(N__44480),
            .I(N__44472));
    LocalMux I__10273 (
            .O(N__44477),
            .I(N__44469));
    LocalMux I__10272 (
            .O(N__44472),
            .I(N__44466));
    Span12Mux_h I__10271 (
            .O(N__44469),
            .I(N__44461));
    Span12Mux_s8_v I__10270 (
            .O(N__44466),
            .I(N__44461));
    Span12Mux_v I__10269 (
            .O(N__44461),
            .I(N__44458));
    Span12Mux_h I__10268 (
            .O(N__44458),
            .I(N__44455));
    Odrv12 I__10267 (
            .O(N__44455),
            .I(dd_pad_i_c_8));
    InMux I__10266 (
            .O(N__44452),
            .I(N__44449));
    LocalMux I__10265 (
            .O(N__44449),
            .I(PIOq_8));
    InMux I__10264 (
            .O(N__44446),
            .I(N__44443));
    LocalMux I__10263 (
            .O(N__44443),
            .I(N__44440));
    Odrv12 I__10262 (
            .O(N__44440),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI6DCMZ0Z_8 ));
    InMux I__10261 (
            .O(N__44437),
            .I(N__44434));
    LocalMux I__10260 (
            .O(N__44434),
            .I(N__44431));
    Span4Mux_v I__10259 (
            .O(N__44431),
            .I(N__44428));
    Span4Mux_v I__10258 (
            .O(N__44428),
            .I(N__44425));
    Span4Mux_h I__10257 (
            .O(N__44425),
            .I(N__44422));
    Odrv4 I__10256 (
            .O(N__44422),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIAT4NZ0Z_8 ));
    CascadeMux I__10255 (
            .O(N__44419),
            .I(\u0.dat_o_i_i_a2_0_0_29_cascade_ ));
    InMux I__10254 (
            .O(N__44416),
            .I(N__44412));
    CascadeMux I__10253 (
            .O(N__44415),
            .I(N__44409));
    LocalMux I__10252 (
            .O(N__44412),
            .I(N__44406));
    InMux I__10251 (
            .O(N__44409),
            .I(N__44403));
    Span4Mux_v I__10250 (
            .O(N__44406),
            .I(N__44400));
    LocalMux I__10249 (
            .O(N__44403),
            .I(N__44397));
    Span4Mux_h I__10248 (
            .O(N__44400),
            .I(N__44394));
    Span4Mux_v I__10247 (
            .O(N__44397),
            .I(N__44391));
    Odrv4 I__10246 (
            .O(N__44394),
            .I(PIO_dport1_Teoc_5));
    Odrv4 I__10245 (
            .O(N__44391),
            .I(PIO_dport1_Teoc_5));
    InMux I__10244 (
            .O(N__44386),
            .I(N__44383));
    LocalMux I__10243 (
            .O(N__44383),
            .I(N__44380));
    Span4Mux_v I__10242 (
            .O(N__44380),
            .I(N__44377));
    Span4Mux_v I__10241 (
            .O(N__44377),
            .I(N__44374));
    Odrv4 I__10240 (
            .O(N__44374),
            .I(\u0.N_1696 ));
    InMux I__10239 (
            .O(N__44371),
            .I(N__44368));
    LocalMux I__10238 (
            .O(N__44368),
            .I(\u0.dat_o_i_i_4_29 ));
    CascadeMux I__10237 (
            .O(N__44365),
            .I(\u0.dat_o_i_i_2_29_cascade_ ));
    IoInMux I__10236 (
            .O(N__44362),
            .I(N__44359));
    LocalMux I__10235 (
            .O(N__44359),
            .I(N__44356));
    IoSpan4Mux I__10234 (
            .O(N__44356),
            .I(N__44353));
    Span4Mux_s0_v I__10233 (
            .O(N__44353),
            .I(N__44350));
    Sp12to4 I__10232 (
            .O(N__44350),
            .I(N__44347));
    Span12Mux_s11_v I__10231 (
            .O(N__44347),
            .I(N__44344));
    Odrv12 I__10230 (
            .O(N__44344),
            .I(N_273));
    InMux I__10229 (
            .O(N__44341),
            .I(N__44338));
    LocalMux I__10228 (
            .O(N__44338),
            .I(N__44334));
    InMux I__10227 (
            .O(N__44337),
            .I(N__44331));
    Span4Mux_v I__10226 (
            .O(N__44334),
            .I(N__44328));
    LocalMux I__10225 (
            .O(N__44331),
            .I(N__44325));
    Sp12to4 I__10224 (
            .O(N__44328),
            .I(N__44322));
    Span4Mux_v I__10223 (
            .O(N__44325),
            .I(N__44319));
    Span12Mux_h I__10222 (
            .O(N__44322),
            .I(N__44316));
    Span4Mux_h I__10221 (
            .O(N__44319),
            .I(N__44313));
    Odrv12 I__10220 (
            .O(N__44316),
            .I(DMA_dev1_Teoc_2));
    Odrv4 I__10219 (
            .O(N__44313),
            .I(DMA_dev1_Teoc_2));
    CascadeMux I__10218 (
            .O(N__44308),
            .I(\u0.N_1675_cascade_ ));
    InMux I__10217 (
            .O(N__44305),
            .I(N__44302));
    LocalMux I__10216 (
            .O(N__44302),
            .I(N__44298));
    InMux I__10215 (
            .O(N__44301),
            .I(N__44295));
    Span4Mux_v I__10214 (
            .O(N__44298),
            .I(N__44292));
    LocalMux I__10213 (
            .O(N__44295),
            .I(N__44289));
    Odrv4 I__10212 (
            .O(N__44292),
            .I(PIO_dport0_Teoc_2));
    Odrv12 I__10211 (
            .O(N__44289),
            .I(PIO_dport0_Teoc_2));
    CascadeMux I__10210 (
            .O(N__44284),
            .I(\u0.dat_o_i_i_4_26_cascade_ ));
    InMux I__10209 (
            .O(N__44281),
            .I(N__44277));
    InMux I__10208 (
            .O(N__44280),
            .I(N__44274));
    LocalMux I__10207 (
            .O(N__44277),
            .I(N__44271));
    LocalMux I__10206 (
            .O(N__44274),
            .I(N__44268));
    Span4Mux_v I__10205 (
            .O(N__44271),
            .I(N__44263));
    Span4Mux_h I__10204 (
            .O(N__44268),
            .I(N__44263));
    Odrv4 I__10203 (
            .O(N__44263),
            .I(PIO_dport1_Teoc_2));
    IoInMux I__10202 (
            .O(N__44260),
            .I(N__44257));
    LocalMux I__10201 (
            .O(N__44257),
            .I(N__44254));
    Span4Mux_s2_v I__10200 (
            .O(N__44254),
            .I(N__44251));
    Span4Mux_h I__10199 (
            .O(N__44251),
            .I(N__44248));
    Span4Mux_v I__10198 (
            .O(N__44248),
            .I(N__44245));
    Span4Mux_v I__10197 (
            .O(N__44245),
            .I(N__44242));
    Odrv4 I__10196 (
            .O(N__44242),
            .I(N_267));
    InMux I__10195 (
            .O(N__44239),
            .I(N__44234));
    InMux I__10194 (
            .O(N__44238),
            .I(N__44231));
    InMux I__10193 (
            .O(N__44237),
            .I(N__44227));
    LocalMux I__10192 (
            .O(N__44234),
            .I(N__44222));
    LocalMux I__10191 (
            .O(N__44231),
            .I(N__44222));
    InMux I__10190 (
            .O(N__44230),
            .I(N__44219));
    LocalMux I__10189 (
            .O(N__44227),
            .I(N__44215));
    Span4Mux_v I__10188 (
            .O(N__44222),
            .I(N__44210));
    LocalMux I__10187 (
            .O(N__44219),
            .I(N__44210));
    InMux I__10186 (
            .O(N__44218),
            .I(N__44207));
    Span4Mux_v I__10185 (
            .O(N__44215),
            .I(N__44202));
    Span4Mux_h I__10184 (
            .O(N__44210),
            .I(N__44199));
    LocalMux I__10183 (
            .O(N__44207),
            .I(N__44196));
    InMux I__10182 (
            .O(N__44206),
            .I(N__44193));
    InMux I__10181 (
            .O(N__44205),
            .I(N__44190));
    Span4Mux_h I__10180 (
            .O(N__44202),
            .I(N__44187));
    Span4Mux_v I__10179 (
            .O(N__44199),
            .I(N__44182));
    Span4Mux_v I__10178 (
            .O(N__44196),
            .I(N__44182));
    LocalMux I__10177 (
            .O(N__44193),
            .I(N__44179));
    LocalMux I__10176 (
            .O(N__44190),
            .I(N__44176));
    Sp12to4 I__10175 (
            .O(N__44187),
            .I(N__44171));
    Sp12to4 I__10174 (
            .O(N__44182),
            .I(N__44171));
    Span4Mux_h I__10173 (
            .O(N__44179),
            .I(N__44166));
    Span4Mux_v I__10172 (
            .O(N__44176),
            .I(N__44166));
    Odrv12 I__10171 (
            .O(N__44171),
            .I(wb_dat_i_c_26));
    Odrv4 I__10170 (
            .O(N__44166),
            .I(wb_dat_i_c_26));
    InMux I__10169 (
            .O(N__44161),
            .I(N__44158));
    LocalMux I__10168 (
            .O(N__44158),
            .I(N__44155));
    Span12Mux_h I__10167 (
            .O(N__44155),
            .I(N__44152));
    Odrv12 I__10166 (
            .O(N__44152),
            .I(DMAq_26));
    CascadeMux I__10165 (
            .O(N__44149),
            .I(N__44146));
    InMux I__10164 (
            .O(N__44146),
            .I(N__44143));
    LocalMux I__10163 (
            .O(N__44143),
            .I(N__44140));
    Span12Mux_h I__10162 (
            .O(N__44140),
            .I(N__44136));
    InMux I__10161 (
            .O(N__44139),
            .I(N__44133));
    Odrv12 I__10160 (
            .O(N__44136),
            .I(DMA_dev0_Teoc_2));
    LocalMux I__10159 (
            .O(N__44133),
            .I(DMA_dev0_Teoc_2));
    InMux I__10158 (
            .O(N__44128),
            .I(N__44125));
    LocalMux I__10157 (
            .O(N__44125),
            .I(\u0.dat_o_i_i_0_26 ));
    InMux I__10156 (
            .O(N__44122),
            .I(N__44118));
    InMux I__10155 (
            .O(N__44121),
            .I(N__44115));
    LocalMux I__10154 (
            .O(N__44118),
            .I(N__44112));
    LocalMux I__10153 (
            .O(N__44115),
            .I(N__44109));
    Span4Mux_h I__10152 (
            .O(N__44112),
            .I(N__44106));
    Span12Mux_h I__10151 (
            .O(N__44109),
            .I(N__44103));
    Span4Mux_h I__10150 (
            .O(N__44106),
            .I(N__44100));
    Odrv12 I__10149 (
            .O(N__44103),
            .I(DMA_dev0_Td_6));
    Odrv4 I__10148 (
            .O(N__44100),
            .I(DMA_dev0_Td_6));
    CascadeMux I__10147 (
            .O(N__44095),
            .I(N__44091));
    InMux I__10146 (
            .O(N__44094),
            .I(N__44088));
    InMux I__10145 (
            .O(N__44091),
            .I(N__44085));
    LocalMux I__10144 (
            .O(N__44088),
            .I(N__44082));
    LocalMux I__10143 (
            .O(N__44085),
            .I(N__44079));
    Span4Mux_h I__10142 (
            .O(N__44082),
            .I(N__44076));
    Odrv12 I__10141 (
            .O(N__44079),
            .I(PIO_dport1_T2_6));
    Odrv4 I__10140 (
            .O(N__44076),
            .I(PIO_dport1_T2_6));
    InMux I__10139 (
            .O(N__44071),
            .I(N__44068));
    LocalMux I__10138 (
            .O(N__44068),
            .I(\u0.dat_o_0_0_0_14 ));
    InMux I__10137 (
            .O(N__44065),
            .I(N__44062));
    LocalMux I__10136 (
            .O(N__44062),
            .I(N__44055));
    InMux I__10135 (
            .O(N__44061),
            .I(N__44052));
    InMux I__10134 (
            .O(N__44060),
            .I(N__44049));
    InMux I__10133 (
            .O(N__44059),
            .I(N__44046));
    InMux I__10132 (
            .O(N__44058),
            .I(N__44043));
    Span4Mux_h I__10131 (
            .O(N__44055),
            .I(N__44036));
    LocalMux I__10130 (
            .O(N__44052),
            .I(N__44036));
    LocalMux I__10129 (
            .O(N__44049),
            .I(N__44036));
    LocalMux I__10128 (
            .O(N__44046),
            .I(N__44032));
    LocalMux I__10127 (
            .O(N__44043),
            .I(N__44029));
    Span4Mux_h I__10126 (
            .O(N__44036),
            .I(N__44025));
    InMux I__10125 (
            .O(N__44035),
            .I(N__44022));
    Span4Mux_v I__10124 (
            .O(N__44032),
            .I(N__44019));
    Span4Mux_v I__10123 (
            .O(N__44029),
            .I(N__44016));
    InMux I__10122 (
            .O(N__44028),
            .I(N__44012));
    Span4Mux_h I__10121 (
            .O(N__44025),
            .I(N__44007));
    LocalMux I__10120 (
            .O(N__44022),
            .I(N__44007));
    Span4Mux_v I__10119 (
            .O(N__44019),
            .I(N__44003));
    Span4Mux_v I__10118 (
            .O(N__44016),
            .I(N__44000));
    InMux I__10117 (
            .O(N__44015),
            .I(N__43997));
    LocalMux I__10116 (
            .O(N__44012),
            .I(N__43994));
    Span4Mux_h I__10115 (
            .O(N__44007),
            .I(N__43991));
    InMux I__10114 (
            .O(N__44006),
            .I(N__43988));
    Sp12to4 I__10113 (
            .O(N__44003),
            .I(N__43983));
    Sp12to4 I__10112 (
            .O(N__44000),
            .I(N__43983));
    LocalMux I__10111 (
            .O(N__43997),
            .I(N__43980));
    Span4Mux_v I__10110 (
            .O(N__43994),
            .I(N__43977));
    Span4Mux_v I__10109 (
            .O(N__43991),
            .I(N__43972));
    LocalMux I__10108 (
            .O(N__43988),
            .I(N__43972));
    Span12Mux_h I__10107 (
            .O(N__43983),
            .I(N__43967));
    Span12Mux_v I__10106 (
            .O(N__43980),
            .I(N__43967));
    Span4Mux_h I__10105 (
            .O(N__43977),
            .I(N__43964));
    Span4Mux_v I__10104 (
            .O(N__43972),
            .I(N__43961));
    Odrv12 I__10103 (
            .O(N__43967),
            .I(wb_dat_i_c_14));
    Odrv4 I__10102 (
            .O(N__43964),
            .I(wb_dat_i_c_14));
    Odrv4 I__10101 (
            .O(N__43961),
            .I(wb_dat_i_c_14));
    InMux I__10100 (
            .O(N__43954),
            .I(N__43951));
    LocalMux I__10099 (
            .O(N__43951),
            .I(\u0.CtrlRegZ0Z_14 ));
    InMux I__10098 (
            .O(N__43948),
            .I(N__43945));
    LocalMux I__10097 (
            .O(N__43945),
            .I(N__43941));
    InMux I__10096 (
            .O(N__43944),
            .I(N__43938));
    Odrv12 I__10095 (
            .O(N__43941),
            .I(PIO_cmdport_T2_6));
    LocalMux I__10094 (
            .O(N__43938),
            .I(PIO_cmdport_T2_6));
    InMux I__10093 (
            .O(N__43933),
            .I(N__43930));
    LocalMux I__10092 (
            .O(N__43930),
            .I(\u0.dat_o_0_0_2_14 ));
    InMux I__10091 (
            .O(N__43927),
            .I(N__43924));
    LocalMux I__10090 (
            .O(N__43924),
            .I(N__43921));
    Span4Mux_v I__10089 (
            .O(N__43921),
            .I(N__43918));
    Span4Mux_h I__10088 (
            .O(N__43918),
            .I(N__43915));
    Odrv4 I__10087 (
            .O(N__43915),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI7SA71Z0Z_14 ));
    InMux I__10086 (
            .O(N__43912),
            .I(N__43909));
    LocalMux I__10085 (
            .O(N__43909),
            .I(N__43906));
    Span4Mux_h I__10084 (
            .O(N__43906),
            .I(N__43903));
    Span4Mux_v I__10083 (
            .O(N__43903),
            .I(N__43900));
    Span4Mux_v I__10082 (
            .O(N__43900),
            .I(N__43897));
    Odrv4 I__10081 (
            .O(N__43897),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIMCDM1Z0Z_2 ));
    InMux I__10080 (
            .O(N__43894),
            .I(N__43891));
    LocalMux I__10079 (
            .O(N__43891),
            .I(DMAq_14));
    InMux I__10078 (
            .O(N__43888),
            .I(N__43884));
    CascadeMux I__10077 (
            .O(N__43887),
            .I(N__43881));
    LocalMux I__10076 (
            .O(N__43884),
            .I(N__43878));
    InMux I__10075 (
            .O(N__43881),
            .I(N__43875));
    Span4Mux_h I__10074 (
            .O(N__43878),
            .I(N__43872));
    LocalMux I__10073 (
            .O(N__43875),
            .I(N__43869));
    Span4Mux_h I__10072 (
            .O(N__43872),
            .I(N__43866));
    Span4Mux_v I__10071 (
            .O(N__43869),
            .I(N__43863));
    Span4Mux_h I__10070 (
            .O(N__43866),
            .I(N__43860));
    Odrv4 I__10069 (
            .O(N__43863),
            .I(DMA_dev1_Teoc_5));
    Odrv4 I__10068 (
            .O(N__43860),
            .I(DMA_dev1_Teoc_5));
    CascadeMux I__10067 (
            .O(N__43855),
            .I(N__43851));
    InMux I__10066 (
            .O(N__43854),
            .I(N__43848));
    InMux I__10065 (
            .O(N__43851),
            .I(N__43845));
    LocalMux I__10064 (
            .O(N__43848),
            .I(N__43842));
    LocalMux I__10063 (
            .O(N__43845),
            .I(N__43839));
    Span12Mux_v I__10062 (
            .O(N__43842),
            .I(N__43836));
    Span4Mux_v I__10061 (
            .O(N__43839),
            .I(N__43833));
    Span12Mux_h I__10060 (
            .O(N__43836),
            .I(N__43830));
    Odrv4 I__10059 (
            .O(N__43833),
            .I(DMA_dev0_Teoc_5));
    Odrv12 I__10058 (
            .O(N__43830),
            .I(DMA_dev0_Teoc_5));
    InMux I__10057 (
            .O(N__43825),
            .I(N__43822));
    LocalMux I__10056 (
            .O(N__43822),
            .I(\u0.dat_o_i_i_0_29 ));
    InMux I__10055 (
            .O(N__43819),
            .I(N__43815));
    InMux I__10054 (
            .O(N__43818),
            .I(N__43812));
    LocalMux I__10053 (
            .O(N__43815),
            .I(N__43809));
    LocalMux I__10052 (
            .O(N__43812),
            .I(N__43806));
    Span4Mux_h I__10051 (
            .O(N__43809),
            .I(N__43803));
    Odrv12 I__10050 (
            .O(N__43806),
            .I(PIO_dport0_Teoc_5));
    Odrv4 I__10049 (
            .O(N__43803),
            .I(PIO_dport0_Teoc_5));
    IoInMux I__10048 (
            .O(N__43798),
            .I(N__43795));
    LocalMux I__10047 (
            .O(N__43795),
            .I(N__43792));
    IoSpan4Mux I__10046 (
            .O(N__43792),
            .I(N__43789));
    Span4Mux_s3_v I__10045 (
            .O(N__43789),
            .I(N__43786));
    Sp12to4 I__10044 (
            .O(N__43786),
            .I(N__43783));
    Odrv12 I__10043 (
            .O(N__43783),
            .I(N_448));
    InMux I__10042 (
            .O(N__43780),
            .I(N__43776));
    InMux I__10041 (
            .O(N__43779),
            .I(N__43773));
    LocalMux I__10040 (
            .O(N__43776),
            .I(N__43768));
    LocalMux I__10039 (
            .O(N__43773),
            .I(N__43768));
    Odrv12 I__10038 (
            .O(N__43768),
            .I(PIO_dport1_T2_3));
    InMux I__10037 (
            .O(N__43765),
            .I(N__43762));
    LocalMux I__10036 (
            .O(N__43762),
            .I(N__43759));
    Span4Mux_v I__10035 (
            .O(N__43759),
            .I(N__43756));
    Span4Mux_h I__10034 (
            .O(N__43756),
            .I(N__43753));
    Span4Mux_h I__10033 (
            .O(N__43753),
            .I(N__43749));
    InMux I__10032 (
            .O(N__43752),
            .I(N__43746));
    Odrv4 I__10031 (
            .O(N__43749),
            .I(DMA_dev0_Td_3));
    LocalMux I__10030 (
            .O(N__43746),
            .I(DMA_dev0_Td_3));
    CascadeMux I__10029 (
            .O(N__43741),
            .I(\u0.dat_o_0_0_0_11_cascade_ ));
    InMux I__10028 (
            .O(N__43738),
            .I(N__43735));
    LocalMux I__10027 (
            .O(N__43735),
            .I(N__43732));
    Span4Mux_h I__10026 (
            .O(N__43732),
            .I(N__43729));
    Span4Mux_h I__10025 (
            .O(N__43729),
            .I(N__43726));
    Odrv4 I__10024 (
            .O(N__43726),
            .I(\u0.dat_o_0_0_3_11 ));
    IoInMux I__10023 (
            .O(N__43723),
            .I(N__43720));
    LocalMux I__10022 (
            .O(N__43720),
            .I(N__43717));
    Span4Mux_s3_h I__10021 (
            .O(N__43717),
            .I(N__43714));
    Sp12to4 I__10020 (
            .O(N__43714),
            .I(N__43711));
    Span12Mux_v I__10019 (
            .O(N__43711),
            .I(N__43708));
    Span12Mux_h I__10018 (
            .O(N__43708),
            .I(N__43705));
    Odrv12 I__10017 (
            .O(N__43705),
            .I(wb_dat_o_c_11));
    InMux I__10016 (
            .O(N__43702),
            .I(N__43696));
    InMux I__10015 (
            .O(N__43701),
            .I(N__43693));
    InMux I__10014 (
            .O(N__43700),
            .I(N__43690));
    InMux I__10013 (
            .O(N__43699),
            .I(N__43687));
    LocalMux I__10012 (
            .O(N__43696),
            .I(N__43682));
    LocalMux I__10011 (
            .O(N__43693),
            .I(N__43682));
    LocalMux I__10010 (
            .O(N__43690),
            .I(N__43677));
    LocalMux I__10009 (
            .O(N__43687),
            .I(N__43677));
    Span4Mux_v I__10008 (
            .O(N__43682),
            .I(N__43673));
    Span4Mux_h I__10007 (
            .O(N__43677),
            .I(N__43668));
    InMux I__10006 (
            .O(N__43676),
            .I(N__43665));
    Span4Mux_h I__10005 (
            .O(N__43673),
            .I(N__43662));
    InMux I__10004 (
            .O(N__43672),
            .I(N__43659));
    InMux I__10003 (
            .O(N__43671),
            .I(N__43656));
    Span4Mux_v I__10002 (
            .O(N__43668),
            .I(N__43653));
    LocalMux I__10001 (
            .O(N__43665),
            .I(N__43650));
    Span4Mux_v I__10000 (
            .O(N__43662),
            .I(N__43643));
    LocalMux I__9999 (
            .O(N__43659),
            .I(N__43643));
    LocalMux I__9998 (
            .O(N__43656),
            .I(N__43643));
    Span4Mux_v I__9997 (
            .O(N__43653),
            .I(N__43640));
    Span4Mux_v I__9996 (
            .O(N__43650),
            .I(N__43634));
    Span4Mux_h I__9995 (
            .O(N__43643),
            .I(N__43634));
    Span4Mux_h I__9994 (
            .O(N__43640),
            .I(N__43631));
    InMux I__9993 (
            .O(N__43639),
            .I(N__43628));
    Span4Mux_v I__9992 (
            .O(N__43634),
            .I(N__43624));
    Span4Mux_h I__9991 (
            .O(N__43631),
            .I(N__43619));
    LocalMux I__9990 (
            .O(N__43628),
            .I(N__43619));
    InMux I__9989 (
            .O(N__43627),
            .I(N__43616));
    Span4Mux_v I__9988 (
            .O(N__43624),
            .I(N__43613));
    Span4Mux_h I__9987 (
            .O(N__43619),
            .I(N__43610));
    LocalMux I__9986 (
            .O(N__43616),
            .I(N__43607));
    Span4Mux_v I__9985 (
            .O(N__43613),
            .I(N__43604));
    Span4Mux_v I__9984 (
            .O(N__43610),
            .I(N__43599));
    Span4Mux_h I__9983 (
            .O(N__43607),
            .I(N__43599));
    IoSpan4Mux I__9982 (
            .O(N__43604),
            .I(N__43594));
    IoSpan4Mux I__9981 (
            .O(N__43599),
            .I(N__43594));
    Odrv4 I__9980 (
            .O(N__43594),
            .I(wb_dat_i_c_11));
    InMux I__9979 (
            .O(N__43591),
            .I(N__43588));
    LocalMux I__9978 (
            .O(N__43588),
            .I(\u0.CtrlRegZ0Z_11 ));
    InMux I__9977 (
            .O(N__43585),
            .I(N__43581));
    InMux I__9976 (
            .O(N__43584),
            .I(N__43578));
    LocalMux I__9975 (
            .O(N__43581),
            .I(N__43575));
    LocalMux I__9974 (
            .O(N__43578),
            .I(N__43572));
    Odrv12 I__9973 (
            .O(N__43575),
            .I(PIO_cmdport_T2_3));
    Odrv12 I__9972 (
            .O(N__43572),
            .I(PIO_cmdport_T2_3));
    InMux I__9971 (
            .O(N__43567),
            .I(N__43564));
    LocalMux I__9970 (
            .O(N__43564),
            .I(\u0.dat_o_0_0_2_11 ));
    CascadeMux I__9969 (
            .O(N__43561),
            .I(N__43557));
    InMux I__9968 (
            .O(N__43560),
            .I(N__43554));
    InMux I__9967 (
            .O(N__43557),
            .I(N__43551));
    LocalMux I__9966 (
            .O(N__43554),
            .I(N__43548));
    LocalMux I__9965 (
            .O(N__43551),
            .I(N__43543));
    Span12Mux_v I__9964 (
            .O(N__43548),
            .I(N__43543));
    Odrv12 I__9963 (
            .O(N__43543),
            .I(DMA_dev1_Td_2));
    InMux I__9962 (
            .O(N__43540),
            .I(N__43537));
    LocalMux I__9961 (
            .O(N__43537),
            .I(N__43533));
    InMux I__9960 (
            .O(N__43536),
            .I(N__43530));
    Span4Mux_v I__9959 (
            .O(N__43533),
            .I(N__43527));
    LocalMux I__9958 (
            .O(N__43530),
            .I(N__43524));
    Odrv4 I__9957 (
            .O(N__43527),
            .I(PIO_dport1_T2_2));
    Odrv4 I__9956 (
            .O(N__43524),
            .I(PIO_dport1_T2_2));
    InMux I__9955 (
            .O(N__43519),
            .I(N__43516));
    LocalMux I__9954 (
            .O(N__43516),
            .I(N__43513));
    Odrv4 I__9953 (
            .O(N__43513),
            .I(\u0.dat_o_i_i_0_10 ));
    CascadeMux I__9952 (
            .O(N__43510),
            .I(N__43506));
    InMux I__9951 (
            .O(N__43509),
            .I(N__43503));
    InMux I__9950 (
            .O(N__43506),
            .I(N__43500));
    LocalMux I__9949 (
            .O(N__43503),
            .I(N__43497));
    LocalMux I__9948 (
            .O(N__43500),
            .I(N__43494));
    Span4Mux_h I__9947 (
            .O(N__43497),
            .I(N__43491));
    Odrv12 I__9946 (
            .O(N__43494),
            .I(PIO_dport0_T2_6));
    Odrv4 I__9945 (
            .O(N__43491),
            .I(PIO_dport0_T2_6));
    InMux I__9944 (
            .O(N__43486),
            .I(N__43482));
    InMux I__9943 (
            .O(N__43485),
            .I(N__43479));
    LocalMux I__9942 (
            .O(N__43482),
            .I(N__43476));
    LocalMux I__9941 (
            .O(N__43479),
            .I(N__43473));
    Odrv12 I__9940 (
            .O(N__43476),
            .I(DMA_dev1_Td_6));
    Odrv4 I__9939 (
            .O(N__43473),
            .I(DMA_dev1_Td_6));
    CascadeMux I__9938 (
            .O(N__43468),
            .I(\u0.dat_o_0_0_3_14_cascade_ ));
    IoInMux I__9937 (
            .O(N__43465),
            .I(N__43462));
    LocalMux I__9936 (
            .O(N__43462),
            .I(N__43459));
    Span12Mux_s3_h I__9935 (
            .O(N__43459),
            .I(N__43456));
    Span12Mux_h I__9934 (
            .O(N__43456),
            .I(N__43453));
    Odrv12 I__9933 (
            .O(N__43453),
            .I(wb_dat_o_c_14));
    InMux I__9932 (
            .O(N__43450),
            .I(N__43447));
    LocalMux I__9931 (
            .O(N__43447),
            .I(N__43444));
    Span4Mux_v I__9930 (
            .O(N__43444),
            .I(N__43441));
    Span4Mux_h I__9929 (
            .O(N__43441),
            .I(N__43438));
    Sp12to4 I__9928 (
            .O(N__43438),
            .I(N__43435));
    Span12Mux_h I__9927 (
            .O(N__43435),
            .I(N__43432));
    Odrv12 I__9926 (
            .O(N__43432),
            .I(PIOq_14));
    InMux I__9925 (
            .O(N__43429),
            .I(N__43426));
    LocalMux I__9924 (
            .O(N__43426),
            .I(\u0.dat_o_0_0_1Z0Z_14 ));
    InMux I__9923 (
            .O(N__43423),
            .I(N__43420));
    LocalMux I__9922 (
            .O(N__43420),
            .I(N__43417));
    Span4Mux_v I__9921 (
            .O(N__43417),
            .I(N__43414));
    Span4Mux_v I__9920 (
            .O(N__43414),
            .I(N__43411));
    Odrv4 I__9919 (
            .O(N__43411),
            .I(\u0.dat_o_0_0_6_0 ));
    CascadeMux I__9918 (
            .O(N__43408),
            .I(\u0.N_1938_cascade_ ));
    IoInMux I__9917 (
            .O(N__43405),
            .I(N__43402));
    LocalMux I__9916 (
            .O(N__43402),
            .I(N__43399));
    Span4Mux_s3_v I__9915 (
            .O(N__43399),
            .I(N__43396));
    Sp12to4 I__9914 (
            .O(N__43396),
            .I(N__43393));
    Span12Mux_h I__9913 (
            .O(N__43393),
            .I(N__43390));
    Odrv12 I__9912 (
            .O(N__43390),
            .I(wb_dat_o_c_0));
    InMux I__9911 (
            .O(N__43387),
            .I(N__43384));
    LocalMux I__9910 (
            .O(N__43384),
            .I(N__43381));
    Span4Mux_v I__9909 (
            .O(N__43381),
            .I(N__43376));
    InMux I__9908 (
            .O(N__43380),
            .I(N__43371));
    InMux I__9907 (
            .O(N__43379),
            .I(N__43371));
    Span4Mux_v I__9906 (
            .O(N__43376),
            .I(N__43368));
    LocalMux I__9905 (
            .O(N__43371),
            .I(N__43365));
    Sp12to4 I__9904 (
            .O(N__43368),
            .I(N__43362));
    Span12Mux_s9_v I__9903 (
            .O(N__43365),
            .I(N__43359));
    Span12Mux_h I__9902 (
            .O(N__43362),
            .I(N__43356));
    Span12Mux_h I__9901 (
            .O(N__43359),
            .I(N__43353));
    Span12Mux_v I__9900 (
            .O(N__43356),
            .I(N__43350));
    Span12Mux_v I__9899 (
            .O(N__43353),
            .I(N__43347));
    Odrv12 I__9898 (
            .O(N__43350),
            .I(dd_pad_i_c_0));
    Odrv12 I__9897 (
            .O(N__43347),
            .I(dd_pad_i_c_0));
    InMux I__9896 (
            .O(N__43342),
            .I(N__43339));
    LocalMux I__9895 (
            .O(N__43339),
            .I(N__43336));
    Span4Mux_h I__9894 (
            .O(N__43336),
            .I(N__43333));
    Odrv4 I__9893 (
            .O(N__43333),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIMSBMZ0Z_0 ));
    InMux I__9892 (
            .O(N__43330),
            .I(N__43327));
    LocalMux I__9891 (
            .O(N__43327),
            .I(N__43324));
    Span4Mux_v I__9890 (
            .O(N__43324),
            .I(N__43321));
    Span4Mux_h I__9889 (
            .O(N__43321),
            .I(N__43318));
    Odrv4 I__9888 (
            .O(N__43318),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIQC4NZ0Z_0 ));
    CascadeMux I__9887 (
            .O(N__43315),
            .I(iQ_RNI2KNK1_2_cascade_));
    InMux I__9886 (
            .O(N__43312),
            .I(N__43309));
    LocalMux I__9885 (
            .O(N__43309),
            .I(\u0.N_1937 ));
    InMux I__9884 (
            .O(N__43306),
            .I(N__43303));
    LocalMux I__9883 (
            .O(N__43303),
            .I(PIOq_0));
    InMux I__9882 (
            .O(N__43300),
            .I(N__43297));
    LocalMux I__9881 (
            .O(N__43297),
            .I(N__43294));
    Span4Mux_v I__9880 (
            .O(N__43294),
            .I(N__43291));
    Span4Mux_h I__9879 (
            .O(N__43291),
            .I(N__43287));
    InMux I__9878 (
            .O(N__43290),
            .I(N__43282));
    Span4Mux_h I__9877 (
            .O(N__43287),
            .I(N__43279));
    InMux I__9876 (
            .O(N__43286),
            .I(N__43276));
    InMux I__9875 (
            .O(N__43285),
            .I(N__43273));
    LocalMux I__9874 (
            .O(N__43282),
            .I(N__43270));
    Odrv4 I__9873 (
            .O(N__43279),
            .I(IDEctrl_rst));
    LocalMux I__9872 (
            .O(N__43276),
            .I(IDEctrl_rst));
    LocalMux I__9871 (
            .O(N__43273),
            .I(IDEctrl_rst));
    Odrv4 I__9870 (
            .O(N__43270),
            .I(IDEctrl_rst));
    InMux I__9869 (
            .O(N__43261),
            .I(N__43258));
    LocalMux I__9868 (
            .O(N__43258),
            .I(\u0.dat_o_0_0_2_0 ));
    InMux I__9867 (
            .O(N__43255),
            .I(N__43252));
    LocalMux I__9866 (
            .O(N__43252),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_0 ));
    InMux I__9865 (
            .O(N__43249),
            .I(N__43246));
    LocalMux I__9864 (
            .O(N__43246),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNIUSSNZ0Z_0 ));
    InMux I__9863 (
            .O(N__43243),
            .I(N__43240));
    LocalMux I__9862 (
            .O(N__43240),
            .I(mem_mem_ram6__RNI87OD1_0));
    CascadeMux I__9861 (
            .O(N__43237),
            .I(N__43233));
    CascadeMux I__9860 (
            .O(N__43236),
            .I(N__43226));
    InMux I__9859 (
            .O(N__43233),
            .I(N__43220));
    InMux I__9858 (
            .O(N__43232),
            .I(N__43220));
    InMux I__9857 (
            .O(N__43231),
            .I(N__43217));
    InMux I__9856 (
            .O(N__43230),
            .I(N__43212));
    InMux I__9855 (
            .O(N__43229),
            .I(N__43212));
    InMux I__9854 (
            .O(N__43226),
            .I(N__43207));
    InMux I__9853 (
            .O(N__43225),
            .I(N__43207));
    LocalMux I__9852 (
            .O(N__43220),
            .I(N__43199));
    LocalMux I__9851 (
            .O(N__43217),
            .I(N__43194));
    LocalMux I__9850 (
            .O(N__43212),
            .I(N__43194));
    LocalMux I__9849 (
            .O(N__43207),
            .I(N__43191));
    InMux I__9848 (
            .O(N__43206),
            .I(N__43186));
    InMux I__9847 (
            .O(N__43205),
            .I(N__43186));
    InMux I__9846 (
            .O(N__43204),
            .I(N__43183));
    InMux I__9845 (
            .O(N__43203),
            .I(N__43178));
    InMux I__9844 (
            .O(N__43202),
            .I(N__43178));
    Span4Mux_h I__9843 (
            .O(N__43199),
            .I(N__43173));
    Span12Mux_s6_v I__9842 (
            .O(N__43194),
            .I(N__43170));
    Span4Mux_h I__9841 (
            .O(N__43191),
            .I(N__43165));
    LocalMux I__9840 (
            .O(N__43186),
            .I(N__43165));
    LocalMux I__9839 (
            .O(N__43183),
            .I(N__43160));
    LocalMux I__9838 (
            .O(N__43178),
            .I(N__43160));
    InMux I__9837 (
            .O(N__43177),
            .I(N__43157));
    InMux I__9836 (
            .O(N__43176),
            .I(N__43154));
    Odrv4 I__9835 (
            .O(N__43173),
            .I(\u1.DMA_control.readDfw_11 ));
    Odrv12 I__9834 (
            .O(N__43170),
            .I(\u1.DMA_control.readDfw_11 ));
    Odrv4 I__9833 (
            .O(N__43165),
            .I(\u1.DMA_control.readDfw_11 ));
    Odrv4 I__9832 (
            .O(N__43160),
            .I(\u1.DMA_control.readDfw_11 ));
    LocalMux I__9831 (
            .O(N__43157),
            .I(\u1.DMA_control.readDfw_11 ));
    LocalMux I__9830 (
            .O(N__43154),
            .I(\u1.DMA_control.readDfw_11 ));
    CascadeMux I__9829 (
            .O(N__43141),
            .I(N__43131));
    InMux I__9828 (
            .O(N__43140),
            .I(N__43126));
    InMux I__9827 (
            .O(N__43139),
            .I(N__43126));
    InMux I__9826 (
            .O(N__43138),
            .I(N__43121));
    InMux I__9825 (
            .O(N__43137),
            .I(N__43121));
    CascadeMux I__9824 (
            .O(N__43136),
            .I(N__43118));
    InMux I__9823 (
            .O(N__43135),
            .I(N__43114));
    InMux I__9822 (
            .O(N__43134),
            .I(N__43109));
    InMux I__9821 (
            .O(N__43131),
            .I(N__43109));
    LocalMux I__9820 (
            .O(N__43126),
            .I(N__43103));
    LocalMux I__9819 (
            .O(N__43121),
            .I(N__43103));
    InMux I__9818 (
            .O(N__43118),
            .I(N__43098));
    InMux I__9817 (
            .O(N__43117),
            .I(N__43098));
    LocalMux I__9816 (
            .O(N__43114),
            .I(N__43089));
    LocalMux I__9815 (
            .O(N__43109),
            .I(N__43089));
    InMux I__9814 (
            .O(N__43108),
            .I(N__43086));
    Span4Mux_v I__9813 (
            .O(N__43103),
            .I(N__43081));
    LocalMux I__9812 (
            .O(N__43098),
            .I(N__43081));
    InMux I__9811 (
            .O(N__43097),
            .I(N__43078));
    InMux I__9810 (
            .O(N__43096),
            .I(N__43075));
    CascadeMux I__9809 (
            .O(N__43095),
            .I(N__43071));
    InMux I__9808 (
            .O(N__43094),
            .I(N__43068));
    Span4Mux_v I__9807 (
            .O(N__43089),
            .I(N__43065));
    LocalMux I__9806 (
            .O(N__43086),
            .I(N__43056));
    Span4Mux_h I__9805 (
            .O(N__43081),
            .I(N__43056));
    LocalMux I__9804 (
            .O(N__43078),
            .I(N__43056));
    LocalMux I__9803 (
            .O(N__43075),
            .I(N__43056));
    InMux I__9802 (
            .O(N__43074),
            .I(N__43053));
    InMux I__9801 (
            .O(N__43071),
            .I(N__43050));
    LocalMux I__9800 (
            .O(N__43068),
            .I(\u1.DMA_control.readDlw_11 ));
    Odrv4 I__9799 (
            .O(N__43065),
            .I(\u1.DMA_control.readDlw_11 ));
    Odrv4 I__9798 (
            .O(N__43056),
            .I(\u1.DMA_control.readDlw_11 ));
    LocalMux I__9797 (
            .O(N__43053),
            .I(\u1.DMA_control.readDlw_11 ));
    LocalMux I__9796 (
            .O(N__43050),
            .I(\u1.DMA_control.readDlw_11 ));
    InMux I__9795 (
            .O(N__43039),
            .I(N__42997));
    InMux I__9794 (
            .O(N__43038),
            .I(N__42997));
    InMux I__9793 (
            .O(N__43037),
            .I(N__42997));
    InMux I__9792 (
            .O(N__43036),
            .I(N__42997));
    InMux I__9791 (
            .O(N__43035),
            .I(N__42988));
    InMux I__9790 (
            .O(N__43034),
            .I(N__42988));
    InMux I__9789 (
            .O(N__43033),
            .I(N__42988));
    InMux I__9788 (
            .O(N__43032),
            .I(N__42988));
    InMux I__9787 (
            .O(N__43031),
            .I(N__42918));
    InMux I__9786 (
            .O(N__43030),
            .I(N__42918));
    InMux I__9785 (
            .O(N__43029),
            .I(N__42918));
    InMux I__9784 (
            .O(N__43028),
            .I(N__42915));
    InMux I__9783 (
            .O(N__43027),
            .I(N__42910));
    InMux I__9782 (
            .O(N__43026),
            .I(N__42910));
    InMux I__9781 (
            .O(N__43025),
            .I(N__42893));
    InMux I__9780 (
            .O(N__43024),
            .I(N__42876));
    InMux I__9779 (
            .O(N__43023),
            .I(N__42876));
    InMux I__9778 (
            .O(N__43022),
            .I(N__42876));
    InMux I__9777 (
            .O(N__43021),
            .I(N__42876));
    InMux I__9776 (
            .O(N__43020),
            .I(N__42876));
    InMux I__9775 (
            .O(N__43019),
            .I(N__42876));
    InMux I__9774 (
            .O(N__43018),
            .I(N__42876));
    InMux I__9773 (
            .O(N__43017),
            .I(N__42876));
    InMux I__9772 (
            .O(N__43016),
            .I(N__42859));
    InMux I__9771 (
            .O(N__43015),
            .I(N__42859));
    InMux I__9770 (
            .O(N__43014),
            .I(N__42859));
    InMux I__9769 (
            .O(N__43013),
            .I(N__42859));
    InMux I__9768 (
            .O(N__43012),
            .I(N__42859));
    InMux I__9767 (
            .O(N__43011),
            .I(N__42859));
    InMux I__9766 (
            .O(N__43010),
            .I(N__42859));
    InMux I__9765 (
            .O(N__43009),
            .I(N__42859));
    InMux I__9764 (
            .O(N__43008),
            .I(N__42856));
    CascadeMux I__9763 (
            .O(N__43007),
            .I(N__42839));
    CascadeMux I__9762 (
            .O(N__43006),
            .I(N__42836));
    LocalMux I__9761 (
            .O(N__42997),
            .I(N__42825));
    LocalMux I__9760 (
            .O(N__42988),
            .I(N__42825));
    InMux I__9759 (
            .O(N__42987),
            .I(N__42818));
    InMux I__9758 (
            .O(N__42986),
            .I(N__42818));
    InMux I__9757 (
            .O(N__42985),
            .I(N__42818));
    CascadeMux I__9756 (
            .O(N__42984),
            .I(N__42813));
    InMux I__9755 (
            .O(N__42983),
            .I(N__42790));
    InMux I__9754 (
            .O(N__42982),
            .I(N__42790));
    InMux I__9753 (
            .O(N__42981),
            .I(N__42790));
    InMux I__9752 (
            .O(N__42980),
            .I(N__42790));
    InMux I__9751 (
            .O(N__42979),
            .I(N__42790));
    InMux I__9750 (
            .O(N__42978),
            .I(N__42790));
    InMux I__9749 (
            .O(N__42977),
            .I(N__42790));
    InMux I__9748 (
            .O(N__42976),
            .I(N__42790));
    InMux I__9747 (
            .O(N__42975),
            .I(N__42785));
    InMux I__9746 (
            .O(N__42974),
            .I(N__42785));
    InMux I__9745 (
            .O(N__42973),
            .I(N__42777));
    InMux I__9744 (
            .O(N__42972),
            .I(N__42777));
    InMux I__9743 (
            .O(N__42971),
            .I(N__42777));
    InMux I__9742 (
            .O(N__42970),
            .I(N__42768));
    InMux I__9741 (
            .O(N__42969),
            .I(N__42768));
    InMux I__9740 (
            .O(N__42968),
            .I(N__42768));
    InMux I__9739 (
            .O(N__42967),
            .I(N__42768));
    CascadeMux I__9738 (
            .O(N__42966),
            .I(N__42764));
    InMux I__9737 (
            .O(N__42965),
            .I(N__42753));
    CascadeMux I__9736 (
            .O(N__42964),
            .I(N__42750));
    CascadeMux I__9735 (
            .O(N__42963),
            .I(N__42747));
    InMux I__9734 (
            .O(N__42962),
            .I(N__42743));
    InMux I__9733 (
            .O(N__42961),
            .I(N__42716));
    InMux I__9732 (
            .O(N__42960),
            .I(N__42713));
    InMux I__9731 (
            .O(N__42959),
            .I(N__42694));
    InMux I__9730 (
            .O(N__42958),
            .I(N__42694));
    InMux I__9729 (
            .O(N__42957),
            .I(N__42694));
    InMux I__9728 (
            .O(N__42956),
            .I(N__42694));
    InMux I__9727 (
            .O(N__42955),
            .I(N__42677));
    InMux I__9726 (
            .O(N__42954),
            .I(N__42677));
    InMux I__9725 (
            .O(N__42953),
            .I(N__42677));
    InMux I__9724 (
            .O(N__42952),
            .I(N__42677));
    InMux I__9723 (
            .O(N__42951),
            .I(N__42677));
    InMux I__9722 (
            .O(N__42950),
            .I(N__42677));
    InMux I__9721 (
            .O(N__42949),
            .I(N__42677));
    InMux I__9720 (
            .O(N__42948),
            .I(N__42677));
    InMux I__9719 (
            .O(N__42947),
            .I(N__42664));
    InMux I__9718 (
            .O(N__42946),
            .I(N__42664));
    InMux I__9717 (
            .O(N__42945),
            .I(N__42664));
    InMux I__9716 (
            .O(N__42944),
            .I(N__42664));
    InMux I__9715 (
            .O(N__42943),
            .I(N__42664));
    InMux I__9714 (
            .O(N__42942),
            .I(N__42664));
    InMux I__9713 (
            .O(N__42941),
            .I(N__42655));
    InMux I__9712 (
            .O(N__42940),
            .I(N__42655));
    InMux I__9711 (
            .O(N__42939),
            .I(N__42655));
    InMux I__9710 (
            .O(N__42938),
            .I(N__42655));
    InMux I__9709 (
            .O(N__42937),
            .I(N__42644));
    InMux I__9708 (
            .O(N__42936),
            .I(N__42644));
    InMux I__9707 (
            .O(N__42935),
            .I(N__42644));
    InMux I__9706 (
            .O(N__42934),
            .I(N__42644));
    InMux I__9705 (
            .O(N__42933),
            .I(N__42644));
    InMux I__9704 (
            .O(N__42932),
            .I(N__42627));
    InMux I__9703 (
            .O(N__42931),
            .I(N__42627));
    InMux I__9702 (
            .O(N__42930),
            .I(N__42627));
    InMux I__9701 (
            .O(N__42929),
            .I(N__42627));
    InMux I__9700 (
            .O(N__42928),
            .I(N__42627));
    InMux I__9699 (
            .O(N__42927),
            .I(N__42627));
    InMux I__9698 (
            .O(N__42926),
            .I(N__42627));
    InMux I__9697 (
            .O(N__42925),
            .I(N__42627));
    LocalMux I__9696 (
            .O(N__42918),
            .I(N__42620));
    LocalMux I__9695 (
            .O(N__42915),
            .I(N__42620));
    LocalMux I__9694 (
            .O(N__42910),
            .I(N__42620));
    InMux I__9693 (
            .O(N__42909),
            .I(N__42615));
    InMux I__9692 (
            .O(N__42908),
            .I(N__42615));
    InMux I__9691 (
            .O(N__42907),
            .I(N__42610));
    InMux I__9690 (
            .O(N__42906),
            .I(N__42610));
    InMux I__9689 (
            .O(N__42905),
            .I(N__42601));
    InMux I__9688 (
            .O(N__42904),
            .I(N__42601));
    InMux I__9687 (
            .O(N__42903),
            .I(N__42601));
    InMux I__9686 (
            .O(N__42902),
            .I(N__42601));
    InMux I__9685 (
            .O(N__42901),
            .I(N__42592));
    InMux I__9684 (
            .O(N__42900),
            .I(N__42592));
    InMux I__9683 (
            .O(N__42899),
            .I(N__42592));
    InMux I__9682 (
            .O(N__42898),
            .I(N__42592));
    InMux I__9681 (
            .O(N__42897),
            .I(N__42587));
    InMux I__9680 (
            .O(N__42896),
            .I(N__42587));
    LocalMux I__9679 (
            .O(N__42893),
            .I(N__42570));
    LocalMux I__9678 (
            .O(N__42876),
            .I(N__42570));
    LocalMux I__9677 (
            .O(N__42859),
            .I(N__42570));
    LocalMux I__9676 (
            .O(N__42856),
            .I(N__42570));
    InMux I__9675 (
            .O(N__42855),
            .I(N__42561));
    InMux I__9674 (
            .O(N__42854),
            .I(N__42561));
    InMux I__9673 (
            .O(N__42853),
            .I(N__42561));
    InMux I__9672 (
            .O(N__42852),
            .I(N__42561));
    InMux I__9671 (
            .O(N__42851),
            .I(N__42544));
    InMux I__9670 (
            .O(N__42850),
            .I(N__42544));
    InMux I__9669 (
            .O(N__42849),
            .I(N__42544));
    InMux I__9668 (
            .O(N__42848),
            .I(N__42544));
    InMux I__9667 (
            .O(N__42847),
            .I(N__42544));
    InMux I__9666 (
            .O(N__42846),
            .I(N__42544));
    InMux I__9665 (
            .O(N__42845),
            .I(N__42544));
    InMux I__9664 (
            .O(N__42844),
            .I(N__42544));
    InMux I__9663 (
            .O(N__42843),
            .I(N__42539));
    InMux I__9662 (
            .O(N__42842),
            .I(N__42539));
    InMux I__9661 (
            .O(N__42839),
            .I(N__42530));
    InMux I__9660 (
            .O(N__42836),
            .I(N__42530));
    InMux I__9659 (
            .O(N__42835),
            .I(N__42530));
    InMux I__9658 (
            .O(N__42834),
            .I(N__42530));
    InMux I__9657 (
            .O(N__42833),
            .I(N__42525));
    InMux I__9656 (
            .O(N__42832),
            .I(N__42525));
    InMux I__9655 (
            .O(N__42831),
            .I(N__42520));
    InMux I__9654 (
            .O(N__42830),
            .I(N__42520));
    Span4Mux_v I__9653 (
            .O(N__42825),
            .I(N__42515));
    LocalMux I__9652 (
            .O(N__42818),
            .I(N__42515));
    InMux I__9651 (
            .O(N__42817),
            .I(N__42510));
    InMux I__9650 (
            .O(N__42816),
            .I(N__42510));
    InMux I__9649 (
            .O(N__42813),
            .I(N__42474));
    InMux I__9648 (
            .O(N__42812),
            .I(N__42461));
    InMux I__9647 (
            .O(N__42811),
            .I(N__42461));
    InMux I__9646 (
            .O(N__42810),
            .I(N__42461));
    InMux I__9645 (
            .O(N__42809),
            .I(N__42461));
    InMux I__9644 (
            .O(N__42808),
            .I(N__42461));
    InMux I__9643 (
            .O(N__42807),
            .I(N__42461));
    LocalMux I__9642 (
            .O(N__42790),
            .I(N__42456));
    LocalMux I__9641 (
            .O(N__42785),
            .I(N__42456));
    InMux I__9640 (
            .O(N__42784),
            .I(N__42453));
    LocalMux I__9639 (
            .O(N__42777),
            .I(N__42448));
    LocalMux I__9638 (
            .O(N__42768),
            .I(N__42448));
    InMux I__9637 (
            .O(N__42767),
            .I(N__42445));
    InMux I__9636 (
            .O(N__42764),
            .I(N__42440));
    InMux I__9635 (
            .O(N__42763),
            .I(N__42440));
    InMux I__9634 (
            .O(N__42762),
            .I(N__42435));
    InMux I__9633 (
            .O(N__42761),
            .I(N__42435));
    InMux I__9632 (
            .O(N__42760),
            .I(N__42424));
    InMux I__9631 (
            .O(N__42759),
            .I(N__42424));
    InMux I__9630 (
            .O(N__42758),
            .I(N__42424));
    InMux I__9629 (
            .O(N__42757),
            .I(N__42424));
    InMux I__9628 (
            .O(N__42756),
            .I(N__42424));
    LocalMux I__9627 (
            .O(N__42753),
            .I(N__42421));
    InMux I__9626 (
            .O(N__42750),
            .I(N__42414));
    InMux I__9625 (
            .O(N__42747),
            .I(N__42414));
    InMux I__9624 (
            .O(N__42746),
            .I(N__42414));
    LocalMux I__9623 (
            .O(N__42743),
            .I(N__42411));
    InMux I__9622 (
            .O(N__42742),
            .I(N__42400));
    InMux I__9621 (
            .O(N__42741),
            .I(N__42400));
    InMux I__9620 (
            .O(N__42740),
            .I(N__42400));
    InMux I__9619 (
            .O(N__42739),
            .I(N__42400));
    InMux I__9618 (
            .O(N__42738),
            .I(N__42400));
    InMux I__9617 (
            .O(N__42737),
            .I(N__42334));
    InMux I__9616 (
            .O(N__42736),
            .I(N__42334));
    InMux I__9615 (
            .O(N__42735),
            .I(N__42334));
    InMux I__9614 (
            .O(N__42734),
            .I(N__42334));
    InMux I__9613 (
            .O(N__42733),
            .I(N__42334));
    InMux I__9612 (
            .O(N__42732),
            .I(N__42323));
    InMux I__9611 (
            .O(N__42731),
            .I(N__42323));
    InMux I__9610 (
            .O(N__42730),
            .I(N__42323));
    InMux I__9609 (
            .O(N__42729),
            .I(N__42323));
    InMux I__9608 (
            .O(N__42728),
            .I(N__42323));
    InMux I__9607 (
            .O(N__42727),
            .I(N__42314));
    InMux I__9606 (
            .O(N__42726),
            .I(N__42314));
    InMux I__9605 (
            .O(N__42725),
            .I(N__42314));
    InMux I__9604 (
            .O(N__42724),
            .I(N__42314));
    InMux I__9603 (
            .O(N__42723),
            .I(N__42303));
    InMux I__9602 (
            .O(N__42722),
            .I(N__42303));
    InMux I__9601 (
            .O(N__42721),
            .I(N__42303));
    InMux I__9600 (
            .O(N__42720),
            .I(N__42303));
    InMux I__9599 (
            .O(N__42719),
            .I(N__42303));
    LocalMux I__9598 (
            .O(N__42716),
            .I(N__42300));
    LocalMux I__9597 (
            .O(N__42713),
            .I(N__42297));
    InMux I__9596 (
            .O(N__42712),
            .I(N__42292));
    InMux I__9595 (
            .O(N__42711),
            .I(N__42292));
    InMux I__9594 (
            .O(N__42710),
            .I(N__42275));
    InMux I__9593 (
            .O(N__42709),
            .I(N__42275));
    InMux I__9592 (
            .O(N__42708),
            .I(N__42275));
    InMux I__9591 (
            .O(N__42707),
            .I(N__42275));
    InMux I__9590 (
            .O(N__42706),
            .I(N__42275));
    InMux I__9589 (
            .O(N__42705),
            .I(N__42275));
    InMux I__9588 (
            .O(N__42704),
            .I(N__42275));
    InMux I__9587 (
            .O(N__42703),
            .I(N__42275));
    LocalMux I__9586 (
            .O(N__42694),
            .I(N__42272));
    LocalMux I__9585 (
            .O(N__42677),
            .I(N__42269));
    LocalMux I__9584 (
            .O(N__42664),
            .I(N__42260));
    LocalMux I__9583 (
            .O(N__42655),
            .I(N__42260));
    LocalMux I__9582 (
            .O(N__42644),
            .I(N__42260));
    LocalMux I__9581 (
            .O(N__42627),
            .I(N__42260));
    Span4Mux_h I__9580 (
            .O(N__42620),
            .I(N__42251));
    LocalMux I__9579 (
            .O(N__42615),
            .I(N__42251));
    LocalMux I__9578 (
            .O(N__42610),
            .I(N__42251));
    LocalMux I__9577 (
            .O(N__42601),
            .I(N__42251));
    LocalMux I__9576 (
            .O(N__42592),
            .I(N__42246));
    LocalMux I__9575 (
            .O(N__42587),
            .I(N__42246));
    InMux I__9574 (
            .O(N__42586),
            .I(N__42221));
    InMux I__9573 (
            .O(N__42585),
            .I(N__42221));
    InMux I__9572 (
            .O(N__42584),
            .I(N__42221));
    InMux I__9571 (
            .O(N__42583),
            .I(N__42221));
    InMux I__9570 (
            .O(N__42582),
            .I(N__42221));
    InMux I__9569 (
            .O(N__42581),
            .I(N__42221));
    InMux I__9568 (
            .O(N__42580),
            .I(N__42221));
    InMux I__9567 (
            .O(N__42579),
            .I(N__42221));
    Span4Mux_v I__9566 (
            .O(N__42570),
            .I(N__42216));
    LocalMux I__9565 (
            .O(N__42561),
            .I(N__42216));
    LocalMux I__9564 (
            .O(N__42544),
            .I(N__42209));
    LocalMux I__9563 (
            .O(N__42539),
            .I(N__42209));
    LocalMux I__9562 (
            .O(N__42530),
            .I(N__42209));
    LocalMux I__9561 (
            .O(N__42525),
            .I(N__42200));
    LocalMux I__9560 (
            .O(N__42520),
            .I(N__42200));
    Span4Mux_v I__9559 (
            .O(N__42515),
            .I(N__42200));
    LocalMux I__9558 (
            .O(N__42510),
            .I(N__42200));
    InMux I__9557 (
            .O(N__42509),
            .I(N__42183));
    InMux I__9556 (
            .O(N__42508),
            .I(N__42183));
    InMux I__9555 (
            .O(N__42507),
            .I(N__42183));
    InMux I__9554 (
            .O(N__42506),
            .I(N__42183));
    InMux I__9553 (
            .O(N__42505),
            .I(N__42183));
    InMux I__9552 (
            .O(N__42504),
            .I(N__42183));
    InMux I__9551 (
            .O(N__42503),
            .I(N__42183));
    InMux I__9550 (
            .O(N__42502),
            .I(N__42183));
    InMux I__9549 (
            .O(N__42501),
            .I(N__42174));
    InMux I__9548 (
            .O(N__42500),
            .I(N__42174));
    InMux I__9547 (
            .O(N__42499),
            .I(N__42174));
    InMux I__9546 (
            .O(N__42498),
            .I(N__42174));
    InMux I__9545 (
            .O(N__42497),
            .I(N__42159));
    InMux I__9544 (
            .O(N__42496),
            .I(N__42159));
    InMux I__9543 (
            .O(N__42495),
            .I(N__42159));
    InMux I__9542 (
            .O(N__42494),
            .I(N__42159));
    InMux I__9541 (
            .O(N__42493),
            .I(N__42159));
    InMux I__9540 (
            .O(N__42492),
            .I(N__42159));
    InMux I__9539 (
            .O(N__42491),
            .I(N__42159));
    InMux I__9538 (
            .O(N__42490),
            .I(N__42142));
    InMux I__9537 (
            .O(N__42489),
            .I(N__42142));
    InMux I__9536 (
            .O(N__42488),
            .I(N__42142));
    InMux I__9535 (
            .O(N__42487),
            .I(N__42142));
    InMux I__9534 (
            .O(N__42486),
            .I(N__42142));
    InMux I__9533 (
            .O(N__42485),
            .I(N__42142));
    InMux I__9532 (
            .O(N__42484),
            .I(N__42142));
    InMux I__9531 (
            .O(N__42483),
            .I(N__42142));
    InMux I__9530 (
            .O(N__42482),
            .I(N__42129));
    InMux I__9529 (
            .O(N__42481),
            .I(N__42129));
    InMux I__9528 (
            .O(N__42480),
            .I(N__42129));
    InMux I__9527 (
            .O(N__42479),
            .I(N__42129));
    InMux I__9526 (
            .O(N__42478),
            .I(N__42129));
    InMux I__9525 (
            .O(N__42477),
            .I(N__42129));
    LocalMux I__9524 (
            .O(N__42474),
            .I(N__42120));
    LocalMux I__9523 (
            .O(N__42461),
            .I(N__42120));
    Span4Mux_v I__9522 (
            .O(N__42456),
            .I(N__42120));
    LocalMux I__9521 (
            .O(N__42453),
            .I(N__42120));
    Span4Mux_h I__9520 (
            .O(N__42448),
            .I(N__42115));
    LocalMux I__9519 (
            .O(N__42445),
            .I(N__42115));
    LocalMux I__9518 (
            .O(N__42440),
            .I(N__42112));
    LocalMux I__9517 (
            .O(N__42435),
            .I(N__42105));
    LocalMux I__9516 (
            .O(N__42424),
            .I(N__42105));
    Span4Mux_h I__9515 (
            .O(N__42421),
            .I(N__42105));
    LocalMux I__9514 (
            .O(N__42414),
            .I(N__42098));
    Span4Mux_h I__9513 (
            .O(N__42411),
            .I(N__42098));
    LocalMux I__9512 (
            .O(N__42400),
            .I(N__42098));
    InMux I__9511 (
            .O(N__42399),
            .I(N__42081));
    InMux I__9510 (
            .O(N__42398),
            .I(N__42081));
    InMux I__9509 (
            .O(N__42397),
            .I(N__42081));
    InMux I__9508 (
            .O(N__42396),
            .I(N__42081));
    InMux I__9507 (
            .O(N__42395),
            .I(N__42081));
    InMux I__9506 (
            .O(N__42394),
            .I(N__42081));
    InMux I__9505 (
            .O(N__42393),
            .I(N__42081));
    InMux I__9504 (
            .O(N__42392),
            .I(N__42081));
    InMux I__9503 (
            .O(N__42391),
            .I(N__42064));
    InMux I__9502 (
            .O(N__42390),
            .I(N__42064));
    InMux I__9501 (
            .O(N__42389),
            .I(N__42064));
    InMux I__9500 (
            .O(N__42388),
            .I(N__42064));
    InMux I__9499 (
            .O(N__42387),
            .I(N__42064));
    InMux I__9498 (
            .O(N__42386),
            .I(N__42064));
    InMux I__9497 (
            .O(N__42385),
            .I(N__42064));
    InMux I__9496 (
            .O(N__42384),
            .I(N__42064));
    InMux I__9495 (
            .O(N__42383),
            .I(N__42049));
    InMux I__9494 (
            .O(N__42382),
            .I(N__42049));
    InMux I__9493 (
            .O(N__42381),
            .I(N__42049));
    InMux I__9492 (
            .O(N__42380),
            .I(N__42049));
    InMux I__9491 (
            .O(N__42379),
            .I(N__42049));
    InMux I__9490 (
            .O(N__42378),
            .I(N__42049));
    InMux I__9489 (
            .O(N__42377),
            .I(N__42049));
    InMux I__9488 (
            .O(N__42376),
            .I(N__42032));
    InMux I__9487 (
            .O(N__42375),
            .I(N__42032));
    InMux I__9486 (
            .O(N__42374),
            .I(N__42032));
    InMux I__9485 (
            .O(N__42373),
            .I(N__42032));
    InMux I__9484 (
            .O(N__42372),
            .I(N__42032));
    InMux I__9483 (
            .O(N__42371),
            .I(N__42032));
    InMux I__9482 (
            .O(N__42370),
            .I(N__42032));
    InMux I__9481 (
            .O(N__42369),
            .I(N__42032));
    InMux I__9480 (
            .O(N__42368),
            .I(N__42015));
    InMux I__9479 (
            .O(N__42367),
            .I(N__42015));
    InMux I__9478 (
            .O(N__42366),
            .I(N__42015));
    InMux I__9477 (
            .O(N__42365),
            .I(N__42015));
    InMux I__9476 (
            .O(N__42364),
            .I(N__42015));
    InMux I__9475 (
            .O(N__42363),
            .I(N__42015));
    InMux I__9474 (
            .O(N__42362),
            .I(N__42015));
    InMux I__9473 (
            .O(N__42361),
            .I(N__42015));
    InMux I__9472 (
            .O(N__42360),
            .I(N__41998));
    InMux I__9471 (
            .O(N__42359),
            .I(N__41998));
    InMux I__9470 (
            .O(N__42358),
            .I(N__41998));
    InMux I__9469 (
            .O(N__42357),
            .I(N__41998));
    InMux I__9468 (
            .O(N__42356),
            .I(N__41998));
    InMux I__9467 (
            .O(N__42355),
            .I(N__41998));
    InMux I__9466 (
            .O(N__42354),
            .I(N__41998));
    InMux I__9465 (
            .O(N__42353),
            .I(N__41998));
    InMux I__9464 (
            .O(N__42352),
            .I(N__41981));
    InMux I__9463 (
            .O(N__42351),
            .I(N__41981));
    InMux I__9462 (
            .O(N__42350),
            .I(N__41981));
    InMux I__9461 (
            .O(N__42349),
            .I(N__41981));
    InMux I__9460 (
            .O(N__42348),
            .I(N__41981));
    InMux I__9459 (
            .O(N__42347),
            .I(N__41981));
    InMux I__9458 (
            .O(N__42346),
            .I(N__41981));
    InMux I__9457 (
            .O(N__42345),
            .I(N__41981));
    LocalMux I__9456 (
            .O(N__42334),
            .I(N__41976));
    LocalMux I__9455 (
            .O(N__42323),
            .I(N__41976));
    LocalMux I__9454 (
            .O(N__42314),
            .I(N__41971));
    LocalMux I__9453 (
            .O(N__42303),
            .I(N__41971));
    Span4Mux_h I__9452 (
            .O(N__42300),
            .I(N__41964));
    Span4Mux_v I__9451 (
            .O(N__42297),
            .I(N__41964));
    LocalMux I__9450 (
            .O(N__42292),
            .I(N__41964));
    LocalMux I__9449 (
            .O(N__42275),
            .I(N__41951));
    Span4Mux_v I__9448 (
            .O(N__42272),
            .I(N__41951));
    Span4Mux_h I__9447 (
            .O(N__42269),
            .I(N__41951));
    Span4Mux_h I__9446 (
            .O(N__42260),
            .I(N__41951));
    Span4Mux_v I__9445 (
            .O(N__42251),
            .I(N__41951));
    Span4Mux_v I__9444 (
            .O(N__42246),
            .I(N__41951));
    InMux I__9443 (
            .O(N__42245),
            .I(N__41934));
    InMux I__9442 (
            .O(N__42244),
            .I(N__41934));
    InMux I__9441 (
            .O(N__42243),
            .I(N__41934));
    InMux I__9440 (
            .O(N__42242),
            .I(N__41934));
    InMux I__9439 (
            .O(N__42241),
            .I(N__41934));
    InMux I__9438 (
            .O(N__42240),
            .I(N__41934));
    InMux I__9437 (
            .O(N__42239),
            .I(N__41934));
    InMux I__9436 (
            .O(N__42238),
            .I(N__41934));
    LocalMux I__9435 (
            .O(N__42221),
            .I(N__41925));
    Span4Mux_h I__9434 (
            .O(N__42216),
            .I(N__41925));
    Span4Mux_h I__9433 (
            .O(N__42209),
            .I(N__41925));
    Span4Mux_h I__9432 (
            .O(N__42200),
            .I(N__41925));
    LocalMux I__9431 (
            .O(N__42183),
            .I(N__41922));
    LocalMux I__9430 (
            .O(N__42174),
            .I(N__41909));
    LocalMux I__9429 (
            .O(N__42159),
            .I(N__41909));
    LocalMux I__9428 (
            .O(N__42142),
            .I(N__41909));
    LocalMux I__9427 (
            .O(N__42129),
            .I(N__41909));
    Span4Mux_h I__9426 (
            .O(N__42120),
            .I(N__41909));
    Span4Mux_h I__9425 (
            .O(N__42115),
            .I(N__41909));
    Span4Mux_h I__9424 (
            .O(N__42112),
            .I(N__41902));
    Span4Mux_h I__9423 (
            .O(N__42105),
            .I(N__41902));
    Span4Mux_h I__9422 (
            .O(N__42098),
            .I(N__41902));
    LocalMux I__9421 (
            .O(N__42081),
            .I(\u1.DMA_control.N_1313 ));
    LocalMux I__9420 (
            .O(N__42064),
            .I(\u1.DMA_control.N_1313 ));
    LocalMux I__9419 (
            .O(N__42049),
            .I(\u1.DMA_control.N_1313 ));
    LocalMux I__9418 (
            .O(N__42032),
            .I(\u1.DMA_control.N_1313 ));
    LocalMux I__9417 (
            .O(N__42015),
            .I(\u1.DMA_control.N_1313 ));
    LocalMux I__9416 (
            .O(N__41998),
            .I(\u1.DMA_control.N_1313 ));
    LocalMux I__9415 (
            .O(N__41981),
            .I(\u1.DMA_control.N_1313 ));
    Odrv4 I__9414 (
            .O(N__41976),
            .I(\u1.DMA_control.N_1313 ));
    Odrv12 I__9413 (
            .O(N__41971),
            .I(\u1.DMA_control.N_1313 ));
    Odrv4 I__9412 (
            .O(N__41964),
            .I(\u1.DMA_control.N_1313 ));
    Odrv4 I__9411 (
            .O(N__41951),
            .I(\u1.DMA_control.N_1313 ));
    LocalMux I__9410 (
            .O(N__41934),
            .I(\u1.DMA_control.N_1313 ));
    Odrv4 I__9409 (
            .O(N__41925),
            .I(\u1.DMA_control.N_1313 ));
    Odrv12 I__9408 (
            .O(N__41922),
            .I(\u1.DMA_control.N_1313 ));
    Odrv4 I__9407 (
            .O(N__41909),
            .I(\u1.DMA_control.N_1313 ));
    Odrv4 I__9406 (
            .O(N__41902),
            .I(\u1.DMA_control.N_1313 ));
    InMux I__9405 (
            .O(N__41869),
            .I(N__41866));
    LocalMux I__9404 (
            .O(N__41866),
            .I(N__41863));
    Odrv4 I__9403 (
            .O(N__41863),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_27 ));
    CEMux I__9402 (
            .O(N__41860),
            .I(N__41856));
    CEMux I__9401 (
            .O(N__41859),
            .I(N__41850));
    LocalMux I__9400 (
            .O(N__41856),
            .I(N__41846));
    CEMux I__9399 (
            .O(N__41855),
            .I(N__41843));
    CEMux I__9398 (
            .O(N__41854),
            .I(N__41840));
    CEMux I__9397 (
            .O(N__41853),
            .I(N__41837));
    LocalMux I__9396 (
            .O(N__41850),
            .I(N__41834));
    CEMux I__9395 (
            .O(N__41849),
            .I(N__41830));
    Span4Mux_v I__9394 (
            .O(N__41846),
            .I(N__41827));
    LocalMux I__9393 (
            .O(N__41843),
            .I(N__41822));
    LocalMux I__9392 (
            .O(N__41840),
            .I(N__41822));
    LocalMux I__9391 (
            .O(N__41837),
            .I(N__41819));
    Span4Mux_v I__9390 (
            .O(N__41834),
            .I(N__41815));
    CEMux I__9389 (
            .O(N__41833),
            .I(N__41812));
    LocalMux I__9388 (
            .O(N__41830),
            .I(N__41809));
    Span4Mux_h I__9387 (
            .O(N__41827),
            .I(N__41802));
    Span4Mux_v I__9386 (
            .O(N__41822),
            .I(N__41802));
    Span4Mux_v I__9385 (
            .O(N__41819),
            .I(N__41802));
    CEMux I__9384 (
            .O(N__41818),
            .I(N__41799));
    Span4Mux_h I__9383 (
            .O(N__41815),
            .I(N__41795));
    LocalMux I__9382 (
            .O(N__41812),
            .I(N__41792));
    Span4Mux_h I__9381 (
            .O(N__41809),
            .I(N__41785));
    Span4Mux_h I__9380 (
            .O(N__41802),
            .I(N__41785));
    LocalMux I__9379 (
            .O(N__41799),
            .I(N__41785));
    CEMux I__9378 (
            .O(N__41798),
            .I(N__41782));
    Span4Mux_h I__9377 (
            .O(N__41795),
            .I(N__41777));
    Span4Mux_v I__9376 (
            .O(N__41792),
            .I(N__41777));
    Span4Mux_h I__9375 (
            .O(N__41785),
            .I(N__41774));
    LocalMux I__9374 (
            .O(N__41782),
            .I(N__41771));
    Odrv4 I__9373 (
            .O(N__41777),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_awe4 ));
    Odrv4 I__9372 (
            .O(N__41774),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_awe4 ));
    Odrv12 I__9371 (
            .O(N__41771),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_awe4 ));
    InMux I__9370 (
            .O(N__41764),
            .I(N__41761));
    LocalMux I__9369 (
            .O(N__41761),
            .I(N__41758));
    Odrv12 I__9368 (
            .O(N__41758),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI1SG71Z0Z_30 ));
    InMux I__9367 (
            .O(N__41755),
            .I(N__41752));
    LocalMux I__9366 (
            .O(N__41752),
            .I(N__41749));
    Odrv12 I__9365 (
            .O(N__41749),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIECLM1Z0Z_2 ));
    InMux I__9364 (
            .O(N__41746),
            .I(N__41743));
    LocalMux I__9363 (
            .O(N__41743),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI4RUQZ0Z_16 ));
    InMux I__9362 (
            .O(N__41740),
            .I(N__41734));
    InMux I__9361 (
            .O(N__41739),
            .I(N__41725));
    InMux I__9360 (
            .O(N__41738),
            .I(N__41725));
    InMux I__9359 (
            .O(N__41737),
            .I(N__41722));
    LocalMux I__9358 (
            .O(N__41734),
            .I(N__41719));
    InMux I__9357 (
            .O(N__41733),
            .I(N__41714));
    InMux I__9356 (
            .O(N__41732),
            .I(N__41714));
    InMux I__9355 (
            .O(N__41731),
            .I(N__41709));
    InMux I__9354 (
            .O(N__41730),
            .I(N__41709));
    LocalMux I__9353 (
            .O(N__41725),
            .I(N__41704));
    LocalMux I__9352 (
            .O(N__41722),
            .I(N__41704));
    Span4Mux_v I__9351 (
            .O(N__41719),
            .I(N__41696));
    LocalMux I__9350 (
            .O(N__41714),
            .I(N__41696));
    LocalMux I__9349 (
            .O(N__41709),
            .I(N__41693));
    Span4Mux_h I__9348 (
            .O(N__41704),
            .I(N__41690));
    InMux I__9347 (
            .O(N__41703),
            .I(N__41685));
    InMux I__9346 (
            .O(N__41702),
            .I(N__41685));
    InMux I__9345 (
            .O(N__41701),
            .I(N__41678));
    Span4Mux_h I__9344 (
            .O(N__41696),
            .I(N__41675));
    Span4Mux_h I__9343 (
            .O(N__41693),
            .I(N__41672));
    Sp12to4 I__9342 (
            .O(N__41690),
            .I(N__41667));
    LocalMux I__9341 (
            .O(N__41685),
            .I(N__41667));
    InMux I__9340 (
            .O(N__41684),
            .I(N__41662));
    InMux I__9339 (
            .O(N__41683),
            .I(N__41662));
    InMux I__9338 (
            .O(N__41682),
            .I(N__41657));
    InMux I__9337 (
            .O(N__41681),
            .I(N__41657));
    LocalMux I__9336 (
            .O(N__41678),
            .I(\u1.DMA_control.readDlw_0 ));
    Odrv4 I__9335 (
            .O(N__41675),
            .I(\u1.DMA_control.readDlw_0 ));
    Odrv4 I__9334 (
            .O(N__41672),
            .I(\u1.DMA_control.readDlw_0 ));
    Odrv12 I__9333 (
            .O(N__41667),
            .I(\u1.DMA_control.readDlw_0 ));
    LocalMux I__9332 (
            .O(N__41662),
            .I(\u1.DMA_control.readDlw_0 ));
    LocalMux I__9331 (
            .O(N__41657),
            .I(\u1.DMA_control.readDlw_0 ));
    InMux I__9330 (
            .O(N__41644),
            .I(N__41638));
    InMux I__9329 (
            .O(N__41643),
            .I(N__41633));
    InMux I__9328 (
            .O(N__41642),
            .I(N__41633));
    InMux I__9327 (
            .O(N__41641),
            .I(N__41630));
    LocalMux I__9326 (
            .O(N__41638),
            .I(N__41618));
    LocalMux I__9325 (
            .O(N__41633),
            .I(N__41618));
    LocalMux I__9324 (
            .O(N__41630),
            .I(N__41618));
    InMux I__9323 (
            .O(N__41629),
            .I(N__41615));
    InMux I__9322 (
            .O(N__41628),
            .I(N__41612));
    InMux I__9321 (
            .O(N__41627),
            .I(N__41609));
    InMux I__9320 (
            .O(N__41626),
            .I(N__41606));
    CascadeMux I__9319 (
            .O(N__41625),
            .I(N__41603));
    Span4Mux_v I__9318 (
            .O(N__41618),
            .I(N__41595));
    LocalMux I__9317 (
            .O(N__41615),
            .I(N__41595));
    LocalMux I__9316 (
            .O(N__41612),
            .I(N__41595));
    LocalMux I__9315 (
            .O(N__41609),
            .I(N__41590));
    LocalMux I__9314 (
            .O(N__41606),
            .I(N__41590));
    InMux I__9313 (
            .O(N__41603),
            .I(N__41585));
    InMux I__9312 (
            .O(N__41602),
            .I(N__41585));
    Span4Mux_h I__9311 (
            .O(N__41595),
            .I(N__41578));
    Span4Mux_h I__9310 (
            .O(N__41590),
            .I(N__41575));
    LocalMux I__9309 (
            .O(N__41585),
            .I(N__41572));
    InMux I__9308 (
            .O(N__41584),
            .I(N__41569));
    InMux I__9307 (
            .O(N__41583),
            .I(N__41566));
    InMux I__9306 (
            .O(N__41582),
            .I(N__41563));
    InMux I__9305 (
            .O(N__41581),
            .I(N__41560));
    Odrv4 I__9304 (
            .O(N__41578),
            .I(\u1.DMA_control.readDfw_0 ));
    Odrv4 I__9303 (
            .O(N__41575),
            .I(\u1.DMA_control.readDfw_0 ));
    Odrv12 I__9302 (
            .O(N__41572),
            .I(\u1.DMA_control.readDfw_0 ));
    LocalMux I__9301 (
            .O(N__41569),
            .I(\u1.DMA_control.readDfw_0 ));
    LocalMux I__9300 (
            .O(N__41566),
            .I(\u1.DMA_control.readDfw_0 ));
    LocalMux I__9299 (
            .O(N__41563),
            .I(\u1.DMA_control.readDfw_0 ));
    LocalMux I__9298 (
            .O(N__41560),
            .I(\u1.DMA_control.readDfw_0 ));
    InMux I__9297 (
            .O(N__41545),
            .I(N__41542));
    LocalMux I__9296 (
            .O(N__41542),
            .I(N__41539));
    Odrv4 I__9295 (
            .O(N__41539),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_1 ));
    CascadeMux I__9294 (
            .O(N__41536),
            .I(N__41531));
    InMux I__9293 (
            .O(N__41535),
            .I(N__41528));
    CascadeMux I__9292 (
            .O(N__41534),
            .I(N__41525));
    InMux I__9291 (
            .O(N__41531),
            .I(N__41522));
    LocalMux I__9290 (
            .O(N__41528),
            .I(N__41515));
    InMux I__9289 (
            .O(N__41525),
            .I(N__41506));
    LocalMux I__9288 (
            .O(N__41522),
            .I(N__41503));
    InMux I__9287 (
            .O(N__41521),
            .I(N__41500));
    InMux I__9286 (
            .O(N__41520),
            .I(N__41497));
    InMux I__9285 (
            .O(N__41519),
            .I(N__41492));
    InMux I__9284 (
            .O(N__41518),
            .I(N__41492));
    Span4Mux_h I__9283 (
            .O(N__41515),
            .I(N__41489));
    InMux I__9282 (
            .O(N__41514),
            .I(N__41486));
    InMux I__9281 (
            .O(N__41513),
            .I(N__41481));
    InMux I__9280 (
            .O(N__41512),
            .I(N__41476));
    InMux I__9279 (
            .O(N__41511),
            .I(N__41476));
    InMux I__9278 (
            .O(N__41510),
            .I(N__41471));
    InMux I__9277 (
            .O(N__41509),
            .I(N__41471));
    LocalMux I__9276 (
            .O(N__41506),
            .I(N__41462));
    Span4Mux_h I__9275 (
            .O(N__41503),
            .I(N__41462));
    LocalMux I__9274 (
            .O(N__41500),
            .I(N__41462));
    LocalMux I__9273 (
            .O(N__41497),
            .I(N__41462));
    LocalMux I__9272 (
            .O(N__41492),
            .I(N__41459));
    Span4Mux_v I__9271 (
            .O(N__41489),
            .I(N__41454));
    LocalMux I__9270 (
            .O(N__41486),
            .I(N__41454));
    InMux I__9269 (
            .O(N__41485),
            .I(N__41451));
    InMux I__9268 (
            .O(N__41484),
            .I(N__41448));
    LocalMux I__9267 (
            .O(N__41481),
            .I(N__41445));
    LocalMux I__9266 (
            .O(N__41476),
            .I(N__41442));
    LocalMux I__9265 (
            .O(N__41471),
            .I(N__41435));
    Span4Mux_v I__9264 (
            .O(N__41462),
            .I(N__41435));
    Span4Mux_v I__9263 (
            .O(N__41459),
            .I(N__41435));
    Span4Mux_h I__9262 (
            .O(N__41454),
            .I(N__41432));
    LocalMux I__9261 (
            .O(N__41451),
            .I(\u1.DMA_control.readDlw_1 ));
    LocalMux I__9260 (
            .O(N__41448),
            .I(\u1.DMA_control.readDlw_1 ));
    Odrv4 I__9259 (
            .O(N__41445),
            .I(\u1.DMA_control.readDlw_1 ));
    Odrv4 I__9258 (
            .O(N__41442),
            .I(\u1.DMA_control.readDlw_1 ));
    Odrv4 I__9257 (
            .O(N__41435),
            .I(\u1.DMA_control.readDlw_1 ));
    Odrv4 I__9256 (
            .O(N__41432),
            .I(\u1.DMA_control.readDlw_1 ));
    InMux I__9255 (
            .O(N__41419),
            .I(N__41414));
    InMux I__9254 (
            .O(N__41418),
            .I(N__41406));
    InMux I__9253 (
            .O(N__41417),
            .I(N__41403));
    LocalMux I__9252 (
            .O(N__41414),
            .I(N__41399));
    InMux I__9251 (
            .O(N__41413),
            .I(N__41396));
    InMux I__9250 (
            .O(N__41412),
            .I(N__41393));
    InMux I__9249 (
            .O(N__41411),
            .I(N__41390));
    InMux I__9248 (
            .O(N__41410),
            .I(N__41387));
    InMux I__9247 (
            .O(N__41409),
            .I(N__41384));
    LocalMux I__9246 (
            .O(N__41406),
            .I(N__41379));
    LocalMux I__9245 (
            .O(N__41403),
            .I(N__41376));
    InMux I__9244 (
            .O(N__41402),
            .I(N__41373));
    Span4Mux_h I__9243 (
            .O(N__41399),
            .I(N__41362));
    LocalMux I__9242 (
            .O(N__41396),
            .I(N__41362));
    LocalMux I__9241 (
            .O(N__41393),
            .I(N__41362));
    LocalMux I__9240 (
            .O(N__41390),
            .I(N__41362));
    LocalMux I__9239 (
            .O(N__41387),
            .I(N__41357));
    LocalMux I__9238 (
            .O(N__41384),
            .I(N__41357));
    InMux I__9237 (
            .O(N__41383),
            .I(N__41354));
    InMux I__9236 (
            .O(N__41382),
            .I(N__41351));
    Span4Mux_h I__9235 (
            .O(N__41379),
            .I(N__41345));
    Span4Mux_h I__9234 (
            .O(N__41376),
            .I(N__41345));
    LocalMux I__9233 (
            .O(N__41373),
            .I(N__41342));
    InMux I__9232 (
            .O(N__41372),
            .I(N__41339));
    InMux I__9231 (
            .O(N__41371),
            .I(N__41336));
    Span4Mux_v I__9230 (
            .O(N__41362),
            .I(N__41327));
    Span4Mux_v I__9229 (
            .O(N__41357),
            .I(N__41327));
    LocalMux I__9228 (
            .O(N__41354),
            .I(N__41327));
    LocalMux I__9227 (
            .O(N__41351),
            .I(N__41327));
    InMux I__9226 (
            .O(N__41350),
            .I(N__41324));
    Odrv4 I__9225 (
            .O(N__41345),
            .I(\u1.DMA_control.readDfw_1 ));
    Odrv4 I__9224 (
            .O(N__41342),
            .I(\u1.DMA_control.readDfw_1 ));
    LocalMux I__9223 (
            .O(N__41339),
            .I(\u1.DMA_control.readDfw_1 ));
    LocalMux I__9222 (
            .O(N__41336),
            .I(\u1.DMA_control.readDfw_1 ));
    Odrv4 I__9221 (
            .O(N__41327),
            .I(\u1.DMA_control.readDfw_1 ));
    LocalMux I__9220 (
            .O(N__41324),
            .I(\u1.DMA_control.readDfw_1 ));
    InMux I__9219 (
            .O(N__41311),
            .I(N__41308));
    LocalMux I__9218 (
            .O(N__41308),
            .I(N__41305));
    Span4Mux_v I__9217 (
            .O(N__41305),
            .I(N__41302));
    Odrv4 I__9216 (
            .O(N__41302),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_11 ));
    CEMux I__9215 (
            .O(N__41299),
            .I(N__41292));
    CEMux I__9214 (
            .O(N__41298),
            .I(N__41289));
    CEMux I__9213 (
            .O(N__41297),
            .I(N__41285));
    CEMux I__9212 (
            .O(N__41296),
            .I(N__41282));
    CEMux I__9211 (
            .O(N__41295),
            .I(N__41279));
    LocalMux I__9210 (
            .O(N__41292),
            .I(N__41276));
    LocalMux I__9209 (
            .O(N__41289),
            .I(N__41273));
    CEMux I__9208 (
            .O(N__41288),
            .I(N__41270));
    LocalMux I__9207 (
            .O(N__41285),
            .I(N__41265));
    LocalMux I__9206 (
            .O(N__41282),
            .I(N__41262));
    LocalMux I__9205 (
            .O(N__41279),
            .I(N__41253));
    Span4Mux_h I__9204 (
            .O(N__41276),
            .I(N__41253));
    Span4Mux_h I__9203 (
            .O(N__41273),
            .I(N__41253));
    LocalMux I__9202 (
            .O(N__41270),
            .I(N__41253));
    CEMux I__9201 (
            .O(N__41269),
            .I(N__41250));
    CEMux I__9200 (
            .O(N__41268),
            .I(N__41247));
    Span4Mux_h I__9199 (
            .O(N__41265),
            .I(N__41243));
    Span4Mux_v I__9198 (
            .O(N__41262),
            .I(N__41238));
    Span4Mux_v I__9197 (
            .O(N__41253),
            .I(N__41238));
    LocalMux I__9196 (
            .O(N__41250),
            .I(N__41235));
    LocalMux I__9195 (
            .O(N__41247),
            .I(N__41232));
    CEMux I__9194 (
            .O(N__41246),
            .I(N__41229));
    Span4Mux_h I__9193 (
            .O(N__41243),
            .I(N__41226));
    Span4Mux_h I__9192 (
            .O(N__41238),
            .I(N__41223));
    Span4Mux_h I__9191 (
            .O(N__41235),
            .I(N__41220));
    Span4Mux_h I__9190 (
            .O(N__41232),
            .I(N__41217));
    LocalMux I__9189 (
            .O(N__41229),
            .I(N__41214));
    Odrv4 I__9188 (
            .O(N__41226),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_awe6 ));
    Odrv4 I__9187 (
            .O(N__41223),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_awe6 ));
    Odrv4 I__9186 (
            .O(N__41220),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_awe6 ));
    Odrv4 I__9185 (
            .O(N__41217),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_awe6 ));
    Odrv4 I__9184 (
            .O(N__41214),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_awe6 ));
    InMux I__9183 (
            .O(N__41203),
            .I(N__41200));
    LocalMux I__9182 (
            .O(N__41200),
            .I(N__41197));
    Span4Mux_v I__9181 (
            .O(N__41197),
            .I(N__41194));
    Odrv4 I__9180 (
            .O(N__41194),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIG9ITZ0Z_27 ));
    InMux I__9179 (
            .O(N__41191),
            .I(N__41188));
    LocalMux I__9178 (
            .O(N__41188),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_27 ));
    InMux I__9177 (
            .O(N__41185),
            .I(N__41182));
    LocalMux I__9176 (
            .O(N__41182),
            .I(N__41179));
    Span4Mux_v I__9175 (
            .O(N__41179),
            .I(N__41176));
    Odrv4 I__9174 (
            .O(N__41176),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIJBE71Z0Z_27 ));
    InMux I__9173 (
            .O(N__41173),
            .I(N__41170));
    LocalMux I__9172 (
            .O(N__41170),
            .I(N__41167));
    Span4Mux_h I__9171 (
            .O(N__41167),
            .I(N__41164));
    Span4Mux_h I__9170 (
            .O(N__41164),
            .I(N__41161));
    Span4Mux_h I__9169 (
            .O(N__41161),
            .I(N__41157));
    InMux I__9168 (
            .O(N__41160),
            .I(N__41154));
    Span4Mux_v I__9167 (
            .O(N__41157),
            .I(N__41149));
    LocalMux I__9166 (
            .O(N__41154),
            .I(N__41149));
    Span4Mux_v I__9165 (
            .O(N__41149),
            .I(N__41146));
    Span4Mux_h I__9164 (
            .O(N__41146),
            .I(N__41143));
    Odrv4 I__9163 (
            .O(N__41143),
            .I(DMA_dev0_Tm_0));
    InMux I__9162 (
            .O(N__41140),
            .I(N__41137));
    LocalMux I__9161 (
            .O(N__41137),
            .I(N__41134));
    Span4Mux_v I__9160 (
            .O(N__41134),
            .I(N__41131));
    Odrv4 I__9159 (
            .O(N__41131),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNIEDTNZ0Z_8 ));
    InMux I__9158 (
            .O(N__41128),
            .I(N__41125));
    LocalMux I__9157 (
            .O(N__41125),
            .I(N__41122));
    Span4Mux_v I__9156 (
            .O(N__41122),
            .I(N__41119));
    Odrv4 I__9155 (
            .O(N__41119),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_8 ));
    InMux I__9154 (
            .O(N__41116),
            .I(N__41113));
    LocalMux I__9153 (
            .O(N__41113),
            .I(N__41110));
    Span4Mux_v I__9152 (
            .O(N__41110),
            .I(N__41107));
    Odrv4 I__9151 (
            .O(N__41107),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNI0VSNZ0Z_1 ));
    InMux I__9150 (
            .O(N__41104),
            .I(N__41101));
    LocalMux I__9149 (
            .O(N__41101),
            .I(N__41098));
    Span4Mux_h I__9148 (
            .O(N__41098),
            .I(N__41095));
    Span4Mux_v I__9147 (
            .O(N__41095),
            .I(N__41092));
    Span4Mux_h I__9146 (
            .O(N__41092),
            .I(N__41089));
    Span4Mux_h I__9145 (
            .O(N__41089),
            .I(N__41086));
    Odrv4 I__9144 (
            .O(N__41086),
            .I(\u0.N_1971 ));
    InMux I__9143 (
            .O(N__41083),
            .I(N__41080));
    LocalMux I__9142 (
            .O(N__41080),
            .I(\u0.N_1970 ));
    CascadeMux I__9141 (
            .O(N__41077),
            .I(N__41074));
    InMux I__9140 (
            .O(N__41074),
            .I(N__41071));
    LocalMux I__9139 (
            .O(N__41071),
            .I(\u0.dat_o_0_0_6_6 ));
    InMux I__9138 (
            .O(N__41068),
            .I(N__41065));
    LocalMux I__9137 (
            .O(N__41065),
            .I(\u0.dat_o_0_0_2_6 ));
    IoInMux I__9136 (
            .O(N__41062),
            .I(N__41059));
    LocalMux I__9135 (
            .O(N__41059),
            .I(N__41056));
    Span4Mux_s1_v I__9134 (
            .O(N__41056),
            .I(N__41053));
    Sp12to4 I__9133 (
            .O(N__41053),
            .I(N__41050));
    Span12Mux_h I__9132 (
            .O(N__41050),
            .I(N__41047));
    Odrv12 I__9131 (
            .O(N__41047),
            .I(wb_dat_o_c_6));
    InMux I__9130 (
            .O(N__41044),
            .I(N__41041));
    LocalMux I__9129 (
            .O(N__41041),
            .I(N__41038));
    Span4Mux_v I__9128 (
            .O(N__41038),
            .I(N__41035));
    Span4Mux_h I__9127 (
            .O(N__41035),
            .I(N__41031));
    InMux I__9126 (
            .O(N__41034),
            .I(N__41028));
    Odrv4 I__9125 (
            .O(N__41031),
            .I(PIO_cmdport_T4_0));
    LocalMux I__9124 (
            .O(N__41028),
            .I(PIO_cmdport_T4_0));
    InMux I__9123 (
            .O(N__41023),
            .I(N__41020));
    LocalMux I__9122 (
            .O(N__41020),
            .I(N__41015));
    InMux I__9121 (
            .O(N__41019),
            .I(N__41012));
    InMux I__9120 (
            .O(N__41018),
            .I(N__41009));
    Span4Mux_h I__9119 (
            .O(N__41015),
            .I(N__41006));
    LocalMux I__9118 (
            .O(N__41012),
            .I(N__41001));
    LocalMux I__9117 (
            .O(N__41009),
            .I(N__41001));
    Span4Mux_v I__9116 (
            .O(N__41006),
            .I(N__40995));
    Span4Mux_v I__9115 (
            .O(N__41001),
            .I(N__40995));
    InMux I__9114 (
            .O(N__41000),
            .I(N__40991));
    Span4Mux_h I__9113 (
            .O(N__40995),
            .I(N__40988));
    InMux I__9112 (
            .O(N__40994),
            .I(N__40985));
    LocalMux I__9111 (
            .O(N__40991),
            .I(N__40982));
    Span4Mux_h I__9110 (
            .O(N__40988),
            .I(N__40977));
    LocalMux I__9109 (
            .O(N__40985),
            .I(N__40977));
    Span12Mux_v I__9108 (
            .O(N__40982),
            .I(N__40974));
    Span4Mux_v I__9107 (
            .O(N__40977),
            .I(N__40971));
    Span12Mux_h I__9106 (
            .O(N__40974),
            .I(N__40968));
    Span4Mux_h I__9105 (
            .O(N__40971),
            .I(N__40965));
    Odrv12 I__9104 (
            .O(N__40968),
            .I(wb_dat_i_c_16));
    Odrv4 I__9103 (
            .O(N__40965),
            .I(wb_dat_i_c_16));
    InMux I__9102 (
            .O(N__40960),
            .I(N__40957));
    LocalMux I__9101 (
            .O(N__40957),
            .I(\u0.CtrlRegZ0Z_16 ));
    InMux I__9100 (
            .O(N__40954),
            .I(N__40951));
    LocalMux I__9099 (
            .O(N__40951),
            .I(N__40948));
    Span4Mux_h I__9098 (
            .O(N__40948),
            .I(N__40945));
    Odrv4 I__9097 (
            .O(N__40945),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_16 ));
    InMux I__9096 (
            .O(N__40942),
            .I(N__40939));
    LocalMux I__9095 (
            .O(N__40939),
            .I(N__40936));
    Span12Mux_h I__9094 (
            .O(N__40936),
            .I(N__40933));
    Odrv12 I__9093 (
            .O(N__40933),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_16 ));
    InMux I__9092 (
            .O(N__40930),
            .I(N__40927));
    LocalMux I__9091 (
            .O(N__40927),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIUM0RZ0Z_22 ));
    InMux I__9090 (
            .O(N__40924),
            .I(N__40921));
    LocalMux I__9089 (
            .O(N__40921),
            .I(N__40918));
    Span4Mux_h I__9088 (
            .O(N__40918),
            .I(N__40915));
    Span4Mux_v I__9087 (
            .O(N__40915),
            .I(N__40912));
    Span4Mux_h I__9086 (
            .O(N__40912),
            .I(N__40909));
    Odrv4 I__9085 (
            .O(N__40909),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI2B9KZ0Z_22 ));
    InMux I__9084 (
            .O(N__40906),
            .I(N__40903));
    LocalMux I__9083 (
            .O(N__40903),
            .I(mem_mem_ram6__RNI4SD71_22));
    CascadeMux I__9082 (
            .O(N__40900),
            .I(iQ_RNIICHM1_2_cascade_));
    InMux I__9081 (
            .O(N__40897),
            .I(N__40894));
    LocalMux I__9080 (
            .O(N__40894),
            .I(\u0.N_1719 ));
    InMux I__9079 (
            .O(N__40891),
            .I(N__40888));
    LocalMux I__9078 (
            .O(N__40888),
            .I(N__40885));
    Span4Mux_v I__9077 (
            .O(N__40885),
            .I(N__40882));
    Span4Mux_v I__9076 (
            .O(N__40882),
            .I(N__40879));
    Span4Mux_h I__9075 (
            .O(N__40879),
            .I(N__40876));
    Odrv4 I__9074 (
            .O(N__40876),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI8F7KZ0Z_16 ));
    InMux I__9073 (
            .O(N__40873),
            .I(N__40868));
    InMux I__9072 (
            .O(N__40872),
            .I(N__40864));
    InMux I__9071 (
            .O(N__40871),
            .I(N__40861));
    LocalMux I__9070 (
            .O(N__40868),
            .I(N__40858));
    InMux I__9069 (
            .O(N__40867),
            .I(N__40855));
    LocalMux I__9068 (
            .O(N__40864),
            .I(N__40851));
    LocalMux I__9067 (
            .O(N__40861),
            .I(N__40848));
    Span4Mux_v I__9066 (
            .O(N__40858),
            .I(N__40843));
    LocalMux I__9065 (
            .O(N__40855),
            .I(N__40843));
    InMux I__9064 (
            .O(N__40854),
            .I(N__40840));
    Span4Mux_v I__9063 (
            .O(N__40851),
            .I(N__40834));
    Span4Mux_h I__9062 (
            .O(N__40848),
            .I(N__40834));
    Span4Mux_h I__9061 (
            .O(N__40843),
            .I(N__40831));
    LocalMux I__9060 (
            .O(N__40840),
            .I(N__40828));
    InMux I__9059 (
            .O(N__40839),
            .I(N__40825));
    Span4Mux_h I__9058 (
            .O(N__40834),
            .I(N__40822));
    Sp12to4 I__9057 (
            .O(N__40831),
            .I(N__40819));
    Span4Mux_v I__9056 (
            .O(N__40828),
            .I(N__40816));
    LocalMux I__9055 (
            .O(N__40825),
            .I(N__40813));
    Sp12to4 I__9054 (
            .O(N__40822),
            .I(N__40807));
    Span12Mux_s10_v I__9053 (
            .O(N__40819),
            .I(N__40807));
    Span4Mux_h I__9052 (
            .O(N__40816),
            .I(N__40802));
    Span4Mux_v I__9051 (
            .O(N__40813),
            .I(N__40802));
    InMux I__9050 (
            .O(N__40812),
            .I(N__40799));
    Odrv12 I__9049 (
            .O(N__40807),
            .I(wb_dat_i_c_25));
    Odrv4 I__9048 (
            .O(N__40802),
            .I(wb_dat_i_c_25));
    LocalMux I__9047 (
            .O(N__40799),
            .I(wb_dat_i_c_25));
    InMux I__9046 (
            .O(N__40792),
            .I(N__40789));
    LocalMux I__9045 (
            .O(N__40789),
            .I(\u0.CtrlRegZ0Z_25 ));
    InMux I__9044 (
            .O(N__40786),
            .I(N__40783));
    LocalMux I__9043 (
            .O(N__40783),
            .I(N__40780));
    Span12Mux_v I__9042 (
            .O(N__40780),
            .I(N__40777));
    Odrv12 I__9041 (
            .O(N__40777),
            .I(DMAq_25));
    CascadeMux I__9040 (
            .O(N__40774),
            .I(N__40771));
    InMux I__9039 (
            .O(N__40771),
            .I(N__40768));
    LocalMux I__9038 (
            .O(N__40768),
            .I(N__40765));
    Sp12to4 I__9037 (
            .O(N__40765),
            .I(N__40762));
    Span12Mux_h I__9036 (
            .O(N__40762),
            .I(N__40758));
    InMux I__9035 (
            .O(N__40761),
            .I(N__40755));
    Odrv12 I__9034 (
            .O(N__40758),
            .I(DMA_dev0_Teoc_1));
    LocalMux I__9033 (
            .O(N__40755),
            .I(DMA_dev0_Teoc_1));
    InMux I__9032 (
            .O(N__40750),
            .I(N__40747));
    LocalMux I__9031 (
            .O(N__40747),
            .I(N__40743));
    InMux I__9030 (
            .O(N__40746),
            .I(N__40740));
    Odrv4 I__9029 (
            .O(N__40743),
            .I(DMA_dev0_Tm_6));
    LocalMux I__9028 (
            .O(N__40740),
            .I(DMA_dev0_Tm_6));
    CascadeMux I__9027 (
            .O(N__40735),
            .I(N__40732));
    InMux I__9026 (
            .O(N__40732),
            .I(N__40729));
    LocalMux I__9025 (
            .O(N__40729),
            .I(N__40726));
    Span4Mux_v I__9024 (
            .O(N__40726),
            .I(N__40722));
    CascadeMux I__9023 (
            .O(N__40725),
            .I(N__40719));
    Span4Mux_v I__9022 (
            .O(N__40722),
            .I(N__40716));
    InMux I__9021 (
            .O(N__40719),
            .I(N__40713));
    Odrv4 I__9020 (
            .O(N__40716),
            .I(PIO_dport1_T1_6));
    LocalMux I__9019 (
            .O(N__40713),
            .I(PIO_dport1_T1_6));
    CascadeMux I__9018 (
            .O(N__40708),
            .I(\u0.dat_o_0_0_0_6_cascade_ ));
    InMux I__9017 (
            .O(N__40705),
            .I(N__40702));
    LocalMux I__9016 (
            .O(N__40702),
            .I(N__40698));
    InMux I__9015 (
            .O(N__40701),
            .I(N__40695));
    Span4Mux_h I__9014 (
            .O(N__40698),
            .I(N__40692));
    LocalMux I__9013 (
            .O(N__40695),
            .I(DMA_dev1_Tm_6));
    Odrv4 I__9012 (
            .O(N__40692),
            .I(DMA_dev1_Tm_6));
    InMux I__9011 (
            .O(N__40687),
            .I(N__40684));
    LocalMux I__9010 (
            .O(N__40684),
            .I(N__40679));
    InMux I__9009 (
            .O(N__40683),
            .I(N__40674));
    InMux I__9008 (
            .O(N__40682),
            .I(N__40674));
    Span4Mux_v I__9007 (
            .O(N__40679),
            .I(N__40671));
    LocalMux I__9006 (
            .O(N__40674),
            .I(N__40668));
    Span4Mux_h I__9005 (
            .O(N__40671),
            .I(N__40663));
    Span4Mux_v I__9004 (
            .O(N__40668),
            .I(N__40663));
    Span4Mux_h I__9003 (
            .O(N__40663),
            .I(N__40660));
    Span4Mux_v I__9002 (
            .O(N__40660),
            .I(N__40657));
    Span4Mux_v I__9001 (
            .O(N__40657),
            .I(N__40654));
    Sp12to4 I__9000 (
            .O(N__40654),
            .I(N__40651));
    Odrv12 I__8999 (
            .O(N__40651),
            .I(dd_pad_i_c_6));
    InMux I__8998 (
            .O(N__40648),
            .I(N__40645));
    LocalMux I__8997 (
            .O(N__40645),
            .I(PIOq_6));
    InMux I__8996 (
            .O(N__40642),
            .I(N__40639));
    LocalMux I__8995 (
            .O(N__40639),
            .I(N__40636));
    Span4Mux_v I__8994 (
            .O(N__40636),
            .I(N__40633));
    Sp12to4 I__8993 (
            .O(N__40633),
            .I(N__40630));
    Span12Mux_h I__8992 (
            .O(N__40630),
            .I(N__40627));
    Odrv12 I__8991 (
            .O(N__40627),
            .I(\u0.N_1969 ));
    InMux I__8990 (
            .O(N__40624),
            .I(N__40620));
    InMux I__8989 (
            .O(N__40623),
            .I(N__40616));
    LocalMux I__8988 (
            .O(N__40620),
            .I(N__40613));
    InMux I__8987 (
            .O(N__40619),
            .I(N__40610));
    LocalMux I__8986 (
            .O(N__40616),
            .I(N__40607));
    Span4Mux_h I__8985 (
            .O(N__40613),
            .I(N__40604));
    LocalMux I__8984 (
            .O(N__40610),
            .I(N__40601));
    Span4Mux_h I__8983 (
            .O(N__40607),
            .I(N__40598));
    Span4Mux_h I__8982 (
            .O(N__40604),
            .I(N__40593));
    Span4Mux_v I__8981 (
            .O(N__40601),
            .I(N__40593));
    Odrv4 I__8980 (
            .O(N__40598),
            .I(IDEctrl_FATR1));
    Odrv4 I__8979 (
            .O(N__40593),
            .I(IDEctrl_FATR1));
    InMux I__8978 (
            .O(N__40588),
            .I(N__40585));
    LocalMux I__8977 (
            .O(N__40585),
            .I(N__40582));
    Span4Mux_v I__8976 (
            .O(N__40582),
            .I(N__40579));
    Span4Mux_v I__8975 (
            .O(N__40579),
            .I(N__40575));
    InMux I__8974 (
            .O(N__40578),
            .I(N__40572));
    Span4Mux_h I__8973 (
            .O(N__40575),
            .I(N__40567));
    LocalMux I__8972 (
            .O(N__40572),
            .I(N__40567));
    Span4Mux_v I__8971 (
            .O(N__40567),
            .I(N__40564));
    Odrv4 I__8970 (
            .O(N__40564),
            .I(PIO_cmdport_T1_6));
    InMux I__8969 (
            .O(N__40561),
            .I(N__40558));
    LocalMux I__8968 (
            .O(N__40558),
            .I(N__40554));
    InMux I__8967 (
            .O(N__40557),
            .I(N__40551));
    Span4Mux_h I__8966 (
            .O(N__40554),
            .I(N__40548));
    LocalMux I__8965 (
            .O(N__40551),
            .I(N__40545));
    Span4Mux_h I__8964 (
            .O(N__40548),
            .I(N__40542));
    Odrv12 I__8963 (
            .O(N__40545),
            .I(PIO_dport0_T1_6));
    Odrv4 I__8962 (
            .O(N__40542),
            .I(PIO_dport0_T1_6));
    InMux I__8961 (
            .O(N__40537),
            .I(N__40534));
    LocalMux I__8960 (
            .O(N__40534),
            .I(\u0.dat_o_0_0_3_6 ));
    InMux I__8959 (
            .O(N__40531),
            .I(N__40528));
    LocalMux I__8958 (
            .O(N__40528),
            .I(N__40523));
    InMux I__8957 (
            .O(N__40527),
            .I(N__40520));
    InMux I__8956 (
            .O(N__40526),
            .I(N__40516));
    Span4Mux_h I__8955 (
            .O(N__40523),
            .I(N__40511));
    LocalMux I__8954 (
            .O(N__40520),
            .I(N__40511));
    InMux I__8953 (
            .O(N__40519),
            .I(N__40508));
    LocalMux I__8952 (
            .O(N__40516),
            .I(N__40505));
    Span4Mux_h I__8951 (
            .O(N__40511),
            .I(N__40497));
    LocalMux I__8950 (
            .O(N__40508),
            .I(N__40497));
    Span4Mux_h I__8949 (
            .O(N__40505),
            .I(N__40497));
    InMux I__8948 (
            .O(N__40504),
            .I(N__40494));
    Span4Mux_v I__8947 (
            .O(N__40497),
            .I(N__40489));
    LocalMux I__8946 (
            .O(N__40494),
            .I(N__40489));
    Span4Mux_v I__8945 (
            .O(N__40489),
            .I(N__40484));
    InMux I__8944 (
            .O(N__40488),
            .I(N__40481));
    InMux I__8943 (
            .O(N__40487),
            .I(N__40478));
    Sp12to4 I__8942 (
            .O(N__40484),
            .I(N__40475));
    LocalMux I__8941 (
            .O(N__40481),
            .I(N__40472));
    LocalMux I__8940 (
            .O(N__40478),
            .I(N__40469));
    Span12Mux_h I__8939 (
            .O(N__40475),
            .I(N__40466));
    Span4Mux_v I__8938 (
            .O(N__40472),
            .I(N__40463));
    Span4Mux_v I__8937 (
            .O(N__40469),
            .I(N__40460));
    Odrv12 I__8936 (
            .O(N__40466),
            .I(wb_dat_i_c_31));
    Odrv4 I__8935 (
            .O(N__40463),
            .I(wb_dat_i_c_31));
    Odrv4 I__8934 (
            .O(N__40460),
            .I(wb_dat_i_c_31));
    InMux I__8933 (
            .O(N__40453),
            .I(N__40450));
    LocalMux I__8932 (
            .O(N__40450),
            .I(N__40447));
    Span4Mux_h I__8931 (
            .O(N__40447),
            .I(N__40444));
    Span4Mux_h I__8930 (
            .O(N__40444),
            .I(N__40441));
    Odrv4 I__8929 (
            .O(N__40441),
            .I(DMAq_31));
    InMux I__8928 (
            .O(N__40438),
            .I(N__40435));
    LocalMux I__8927 (
            .O(N__40435),
            .I(N__40431));
    InMux I__8926 (
            .O(N__40434),
            .I(N__40428));
    Span12Mux_h I__8925 (
            .O(N__40431),
            .I(N__40425));
    LocalMux I__8924 (
            .O(N__40428),
            .I(N__40422));
    Span12Mux_h I__8923 (
            .O(N__40425),
            .I(N__40419));
    Span4Mux_h I__8922 (
            .O(N__40422),
            .I(N__40416));
    Odrv12 I__8921 (
            .O(N__40419),
            .I(DMA_dev0_Teoc_7));
    Odrv4 I__8920 (
            .O(N__40416),
            .I(DMA_dev0_Teoc_7));
    CascadeMux I__8919 (
            .O(N__40411),
            .I(\u0.dat_o_i_i_0_31_cascade_ ));
    InMux I__8918 (
            .O(N__40408),
            .I(N__40405));
    LocalMux I__8917 (
            .O(N__40405),
            .I(N__40402));
    Span4Mux_v I__8916 (
            .O(N__40402),
            .I(N__40399));
    Sp12to4 I__8915 (
            .O(N__40399),
            .I(N__40395));
    InMux I__8914 (
            .O(N__40398),
            .I(N__40392));
    Span12Mux_s6_h I__8913 (
            .O(N__40395),
            .I(N__40389));
    LocalMux I__8912 (
            .O(N__40392),
            .I(DMA_dev1_Teoc_7));
    Odrv12 I__8911 (
            .O(N__40389),
            .I(DMA_dev1_Teoc_7));
    IoInMux I__8910 (
            .O(N__40384),
            .I(N__40381));
    LocalMux I__8909 (
            .O(N__40381),
            .I(N__40378));
    IoSpan4Mux I__8908 (
            .O(N__40378),
            .I(N__40375));
    Span4Mux_s3_v I__8907 (
            .O(N__40375),
            .I(N__40372));
    Span4Mux_v I__8906 (
            .O(N__40372),
            .I(N__40369));
    Span4Mux_v I__8905 (
            .O(N__40369),
            .I(N__40366));
    Odrv4 I__8904 (
            .O(N__40366),
            .I(N_277));
    InMux I__8903 (
            .O(N__40363),
            .I(N__40359));
    InMux I__8902 (
            .O(N__40362),
            .I(N__40356));
    LocalMux I__8901 (
            .O(N__40359),
            .I(N__40353));
    LocalMux I__8900 (
            .O(N__40356),
            .I(PIO_dport1_Teoc_7));
    Odrv12 I__8899 (
            .O(N__40353),
            .I(PIO_dport1_Teoc_7));
    InMux I__8898 (
            .O(N__40348),
            .I(N__40345));
    LocalMux I__8897 (
            .O(N__40345),
            .I(\u0.CtrlRegZ0Z_31 ));
    InMux I__8896 (
            .O(N__40342),
            .I(N__40338));
    InMux I__8895 (
            .O(N__40341),
            .I(N__40335));
    LocalMux I__8894 (
            .O(N__40338),
            .I(N__40332));
    LocalMux I__8893 (
            .O(N__40335),
            .I(N__40329));
    Span4Mux_v I__8892 (
            .O(N__40332),
            .I(N__40326));
    Span4Mux_v I__8891 (
            .O(N__40329),
            .I(N__40323));
    Odrv4 I__8890 (
            .O(N__40326),
            .I(PIO_cmdport_Teoc_7));
    Odrv4 I__8889 (
            .O(N__40323),
            .I(PIO_cmdport_Teoc_7));
    InMux I__8888 (
            .O(N__40318),
            .I(N__40315));
    LocalMux I__8887 (
            .O(N__40315),
            .I(\u0.N_1710 ));
    CascadeMux I__8886 (
            .O(N__40312),
            .I(\u0.dat_o_i_i_1_31_cascade_ ));
    InMux I__8885 (
            .O(N__40309),
            .I(N__40306));
    LocalMux I__8884 (
            .O(N__40306),
            .I(N__40302));
    InMux I__8883 (
            .O(N__40305),
            .I(N__40299));
    Span4Mux_v I__8882 (
            .O(N__40302),
            .I(N__40296));
    LocalMux I__8881 (
            .O(N__40299),
            .I(N__40293));
    Odrv4 I__8880 (
            .O(N__40296),
            .I(PIO_dport0_Teoc_7));
    Odrv12 I__8879 (
            .O(N__40293),
            .I(PIO_dport0_Teoc_7));
    InMux I__8878 (
            .O(N__40288),
            .I(N__40285));
    LocalMux I__8877 (
            .O(N__40285),
            .I(\u0.dat_o_i_i_4_31 ));
    InMux I__8876 (
            .O(N__40282),
            .I(N__40279));
    LocalMux I__8875 (
            .O(N__40279),
            .I(N__40276));
    Span4Mux_v I__8874 (
            .O(N__40276),
            .I(N__40272));
    InMux I__8873 (
            .O(N__40275),
            .I(N__40269));
    Odrv4 I__8872 (
            .O(N__40272),
            .I(PIO_cmdport_Teoc_1));
    LocalMux I__8871 (
            .O(N__40269),
            .I(PIO_cmdport_Teoc_1));
    CascadeMux I__8870 (
            .O(N__40264),
            .I(\u0.dat_o_i_i_1_25_cascade_ ));
    InMux I__8869 (
            .O(N__40261),
            .I(N__40257));
    InMux I__8868 (
            .O(N__40260),
            .I(N__40254));
    LocalMux I__8867 (
            .O(N__40257),
            .I(N__40251));
    LocalMux I__8866 (
            .O(N__40254),
            .I(N__40248));
    Span4Mux_v I__8865 (
            .O(N__40251),
            .I(N__40243));
    Span4Mux_v I__8864 (
            .O(N__40248),
            .I(N__40243));
    Odrv4 I__8863 (
            .O(N__40243),
            .I(PIO_dport0_Teoc_1));
    CascadeMux I__8862 (
            .O(N__40240),
            .I(N__40236));
    InMux I__8861 (
            .O(N__40239),
            .I(N__40233));
    InMux I__8860 (
            .O(N__40236),
            .I(N__40230));
    LocalMux I__8859 (
            .O(N__40233),
            .I(N__40227));
    LocalMux I__8858 (
            .O(N__40230),
            .I(N__40224));
    Span4Mux_v I__8857 (
            .O(N__40227),
            .I(N__40221));
    Span4Mux_h I__8856 (
            .O(N__40224),
            .I(N__40218));
    Odrv4 I__8855 (
            .O(N__40221),
            .I(PIO_dport1_Teoc_1));
    Odrv4 I__8854 (
            .O(N__40218),
            .I(PIO_dport1_Teoc_1));
    InMux I__8853 (
            .O(N__40213),
            .I(N__40210));
    LocalMux I__8852 (
            .O(N__40210),
            .I(\u0.N_1668 ));
    CascadeMux I__8851 (
            .O(N__40207),
            .I(\u0.dat_o_i_i_3_10_cascade_ ));
    InMux I__8850 (
            .O(N__40204),
            .I(N__40201));
    LocalMux I__8849 (
            .O(N__40201),
            .I(N__40198));
    Span4Mux_v I__8848 (
            .O(N__40198),
            .I(N__40194));
    InMux I__8847 (
            .O(N__40197),
            .I(N__40191));
    Odrv4 I__8846 (
            .O(N__40194),
            .I(PIO_dport0_T2_2));
    LocalMux I__8845 (
            .O(N__40191),
            .I(PIO_dport0_T2_2));
    InMux I__8844 (
            .O(N__40186),
            .I(N__40182));
    InMux I__8843 (
            .O(N__40185),
            .I(N__40179));
    LocalMux I__8842 (
            .O(N__40182),
            .I(N__40174));
    LocalMux I__8841 (
            .O(N__40179),
            .I(N__40174));
    Span4Mux_v I__8840 (
            .O(N__40174),
            .I(N__40169));
    InMux I__8839 (
            .O(N__40173),
            .I(N__40163));
    InMux I__8838 (
            .O(N__40172),
            .I(N__40160));
    Span4Mux_h I__8837 (
            .O(N__40169),
            .I(N__40157));
    InMux I__8836 (
            .O(N__40168),
            .I(N__40154));
    InMux I__8835 (
            .O(N__40167),
            .I(N__40151));
    InMux I__8834 (
            .O(N__40166),
            .I(N__40148));
    LocalMux I__8833 (
            .O(N__40163),
            .I(N__40145));
    LocalMux I__8832 (
            .O(N__40160),
            .I(N__40142));
    Span4Mux_v I__8831 (
            .O(N__40157),
            .I(N__40135));
    LocalMux I__8830 (
            .O(N__40154),
            .I(N__40135));
    LocalMux I__8829 (
            .O(N__40151),
            .I(N__40135));
    LocalMux I__8828 (
            .O(N__40148),
            .I(N__40132));
    Span4Mux_v I__8827 (
            .O(N__40145),
            .I(N__40129));
    Span4Mux_v I__8826 (
            .O(N__40142),
            .I(N__40123));
    Span4Mux_h I__8825 (
            .O(N__40135),
            .I(N__40123));
    Span4Mux_v I__8824 (
            .O(N__40132),
            .I(N__40119));
    Sp12to4 I__8823 (
            .O(N__40129),
            .I(N__40116));
    InMux I__8822 (
            .O(N__40128),
            .I(N__40113));
    Span4Mux_v I__8821 (
            .O(N__40123),
            .I(N__40110));
    InMux I__8820 (
            .O(N__40122),
            .I(N__40107));
    Sp12to4 I__8819 (
            .O(N__40119),
            .I(N__40100));
    Span12Mux_h I__8818 (
            .O(N__40116),
            .I(N__40100));
    LocalMux I__8817 (
            .O(N__40113),
            .I(N__40100));
    Span4Mux_v I__8816 (
            .O(N__40110),
            .I(N__40097));
    LocalMux I__8815 (
            .O(N__40107),
            .I(N__40094));
    Span12Mux_h I__8814 (
            .O(N__40100),
            .I(N__40091));
    Span4Mux_v I__8813 (
            .O(N__40097),
            .I(N__40088));
    Span4Mux_v I__8812 (
            .O(N__40094),
            .I(N__40085));
    Span12Mux_v I__8811 (
            .O(N__40091),
            .I(N__40082));
    Span4Mux_h I__8810 (
            .O(N__40088),
            .I(N__40079));
    IoSpan4Mux I__8809 (
            .O(N__40085),
            .I(N__40076));
    Odrv12 I__8808 (
            .O(N__40082),
            .I(wb_dat_i_c_10));
    Odrv4 I__8807 (
            .O(N__40079),
            .I(wb_dat_i_c_10));
    Odrv4 I__8806 (
            .O(N__40076),
            .I(wb_dat_i_c_10));
    InMux I__8805 (
            .O(N__40069),
            .I(N__40066));
    LocalMux I__8804 (
            .O(N__40066),
            .I(\u0.CtrlRegZ0Z_10 ));
    InMux I__8803 (
            .O(N__40063),
            .I(N__40060));
    LocalMux I__8802 (
            .O(N__40060),
            .I(N__40057));
    Span12Mux_h I__8801 (
            .O(N__40057),
            .I(N__40053));
    InMux I__8800 (
            .O(N__40056),
            .I(N__40050));
    Odrv12 I__8799 (
            .O(N__40053),
            .I(DMA_dev0_Td_2));
    LocalMux I__8798 (
            .O(N__40050),
            .I(DMA_dev0_Td_2));
    InMux I__8797 (
            .O(N__40045),
            .I(N__40042));
    LocalMux I__8796 (
            .O(N__40042),
            .I(N__40039));
    Span12Mux_v I__8795 (
            .O(N__40039),
            .I(N__40036));
    Odrv12 I__8794 (
            .O(N__40036),
            .I(\u0.N_1989 ));
    InMux I__8793 (
            .O(N__40033),
            .I(N__40030));
    LocalMux I__8792 (
            .O(N__40030),
            .I(N__40027));
    Span12Mux_h I__8791 (
            .O(N__40027),
            .I(N__40024));
    Odrv12 I__8790 (
            .O(N__40024),
            .I(\u0.dat_o_i_i_2Z0Z_10 ));
    CascadeMux I__8789 (
            .O(N__40021),
            .I(\u0.N_1990_cascade_ ));
    InMux I__8788 (
            .O(N__40018),
            .I(N__40015));
    LocalMux I__8787 (
            .O(N__40015),
            .I(\u0.dat_o_i_i_6_10 ));
    IoInMux I__8786 (
            .O(N__40012),
            .I(N__40009));
    LocalMux I__8785 (
            .O(N__40009),
            .I(N__40006));
    Span4Mux_s2_v I__8784 (
            .O(N__40006),
            .I(N__40003));
    Span4Mux_v I__8783 (
            .O(N__40003),
            .I(N__40000));
    Span4Mux_v I__8782 (
            .O(N__40000),
            .I(N__39997));
    Odrv4 I__8781 (
            .O(N__39997),
            .I(N_1097));
    InMux I__8780 (
            .O(N__39994),
            .I(N__39990));
    InMux I__8779 (
            .O(N__39993),
            .I(N__39987));
    LocalMux I__8778 (
            .O(N__39990),
            .I(N__39984));
    LocalMux I__8777 (
            .O(N__39987),
            .I(N__39981));
    Span4Mux_h I__8776 (
            .O(N__39984),
            .I(N__39976));
    Span4Mux_h I__8775 (
            .O(N__39981),
            .I(N__39976));
    Odrv4 I__8774 (
            .O(N__39976),
            .I(PIO_dport1_Teoc_0));
    CascadeMux I__8773 (
            .O(N__39973),
            .I(\u0.N_1661_cascade_ ));
    InMux I__8772 (
            .O(N__39970),
            .I(N__39967));
    LocalMux I__8771 (
            .O(N__39967),
            .I(N__39964));
    Span4Mux_v I__8770 (
            .O(N__39964),
            .I(N__39960));
    InMux I__8769 (
            .O(N__39963),
            .I(N__39957));
    Span4Mux_h I__8768 (
            .O(N__39960),
            .I(N__39952));
    LocalMux I__8767 (
            .O(N__39957),
            .I(N__39952));
    Odrv4 I__8766 (
            .O(N__39952),
            .I(PIO_dport0_Teoc_0));
    InMux I__8765 (
            .O(N__39949),
            .I(N__39945));
    InMux I__8764 (
            .O(N__39948),
            .I(N__39942));
    LocalMux I__8763 (
            .O(N__39945),
            .I(N__39939));
    LocalMux I__8762 (
            .O(N__39942),
            .I(N__39936));
    Span4Mux_h I__8761 (
            .O(N__39939),
            .I(N__39933));
    Odrv4 I__8760 (
            .O(N__39936),
            .I(PIO_cmdport_Teoc_0));
    Odrv4 I__8759 (
            .O(N__39933),
            .I(PIO_cmdport_Teoc_0));
    InMux I__8758 (
            .O(N__39928),
            .I(N__39925));
    LocalMux I__8757 (
            .O(N__39925),
            .I(\u0.dat_o_i_i_1_24 ));
    InMux I__8756 (
            .O(N__39922),
            .I(N__39917));
    InMux I__8755 (
            .O(N__39921),
            .I(N__39914));
    InMux I__8754 (
            .O(N__39920),
            .I(N__39911));
    LocalMux I__8753 (
            .O(N__39917),
            .I(N__39908));
    LocalMux I__8752 (
            .O(N__39914),
            .I(N__39904));
    LocalMux I__8751 (
            .O(N__39911),
            .I(N__39901));
    Span4Mux_v I__8750 (
            .O(N__39908),
            .I(N__39898));
    InMux I__8749 (
            .O(N__39907),
            .I(N__39895));
    Span4Mux_v I__8748 (
            .O(N__39904),
            .I(N__39892));
    Span4Mux_v I__8747 (
            .O(N__39901),
            .I(N__39889));
    Span4Mux_h I__8746 (
            .O(N__39898),
            .I(N__39884));
    LocalMux I__8745 (
            .O(N__39895),
            .I(N__39884));
    Span4Mux_h I__8744 (
            .O(N__39892),
            .I(N__39880));
    Span4Mux_v I__8743 (
            .O(N__39889),
            .I(N__39875));
    Span4Mux_h I__8742 (
            .O(N__39884),
            .I(N__39872));
    InMux I__8741 (
            .O(N__39883),
            .I(N__39869));
    Span4Mux_h I__8740 (
            .O(N__39880),
            .I(N__39866));
    InMux I__8739 (
            .O(N__39879),
            .I(N__39863));
    InMux I__8738 (
            .O(N__39878),
            .I(N__39860));
    Span4Mux_v I__8737 (
            .O(N__39875),
            .I(N__39857));
    Span4Mux_v I__8736 (
            .O(N__39872),
            .I(N__39852));
    LocalMux I__8735 (
            .O(N__39869),
            .I(N__39852));
    Span4Mux_h I__8734 (
            .O(N__39866),
            .I(N__39847));
    LocalMux I__8733 (
            .O(N__39863),
            .I(N__39847));
    LocalMux I__8732 (
            .O(N__39860),
            .I(N__39844));
    Span4Mux_v I__8731 (
            .O(N__39857),
            .I(N__39841));
    Span4Mux_h I__8730 (
            .O(N__39852),
            .I(N__39838));
    Span4Mux_v I__8729 (
            .O(N__39847),
            .I(N__39835));
    Span4Mux_v I__8728 (
            .O(N__39844),
            .I(N__39832));
    Span4Mux_h I__8727 (
            .O(N__39841),
            .I(N__39829));
    Sp12to4 I__8726 (
            .O(N__39838),
            .I(N__39826));
    Span4Mux_h I__8725 (
            .O(N__39835),
            .I(N__39821));
    Span4Mux_v I__8724 (
            .O(N__39832),
            .I(N__39821));
    Sp12to4 I__8723 (
            .O(N__39829),
            .I(N__39818));
    Span12Mux_v I__8722 (
            .O(N__39826),
            .I(N__39815));
    Span4Mux_v I__8721 (
            .O(N__39821),
            .I(N__39812));
    Odrv12 I__8720 (
            .O(N__39818),
            .I(wb_dat_i_c_24));
    Odrv12 I__8719 (
            .O(N__39815),
            .I(wb_dat_i_c_24));
    Odrv4 I__8718 (
            .O(N__39812),
            .I(wb_dat_i_c_24));
    InMux I__8717 (
            .O(N__39805),
            .I(N__39802));
    LocalMux I__8716 (
            .O(N__39802),
            .I(\u0.CtrlRegZ0Z_24 ));
    CascadeMux I__8715 (
            .O(N__39799),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIC5ITZ0Z_25_cascade_ ));
    InMux I__8714 (
            .O(N__39796),
            .I(N__39793));
    LocalMux I__8713 (
            .O(N__39793),
            .I(N__39790));
    Odrv4 I__8712 (
            .O(N__39790),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_25 ));
    InMux I__8711 (
            .O(N__39787),
            .I(N__39784));
    LocalMux I__8710 (
            .O(N__39784),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNID5E71Z0Z_25 ));
    InMux I__8709 (
            .O(N__39781),
            .I(N__39778));
    LocalMux I__8708 (
            .O(N__39778),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI2PFTZ0Z_11 ));
    CascadeMux I__8707 (
            .O(N__39775),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIUIA71Z0Z_11_cascade_ ));
    InMux I__8706 (
            .O(N__39772),
            .I(N__39769));
    LocalMux I__8705 (
            .O(N__39769),
            .I(N__39766));
    Odrv4 I__8704 (
            .O(N__39766),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIA0DM1Z0Z_2 ));
    InMux I__8703 (
            .O(N__39763),
            .I(N__39760));
    LocalMux I__8702 (
            .O(N__39760),
            .I(N__39757));
    Span4Mux_v I__8701 (
            .O(N__39757),
            .I(N__39754));
    Sp12to4 I__8700 (
            .O(N__39754),
            .I(N__39750));
    InMux I__8699 (
            .O(N__39753),
            .I(N__39747));
    Odrv12 I__8698 (
            .O(N__39750),
            .I(DMA_dev0_Tm_7));
    LocalMux I__8697 (
            .O(N__39747),
            .I(DMA_dev0_Tm_7));
    CEMux I__8696 (
            .O(N__39742),
            .I(N__39737));
    CEMux I__8695 (
            .O(N__39741),
            .I(N__39733));
    CEMux I__8694 (
            .O(N__39740),
            .I(N__39730));
    LocalMux I__8693 (
            .O(N__39737),
            .I(N__39727));
    CEMux I__8692 (
            .O(N__39736),
            .I(N__39724));
    LocalMux I__8691 (
            .O(N__39733),
            .I(N__39720));
    LocalMux I__8690 (
            .O(N__39730),
            .I(N__39717));
    Span4Mux_v I__8689 (
            .O(N__39727),
            .I(N__39714));
    LocalMux I__8688 (
            .O(N__39724),
            .I(N__39711));
    CEMux I__8687 (
            .O(N__39723),
            .I(N__39708));
    Span4Mux_v I__8686 (
            .O(N__39720),
            .I(N__39705));
    Span4Mux_v I__8685 (
            .O(N__39717),
            .I(N__39702));
    Span4Mux_h I__8684 (
            .O(N__39714),
            .I(N__39697));
    Span4Mux_v I__8683 (
            .O(N__39711),
            .I(N__39697));
    LocalMux I__8682 (
            .O(N__39708),
            .I(N__39694));
    Span4Mux_h I__8681 (
            .O(N__39705),
            .I(N__39690));
    Span4Mux_v I__8680 (
            .O(N__39702),
            .I(N__39685));
    Span4Mux_v I__8679 (
            .O(N__39697),
            .I(N__39685));
    Span4Mux_v I__8678 (
            .O(N__39694),
            .I(N__39682));
    CEMux I__8677 (
            .O(N__39693),
            .I(N__39679));
    Span4Mux_v I__8676 (
            .O(N__39690),
            .I(N__39676));
    Span4Mux_h I__8675 (
            .O(N__39685),
            .I(N__39671));
    Span4Mux_h I__8674 (
            .O(N__39682),
            .I(N__39671));
    LocalMux I__8673 (
            .O(N__39679),
            .I(N__39668));
    Odrv4 I__8672 (
            .O(N__39676),
            .I(\u0.N_444 ));
    Odrv4 I__8671 (
            .O(N__39671),
            .I(\u0.N_444 ));
    Odrv4 I__8670 (
            .O(N__39668),
            .I(\u0.N_444 ));
    InMux I__8669 (
            .O(N__39661),
            .I(N__39658));
    LocalMux I__8668 (
            .O(N__39658),
            .I(N__39654));
    InMux I__8667 (
            .O(N__39657),
            .I(N__39651));
    Span4Mux_v I__8666 (
            .O(N__39654),
            .I(N__39644));
    LocalMux I__8665 (
            .O(N__39651),
            .I(N__39644));
    InMux I__8664 (
            .O(N__39650),
            .I(N__39641));
    InMux I__8663 (
            .O(N__39649),
            .I(N__39637));
    Span4Mux_h I__8662 (
            .O(N__39644),
            .I(N__39632));
    LocalMux I__8661 (
            .O(N__39641),
            .I(N__39632));
    InMux I__8660 (
            .O(N__39640),
            .I(N__39629));
    LocalMux I__8659 (
            .O(N__39637),
            .I(N__39625));
    Sp12to4 I__8658 (
            .O(N__39632),
            .I(N__39621));
    LocalMux I__8657 (
            .O(N__39629),
            .I(N__39618));
    InMux I__8656 (
            .O(N__39628),
            .I(N__39615));
    Span4Mux_v I__8655 (
            .O(N__39625),
            .I(N__39611));
    InMux I__8654 (
            .O(N__39624),
            .I(N__39608));
    Span12Mux_v I__8653 (
            .O(N__39621),
            .I(N__39604));
    Span4Mux_v I__8652 (
            .O(N__39618),
            .I(N__39601));
    LocalMux I__8651 (
            .O(N__39615),
            .I(N__39598));
    InMux I__8650 (
            .O(N__39614),
            .I(N__39595));
    Sp12to4 I__8649 (
            .O(N__39611),
            .I(N__39592));
    LocalMux I__8648 (
            .O(N__39608),
            .I(N__39589));
    InMux I__8647 (
            .O(N__39607),
            .I(N__39586));
    Span12Mux_h I__8646 (
            .O(N__39604),
            .I(N__39583));
    Sp12to4 I__8645 (
            .O(N__39601),
            .I(N__39576));
    Span12Mux_v I__8644 (
            .O(N__39598),
            .I(N__39576));
    LocalMux I__8643 (
            .O(N__39595),
            .I(N__39576));
    Span12Mux_h I__8642 (
            .O(N__39592),
            .I(N__39569));
    Span12Mux_v I__8641 (
            .O(N__39589),
            .I(N__39569));
    LocalMux I__8640 (
            .O(N__39586),
            .I(N__39569));
    Span12Mux_h I__8639 (
            .O(N__39583),
            .I(N__39566));
    Span12Mux_h I__8638 (
            .O(N__39576),
            .I(N__39563));
    Span12Mux_h I__8637 (
            .O(N__39569),
            .I(N__39560));
    Odrv12 I__8636 (
            .O(N__39566),
            .I(wb_dat_i_c_7));
    Odrv12 I__8635 (
            .O(N__39563),
            .I(wb_dat_i_c_7));
    Odrv12 I__8634 (
            .O(N__39560),
            .I(wb_dat_i_c_7));
    InMux I__8633 (
            .O(N__39553),
            .I(N__39547));
    InMux I__8632 (
            .O(N__39552),
            .I(N__39547));
    LocalMux I__8631 (
            .O(N__39547),
            .I(DMA_dev1_Tm_7));
    CEMux I__8630 (
            .O(N__39544),
            .I(N__39539));
    CEMux I__8629 (
            .O(N__39543),
            .I(N__39536));
    CEMux I__8628 (
            .O(N__39542),
            .I(N__39533));
    LocalMux I__8627 (
            .O(N__39539),
            .I(N__39529));
    LocalMux I__8626 (
            .O(N__39536),
            .I(N__39526));
    LocalMux I__8625 (
            .O(N__39533),
            .I(N__39523));
    CEMux I__8624 (
            .O(N__39532),
            .I(N__39520));
    Span4Mux_v I__8623 (
            .O(N__39529),
            .I(N__39517));
    Span4Mux_h I__8622 (
            .O(N__39526),
            .I(N__39512));
    Span4Mux_v I__8621 (
            .O(N__39523),
            .I(N__39512));
    LocalMux I__8620 (
            .O(N__39520),
            .I(N__39509));
    Span4Mux_h I__8619 (
            .O(N__39517),
            .I(N__39506));
    Span4Mux_v I__8618 (
            .O(N__39512),
            .I(N__39503));
    Span4Mux_v I__8617 (
            .O(N__39509),
            .I(N__39500));
    Span4Mux_v I__8616 (
            .O(N__39506),
            .I(N__39495));
    Span4Mux_h I__8615 (
            .O(N__39503),
            .I(N__39495));
    Span4Mux_v I__8614 (
            .O(N__39500),
            .I(N__39492));
    Odrv4 I__8613 (
            .O(N__39495),
            .I(\u0.N_442 ));
    Odrv4 I__8612 (
            .O(N__39492),
            .I(\u0.N_442 ));
    InMux I__8611 (
            .O(N__39487),
            .I(N__39484));
    LocalMux I__8610 (
            .O(N__39484),
            .I(N__39481));
    Span4Mux_v I__8609 (
            .O(N__39481),
            .I(N__39477));
    InMux I__8608 (
            .O(N__39480),
            .I(N__39472));
    Span4Mux_v I__8607 (
            .O(N__39477),
            .I(N__39468));
    InMux I__8606 (
            .O(N__39476),
            .I(N__39465));
    InMux I__8605 (
            .O(N__39475),
            .I(N__39462));
    LocalMux I__8604 (
            .O(N__39472),
            .I(N__39459));
    InMux I__8603 (
            .O(N__39471),
            .I(N__39456));
    Span4Mux_h I__8602 (
            .O(N__39468),
            .I(N__39450));
    LocalMux I__8601 (
            .O(N__39465),
            .I(N__39450));
    LocalMux I__8600 (
            .O(N__39462),
            .I(N__39446));
    Span4Mux_v I__8599 (
            .O(N__39459),
            .I(N__39443));
    LocalMux I__8598 (
            .O(N__39456),
            .I(N__39440));
    InMux I__8597 (
            .O(N__39455),
            .I(N__39437));
    Span4Mux_v I__8596 (
            .O(N__39450),
            .I(N__39434));
    InMux I__8595 (
            .O(N__39449),
            .I(N__39431));
    Span4Mux_v I__8594 (
            .O(N__39446),
            .I(N__39427));
    Span4Mux_h I__8593 (
            .O(N__39443),
            .I(N__39422));
    Span4Mux_v I__8592 (
            .O(N__39440),
            .I(N__39422));
    LocalMux I__8591 (
            .O(N__39437),
            .I(N__39418));
    Span4Mux_h I__8590 (
            .O(N__39434),
            .I(N__39415));
    LocalMux I__8589 (
            .O(N__39431),
            .I(N__39412));
    InMux I__8588 (
            .O(N__39430),
            .I(N__39409));
    Span4Mux_h I__8587 (
            .O(N__39427),
            .I(N__39406));
    Span4Mux_h I__8586 (
            .O(N__39422),
            .I(N__39403));
    InMux I__8585 (
            .O(N__39421),
            .I(N__39400));
    Span4Mux_v I__8584 (
            .O(N__39418),
            .I(N__39397));
    Span4Mux_h I__8583 (
            .O(N__39415),
            .I(N__39390));
    Span4Mux_v I__8582 (
            .O(N__39412),
            .I(N__39390));
    LocalMux I__8581 (
            .O(N__39409),
            .I(N__39390));
    Span4Mux_h I__8580 (
            .O(N__39406),
            .I(N__39387));
    Sp12to4 I__8579 (
            .O(N__39403),
            .I(N__39382));
    LocalMux I__8578 (
            .O(N__39400),
            .I(N__39382));
    Span4Mux_v I__8577 (
            .O(N__39397),
            .I(N__39377));
    Span4Mux_v I__8576 (
            .O(N__39390),
            .I(N__39377));
    Sp12to4 I__8575 (
            .O(N__39387),
            .I(N__39372));
    Span12Mux_h I__8574 (
            .O(N__39382),
            .I(N__39372));
    Sp12to4 I__8573 (
            .O(N__39377),
            .I(N__39369));
    Span12Mux_v I__8572 (
            .O(N__39372),
            .I(N__39366));
    Span12Mux_h I__8571 (
            .O(N__39369),
            .I(N__39363));
    Odrv12 I__8570 (
            .O(N__39366),
            .I(wb_dat_i_c_6));
    Odrv12 I__8569 (
            .O(N__39363),
            .I(wb_dat_i_c_6));
    InMux I__8568 (
            .O(N__39358),
            .I(N__39355));
    LocalMux I__8567 (
            .O(N__39355),
            .I(N__39349));
    InMux I__8566 (
            .O(N__39354),
            .I(N__39346));
    InMux I__8565 (
            .O(N__39353),
            .I(N__39342));
    InMux I__8564 (
            .O(N__39352),
            .I(N__39338));
    Span4Mux_v I__8563 (
            .O(N__39349),
            .I(N__39334));
    LocalMux I__8562 (
            .O(N__39346),
            .I(N__39331));
    InMux I__8561 (
            .O(N__39345),
            .I(N__39328));
    LocalMux I__8560 (
            .O(N__39342),
            .I(N__39325));
    InMux I__8559 (
            .O(N__39341),
            .I(N__39322));
    LocalMux I__8558 (
            .O(N__39338),
            .I(N__39319));
    InMux I__8557 (
            .O(N__39337),
            .I(N__39316));
    Span4Mux_h I__8556 (
            .O(N__39334),
            .I(N__39309));
    Span4Mux_v I__8555 (
            .O(N__39331),
            .I(N__39309));
    LocalMux I__8554 (
            .O(N__39328),
            .I(N__39309));
    Span4Mux_h I__8553 (
            .O(N__39325),
            .I(N__39305));
    LocalMux I__8552 (
            .O(N__39322),
            .I(N__39302));
    Span4Mux_h I__8551 (
            .O(N__39319),
            .I(N__39299));
    LocalMux I__8550 (
            .O(N__39316),
            .I(N__39296));
    Span4Mux_v I__8549 (
            .O(N__39309),
            .I(N__39292));
    InMux I__8548 (
            .O(N__39308),
            .I(N__39289));
    Span4Mux_v I__8547 (
            .O(N__39305),
            .I(N__39286));
    Span4Mux_v I__8546 (
            .O(N__39302),
            .I(N__39279));
    Span4Mux_v I__8545 (
            .O(N__39299),
            .I(N__39279));
    Span4Mux_h I__8544 (
            .O(N__39296),
            .I(N__39279));
    InMux I__8543 (
            .O(N__39295),
            .I(N__39276));
    Sp12to4 I__8542 (
            .O(N__39292),
            .I(N__39273));
    LocalMux I__8541 (
            .O(N__39289),
            .I(N__39270));
    Sp12to4 I__8540 (
            .O(N__39286),
            .I(N__39263));
    Sp12to4 I__8539 (
            .O(N__39279),
            .I(N__39263));
    LocalMux I__8538 (
            .O(N__39276),
            .I(N__39263));
    Span12Mux_h I__8537 (
            .O(N__39273),
            .I(N__39258));
    Span12Mux_v I__8536 (
            .O(N__39270),
            .I(N__39258));
    Span12Mux_v I__8535 (
            .O(N__39263),
            .I(N__39255));
    Span12Mux_v I__8534 (
            .O(N__39258),
            .I(N__39252));
    Span12Mux_h I__8533 (
            .O(N__39255),
            .I(N__39249));
    Span12Mux_h I__8532 (
            .O(N__39252),
            .I(N__39246));
    Odrv12 I__8531 (
            .O(N__39249),
            .I(wb_dat_i_c_1));
    Odrv12 I__8530 (
            .O(N__39246),
            .I(wb_dat_i_c_1));
    CascadeMux I__8529 (
            .O(N__39241),
            .I(N__39238));
    InMux I__8528 (
            .O(N__39238),
            .I(N__39234));
    InMux I__8527 (
            .O(N__39237),
            .I(N__39231));
    LocalMux I__8526 (
            .O(N__39234),
            .I(N__39228));
    LocalMux I__8525 (
            .O(N__39231),
            .I(N__39225));
    Span4Mux_h I__8524 (
            .O(N__39228),
            .I(N__39222));
    Span4Mux_h I__8523 (
            .O(N__39225),
            .I(N__39219));
    Span4Mux_v I__8522 (
            .O(N__39222),
            .I(N__39216));
    Span4Mux_h I__8521 (
            .O(N__39219),
            .I(N__39213));
    Odrv4 I__8520 (
            .O(N__39216),
            .I(PIO_cmdport_IORDYen));
    Odrv4 I__8519 (
            .O(N__39213),
            .I(PIO_cmdport_IORDYen));
    CEMux I__8518 (
            .O(N__39208),
            .I(N__39202));
    CEMux I__8517 (
            .O(N__39207),
            .I(N__39198));
    CEMux I__8516 (
            .O(N__39206),
            .I(N__39195));
    CEMux I__8515 (
            .O(N__39205),
            .I(N__39192));
    LocalMux I__8514 (
            .O(N__39202),
            .I(N__39189));
    CEMux I__8513 (
            .O(N__39201),
            .I(N__39185));
    LocalMux I__8512 (
            .O(N__39198),
            .I(N__39180));
    LocalMux I__8511 (
            .O(N__39195),
            .I(N__39180));
    LocalMux I__8510 (
            .O(N__39192),
            .I(N__39177));
    Span4Mux_v I__8509 (
            .O(N__39189),
            .I(N__39174));
    CEMux I__8508 (
            .O(N__39188),
            .I(N__39171));
    LocalMux I__8507 (
            .O(N__39185),
            .I(N__39168));
    Span4Mux_h I__8506 (
            .O(N__39180),
            .I(N__39165));
    Span4Mux_v I__8505 (
            .O(N__39177),
            .I(N__39162));
    Span4Mux_v I__8504 (
            .O(N__39174),
            .I(N__39159));
    LocalMux I__8503 (
            .O(N__39171),
            .I(N__39156));
    Span12Mux_v I__8502 (
            .O(N__39168),
            .I(N__39151));
    Span4Mux_v I__8501 (
            .O(N__39165),
            .I(N__39148));
    Span4Mux_h I__8500 (
            .O(N__39162),
            .I(N__39145));
    Span4Mux_h I__8499 (
            .O(N__39159),
            .I(N__39140));
    Span4Mux_v I__8498 (
            .O(N__39156),
            .I(N__39140));
    CEMux I__8497 (
            .O(N__39155),
            .I(N__39137));
    CEMux I__8496 (
            .O(N__39154),
            .I(N__39134));
    Odrv12 I__8495 (
            .O(N__39151),
            .I(\u0.N_446 ));
    Odrv4 I__8494 (
            .O(N__39148),
            .I(\u0.N_446 ));
    Odrv4 I__8493 (
            .O(N__39145),
            .I(\u0.N_446 ));
    Odrv4 I__8492 (
            .O(N__39140),
            .I(\u0.N_446 ));
    LocalMux I__8491 (
            .O(N__39137),
            .I(\u0.N_446 ));
    LocalMux I__8490 (
            .O(N__39134),
            .I(\u0.N_446 ));
    InMux I__8489 (
            .O(N__39121),
            .I(N__39117));
    InMux I__8488 (
            .O(N__39120),
            .I(N__39114));
    LocalMux I__8487 (
            .O(N__39117),
            .I(N__39111));
    LocalMux I__8486 (
            .O(N__39114),
            .I(PIO_cmdport_T2_2));
    Odrv12 I__8485 (
            .O(N__39111),
            .I(PIO_cmdport_T2_2));
    InMux I__8484 (
            .O(N__39106),
            .I(N__39103));
    LocalMux I__8483 (
            .O(N__39103),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_23 ));
    InMux I__8482 (
            .O(N__39100),
            .I(N__39097));
    LocalMux I__8481 (
            .O(N__39097),
            .I(N__39094));
    Span4Mux_v I__8480 (
            .O(N__39094),
            .I(N__39091));
    Span4Mux_h I__8479 (
            .O(N__39091),
            .I(N__39088));
    Odrv4 I__8478 (
            .O(N__39088),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_23 ));
    InMux I__8477 (
            .O(N__39085),
            .I(N__39082));
    LocalMux I__8476 (
            .O(N__39082),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI81ITZ0Z_23 ));
    InMux I__8475 (
            .O(N__39079),
            .I(N__39076));
    LocalMux I__8474 (
            .O(N__39076),
            .I(N__39073));
    Odrv12 I__8473 (
            .O(N__39073),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_9 ));
    InMux I__8472 (
            .O(N__39070),
            .I(N__39067));
    LocalMux I__8471 (
            .O(N__39067),
            .I(N__39064));
    Span4Mux_v I__8470 (
            .O(N__39064),
            .I(N__39061));
    Odrv4 I__8469 (
            .O(N__39061),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_9 ));
    CascadeMux I__8468 (
            .O(N__39058),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNIGFTNZ0Z_9_cascade_ ));
    InMux I__8467 (
            .O(N__39055),
            .I(N__39052));
    LocalMux I__8466 (
            .O(N__39052),
            .I(N__39049));
    Span4Mux_v I__8465 (
            .O(N__39049),
            .I(N__39046));
    Odrv4 I__8464 (
            .O(N__39046),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_9 ));
    InMux I__8463 (
            .O(N__39043),
            .I(N__39040));
    LocalMux I__8462 (
            .O(N__39040),
            .I(N__39037));
    Span4Mux_h I__8461 (
            .O(N__39037),
            .I(N__39034));
    Odrv4 I__8460 (
            .O(N__39034),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_0 ));
    InMux I__8459 (
            .O(N__39031),
            .I(N__39028));
    LocalMux I__8458 (
            .O(N__39028),
            .I(N__39025));
    Span4Mux_v I__8457 (
            .O(N__39025),
            .I(N__39022));
    Odrv4 I__8456 (
            .O(N__39022),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_0 ));
    InMux I__8455 (
            .O(N__39019),
            .I(N__39016));
    LocalMux I__8454 (
            .O(N__39016),
            .I(N__39013));
    Span4Mux_h I__8453 (
            .O(N__39013),
            .I(N__39010));
    Odrv4 I__8452 (
            .O(N__39010),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIUOHM1Z0Z_2 ));
    InMux I__8451 (
            .O(N__39007),
            .I(N__39004));
    LocalMux I__8450 (
            .O(N__39004),
            .I(N__39001));
    Span4Mux_h I__8449 (
            .O(N__39001),
            .I(N__38998));
    Odrv4 I__8448 (
            .O(N__38998),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI4D9KZ0Z_23 ));
    InMux I__8447 (
            .O(N__38995),
            .I(N__38992));
    LocalMux I__8446 (
            .O(N__38992),
            .I(N__38989));
    Span4Mux_h I__8445 (
            .O(N__38989),
            .I(N__38986));
    Odrv4 I__8444 (
            .O(N__38986),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_23 ));
    InMux I__8443 (
            .O(N__38983),
            .I(N__38980));
    LocalMux I__8442 (
            .O(N__38980),
            .I(N__38977));
    Span4Mux_h I__8441 (
            .O(N__38977),
            .I(N__38974));
    Odrv4 I__8440 (
            .O(N__38974),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_23 ));
    InMux I__8439 (
            .O(N__38971),
            .I(N__38968));
    LocalMux I__8438 (
            .O(N__38968),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI0P0RZ0Z_23 ));
    InMux I__8437 (
            .O(N__38965),
            .I(N__38962));
    LocalMux I__8436 (
            .O(N__38962),
            .I(N__38959));
    Odrv12 I__8435 (
            .O(N__38959),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_25 ));
    InMux I__8434 (
            .O(N__38956),
            .I(N__38953));
    LocalMux I__8433 (
            .O(N__38953),
            .I(N__38950));
    Span4Mux_v I__8432 (
            .O(N__38950),
            .I(N__38947));
    Odrv4 I__8431 (
            .O(N__38947),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_25 ));
    InMux I__8430 (
            .O(N__38944),
            .I(N__38941));
    LocalMux I__8429 (
            .O(N__38941),
            .I(\u0.CtrlRegZ0Z_22 ));
    InMux I__8428 (
            .O(N__38938),
            .I(N__38935));
    LocalMux I__8427 (
            .O(N__38935),
            .I(N__38932));
    Span4Mux_h I__8426 (
            .O(N__38932),
            .I(N__38929));
    Span4Mux_v I__8425 (
            .O(N__38929),
            .I(N__38925));
    InMux I__8424 (
            .O(N__38928),
            .I(N__38922));
    Odrv4 I__8423 (
            .O(N__38925),
            .I(PIO_cmdport_T4_6));
    LocalMux I__8422 (
            .O(N__38922),
            .I(PIO_cmdport_T4_6));
    CascadeMux I__8421 (
            .O(N__38917),
            .I(\u0.dat_o_i_0_2_22_cascade_ ));
    InMux I__8420 (
            .O(N__38914),
            .I(N__38911));
    LocalMux I__8419 (
            .O(N__38911),
            .I(N__38908));
    Odrv12 I__8418 (
            .O(N__38908),
            .I(\u0.dat_o_i_0_0_22 ));
    IoInMux I__8417 (
            .O(N__38905),
            .I(N__38902));
    LocalMux I__8416 (
            .O(N__38902),
            .I(N__38899));
    IoSpan4Mux I__8415 (
            .O(N__38899),
            .I(N__38896));
    Sp12to4 I__8414 (
            .O(N__38896),
            .I(N__38893));
    Span12Mux_s7_h I__8413 (
            .O(N__38893),
            .I(N__38890));
    Odrv12 I__8412 (
            .O(N__38890),
            .I(N_330_i));
    InMux I__8411 (
            .O(N__38887),
            .I(N__38884));
    LocalMux I__8410 (
            .O(N__38884),
            .I(N__38881));
    Span4Mux_h I__8409 (
            .O(N__38881),
            .I(N__38878));
    Span4Mux_h I__8408 (
            .O(N__38878),
            .I(N__38875));
    Odrv4 I__8407 (
            .O(N__38875),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_7 ));
    InMux I__8406 (
            .O(N__38872),
            .I(N__38869));
    LocalMux I__8405 (
            .O(N__38869),
            .I(N__38866));
    Odrv4 I__8404 (
            .O(N__38866),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNICBTNZ0Z_7 ));
    InMux I__8403 (
            .O(N__38863),
            .I(N__38860));
    LocalMux I__8402 (
            .O(N__38860),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_7 ));
    CascadeMux I__8401 (
            .O(N__38857),
            .I(N__38852));
    CascadeMux I__8400 (
            .O(N__38856),
            .I(N__38846));
    CascadeMux I__8399 (
            .O(N__38855),
            .I(N__38842));
    InMux I__8398 (
            .O(N__38852),
            .I(N__38834));
    InMux I__8397 (
            .O(N__38851),
            .I(N__38834));
    InMux I__8396 (
            .O(N__38850),
            .I(N__38831));
    InMux I__8395 (
            .O(N__38849),
            .I(N__38826));
    InMux I__8394 (
            .O(N__38846),
            .I(N__38821));
    InMux I__8393 (
            .O(N__38845),
            .I(N__38821));
    InMux I__8392 (
            .O(N__38842),
            .I(N__38816));
    InMux I__8391 (
            .O(N__38841),
            .I(N__38816));
    InMux I__8390 (
            .O(N__38840),
            .I(N__38811));
    InMux I__8389 (
            .O(N__38839),
            .I(N__38811));
    LocalMux I__8388 (
            .O(N__38834),
            .I(N__38808));
    LocalMux I__8387 (
            .O(N__38831),
            .I(N__38805));
    InMux I__8386 (
            .O(N__38830),
            .I(N__38797));
    InMux I__8385 (
            .O(N__38829),
            .I(N__38797));
    LocalMux I__8384 (
            .O(N__38826),
            .I(N__38792));
    LocalMux I__8383 (
            .O(N__38821),
            .I(N__38792));
    LocalMux I__8382 (
            .O(N__38816),
            .I(N__38789));
    LocalMux I__8381 (
            .O(N__38811),
            .I(N__38786));
    Span4Mux_s3_v I__8380 (
            .O(N__38808),
            .I(N__38781));
    Span4Mux_h I__8379 (
            .O(N__38805),
            .I(N__38781));
    InMux I__8378 (
            .O(N__38804),
            .I(N__38778));
    InMux I__8377 (
            .O(N__38803),
            .I(N__38773));
    InMux I__8376 (
            .O(N__38802),
            .I(N__38773));
    LocalMux I__8375 (
            .O(N__38797),
            .I(N__38768));
    Span4Mux_h I__8374 (
            .O(N__38792),
            .I(N__38768));
    Span4Mux_v I__8373 (
            .O(N__38789),
            .I(N__38765));
    Span4Mux_v I__8372 (
            .O(N__38786),
            .I(N__38760));
    Span4Mux_v I__8371 (
            .O(N__38781),
            .I(N__38760));
    LocalMux I__8370 (
            .O(N__38778),
            .I(\u1.DMA_control.readDlw_7 ));
    LocalMux I__8369 (
            .O(N__38773),
            .I(\u1.DMA_control.readDlw_7 ));
    Odrv4 I__8368 (
            .O(N__38768),
            .I(\u1.DMA_control.readDlw_7 ));
    Odrv4 I__8367 (
            .O(N__38765),
            .I(\u1.DMA_control.readDlw_7 ));
    Odrv4 I__8366 (
            .O(N__38760),
            .I(\u1.DMA_control.readDlw_7 ));
    InMux I__8365 (
            .O(N__38749),
            .I(N__38746));
    LocalMux I__8364 (
            .O(N__38746),
            .I(N__38736));
    InMux I__8363 (
            .O(N__38745),
            .I(N__38731));
    InMux I__8362 (
            .O(N__38744),
            .I(N__38731));
    InMux I__8361 (
            .O(N__38743),
            .I(N__38728));
    InMux I__8360 (
            .O(N__38742),
            .I(N__38725));
    InMux I__8359 (
            .O(N__38741),
            .I(N__38722));
    InMux I__8358 (
            .O(N__38740),
            .I(N__38717));
    InMux I__8357 (
            .O(N__38739),
            .I(N__38717));
    Sp12to4 I__8356 (
            .O(N__38736),
            .I(N__38710));
    LocalMux I__8355 (
            .O(N__38731),
            .I(N__38710));
    LocalMux I__8354 (
            .O(N__38728),
            .I(N__38707));
    LocalMux I__8353 (
            .O(N__38725),
            .I(N__38702));
    LocalMux I__8352 (
            .O(N__38722),
            .I(N__38702));
    LocalMux I__8351 (
            .O(N__38717),
            .I(N__38699));
    InMux I__8350 (
            .O(N__38716),
            .I(N__38694));
    InMux I__8349 (
            .O(N__38715),
            .I(N__38694));
    Span12Mux_s7_v I__8348 (
            .O(N__38710),
            .I(N__38687));
    Span4Mux_h I__8347 (
            .O(N__38707),
            .I(N__38682));
    Span4Mux_h I__8346 (
            .O(N__38702),
            .I(N__38682));
    Span4Mux_v I__8345 (
            .O(N__38699),
            .I(N__38677));
    LocalMux I__8344 (
            .O(N__38694),
            .I(N__38677));
    InMux I__8343 (
            .O(N__38693),
            .I(N__38674));
    InMux I__8342 (
            .O(N__38692),
            .I(N__38671));
    InMux I__8341 (
            .O(N__38691),
            .I(N__38668));
    InMux I__8340 (
            .O(N__38690),
            .I(N__38665));
    Odrv12 I__8339 (
            .O(N__38687),
            .I(\u1.DMA_control.readDfw_7 ));
    Odrv4 I__8338 (
            .O(N__38682),
            .I(\u1.DMA_control.readDfw_7 ));
    Odrv4 I__8337 (
            .O(N__38677),
            .I(\u1.DMA_control.readDfw_7 ));
    LocalMux I__8336 (
            .O(N__38674),
            .I(\u1.DMA_control.readDfw_7 ));
    LocalMux I__8335 (
            .O(N__38671),
            .I(\u1.DMA_control.readDfw_7 ));
    LocalMux I__8334 (
            .O(N__38668),
            .I(\u1.DMA_control.readDfw_7 ));
    LocalMux I__8333 (
            .O(N__38665),
            .I(\u1.DMA_control.readDfw_7 ));
    InMux I__8332 (
            .O(N__38650),
            .I(N__38647));
    LocalMux I__8331 (
            .O(N__38647),
            .I(N__38644));
    Span4Mux_v I__8330 (
            .O(N__38644),
            .I(N__38641));
    Span4Mux_h I__8329 (
            .O(N__38641),
            .I(N__38638));
    Odrv4 I__8328 (
            .O(N__38638),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_8 ));
    InMux I__8327 (
            .O(N__38635),
            .I(N__38632));
    LocalMux I__8326 (
            .O(N__38632),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_8 ));
    InMux I__8325 (
            .O(N__38629),
            .I(N__38620));
    InMux I__8324 (
            .O(N__38628),
            .I(N__38615));
    InMux I__8323 (
            .O(N__38627),
            .I(N__38610));
    InMux I__8322 (
            .O(N__38626),
            .I(N__38610));
    InMux I__8321 (
            .O(N__38625),
            .I(N__38606));
    InMux I__8320 (
            .O(N__38624),
            .I(N__38601));
    InMux I__8319 (
            .O(N__38623),
            .I(N__38601));
    LocalMux I__8318 (
            .O(N__38620),
            .I(N__38598));
    InMux I__8317 (
            .O(N__38619),
            .I(N__38595));
    InMux I__8316 (
            .O(N__38618),
            .I(N__38592));
    LocalMux I__8315 (
            .O(N__38615),
            .I(N__38587));
    LocalMux I__8314 (
            .O(N__38610),
            .I(N__38587));
    InMux I__8313 (
            .O(N__38609),
            .I(N__38580));
    LocalMux I__8312 (
            .O(N__38606),
            .I(N__38577));
    LocalMux I__8311 (
            .O(N__38601),
            .I(N__38574));
    Span4Mux_v I__8310 (
            .O(N__38598),
            .I(N__38565));
    LocalMux I__8309 (
            .O(N__38595),
            .I(N__38565));
    LocalMux I__8308 (
            .O(N__38592),
            .I(N__38565));
    Span4Mux_s2_v I__8307 (
            .O(N__38587),
            .I(N__38565));
    InMux I__8306 (
            .O(N__38586),
            .I(N__38560));
    InMux I__8305 (
            .O(N__38585),
            .I(N__38560));
    InMux I__8304 (
            .O(N__38584),
            .I(N__38555));
    InMux I__8303 (
            .O(N__38583),
            .I(N__38555));
    LocalMux I__8302 (
            .O(N__38580),
            .I(N__38552));
    Span12Mux_h I__8301 (
            .O(N__38577),
            .I(N__38549));
    Span4Mux_v I__8300 (
            .O(N__38574),
            .I(N__38544));
    Span4Mux_v I__8299 (
            .O(N__38565),
            .I(N__38544));
    LocalMux I__8298 (
            .O(N__38560),
            .I(\u1.DMA_control.readDfw_8 ));
    LocalMux I__8297 (
            .O(N__38555),
            .I(\u1.DMA_control.readDfw_8 ));
    Odrv12 I__8296 (
            .O(N__38552),
            .I(\u1.DMA_control.readDfw_8 ));
    Odrv12 I__8295 (
            .O(N__38549),
            .I(\u1.DMA_control.readDfw_8 ));
    Odrv4 I__8294 (
            .O(N__38544),
            .I(\u1.DMA_control.readDfw_8 ));
    InMux I__8293 (
            .O(N__38533),
            .I(N__38523));
    InMux I__8292 (
            .O(N__38532),
            .I(N__38520));
    InMux I__8291 (
            .O(N__38531),
            .I(N__38517));
    InMux I__8290 (
            .O(N__38530),
            .I(N__38514));
    InMux I__8289 (
            .O(N__38529),
            .I(N__38509));
    InMux I__8288 (
            .O(N__38528),
            .I(N__38509));
    InMux I__8287 (
            .O(N__38527),
            .I(N__38505));
    InMux I__8286 (
            .O(N__38526),
            .I(N__38502));
    LocalMux I__8285 (
            .O(N__38523),
            .I(N__38495));
    LocalMux I__8284 (
            .O(N__38520),
            .I(N__38495));
    LocalMux I__8283 (
            .O(N__38517),
            .I(N__38495));
    LocalMux I__8282 (
            .O(N__38514),
            .I(N__38492));
    LocalMux I__8281 (
            .O(N__38509),
            .I(N__38489));
    InMux I__8280 (
            .O(N__38508),
            .I(N__38486));
    LocalMux I__8279 (
            .O(N__38505),
            .I(N__38478));
    LocalMux I__8278 (
            .O(N__38502),
            .I(N__38478));
    Span4Mux_s3_v I__8277 (
            .O(N__38495),
            .I(N__38473));
    Span4Mux_h I__8276 (
            .O(N__38492),
            .I(N__38473));
    Span4Mux_v I__8275 (
            .O(N__38489),
            .I(N__38468));
    LocalMux I__8274 (
            .O(N__38486),
            .I(N__38468));
    InMux I__8273 (
            .O(N__38485),
            .I(N__38465));
    CascadeMux I__8272 (
            .O(N__38484),
            .I(N__38462));
    InMux I__8271 (
            .O(N__38483),
            .I(N__38456));
    Span4Mux_v I__8270 (
            .O(N__38478),
            .I(N__38453));
    Span4Mux_h I__8269 (
            .O(N__38473),
            .I(N__38448));
    Span4Mux_h I__8268 (
            .O(N__38468),
            .I(N__38448));
    LocalMux I__8267 (
            .O(N__38465),
            .I(N__38445));
    InMux I__8266 (
            .O(N__38462),
            .I(N__38440));
    InMux I__8265 (
            .O(N__38461),
            .I(N__38440));
    InMux I__8264 (
            .O(N__38460),
            .I(N__38437));
    InMux I__8263 (
            .O(N__38459),
            .I(N__38434));
    LocalMux I__8262 (
            .O(N__38456),
            .I(\u1.DMA_control.readDlw_8 ));
    Odrv4 I__8261 (
            .O(N__38453),
            .I(\u1.DMA_control.readDlw_8 ));
    Odrv4 I__8260 (
            .O(N__38448),
            .I(\u1.DMA_control.readDlw_8 ));
    Odrv12 I__8259 (
            .O(N__38445),
            .I(\u1.DMA_control.readDlw_8 ));
    LocalMux I__8258 (
            .O(N__38440),
            .I(\u1.DMA_control.readDlw_8 ));
    LocalMux I__8257 (
            .O(N__38437),
            .I(\u1.DMA_control.readDlw_8 ));
    LocalMux I__8256 (
            .O(N__38434),
            .I(\u1.DMA_control.readDlw_8 ));
    InMux I__8255 (
            .O(N__38419),
            .I(N__38416));
    LocalMux I__8254 (
            .O(N__38416),
            .I(N__38413));
    Span4Mux_v I__8253 (
            .O(N__38413),
            .I(N__38410));
    Odrv4 I__8252 (
            .O(N__38410),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_24 ));
    InMux I__8251 (
            .O(N__38407),
            .I(N__38404));
    LocalMux I__8250 (
            .O(N__38404),
            .I(N__38401));
    Span4Mux_v I__8249 (
            .O(N__38401),
            .I(N__38398));
    Odrv4 I__8248 (
            .O(N__38398),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_23 ));
    InMux I__8247 (
            .O(N__38395),
            .I(N__38392));
    LocalMux I__8246 (
            .O(N__38392),
            .I(N__38387));
    InMux I__8245 (
            .O(N__38391),
            .I(N__38382));
    InMux I__8244 (
            .O(N__38390),
            .I(N__38382));
    Span4Mux_v I__8243 (
            .O(N__38387),
            .I(N__38379));
    LocalMux I__8242 (
            .O(N__38382),
            .I(N__38376));
    Span4Mux_v I__8241 (
            .O(N__38379),
            .I(N__38373));
    Span4Mux_v I__8240 (
            .O(N__38376),
            .I(N__38370));
    Span4Mux_v I__8239 (
            .O(N__38373),
            .I(N__38367));
    Sp12to4 I__8238 (
            .O(N__38370),
            .I(N__38364));
    Sp12to4 I__8237 (
            .O(N__38367),
            .I(N__38359));
    Span12Mux_v I__8236 (
            .O(N__38364),
            .I(N__38359));
    Span12Mux_h I__8235 (
            .O(N__38359),
            .I(N__38356));
    Odrv12 I__8234 (
            .O(N__38356),
            .I(dd_pad_i_c_7));
    InMux I__8233 (
            .O(N__38353),
            .I(N__38350));
    LocalMux I__8232 (
            .O(N__38350),
            .I(PIOq_7));
    CascadeMux I__8231 (
            .O(N__38347),
            .I(N__38344));
    InMux I__8230 (
            .O(N__38344),
            .I(N__38341));
    LocalMux I__8229 (
            .O(N__38341),
            .I(N__38336));
    InMux I__8228 (
            .O(N__38340),
            .I(N__38330));
    InMux I__8227 (
            .O(N__38339),
            .I(N__38330));
    Span4Mux_h I__8226 (
            .O(N__38336),
            .I(N__38327));
    InMux I__8225 (
            .O(N__38335),
            .I(N__38323));
    LocalMux I__8224 (
            .O(N__38330),
            .I(N__38320));
    Span4Mux_h I__8223 (
            .O(N__38327),
            .I(N__38317));
    InMux I__8222 (
            .O(N__38326),
            .I(N__38314));
    LocalMux I__8221 (
            .O(N__38323),
            .I(N__38311));
    Span4Mux_h I__8220 (
            .O(N__38320),
            .I(N__38308));
    Odrv4 I__8219 (
            .O(N__38317),
            .I(IDEctrl_IDEen));
    LocalMux I__8218 (
            .O(N__38314),
            .I(IDEctrl_IDEen));
    Odrv12 I__8217 (
            .O(N__38311),
            .I(IDEctrl_IDEen));
    Odrv4 I__8216 (
            .O(N__38308),
            .I(IDEctrl_IDEen));
    InMux I__8215 (
            .O(N__38299),
            .I(N__38296));
    LocalMux I__8214 (
            .O(N__38296),
            .I(\u0.dat_o_0_0_2_7 ));
    InMux I__8213 (
            .O(N__38293),
            .I(N__38290));
    LocalMux I__8212 (
            .O(N__38290),
            .I(N__38287));
    Span4Mux_v I__8211 (
            .O(N__38287),
            .I(N__38284));
    Odrv4 I__8210 (
            .O(N__38284),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI8R4NZ0Z_7 ));
    InMux I__8209 (
            .O(N__38281),
            .I(N__38278));
    LocalMux I__8208 (
            .O(N__38278),
            .I(N__38275));
    Span4Mux_v I__8207 (
            .O(N__38275),
            .I(N__38272));
    Span4Mux_h I__8206 (
            .O(N__38272),
            .I(N__38269));
    Odrv4 I__8205 (
            .O(N__38269),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI4BCMZ0Z_7 ));
    InMux I__8204 (
            .O(N__38266),
            .I(N__38263));
    LocalMux I__8203 (
            .O(N__38263),
            .I(iQ_RNIUGOK1_2));
    InMux I__8202 (
            .O(N__38260),
            .I(N__38257));
    LocalMux I__8201 (
            .O(N__38257),
            .I(\u0.N_1980 ));
    InMux I__8200 (
            .O(N__38254),
            .I(N__38251));
    LocalMux I__8199 (
            .O(N__38251),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_7 ));
    InMux I__8198 (
            .O(N__38248),
            .I(N__38245));
    LocalMux I__8197 (
            .O(N__38245),
            .I(mem_mem_ram6__RNITSOD1_7));
    InMux I__8196 (
            .O(N__38242),
            .I(N__38239));
    LocalMux I__8195 (
            .O(N__38239),
            .I(N__38236));
    Span4Mux_v I__8194 (
            .O(N__38236),
            .I(N__38233));
    Span4Mux_h I__8193 (
            .O(N__38233),
            .I(N__38230));
    Odrv4 I__8192 (
            .O(N__38230),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI6VHTZ0Z_22 ));
    InMux I__8191 (
            .O(N__38227),
            .I(N__38224));
    LocalMux I__8190 (
            .O(N__38224),
            .I(N__38221));
    Span4Mux_v I__8189 (
            .O(N__38221),
            .I(N__38218));
    Sp12to4 I__8188 (
            .O(N__38218),
            .I(N__38215));
    Odrv12 I__8187 (
            .O(N__38215),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_22 ));
    InMux I__8186 (
            .O(N__38212),
            .I(N__38209));
    LocalMux I__8185 (
            .O(N__38209),
            .I(N__38206));
    Span4Mux_v I__8184 (
            .O(N__38206),
            .I(N__38203));
    Odrv4 I__8183 (
            .O(N__38203),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_22 ));
    InMux I__8182 (
            .O(N__38200),
            .I(N__38197));
    LocalMux I__8181 (
            .O(N__38197),
            .I(N__38194));
    Span4Mux_v I__8180 (
            .O(N__38194),
            .I(N__38191));
    Odrv4 I__8179 (
            .O(N__38191),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_22 ));
    CascadeMux I__8178 (
            .O(N__38188),
            .I(N__38185));
    InMux I__8177 (
            .O(N__38185),
            .I(N__38179));
    InMux I__8176 (
            .O(N__38184),
            .I(N__38176));
    InMux I__8175 (
            .O(N__38183),
            .I(N__38173));
    InMux I__8174 (
            .O(N__38182),
            .I(N__38170));
    LocalMux I__8173 (
            .O(N__38179),
            .I(N__38165));
    LocalMux I__8172 (
            .O(N__38176),
            .I(N__38165));
    LocalMux I__8171 (
            .O(N__38173),
            .I(N__38162));
    LocalMux I__8170 (
            .O(N__38170),
            .I(N__38159));
    Span4Mux_v I__8169 (
            .O(N__38165),
            .I(N__38156));
    Span4Mux_v I__8168 (
            .O(N__38162),
            .I(N__38153));
    Span4Mux_v I__8167 (
            .O(N__38159),
            .I(N__38150));
    Span4Mux_v I__8166 (
            .O(N__38156),
            .I(N__38146));
    Span4Mux_v I__8165 (
            .O(N__38153),
            .I(N__38143));
    Span4Mux_h I__8164 (
            .O(N__38150),
            .I(N__38140));
    InMux I__8163 (
            .O(N__38149),
            .I(N__38137));
    Sp12to4 I__8162 (
            .O(N__38146),
            .I(N__38134));
    Span4Mux_h I__8161 (
            .O(N__38143),
            .I(N__38129));
    Span4Mux_h I__8160 (
            .O(N__38140),
            .I(N__38129));
    LocalMux I__8159 (
            .O(N__38137),
            .I(N__38126));
    Span12Mux_h I__8158 (
            .O(N__38134),
            .I(N__38123));
    Span4Mux_h I__8157 (
            .O(N__38129),
            .I(N__38118));
    Span4Mux_v I__8156 (
            .O(N__38126),
            .I(N__38118));
    Odrv12 I__8155 (
            .O(N__38123),
            .I(wb_dat_i_c_22));
    Odrv4 I__8154 (
            .O(N__38118),
            .I(wb_dat_i_c_22));
    CascadeMux I__8153 (
            .O(N__38113),
            .I(\u0.N_1636_cascade_ ));
    InMux I__8152 (
            .O(N__38110),
            .I(N__38107));
    LocalMux I__8151 (
            .O(N__38107),
            .I(N__38104));
    Odrv4 I__8150 (
            .O(N__38104),
            .I(\u0.dat_o_i_0_21 ));
    IoInMux I__8149 (
            .O(N__38101),
            .I(N__38098));
    LocalMux I__8148 (
            .O(N__38098),
            .I(N__38095));
    Span4Mux_s1_h I__8147 (
            .O(N__38095),
            .I(N__38092));
    Span4Mux_h I__8146 (
            .O(N__38092),
            .I(N__38089));
    Sp12to4 I__8145 (
            .O(N__38089),
            .I(N__38086));
    Span12Mux_s11_v I__8144 (
            .O(N__38086),
            .I(N__38083));
    Span12Mux_h I__8143 (
            .O(N__38083),
            .I(N__38080));
    Odrv12 I__8142 (
            .O(N__38080),
            .I(N_259_i));
    InMux I__8141 (
            .O(N__38077),
            .I(N__38073));
    InMux I__8140 (
            .O(N__38076),
            .I(N__38070));
    LocalMux I__8139 (
            .O(N__38073),
            .I(N__38066));
    LocalMux I__8138 (
            .O(N__38070),
            .I(N__38063));
    InMux I__8137 (
            .O(N__38069),
            .I(N__38060));
    Span4Mux_h I__8136 (
            .O(N__38066),
            .I(N__38057));
    Span4Mux_v I__8135 (
            .O(N__38063),
            .I(N__38051));
    LocalMux I__8134 (
            .O(N__38060),
            .I(N__38051));
    Span4Mux_h I__8133 (
            .O(N__38057),
            .I(N__38048));
    InMux I__8132 (
            .O(N__38056),
            .I(N__38044));
    Sp12to4 I__8131 (
            .O(N__38051),
            .I(N__38041));
    Span4Mux_v I__8130 (
            .O(N__38048),
            .I(N__38038));
    InMux I__8129 (
            .O(N__38047),
            .I(N__38035));
    LocalMux I__8128 (
            .O(N__38044),
            .I(N__38032));
    Span12Mux_v I__8127 (
            .O(N__38041),
            .I(N__38029));
    Span4Mux_h I__8126 (
            .O(N__38038),
            .I(N__38024));
    LocalMux I__8125 (
            .O(N__38035),
            .I(N__38024));
    Span12Mux_v I__8124 (
            .O(N__38032),
            .I(N__38021));
    Span12Mux_h I__8123 (
            .O(N__38029),
            .I(N__38018));
    Span4Mux_v I__8122 (
            .O(N__38024),
            .I(N__38015));
    Odrv12 I__8121 (
            .O(N__38021),
            .I(wb_dat_i_c_21));
    Odrv12 I__8120 (
            .O(N__38018),
            .I(wb_dat_i_c_21));
    Odrv4 I__8119 (
            .O(N__38015),
            .I(wb_dat_i_c_21));
    InMux I__8118 (
            .O(N__38008),
            .I(N__38005));
    LocalMux I__8117 (
            .O(N__38005),
            .I(N__38002));
    Span4Mux_h I__8116 (
            .O(N__38002),
            .I(N__37999));
    Span4Mux_h I__8115 (
            .O(N__37999),
            .I(N__37996));
    Odrv4 I__8114 (
            .O(N__37996),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_21 ));
    InMux I__8113 (
            .O(N__37993),
            .I(N__37990));
    LocalMux I__8112 (
            .O(N__37990),
            .I(N__37987));
    Span4Mux_v I__8111 (
            .O(N__37987),
            .I(N__37984));
    Odrv4 I__8110 (
            .O(N__37984),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_21 ));
    CascadeMux I__8109 (
            .O(N__37981),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNISK0RZ0Z_21_cascade_ ));
    InMux I__8108 (
            .O(N__37978),
            .I(N__37975));
    LocalMux I__8107 (
            .O(N__37975),
            .I(N__37972));
    Span12Mux_v I__8106 (
            .O(N__37972),
            .I(N__37969));
    Odrv12 I__8105 (
            .O(N__37969),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI099KZ0Z_21 ));
    InMux I__8104 (
            .O(N__37966),
            .I(N__37963));
    LocalMux I__8103 (
            .O(N__37963),
            .I(iQ_RNIE8HM1_2));
    InMux I__8102 (
            .O(N__37960),
            .I(N__37957));
    LocalMux I__8101 (
            .O(N__37957),
            .I(N__37954));
    Sp12to4 I__8100 (
            .O(N__37954),
            .I(N__37951));
    Span12Mux_h I__8099 (
            .O(N__37951),
            .I(N__37948));
    Odrv12 I__8098 (
            .O(N__37948),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI4THTZ0Z_21 ));
    InMux I__8097 (
            .O(N__37945),
            .I(N__37942));
    LocalMux I__8096 (
            .O(N__37942),
            .I(N__37939));
    Span12Mux_h I__8095 (
            .O(N__37939),
            .I(N__37936));
    Odrv12 I__8094 (
            .O(N__37936),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_21 ));
    CascadeMux I__8093 (
            .O(N__37933),
            .I(N__37930));
    InMux I__8092 (
            .O(N__37930),
            .I(N__37927));
    LocalMux I__8091 (
            .O(N__37927),
            .I(mem_mem_ram6__RNI1PD71_21));
    InMux I__8090 (
            .O(N__37924),
            .I(N__37921));
    LocalMux I__8089 (
            .O(N__37921),
            .I(N__37918));
    Odrv4 I__8088 (
            .O(N__37918),
            .I(\u0.CtrlRegZ0Z_21 ));
    InMux I__8087 (
            .O(N__37915),
            .I(N__37912));
    LocalMux I__8086 (
            .O(N__37912),
            .I(N__37908));
    InMux I__8085 (
            .O(N__37911),
            .I(N__37905));
    Span4Mux_v I__8084 (
            .O(N__37908),
            .I(N__37902));
    LocalMux I__8083 (
            .O(N__37905),
            .I(N__37899));
    Odrv4 I__8082 (
            .O(N__37902),
            .I(PIO_cmdport_T4_5));
    Odrv4 I__8081 (
            .O(N__37899),
            .I(PIO_cmdport_T4_5));
    InMux I__8080 (
            .O(N__37894),
            .I(N__37891));
    LocalMux I__8079 (
            .O(N__37891),
            .I(\u0.dat_o_i_2_21 ));
    InMux I__8078 (
            .O(N__37888),
            .I(N__37885));
    LocalMux I__8077 (
            .O(N__37885),
            .I(N__37882));
    Odrv12 I__8076 (
            .O(N__37882),
            .I(\u0.dat_o_0_0_6_7 ));
    CascadeMux I__8075 (
            .O(N__37879),
            .I(\u0.N_1979_cascade_ ));
    IoInMux I__8074 (
            .O(N__37876),
            .I(N__37873));
    LocalMux I__8073 (
            .O(N__37873),
            .I(N__37870));
    IoSpan4Mux I__8072 (
            .O(N__37870),
            .I(N__37867));
    Sp12to4 I__8071 (
            .O(N__37867),
            .I(N__37864));
    Span12Mux_s6_v I__8070 (
            .O(N__37864),
            .I(N__37861));
    Span12Mux_h I__8069 (
            .O(N__37861),
            .I(N__37858));
    Odrv12 I__8068 (
            .O(N__37858),
            .I(wb_dat_o_c_7));
    CascadeMux I__8067 (
            .O(N__37855),
            .I(N__37851));
    CascadeMux I__8066 (
            .O(N__37854),
            .I(N__37848));
    InMux I__8065 (
            .O(N__37851),
            .I(N__37845));
    InMux I__8064 (
            .O(N__37848),
            .I(N__37842));
    LocalMux I__8063 (
            .O(N__37845),
            .I(N__37839));
    LocalMux I__8062 (
            .O(N__37842),
            .I(N__37836));
    Span4Mux_v I__8061 (
            .O(N__37839),
            .I(N__37833));
    Odrv4 I__8060 (
            .O(N__37836),
            .I(DMA_dev1_Tm_4));
    Odrv4 I__8059 (
            .O(N__37833),
            .I(DMA_dev1_Tm_4));
    InMux I__8058 (
            .O(N__37828),
            .I(N__37824));
    InMux I__8057 (
            .O(N__37827),
            .I(N__37821));
    LocalMux I__8056 (
            .O(N__37824),
            .I(N__37818));
    LocalMux I__8055 (
            .O(N__37821),
            .I(N__37815));
    Span4Mux_v I__8054 (
            .O(N__37818),
            .I(N__37812));
    Span4Mux_h I__8053 (
            .O(N__37815),
            .I(N__37809));
    Odrv4 I__8052 (
            .O(N__37812),
            .I(DMA_dev1_Tm_5));
    Odrv4 I__8051 (
            .O(N__37809),
            .I(DMA_dev1_Tm_5));
    InMux I__8050 (
            .O(N__37804),
            .I(N__37801));
    LocalMux I__8049 (
            .O(N__37801),
            .I(N__37797));
    InMux I__8048 (
            .O(N__37800),
            .I(N__37794));
    Span4Mux_v I__8047 (
            .O(N__37797),
            .I(N__37791));
    LocalMux I__8046 (
            .O(N__37794),
            .I(N__37788));
    Odrv4 I__8045 (
            .O(N__37791),
            .I(PIO_cmdport_Teoc_3));
    Odrv4 I__8044 (
            .O(N__37788),
            .I(PIO_cmdport_Teoc_3));
    CascadeMux I__8043 (
            .O(N__37783),
            .I(\u0.dat_o_i_i_1_27_cascade_ ));
    InMux I__8042 (
            .O(N__37780),
            .I(N__37776));
    InMux I__8041 (
            .O(N__37779),
            .I(N__37773));
    LocalMux I__8040 (
            .O(N__37776),
            .I(N__37770));
    LocalMux I__8039 (
            .O(N__37773),
            .I(N__37767));
    Span4Mux_h I__8038 (
            .O(N__37770),
            .I(N__37762));
    Span4Mux_h I__8037 (
            .O(N__37767),
            .I(N__37762));
    Odrv4 I__8036 (
            .O(N__37762),
            .I(PIO_dport0_Teoc_3));
    CascadeMux I__8035 (
            .O(N__37759),
            .I(\u0.dat_o_i_i_4_27_cascade_ ));
    InMux I__8034 (
            .O(N__37756),
            .I(N__37753));
    LocalMux I__8033 (
            .O(N__37753),
            .I(N__37750));
    Span4Mux_v I__8032 (
            .O(N__37750),
            .I(N__37746));
    InMux I__8031 (
            .O(N__37749),
            .I(N__37743));
    Span4Mux_h I__8030 (
            .O(N__37746),
            .I(N__37740));
    LocalMux I__8029 (
            .O(N__37743),
            .I(DMA_dev1_Teoc_3));
    Odrv4 I__8028 (
            .O(N__37740),
            .I(DMA_dev1_Teoc_3));
    IoInMux I__8027 (
            .O(N__37735),
            .I(N__37732));
    LocalMux I__8026 (
            .O(N__37732),
            .I(N__37729));
    Span4Mux_s1_v I__8025 (
            .O(N__37729),
            .I(N__37726));
    Span4Mux_v I__8024 (
            .O(N__37726),
            .I(N__37723));
    Span4Mux_v I__8023 (
            .O(N__37723),
            .I(N__37720));
    Odrv4 I__8022 (
            .O(N__37720),
            .I(N_269));
    InMux I__8021 (
            .O(N__37717),
            .I(N__37711));
    InMux I__8020 (
            .O(N__37716),
            .I(N__37708));
    InMux I__8019 (
            .O(N__37715),
            .I(N__37704));
    InMux I__8018 (
            .O(N__37714),
            .I(N__37701));
    LocalMux I__8017 (
            .O(N__37711),
            .I(N__37696));
    LocalMux I__8016 (
            .O(N__37708),
            .I(N__37696));
    InMux I__8015 (
            .O(N__37707),
            .I(N__37693));
    LocalMux I__8014 (
            .O(N__37704),
            .I(N__37688));
    LocalMux I__8013 (
            .O(N__37701),
            .I(N__37688));
    Span4Mux_v I__8012 (
            .O(N__37696),
            .I(N__37684));
    LocalMux I__8011 (
            .O(N__37693),
            .I(N__37681));
    Span4Mux_v I__8010 (
            .O(N__37688),
            .I(N__37678));
    InMux I__8009 (
            .O(N__37687),
            .I(N__37675));
    Span4Mux_h I__8008 (
            .O(N__37684),
            .I(N__37669));
    Span4Mux_v I__8007 (
            .O(N__37681),
            .I(N__37669));
    Span4Mux_h I__8006 (
            .O(N__37678),
            .I(N__37666));
    LocalMux I__8005 (
            .O(N__37675),
            .I(N__37663));
    InMux I__8004 (
            .O(N__37674),
            .I(N__37660));
    Span4Mux_h I__8003 (
            .O(N__37669),
            .I(N__37657));
    Span4Mux_h I__8002 (
            .O(N__37666),
            .I(N__37650));
    Span4Mux_v I__8001 (
            .O(N__37663),
            .I(N__37650));
    LocalMux I__8000 (
            .O(N__37660),
            .I(N__37650));
    Span4Mux_v I__7999 (
            .O(N__37657),
            .I(N__37647));
    Span4Mux_h I__7998 (
            .O(N__37650),
            .I(N__37644));
    Span4Mux_h I__7997 (
            .O(N__37647),
            .I(N__37641));
    Span4Mux_v I__7996 (
            .O(N__37644),
            .I(N__37638));
    Odrv4 I__7995 (
            .O(N__37641),
            .I(wb_dat_i_c_27));
    Odrv4 I__7994 (
            .O(N__37638),
            .I(wb_dat_i_c_27));
    CascadeMux I__7993 (
            .O(N__37633),
            .I(N__37630));
    InMux I__7992 (
            .O(N__37630),
            .I(N__37627));
    LocalMux I__7991 (
            .O(N__37627),
            .I(N__37624));
    Odrv4 I__7990 (
            .O(N__37624),
            .I(\u0.CtrlRegZ0Z_27 ));
    InMux I__7989 (
            .O(N__37621),
            .I(N__37617));
    CascadeMux I__7988 (
            .O(N__37620),
            .I(N__37614));
    LocalMux I__7987 (
            .O(N__37617),
            .I(N__37611));
    InMux I__7986 (
            .O(N__37614),
            .I(N__37608));
    Span4Mux_v I__7985 (
            .O(N__37611),
            .I(N__37605));
    LocalMux I__7984 (
            .O(N__37608),
            .I(N__37602));
    Span4Mux_h I__7983 (
            .O(N__37605),
            .I(N__37597));
    Span4Mux_h I__7982 (
            .O(N__37602),
            .I(N__37597));
    Span4Mux_v I__7981 (
            .O(N__37597),
            .I(N__37594));
    Span4Mux_h I__7980 (
            .O(N__37594),
            .I(N__37591));
    Odrv4 I__7979 (
            .O(N__37591),
            .I(PIO_dport1_Teoc_3));
    InMux I__7978 (
            .O(N__37588),
            .I(N__37585));
    LocalMux I__7977 (
            .O(N__37585),
            .I(\u0.N_1682 ));
    InMux I__7976 (
            .O(N__37582),
            .I(N__37579));
    LocalMux I__7975 (
            .O(N__37579),
            .I(N__37575));
    InMux I__7974 (
            .O(N__37578),
            .I(N__37572));
    Span4Mux_v I__7973 (
            .O(N__37575),
            .I(N__37569));
    LocalMux I__7972 (
            .O(N__37572),
            .I(DMA_dev0_Teoc_3));
    Odrv4 I__7971 (
            .O(N__37569),
            .I(DMA_dev0_Teoc_3));
    InMux I__7970 (
            .O(N__37564),
            .I(N__37561));
    LocalMux I__7969 (
            .O(N__37561),
            .I(N__37558));
    Span4Mux_v I__7968 (
            .O(N__37558),
            .I(N__37555));
    Odrv4 I__7967 (
            .O(N__37555),
            .I(DMAq_27));
    InMux I__7966 (
            .O(N__37552),
            .I(N__37549));
    LocalMux I__7965 (
            .O(N__37549),
            .I(\u0.dat_o_i_i_0_27 ));
    InMux I__7964 (
            .O(N__37546),
            .I(N__37543));
    LocalMux I__7963 (
            .O(N__37543),
            .I(N__37539));
    InMux I__7962 (
            .O(N__37542),
            .I(N__37536));
    Span4Mux_h I__7961 (
            .O(N__37539),
            .I(N__37533));
    LocalMux I__7960 (
            .O(N__37536),
            .I(PIO_dport0_T4_2));
    Odrv4 I__7959 (
            .O(N__37533),
            .I(PIO_dport0_T4_2));
    CascadeMux I__7958 (
            .O(N__37528),
            .I(N__37525));
    InMux I__7957 (
            .O(N__37525),
            .I(N__37521));
    InMux I__7956 (
            .O(N__37524),
            .I(N__37518));
    LocalMux I__7955 (
            .O(N__37521),
            .I(N__37515));
    LocalMux I__7954 (
            .O(N__37518),
            .I(N__37512));
    Span4Mux_h I__7953 (
            .O(N__37515),
            .I(N__37507));
    Span4Mux_h I__7952 (
            .O(N__37512),
            .I(N__37507));
    Odrv4 I__7951 (
            .O(N__37507),
            .I(PIO_dport1_T4_4));
    CascadeMux I__7950 (
            .O(N__37504),
            .I(N__37501));
    InMux I__7949 (
            .O(N__37501),
            .I(N__37497));
    InMux I__7948 (
            .O(N__37500),
            .I(N__37494));
    LocalMux I__7947 (
            .O(N__37497),
            .I(N__37491));
    LocalMux I__7946 (
            .O(N__37494),
            .I(N__37486));
    Span4Mux_h I__7945 (
            .O(N__37491),
            .I(N__37486));
    Odrv4 I__7944 (
            .O(N__37486),
            .I(PIO_dport0_T4_4));
    InMux I__7943 (
            .O(N__37483),
            .I(N__37480));
    LocalMux I__7942 (
            .O(N__37480),
            .I(N__37477));
    Span4Mux_v I__7941 (
            .O(N__37477),
            .I(N__37474));
    Span4Mux_h I__7940 (
            .O(N__37474),
            .I(N__37471));
    Odrv4 I__7939 (
            .O(N__37471),
            .I(\u0.dat_o_0_a2_i_0_20 ));
    InMux I__7938 (
            .O(N__37468),
            .I(N__37465));
    LocalMux I__7937 (
            .O(N__37465),
            .I(N__37461));
    CascadeMux I__7936 (
            .O(N__37464),
            .I(N__37458));
    Span4Mux_h I__7935 (
            .O(N__37461),
            .I(N__37455));
    InMux I__7934 (
            .O(N__37458),
            .I(N__37452));
    Span4Mux_h I__7933 (
            .O(N__37455),
            .I(N__37449));
    LocalMux I__7932 (
            .O(N__37452),
            .I(PIO_dport1_T4_5));
    Odrv4 I__7931 (
            .O(N__37449),
            .I(PIO_dport1_T4_5));
    CascadeMux I__7930 (
            .O(N__37444),
            .I(N__37441));
    InMux I__7929 (
            .O(N__37441),
            .I(N__37437));
    InMux I__7928 (
            .O(N__37440),
            .I(N__37434));
    LocalMux I__7927 (
            .O(N__37437),
            .I(N__37431));
    LocalMux I__7926 (
            .O(N__37434),
            .I(N__37426));
    Span4Mux_h I__7925 (
            .O(N__37431),
            .I(N__37426));
    Span4Mux_h I__7924 (
            .O(N__37426),
            .I(N__37423));
    Odrv4 I__7923 (
            .O(N__37423),
            .I(PIO_dport0_T4_5));
    CascadeMux I__7922 (
            .O(N__37420),
            .I(N__37417));
    InMux I__7921 (
            .O(N__37417),
            .I(N__37414));
    LocalMux I__7920 (
            .O(N__37414),
            .I(N__37410));
    InMux I__7919 (
            .O(N__37413),
            .I(N__37407));
    Span4Mux_h I__7918 (
            .O(N__37410),
            .I(N__37404));
    LocalMux I__7917 (
            .O(N__37407),
            .I(PIO_dport1_T4_6));
    Odrv4 I__7916 (
            .O(N__37404),
            .I(PIO_dport1_T4_6));
    CascadeMux I__7915 (
            .O(N__37399),
            .I(N__37395));
    InMux I__7914 (
            .O(N__37398),
            .I(N__37392));
    InMux I__7913 (
            .O(N__37395),
            .I(N__37389));
    LocalMux I__7912 (
            .O(N__37392),
            .I(N__37386));
    LocalMux I__7911 (
            .O(N__37389),
            .I(N__37381));
    Span4Mux_v I__7910 (
            .O(N__37386),
            .I(N__37381));
    Odrv4 I__7909 (
            .O(N__37381),
            .I(PIO_dport0_T4_6));
    InMux I__7908 (
            .O(N__37378),
            .I(N__37374));
    InMux I__7907 (
            .O(N__37377),
            .I(N__37371));
    LocalMux I__7906 (
            .O(N__37374),
            .I(N__37365));
    LocalMux I__7905 (
            .O(N__37371),
            .I(N__37360));
    InMux I__7904 (
            .O(N__37370),
            .I(N__37357));
    InMux I__7903 (
            .O(N__37369),
            .I(N__37354));
    InMux I__7902 (
            .O(N__37368),
            .I(N__37351));
    Span4Mux_v I__7901 (
            .O(N__37365),
            .I(N__37348));
    InMux I__7900 (
            .O(N__37364),
            .I(N__37345));
    InMux I__7899 (
            .O(N__37363),
            .I(N__37342));
    Span4Mux_v I__7898 (
            .O(N__37360),
            .I(N__37338));
    LocalMux I__7897 (
            .O(N__37357),
            .I(N__37333));
    LocalMux I__7896 (
            .O(N__37354),
            .I(N__37333));
    LocalMux I__7895 (
            .O(N__37351),
            .I(N__37330));
    Span4Mux_h I__7894 (
            .O(N__37348),
            .I(N__37327));
    LocalMux I__7893 (
            .O(N__37345),
            .I(N__37322));
    LocalMux I__7892 (
            .O(N__37342),
            .I(N__37322));
    InMux I__7891 (
            .O(N__37341),
            .I(N__37319));
    Sp12to4 I__7890 (
            .O(N__37338),
            .I(N__37313));
    Span12Mux_v I__7889 (
            .O(N__37333),
            .I(N__37313));
    Span4Mux_v I__7888 (
            .O(N__37330),
            .I(N__37310));
    Span4Mux_v I__7887 (
            .O(N__37327),
            .I(N__37303));
    Span4Mux_v I__7886 (
            .O(N__37322),
            .I(N__37303));
    LocalMux I__7885 (
            .O(N__37319),
            .I(N__37303));
    InMux I__7884 (
            .O(N__37318),
            .I(N__37300));
    Span12Mux_h I__7883 (
            .O(N__37313),
            .I(N__37297));
    Span4Mux_h I__7882 (
            .O(N__37310),
            .I(N__37292));
    Span4Mux_v I__7881 (
            .O(N__37303),
            .I(N__37292));
    LocalMux I__7880 (
            .O(N__37300),
            .I(N__37289));
    Span12Mux_v I__7879 (
            .O(N__37297),
            .I(N__37284));
    Sp12to4 I__7878 (
            .O(N__37292),
            .I(N__37284));
    Span12Mux_h I__7877 (
            .O(N__37289),
            .I(N__37281));
    Span12Mux_h I__7876 (
            .O(N__37284),
            .I(N__37278));
    Odrv12 I__7875 (
            .O(N__37281),
            .I(wb_dat_i_c_3));
    Odrv12 I__7874 (
            .O(N__37278),
            .I(wb_dat_i_c_3));
    CascadeMux I__7873 (
            .O(N__37273),
            .I(N__37270));
    InMux I__7872 (
            .O(N__37270),
            .I(N__37266));
    InMux I__7871 (
            .O(N__37269),
            .I(N__37263));
    LocalMux I__7870 (
            .O(N__37266),
            .I(N__37260));
    LocalMux I__7869 (
            .O(N__37263),
            .I(N__37257));
    Span4Mux_v I__7868 (
            .O(N__37260),
            .I(N__37254));
    Span4Mux_h I__7867 (
            .O(N__37257),
            .I(N__37251));
    Odrv4 I__7866 (
            .O(N__37254),
            .I(DMA_dev1_Tm_3));
    Odrv4 I__7865 (
            .O(N__37251),
            .I(DMA_dev1_Tm_3));
    InMux I__7864 (
            .O(N__37246),
            .I(N__37242));
    InMux I__7863 (
            .O(N__37245),
            .I(N__37238));
    LocalMux I__7862 (
            .O(N__37242),
            .I(N__37234));
    InMux I__7861 (
            .O(N__37241),
            .I(N__37230));
    LocalMux I__7860 (
            .O(N__37238),
            .I(N__37227));
    InMux I__7859 (
            .O(N__37237),
            .I(N__37222));
    Span4Mux_h I__7858 (
            .O(N__37234),
            .I(N__37218));
    InMux I__7857 (
            .O(N__37233),
            .I(N__37215));
    LocalMux I__7856 (
            .O(N__37230),
            .I(N__37212));
    Span4Mux_v I__7855 (
            .O(N__37227),
            .I(N__37209));
    InMux I__7854 (
            .O(N__37226),
            .I(N__37206));
    InMux I__7853 (
            .O(N__37225),
            .I(N__37203));
    LocalMux I__7852 (
            .O(N__37222),
            .I(N__37200));
    InMux I__7851 (
            .O(N__37221),
            .I(N__37197));
    Span4Mux_v I__7850 (
            .O(N__37218),
            .I(N__37194));
    LocalMux I__7849 (
            .O(N__37215),
            .I(N__37191));
    Span4Mux_v I__7848 (
            .O(N__37212),
            .I(N__37187));
    Sp12to4 I__7847 (
            .O(N__37209),
            .I(N__37182));
    LocalMux I__7846 (
            .O(N__37206),
            .I(N__37182));
    LocalMux I__7845 (
            .O(N__37203),
            .I(N__37179));
    Span4Mux_h I__7844 (
            .O(N__37200),
            .I(N__37176));
    LocalMux I__7843 (
            .O(N__37197),
            .I(N__37173));
    Sp12to4 I__7842 (
            .O(N__37194),
            .I(N__37168));
    Sp12to4 I__7841 (
            .O(N__37191),
            .I(N__37168));
    InMux I__7840 (
            .O(N__37190),
            .I(N__37165));
    Sp12to4 I__7839 (
            .O(N__37187),
            .I(N__37162));
    Span12Mux_v I__7838 (
            .O(N__37182),
            .I(N__37159));
    Sp12to4 I__7837 (
            .O(N__37179),
            .I(N__37152));
    Sp12to4 I__7836 (
            .O(N__37176),
            .I(N__37152));
    Sp12to4 I__7835 (
            .O(N__37173),
            .I(N__37152));
    Span12Mux_v I__7834 (
            .O(N__37168),
            .I(N__37147));
    LocalMux I__7833 (
            .O(N__37165),
            .I(N__37147));
    Span12Mux_h I__7832 (
            .O(N__37162),
            .I(N__37144));
    Span12Mux_h I__7831 (
            .O(N__37159),
            .I(N__37139));
    Span12Mux_v I__7830 (
            .O(N__37152),
            .I(N__37139));
    Span12Mux_h I__7829 (
            .O(N__37147),
            .I(N__37136));
    Span12Mux_v I__7828 (
            .O(N__37144),
            .I(N__37131));
    Span12Mux_h I__7827 (
            .O(N__37139),
            .I(N__37131));
    Span12Mux_h I__7826 (
            .O(N__37136),
            .I(N__37128));
    Odrv12 I__7825 (
            .O(N__37131),
            .I(wb_dat_i_c_4));
    Odrv12 I__7824 (
            .O(N__37128),
            .I(wb_dat_i_c_4));
    InMux I__7823 (
            .O(N__37123),
            .I(N__37120));
    LocalMux I__7822 (
            .O(N__37120),
            .I(N__37117));
    Span4Mux_v I__7821 (
            .O(N__37117),
            .I(N__37114));
    Span4Mux_h I__7820 (
            .O(N__37114),
            .I(N__37111));
    Span4Mux_h I__7819 (
            .O(N__37111),
            .I(N__37108));
    Span4Mux_h I__7818 (
            .O(N__37108),
            .I(N__37105));
    Odrv4 I__7817 (
            .O(N__37105),
            .I(\u0.dat_o_0_0_0_0 ));
    CascadeMux I__7816 (
            .O(N__37102),
            .I(\u0.dat_o_0_0_3_0_cascade_ ));
    InMux I__7815 (
            .O(N__37099),
            .I(N__37096));
    LocalMux I__7814 (
            .O(N__37096),
            .I(N__37092));
    IoInMux I__7813 (
            .O(N__37095),
            .I(N__37089));
    Span4Mux_h I__7812 (
            .O(N__37092),
            .I(N__37086));
    LocalMux I__7811 (
            .O(N__37089),
            .I(N__37083));
    Span4Mux_v I__7810 (
            .O(N__37086),
            .I(N__37080));
    Span12Mux_s3_h I__7809 (
            .O(N__37083),
            .I(N__37076));
    Span4Mux_h I__7808 (
            .O(N__37080),
            .I(N__37073));
    InMux I__7807 (
            .O(N__37079),
            .I(N__37070));
    Odrv12 I__7806 (
            .O(N__37076),
            .I(wb_inta_o_c));
    Odrv4 I__7805 (
            .O(N__37073),
            .I(wb_inta_o_c));
    LocalMux I__7804 (
            .O(N__37070),
            .I(wb_inta_o_c));
    CascadeMux I__7803 (
            .O(N__37063),
            .I(N__37060));
    InMux I__7802 (
            .O(N__37060),
            .I(N__37056));
    InMux I__7801 (
            .O(N__37059),
            .I(N__37053));
    LocalMux I__7800 (
            .O(N__37056),
            .I(N__37050));
    LocalMux I__7799 (
            .O(N__37053),
            .I(N__37047));
    Odrv4 I__7798 (
            .O(N__37050),
            .I(PIO_dport0_T4_0));
    Odrv4 I__7797 (
            .O(N__37047),
            .I(PIO_dport0_T4_0));
    InMux I__7796 (
            .O(N__37042),
            .I(N__37038));
    InMux I__7795 (
            .O(N__37041),
            .I(N__37035));
    LocalMux I__7794 (
            .O(N__37038),
            .I(N__37032));
    LocalMux I__7793 (
            .O(N__37035),
            .I(N__37029));
    Span4Mux_v I__7792 (
            .O(N__37032),
            .I(N__37026));
    Span4Mux_h I__7791 (
            .O(N__37029),
            .I(N__37023));
    Odrv4 I__7790 (
            .O(N__37026),
            .I(PIO_dport1_T4_0));
    Odrv4 I__7789 (
            .O(N__37023),
            .I(PIO_dport1_T4_0));
    CascadeMux I__7788 (
            .O(N__37018),
            .I(N__37014));
    CascadeMux I__7787 (
            .O(N__37017),
            .I(N__37011));
    InMux I__7786 (
            .O(N__37014),
            .I(N__37008));
    InMux I__7785 (
            .O(N__37011),
            .I(N__37005));
    LocalMux I__7784 (
            .O(N__37008),
            .I(N__37002));
    LocalMux I__7783 (
            .O(N__37005),
            .I(N__36999));
    Span4Mux_v I__7782 (
            .O(N__37002),
            .I(N__36994));
    Span4Mux_v I__7781 (
            .O(N__36999),
            .I(N__36994));
    Odrv4 I__7780 (
            .O(N__36994),
            .I(PIO_dport1_T4_2));
    InMux I__7779 (
            .O(N__36991),
            .I(N__36986));
    InMux I__7778 (
            .O(N__36990),
            .I(N__36982));
    InMux I__7777 (
            .O(N__36989),
            .I(N__36978));
    LocalMux I__7776 (
            .O(N__36986),
            .I(N__36975));
    InMux I__7775 (
            .O(N__36985),
            .I(N__36972));
    LocalMux I__7774 (
            .O(N__36982),
            .I(N__36968));
    InMux I__7773 (
            .O(N__36981),
            .I(N__36965));
    LocalMux I__7772 (
            .O(N__36978),
            .I(N__36962));
    Span4Mux_v I__7771 (
            .O(N__36975),
            .I(N__36958));
    LocalMux I__7770 (
            .O(N__36972),
            .I(N__36955));
    InMux I__7769 (
            .O(N__36971),
            .I(N__36952));
    Span4Mux_v I__7768 (
            .O(N__36968),
            .I(N__36948));
    LocalMux I__7767 (
            .O(N__36965),
            .I(N__36945));
    Span4Mux_h I__7766 (
            .O(N__36962),
            .I(N__36942));
    InMux I__7765 (
            .O(N__36961),
            .I(N__36939));
    Sp12to4 I__7764 (
            .O(N__36958),
            .I(N__36935));
    Span4Mux_v I__7763 (
            .O(N__36955),
            .I(N__36930));
    LocalMux I__7762 (
            .O(N__36952),
            .I(N__36930));
    InMux I__7761 (
            .O(N__36951),
            .I(N__36927));
    Span4Mux_h I__7760 (
            .O(N__36948),
            .I(N__36922));
    Span4Mux_v I__7759 (
            .O(N__36945),
            .I(N__36922));
    Span4Mux_v I__7758 (
            .O(N__36942),
            .I(N__36917));
    LocalMux I__7757 (
            .O(N__36939),
            .I(N__36917));
    InMux I__7756 (
            .O(N__36938),
            .I(N__36914));
    Span12Mux_h I__7755 (
            .O(N__36935),
            .I(N__36905));
    Sp12to4 I__7754 (
            .O(N__36930),
            .I(N__36905));
    LocalMux I__7753 (
            .O(N__36927),
            .I(N__36905));
    Sp12to4 I__7752 (
            .O(N__36922),
            .I(N__36905));
    Span4Mux_h I__7751 (
            .O(N__36917),
            .I(N__36900));
    LocalMux I__7750 (
            .O(N__36914),
            .I(N__36900));
    Span12Mux_h I__7749 (
            .O(N__36905),
            .I(N__36897));
    Span4Mux_h I__7748 (
            .O(N__36900),
            .I(N__36894));
    Span12Mux_v I__7747 (
            .O(N__36897),
            .I(N__36891));
    Span4Mux_v I__7746 (
            .O(N__36894),
            .I(N__36888));
    Odrv12 I__7745 (
            .O(N__36891),
            .I(wb_dat_i_c_12));
    Odrv4 I__7744 (
            .O(N__36888),
            .I(wb_dat_i_c_12));
    CascadeMux I__7743 (
            .O(N__36883),
            .I(N__36880));
    InMux I__7742 (
            .O(N__36880),
            .I(N__36876));
    InMux I__7741 (
            .O(N__36879),
            .I(N__36873));
    LocalMux I__7740 (
            .O(N__36876),
            .I(N__36870));
    LocalMux I__7739 (
            .O(N__36873),
            .I(N__36867));
    Span4Mux_v I__7738 (
            .O(N__36870),
            .I(N__36864));
    Span4Mux_h I__7737 (
            .O(N__36867),
            .I(N__36861));
    Odrv4 I__7736 (
            .O(N__36864),
            .I(PIO_cmdport_T2_4));
    Odrv4 I__7735 (
            .O(N__36861),
            .I(PIO_cmdport_T2_4));
    InMux I__7734 (
            .O(N__36856),
            .I(N__36853));
    LocalMux I__7733 (
            .O(N__36853),
            .I(N__36849));
    InMux I__7732 (
            .O(N__36852),
            .I(N__36846));
    Span4Mux_v I__7731 (
            .O(N__36849),
            .I(N__36843));
    LocalMux I__7730 (
            .O(N__36846),
            .I(N__36840));
    Span4Mux_h I__7729 (
            .O(N__36843),
            .I(N__36837));
    Span4Mux_v I__7728 (
            .O(N__36840),
            .I(N__36834));
    Span4Mux_h I__7727 (
            .O(N__36837),
            .I(N__36829));
    Span4Mux_h I__7726 (
            .O(N__36834),
            .I(N__36829));
    Odrv4 I__7725 (
            .O(N__36829),
            .I(DMA_dev1_Teoc_4));
    InMux I__7724 (
            .O(N__36826),
            .I(N__36823));
    LocalMux I__7723 (
            .O(N__36823),
            .I(N__36819));
    InMux I__7722 (
            .O(N__36822),
            .I(N__36816));
    Span4Mux_h I__7721 (
            .O(N__36819),
            .I(N__36811));
    LocalMux I__7720 (
            .O(N__36816),
            .I(N__36811));
    Odrv4 I__7719 (
            .O(N__36811),
            .I(PIO_cmdport_Teoc_4));
    CascadeMux I__7718 (
            .O(N__36808),
            .I(N__36805));
    InMux I__7717 (
            .O(N__36805),
            .I(N__36802));
    LocalMux I__7716 (
            .O(N__36802),
            .I(N__36799));
    Span4Mux_v I__7715 (
            .O(N__36799),
            .I(N__36795));
    InMux I__7714 (
            .O(N__36798),
            .I(N__36792));
    Span4Mux_h I__7713 (
            .O(N__36795),
            .I(N__36787));
    LocalMux I__7712 (
            .O(N__36792),
            .I(N__36787));
    Odrv4 I__7711 (
            .O(N__36787),
            .I(PIO_cmdport_T1_7));
    InMux I__7710 (
            .O(N__36784),
            .I(N__36768));
    InMux I__7709 (
            .O(N__36783),
            .I(N__36765));
    InMux I__7708 (
            .O(N__36782),
            .I(N__36760));
    InMux I__7707 (
            .O(N__36781),
            .I(N__36760));
    InMux I__7706 (
            .O(N__36780),
            .I(N__36755));
    InMux I__7705 (
            .O(N__36779),
            .I(N__36755));
    InMux I__7704 (
            .O(N__36778),
            .I(N__36752));
    InMux I__7703 (
            .O(N__36777),
            .I(N__36749));
    InMux I__7702 (
            .O(N__36776),
            .I(N__36746));
    InMux I__7701 (
            .O(N__36775),
            .I(N__36743));
    InMux I__7700 (
            .O(N__36774),
            .I(N__36731));
    InMux I__7699 (
            .O(N__36773),
            .I(N__36731));
    InMux I__7698 (
            .O(N__36772),
            .I(N__36731));
    InMux I__7697 (
            .O(N__36771),
            .I(N__36731));
    LocalMux I__7696 (
            .O(N__36768),
            .I(N__36727));
    LocalMux I__7695 (
            .O(N__36765),
            .I(N__36720));
    LocalMux I__7694 (
            .O(N__36760),
            .I(N__36720));
    LocalMux I__7693 (
            .O(N__36755),
            .I(N__36720));
    LocalMux I__7692 (
            .O(N__36752),
            .I(N__36715));
    LocalMux I__7691 (
            .O(N__36749),
            .I(N__36715));
    LocalMux I__7690 (
            .O(N__36746),
            .I(N__36710));
    LocalMux I__7689 (
            .O(N__36743),
            .I(N__36710));
    InMux I__7688 (
            .O(N__36742),
            .I(N__36707));
    InMux I__7687 (
            .O(N__36741),
            .I(N__36702));
    InMux I__7686 (
            .O(N__36740),
            .I(N__36702));
    LocalMux I__7685 (
            .O(N__36731),
            .I(N__36699));
    InMux I__7684 (
            .O(N__36730),
            .I(N__36695));
    Sp12to4 I__7683 (
            .O(N__36727),
            .I(N__36691));
    Span4Mux_v I__7682 (
            .O(N__36720),
            .I(N__36688));
    Span4Mux_h I__7681 (
            .O(N__36715),
            .I(N__36685));
    Span4Mux_h I__7680 (
            .O(N__36710),
            .I(N__36678));
    LocalMux I__7679 (
            .O(N__36707),
            .I(N__36678));
    LocalMux I__7678 (
            .O(N__36702),
            .I(N__36678));
    Span4Mux_v I__7677 (
            .O(N__36699),
            .I(N__36675));
    InMux I__7676 (
            .O(N__36698),
            .I(N__36672));
    LocalMux I__7675 (
            .O(N__36695),
            .I(N__36669));
    CascadeMux I__7674 (
            .O(N__36694),
            .I(N__36665));
    Span12Mux_h I__7673 (
            .O(N__36691),
            .I(N__36659));
    Span4Mux_v I__7672 (
            .O(N__36688),
            .I(N__36656));
    Span4Mux_v I__7671 (
            .O(N__36685),
            .I(N__36653));
    Span4Mux_v I__7670 (
            .O(N__36678),
            .I(N__36650));
    Span4Mux_h I__7669 (
            .O(N__36675),
            .I(N__36645));
    LocalMux I__7668 (
            .O(N__36672),
            .I(N__36645));
    Span4Mux_h I__7667 (
            .O(N__36669),
            .I(N__36642));
    InMux I__7666 (
            .O(N__36668),
            .I(N__36639));
    InMux I__7665 (
            .O(N__36665),
            .I(N__36630));
    InMux I__7664 (
            .O(N__36664),
            .I(N__36630));
    InMux I__7663 (
            .O(N__36663),
            .I(N__36630));
    InMux I__7662 (
            .O(N__36662),
            .I(N__36630));
    Odrv12 I__7661 (
            .O(N__36659),
            .I(PIOtip));
    Odrv4 I__7660 (
            .O(N__36656),
            .I(PIOtip));
    Odrv4 I__7659 (
            .O(N__36653),
            .I(PIOtip));
    Odrv4 I__7658 (
            .O(N__36650),
            .I(PIOtip));
    Odrv4 I__7657 (
            .O(N__36645),
            .I(PIOtip));
    Odrv4 I__7656 (
            .O(N__36642),
            .I(PIOtip));
    LocalMux I__7655 (
            .O(N__36639),
            .I(PIOtip));
    LocalMux I__7654 (
            .O(N__36630),
            .I(PIOtip));
    InMux I__7653 (
            .O(N__36613),
            .I(N__36610));
    LocalMux I__7652 (
            .O(N__36610),
            .I(N__36606));
    InMux I__7651 (
            .O(N__36609),
            .I(N__36603));
    Span4Mux_v I__7650 (
            .O(N__36606),
            .I(N__36600));
    LocalMux I__7649 (
            .O(N__36603),
            .I(N__36597));
    Span4Mux_h I__7648 (
            .O(N__36600),
            .I(N__36594));
    Odrv12 I__7647 (
            .O(N__36597),
            .I(PIO_dport0_T1_7));
    Odrv4 I__7646 (
            .O(N__36594),
            .I(PIO_dport0_T1_7));
    InMux I__7645 (
            .O(N__36589),
            .I(N__36586));
    LocalMux I__7644 (
            .O(N__36586),
            .I(N__36583));
    Odrv12 I__7643 (
            .O(N__36583),
            .I(\u0.dat_o_0_0_0_7 ));
    CascadeMux I__7642 (
            .O(N__36580),
            .I(\u0.dat_o_0_0_3_7_cascade_ ));
    CascadeMux I__7641 (
            .O(N__36577),
            .I(N__36574));
    InMux I__7640 (
            .O(N__36574),
            .I(N__36571));
    LocalMux I__7639 (
            .O(N__36571),
            .I(N__36567));
    InMux I__7638 (
            .O(N__36570),
            .I(N__36564));
    Span4Mux_v I__7637 (
            .O(N__36567),
            .I(N__36561));
    LocalMux I__7636 (
            .O(N__36564),
            .I(N__36558));
    Odrv4 I__7635 (
            .O(N__36561),
            .I(PIO_cmdport_T1_0));
    Odrv12 I__7634 (
            .O(N__36558),
            .I(PIO_cmdport_T1_0));
    InMux I__7633 (
            .O(N__36553),
            .I(N__36544));
    InMux I__7632 (
            .O(N__36552),
            .I(N__36544));
    InMux I__7631 (
            .O(N__36551),
            .I(N__36539));
    InMux I__7630 (
            .O(N__36550),
            .I(N__36539));
    CascadeMux I__7629 (
            .O(N__36549),
            .I(N__36531));
    LocalMux I__7628 (
            .O(N__36544),
            .I(N__36526));
    LocalMux I__7627 (
            .O(N__36539),
            .I(N__36523));
    InMux I__7626 (
            .O(N__36538),
            .I(N__36520));
    InMux I__7625 (
            .O(N__36537),
            .I(N__36517));
    InMux I__7624 (
            .O(N__36536),
            .I(N__36512));
    InMux I__7623 (
            .O(N__36535),
            .I(N__36512));
    InMux I__7622 (
            .O(N__36534),
            .I(N__36509));
    InMux I__7621 (
            .O(N__36531),
            .I(N__36504));
    InMux I__7620 (
            .O(N__36530),
            .I(N__36504));
    CascadeMux I__7619 (
            .O(N__36529),
            .I(N__36500));
    Span4Mux_h I__7618 (
            .O(N__36526),
            .I(N__36495));
    Span4Mux_h I__7617 (
            .O(N__36523),
            .I(N__36488));
    LocalMux I__7616 (
            .O(N__36520),
            .I(N__36488));
    LocalMux I__7615 (
            .O(N__36517),
            .I(N__36488));
    LocalMux I__7614 (
            .O(N__36512),
            .I(N__36485));
    LocalMux I__7613 (
            .O(N__36509),
            .I(N__36482));
    LocalMux I__7612 (
            .O(N__36504),
            .I(N__36479));
    InMux I__7611 (
            .O(N__36503),
            .I(N__36474));
    InMux I__7610 (
            .O(N__36500),
            .I(N__36474));
    InMux I__7609 (
            .O(N__36499),
            .I(N__36471));
    InMux I__7608 (
            .O(N__36498),
            .I(N__36468));
    Span4Mux_h I__7607 (
            .O(N__36495),
            .I(N__36465));
    Span4Mux_h I__7606 (
            .O(N__36488),
            .I(N__36460));
    Span4Mux_h I__7605 (
            .O(N__36485),
            .I(N__36460));
    Span4Mux_v I__7604 (
            .O(N__36482),
            .I(N__36453));
    Span4Mux_v I__7603 (
            .O(N__36479),
            .I(N__36453));
    LocalMux I__7602 (
            .O(N__36474),
            .I(N__36453));
    LocalMux I__7601 (
            .O(N__36471),
            .I(N__36448));
    LocalMux I__7600 (
            .O(N__36468),
            .I(N__36448));
    Odrv4 I__7599 (
            .O(N__36465),
            .I(\u1.DMA_control.readDlw_3 ));
    Odrv4 I__7598 (
            .O(N__36460),
            .I(\u1.DMA_control.readDlw_3 ));
    Odrv4 I__7597 (
            .O(N__36453),
            .I(\u1.DMA_control.readDlw_3 ));
    Odrv12 I__7596 (
            .O(N__36448),
            .I(\u1.DMA_control.readDlw_3 ));
    CascadeMux I__7595 (
            .O(N__36439),
            .I(N__36432));
    CascadeMux I__7594 (
            .O(N__36438),
            .I(N__36428));
    InMux I__7593 (
            .O(N__36437),
            .I(N__36421));
    InMux I__7592 (
            .O(N__36436),
            .I(N__36421));
    CascadeMux I__7591 (
            .O(N__36435),
            .I(N__36418));
    InMux I__7590 (
            .O(N__36432),
            .I(N__36413));
    InMux I__7589 (
            .O(N__36431),
            .I(N__36413));
    InMux I__7588 (
            .O(N__36428),
            .I(N__36404));
    InMux I__7587 (
            .O(N__36427),
            .I(N__36404));
    InMux I__7586 (
            .O(N__36426),
            .I(N__36399));
    LocalMux I__7585 (
            .O(N__36421),
            .I(N__36396));
    InMux I__7584 (
            .O(N__36418),
            .I(N__36393));
    LocalMux I__7583 (
            .O(N__36413),
            .I(N__36390));
    InMux I__7582 (
            .O(N__36412),
            .I(N__36385));
    InMux I__7581 (
            .O(N__36411),
            .I(N__36385));
    InMux I__7580 (
            .O(N__36410),
            .I(N__36380));
    InMux I__7579 (
            .O(N__36409),
            .I(N__36380));
    LocalMux I__7578 (
            .O(N__36404),
            .I(N__36377));
    InMux I__7577 (
            .O(N__36403),
            .I(N__36374));
    InMux I__7576 (
            .O(N__36402),
            .I(N__36371));
    LocalMux I__7575 (
            .O(N__36399),
            .I(N__36366));
    Span4Mux_h I__7574 (
            .O(N__36396),
            .I(N__36366));
    LocalMux I__7573 (
            .O(N__36393),
            .I(N__36361));
    Span4Mux_h I__7572 (
            .O(N__36390),
            .I(N__36361));
    LocalMux I__7571 (
            .O(N__36385),
            .I(N__36354));
    LocalMux I__7570 (
            .O(N__36380),
            .I(N__36354));
    Span4Mux_v I__7569 (
            .O(N__36377),
            .I(N__36354));
    LocalMux I__7568 (
            .O(N__36374),
            .I(N__36347));
    LocalMux I__7567 (
            .O(N__36371),
            .I(N__36347));
    Span4Mux_v I__7566 (
            .O(N__36366),
            .I(N__36347));
    Span4Mux_h I__7565 (
            .O(N__36361),
            .I(N__36344));
    Span4Mux_h I__7564 (
            .O(N__36354),
            .I(N__36341));
    Span4Mux_h I__7563 (
            .O(N__36347),
            .I(N__36338));
    Odrv4 I__7562 (
            .O(N__36344),
            .I(\u1.DMA_control.readDfw_3 ));
    Odrv4 I__7561 (
            .O(N__36341),
            .I(\u1.DMA_control.readDfw_3 ));
    Odrv4 I__7560 (
            .O(N__36338),
            .I(\u1.DMA_control.readDfw_3 ));
    InMux I__7559 (
            .O(N__36331),
            .I(N__36328));
    LocalMux I__7558 (
            .O(N__36328),
            .I(N__36318));
    CEMux I__7557 (
            .O(N__36327),
            .I(N__36301));
    CEMux I__7556 (
            .O(N__36326),
            .I(N__36301));
    CEMux I__7555 (
            .O(N__36325),
            .I(N__36301));
    CEMux I__7554 (
            .O(N__36324),
            .I(N__36301));
    CEMux I__7553 (
            .O(N__36323),
            .I(N__36301));
    CEMux I__7552 (
            .O(N__36322),
            .I(N__36301));
    CEMux I__7551 (
            .O(N__36321),
            .I(N__36301));
    Glb2LocalMux I__7550 (
            .O(N__36318),
            .I(N__36301));
    GlobalMux I__7549 (
            .O(N__36301),
            .I(N__36298));
    gio2CtrlBuf I__7548 (
            .O(N__36298),
            .I(\u1.DMA_control.rd_dstrb_g ));
    InMux I__7547 (
            .O(N__36295),
            .I(N__36292));
    LocalMux I__7546 (
            .O(N__36292),
            .I(N__36279));
    InMux I__7545 (
            .O(N__36291),
            .I(N__36276));
    InMux I__7544 (
            .O(N__36290),
            .I(N__36273));
    InMux I__7543 (
            .O(N__36289),
            .I(N__36258));
    InMux I__7542 (
            .O(N__36288),
            .I(N__36258));
    InMux I__7541 (
            .O(N__36287),
            .I(N__36258));
    InMux I__7540 (
            .O(N__36286),
            .I(N__36258));
    InMux I__7539 (
            .O(N__36285),
            .I(N__36258));
    InMux I__7538 (
            .O(N__36284),
            .I(N__36258));
    InMux I__7537 (
            .O(N__36283),
            .I(N__36258));
    InMux I__7536 (
            .O(N__36282),
            .I(N__36248));
    Span4Mux_v I__7535 (
            .O(N__36279),
            .I(N__36245));
    LocalMux I__7534 (
            .O(N__36276),
            .I(N__36242));
    LocalMux I__7533 (
            .O(N__36273),
            .I(N__36238));
    LocalMux I__7532 (
            .O(N__36258),
            .I(N__36235));
    InMux I__7531 (
            .O(N__36257),
            .I(N__36232));
    InMux I__7530 (
            .O(N__36256),
            .I(N__36218));
    InMux I__7529 (
            .O(N__36255),
            .I(N__36218));
    InMux I__7528 (
            .O(N__36254),
            .I(N__36218));
    InMux I__7527 (
            .O(N__36253),
            .I(N__36218));
    InMux I__7526 (
            .O(N__36252),
            .I(N__36213));
    CascadeMux I__7525 (
            .O(N__36251),
            .I(N__36210));
    LocalMux I__7524 (
            .O(N__36248),
            .I(N__36205));
    Span4Mux_v I__7523 (
            .O(N__36245),
            .I(N__36202));
    Sp12to4 I__7522 (
            .O(N__36242),
            .I(N__36199));
    InMux I__7521 (
            .O(N__36241),
            .I(N__36196));
    Span4Mux_v I__7520 (
            .O(N__36238),
            .I(N__36191));
    Span4Mux_v I__7519 (
            .O(N__36235),
            .I(N__36191));
    LocalMux I__7518 (
            .O(N__36232),
            .I(N__36188));
    InMux I__7517 (
            .O(N__36231),
            .I(N__36177));
    InMux I__7516 (
            .O(N__36230),
            .I(N__36177));
    InMux I__7515 (
            .O(N__36229),
            .I(N__36177));
    InMux I__7514 (
            .O(N__36228),
            .I(N__36177));
    InMux I__7513 (
            .O(N__36227),
            .I(N__36177));
    LocalMux I__7512 (
            .O(N__36218),
            .I(N__36174));
    InMux I__7511 (
            .O(N__36217),
            .I(N__36171));
    CascadeMux I__7510 (
            .O(N__36216),
            .I(N__36167));
    LocalMux I__7509 (
            .O(N__36213),
            .I(N__36164));
    InMux I__7508 (
            .O(N__36210),
            .I(N__36161));
    InMux I__7507 (
            .O(N__36209),
            .I(N__36158));
    InMux I__7506 (
            .O(N__36208),
            .I(N__36155));
    Span12Mux_v I__7505 (
            .O(N__36205),
            .I(N__36152));
    Sp12to4 I__7504 (
            .O(N__36202),
            .I(N__36145));
    Span12Mux_s11_v I__7503 (
            .O(N__36199),
            .I(N__36145));
    LocalMux I__7502 (
            .O(N__36196),
            .I(N__36145));
    Span4Mux_h I__7501 (
            .O(N__36191),
            .I(N__36138));
    Span4Mux_v I__7500 (
            .O(N__36188),
            .I(N__36138));
    LocalMux I__7499 (
            .O(N__36177),
            .I(N__36138));
    Span4Mux_v I__7498 (
            .O(N__36174),
            .I(N__36133));
    LocalMux I__7497 (
            .O(N__36171),
            .I(N__36133));
    InMux I__7496 (
            .O(N__36170),
            .I(N__36128));
    InMux I__7495 (
            .O(N__36167),
            .I(N__36128));
    Span4Mux_v I__7494 (
            .O(N__36164),
            .I(N__36125));
    LocalMux I__7493 (
            .O(N__36161),
            .I(N__36120));
    LocalMux I__7492 (
            .O(N__36158),
            .I(N__36120));
    LocalMux I__7491 (
            .O(N__36155),
            .I(\u1.SelDev ));
    Odrv12 I__7490 (
            .O(N__36152),
            .I(\u1.SelDev ));
    Odrv12 I__7489 (
            .O(N__36145),
            .I(\u1.SelDev ));
    Odrv4 I__7488 (
            .O(N__36138),
            .I(\u1.SelDev ));
    Odrv4 I__7487 (
            .O(N__36133),
            .I(\u1.SelDev ));
    LocalMux I__7486 (
            .O(N__36128),
            .I(\u1.SelDev ));
    Odrv4 I__7485 (
            .O(N__36125),
            .I(\u1.SelDev ));
    Odrv4 I__7484 (
            .O(N__36120),
            .I(\u1.SelDev ));
    InMux I__7483 (
            .O(N__36103),
            .I(N__36100));
    LocalMux I__7482 (
            .O(N__36100),
            .I(N__36097));
    Span12Mux_v I__7481 (
            .O(N__36097),
            .I(N__36094));
    Odrv12 I__7480 (
            .O(N__36094),
            .I(\u1.DMA_control.Tm_7 ));
    CascadeMux I__7479 (
            .O(N__36091),
            .I(N__36087));
    CascadeMux I__7478 (
            .O(N__36090),
            .I(N__36084));
    InMux I__7477 (
            .O(N__36087),
            .I(N__36081));
    InMux I__7476 (
            .O(N__36084),
            .I(N__36078));
    LocalMux I__7475 (
            .O(N__36081),
            .I(N__36075));
    LocalMux I__7474 (
            .O(N__36078),
            .I(N__36072));
    Span4Mux_v I__7473 (
            .O(N__36075),
            .I(N__36067));
    Span4Mux_v I__7472 (
            .O(N__36072),
            .I(N__36067));
    Odrv4 I__7471 (
            .O(N__36067),
            .I(PIO_dport1_T1_7));
    InMux I__7470 (
            .O(N__36064),
            .I(N__36060));
    InMux I__7469 (
            .O(N__36063),
            .I(N__36057));
    LocalMux I__7468 (
            .O(N__36060),
            .I(N__36054));
    LocalMux I__7467 (
            .O(N__36057),
            .I(N__36051));
    Span4Mux_h I__7466 (
            .O(N__36054),
            .I(N__36048));
    Odrv4 I__7465 (
            .O(N__36051),
            .I(PIO_dport0_T1_4));
    Odrv4 I__7464 (
            .O(N__36048),
            .I(PIO_dport0_T1_4));
    CascadeMux I__7463 (
            .O(N__36043),
            .I(N__36039));
    InMux I__7462 (
            .O(N__36042),
            .I(N__36036));
    InMux I__7461 (
            .O(N__36039),
            .I(N__36033));
    LocalMux I__7460 (
            .O(N__36036),
            .I(N__36030));
    LocalMux I__7459 (
            .O(N__36033),
            .I(N__36027));
    Span4Mux_v I__7458 (
            .O(N__36030),
            .I(N__36022));
    Span4Mux_h I__7457 (
            .O(N__36027),
            .I(N__36022));
    Odrv4 I__7456 (
            .O(N__36022),
            .I(PIO_dport0_T2_0));
    InMux I__7455 (
            .O(N__36019),
            .I(N__36014));
    CascadeMux I__7454 (
            .O(N__36018),
            .I(N__36011));
    InMux I__7453 (
            .O(N__36017),
            .I(N__36007));
    LocalMux I__7452 (
            .O(N__36014),
            .I(N__36004));
    InMux I__7451 (
            .O(N__36011),
            .I(N__36001));
    InMux I__7450 (
            .O(N__36010),
            .I(N__35998));
    LocalMux I__7449 (
            .O(N__36007),
            .I(N__35995));
    Span4Mux_s3_h I__7448 (
            .O(N__36004),
            .I(N__35991));
    LocalMux I__7447 (
            .O(N__36001),
            .I(N__35986));
    LocalMux I__7446 (
            .O(N__35998),
            .I(N__35986));
    Span4Mux_v I__7445 (
            .O(N__35995),
            .I(N__35982));
    InMux I__7444 (
            .O(N__35994),
            .I(N__35979));
    Span4Mux_h I__7443 (
            .O(N__35991),
            .I(N__35974));
    Span4Mux_v I__7442 (
            .O(N__35986),
            .I(N__35974));
    InMux I__7441 (
            .O(N__35985),
            .I(N__35971));
    Span4Mux_v I__7440 (
            .O(N__35982),
            .I(N__35966));
    LocalMux I__7439 (
            .O(N__35979),
            .I(N__35966));
    Span4Mux_h I__7438 (
            .O(N__35974),
            .I(N__35960));
    LocalMux I__7437 (
            .O(N__35971),
            .I(N__35960));
    Span4Mux_h I__7436 (
            .O(N__35966),
            .I(N__35957));
    InMux I__7435 (
            .O(N__35965),
            .I(N__35954));
    Span4Mux_h I__7434 (
            .O(N__35960),
            .I(N__35949));
    Span4Mux_h I__7433 (
            .O(N__35957),
            .I(N__35944));
    LocalMux I__7432 (
            .O(N__35954),
            .I(N__35944));
    InMux I__7431 (
            .O(N__35953),
            .I(N__35941));
    InMux I__7430 (
            .O(N__35952),
            .I(N__35938));
    Span4Mux_v I__7429 (
            .O(N__35949),
            .I(N__35935));
    Span4Mux_v I__7428 (
            .O(N__35944),
            .I(N__35932));
    LocalMux I__7427 (
            .O(N__35941),
            .I(N__35927));
    LocalMux I__7426 (
            .O(N__35938),
            .I(N__35927));
    Sp12to4 I__7425 (
            .O(N__35935),
            .I(N__35924));
    Span4Mux_h I__7424 (
            .O(N__35932),
            .I(N__35921));
    Span4Mux_v I__7423 (
            .O(N__35927),
            .I(N__35918));
    Span12Mux_v I__7422 (
            .O(N__35924),
            .I(N__35911));
    Sp12to4 I__7421 (
            .O(N__35921),
            .I(N__35911));
    Sp12to4 I__7420 (
            .O(N__35918),
            .I(N__35911));
    Span12Mux_h I__7419 (
            .O(N__35911),
            .I(N__35908));
    Odrv12 I__7418 (
            .O(N__35908),
            .I(wb_dat_i_c_9));
    CEMux I__7417 (
            .O(N__35905),
            .I(N__35902));
    LocalMux I__7416 (
            .O(N__35902),
            .I(N__35896));
    CEMux I__7415 (
            .O(N__35901),
            .I(N__35893));
    CEMux I__7414 (
            .O(N__35900),
            .I(N__35887));
    CEMux I__7413 (
            .O(N__35899),
            .I(N__35884));
    Span4Mux_h I__7412 (
            .O(N__35896),
            .I(N__35879));
    LocalMux I__7411 (
            .O(N__35893),
            .I(N__35879));
    CEMux I__7410 (
            .O(N__35892),
            .I(N__35875));
    CEMux I__7409 (
            .O(N__35891),
            .I(N__35872));
    CEMux I__7408 (
            .O(N__35890),
            .I(N__35869));
    LocalMux I__7407 (
            .O(N__35887),
            .I(N__35866));
    LocalMux I__7406 (
            .O(N__35884),
            .I(N__35863));
    Span4Mux_s2_v I__7405 (
            .O(N__35879),
            .I(N__35860));
    CEMux I__7404 (
            .O(N__35878),
            .I(N__35857));
    LocalMux I__7403 (
            .O(N__35875),
            .I(N__35852));
    LocalMux I__7402 (
            .O(N__35872),
            .I(N__35852));
    LocalMux I__7401 (
            .O(N__35869),
            .I(N__35849));
    Span4Mux_v I__7400 (
            .O(N__35866),
            .I(N__35846));
    Span4Mux_v I__7399 (
            .O(N__35863),
            .I(N__35843));
    Span4Mux_h I__7398 (
            .O(N__35860),
            .I(N__35840));
    LocalMux I__7397 (
            .O(N__35857),
            .I(N__35837));
    Span4Mux_h I__7396 (
            .O(N__35852),
            .I(N__35834));
    Span4Mux_v I__7395 (
            .O(N__35849),
            .I(N__35827));
    Span4Mux_h I__7394 (
            .O(N__35846),
            .I(N__35827));
    Span4Mux_h I__7393 (
            .O(N__35843),
            .I(N__35827));
    Span4Mux_v I__7392 (
            .O(N__35840),
            .I(N__35824));
    Odrv12 I__7391 (
            .O(N__35837),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_awe0 ));
    Odrv4 I__7390 (
            .O(N__35834),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_awe0 ));
    Odrv4 I__7389 (
            .O(N__35827),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_awe0 ));
    Odrv4 I__7388 (
            .O(N__35824),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_awe0 ));
    InMux I__7387 (
            .O(N__35815),
            .I(N__35812));
    LocalMux I__7386 (
            .O(N__35812),
            .I(N__35809));
    Span4Mux_h I__7385 (
            .O(N__35809),
            .I(N__35806));
    Odrv4 I__7384 (
            .O(N__35806),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_11 ));
    InMux I__7383 (
            .O(N__35803),
            .I(N__35800));
    LocalMux I__7382 (
            .O(N__35800),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_11 ));
    CascadeMux I__7381 (
            .O(N__35797),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIQGUQZ0Z_11_cascade_ ));
    InMux I__7380 (
            .O(N__35794),
            .I(N__35791));
    LocalMux I__7379 (
            .O(N__35791),
            .I(N__35788));
    Span12Mux_h I__7378 (
            .O(N__35788),
            .I(N__35785));
    Odrv12 I__7377 (
            .O(N__35785),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIU47KZ0Z_11 ));
    InMux I__7376 (
            .O(N__35782),
            .I(N__35779));
    LocalMux I__7375 (
            .O(N__35779),
            .I(N__35776));
    Span4Mux_v I__7374 (
            .O(N__35776),
            .I(N__35773));
    Odrv4 I__7373 (
            .O(N__35773),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_16 ));
    InMux I__7372 (
            .O(N__35770),
            .I(N__35767));
    LocalMux I__7371 (
            .O(N__35767),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_16 ));
    InMux I__7370 (
            .O(N__35764),
            .I(N__35761));
    LocalMux I__7369 (
            .O(N__35761),
            .I(N__35758));
    Odrv12 I__7368 (
            .O(N__35758),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_11 ));
    InMux I__7367 (
            .O(N__35755),
            .I(N__35752));
    LocalMux I__7366 (
            .O(N__35752),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_11 ));
    InMux I__7365 (
            .O(N__35749),
            .I(N__35746));
    LocalMux I__7364 (
            .O(N__35746),
            .I(N__35743));
    Odrv12 I__7363 (
            .O(N__35743),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_27 ));
    InMux I__7362 (
            .O(N__35740),
            .I(N__35737));
    LocalMux I__7361 (
            .O(N__35737),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_0 ));
    InMux I__7360 (
            .O(N__35734),
            .I(N__35731));
    LocalMux I__7359 (
            .O(N__35731),
            .I(N__35728));
    Odrv4 I__7358 (
            .O(N__35728),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_1 ));
    InMux I__7357 (
            .O(N__35725),
            .I(N__35722));
    LocalMux I__7356 (
            .O(N__35722),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_1 ));
    InMux I__7355 (
            .O(N__35719),
            .I(N__35716));
    LocalMux I__7354 (
            .O(N__35716),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_27 ));
    InMux I__7353 (
            .O(N__35713),
            .I(N__35710));
    LocalMux I__7352 (
            .O(N__35710),
            .I(N__35707));
    Odrv12 I__7351 (
            .O(N__35707),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_27 ));
    InMux I__7350 (
            .O(N__35704),
            .I(N__35701));
    LocalMux I__7349 (
            .O(N__35701),
            .I(N__35698));
    Span4Mux_h I__7348 (
            .O(N__35698),
            .I(N__35695));
    Odrv4 I__7347 (
            .O(N__35695),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_27 ));
    InMux I__7346 (
            .O(N__35692),
            .I(N__35689));
    LocalMux I__7345 (
            .O(N__35689),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI811RZ0Z_27 ));
    CascadeMux I__7344 (
            .O(N__35686),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNICL9KZ0Z_27_cascade_ ));
    CascadeMux I__7343 (
            .O(N__35683),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI61IM1Z0Z_2_cascade_ ));
    InMux I__7342 (
            .O(N__35680),
            .I(N__35677));
    LocalMux I__7341 (
            .O(N__35677),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_27 ));
    InMux I__7340 (
            .O(N__35674),
            .I(N__35671));
    LocalMux I__7339 (
            .O(N__35671),
            .I(N__35661));
    InMux I__7338 (
            .O(N__35670),
            .I(N__35658));
    InMux I__7337 (
            .O(N__35669),
            .I(N__35655));
    InMux I__7336 (
            .O(N__35668),
            .I(N__35648));
    InMux I__7335 (
            .O(N__35667),
            .I(N__35648));
    InMux I__7334 (
            .O(N__35666),
            .I(N__35645));
    InMux I__7333 (
            .O(N__35665),
            .I(N__35642));
    CascadeMux I__7332 (
            .O(N__35664),
            .I(N__35639));
    Span4Mux_v I__7331 (
            .O(N__35661),
            .I(N__35634));
    LocalMux I__7330 (
            .O(N__35658),
            .I(N__35629));
    LocalMux I__7329 (
            .O(N__35655),
            .I(N__35629));
    InMux I__7328 (
            .O(N__35654),
            .I(N__35626));
    InMux I__7327 (
            .O(N__35653),
            .I(N__35623));
    LocalMux I__7326 (
            .O(N__35648),
            .I(N__35620));
    LocalMux I__7325 (
            .O(N__35645),
            .I(N__35617));
    LocalMux I__7324 (
            .O(N__35642),
            .I(N__35614));
    InMux I__7323 (
            .O(N__35639),
            .I(N__35609));
    InMux I__7322 (
            .O(N__35638),
            .I(N__35609));
    CascadeMux I__7321 (
            .O(N__35637),
            .I(N__35606));
    Sp12to4 I__7320 (
            .O(N__35634),
            .I(N__35594));
    Span12Mux_s8_v I__7319 (
            .O(N__35629),
            .I(N__35594));
    LocalMux I__7318 (
            .O(N__35626),
            .I(N__35594));
    LocalMux I__7317 (
            .O(N__35623),
            .I(N__35594));
    Span4Mux_h I__7316 (
            .O(N__35620),
            .I(N__35591));
    Span4Mux_v I__7315 (
            .O(N__35617),
            .I(N__35584));
    Span4Mux_v I__7314 (
            .O(N__35614),
            .I(N__35584));
    LocalMux I__7313 (
            .O(N__35609),
            .I(N__35584));
    InMux I__7312 (
            .O(N__35606),
            .I(N__35579));
    InMux I__7311 (
            .O(N__35605),
            .I(N__35579));
    InMux I__7310 (
            .O(N__35604),
            .I(N__35576));
    InMux I__7309 (
            .O(N__35603),
            .I(N__35573));
    Odrv12 I__7308 (
            .O(N__35594),
            .I(\u1.DMA_control.readDlw_5 ));
    Odrv4 I__7307 (
            .O(N__35591),
            .I(\u1.DMA_control.readDlw_5 ));
    Odrv4 I__7306 (
            .O(N__35584),
            .I(\u1.DMA_control.readDlw_5 ));
    LocalMux I__7305 (
            .O(N__35579),
            .I(\u1.DMA_control.readDlw_5 ));
    LocalMux I__7304 (
            .O(N__35576),
            .I(\u1.DMA_control.readDlw_5 ));
    LocalMux I__7303 (
            .O(N__35573),
            .I(\u1.DMA_control.readDlw_5 ));
    InMux I__7302 (
            .O(N__35560),
            .I(N__35553));
    InMux I__7301 (
            .O(N__35559),
            .I(N__35542));
    InMux I__7300 (
            .O(N__35558),
            .I(N__35542));
    InMux I__7299 (
            .O(N__35557),
            .I(N__35537));
    InMux I__7298 (
            .O(N__35556),
            .I(N__35537));
    LocalMux I__7297 (
            .O(N__35553),
            .I(N__35534));
    InMux I__7296 (
            .O(N__35552),
            .I(N__35531));
    InMux I__7295 (
            .O(N__35551),
            .I(N__35526));
    InMux I__7294 (
            .O(N__35550),
            .I(N__35526));
    InMux I__7293 (
            .O(N__35549),
            .I(N__35521));
    InMux I__7292 (
            .O(N__35548),
            .I(N__35521));
    CascadeMux I__7291 (
            .O(N__35547),
            .I(N__35518));
    LocalMux I__7290 (
            .O(N__35542),
            .I(N__35514));
    LocalMux I__7289 (
            .O(N__35537),
            .I(N__35511));
    Span4Mux_s3_v I__7288 (
            .O(N__35534),
            .I(N__35504));
    LocalMux I__7287 (
            .O(N__35531),
            .I(N__35504));
    LocalMux I__7286 (
            .O(N__35526),
            .I(N__35504));
    LocalMux I__7285 (
            .O(N__35521),
            .I(N__35501));
    InMux I__7284 (
            .O(N__35518),
            .I(N__35496));
    InMux I__7283 (
            .O(N__35517),
            .I(N__35496));
    Span4Mux_h I__7282 (
            .O(N__35514),
            .I(N__35491));
    Span4Mux_v I__7281 (
            .O(N__35511),
            .I(N__35482));
    Span4Mux_v I__7280 (
            .O(N__35504),
            .I(N__35482));
    Span4Mux_h I__7279 (
            .O(N__35501),
            .I(N__35482));
    LocalMux I__7278 (
            .O(N__35496),
            .I(N__35482));
    InMux I__7277 (
            .O(N__35495),
            .I(N__35477));
    InMux I__7276 (
            .O(N__35494),
            .I(N__35477));
    Span4Mux_h I__7275 (
            .O(N__35491),
            .I(N__35474));
    Span4Mux_h I__7274 (
            .O(N__35482),
            .I(N__35471));
    LocalMux I__7273 (
            .O(N__35477),
            .I(N__35468));
    Odrv4 I__7272 (
            .O(N__35474),
            .I(\u1.DMA_control.readDfw_5 ));
    Odrv4 I__7271 (
            .O(N__35471),
            .I(\u1.DMA_control.readDfw_5 ));
    Odrv4 I__7270 (
            .O(N__35468),
            .I(\u1.DMA_control.readDfw_5 ));
    InMux I__7269 (
            .O(N__35461),
            .I(N__35458));
    LocalMux I__7268 (
            .O(N__35458),
            .I(N__35455));
    Span4Mux_h I__7267 (
            .O(N__35455),
            .I(N__35452));
    Odrv4 I__7266 (
            .O(N__35452),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_9 ));
    InMux I__7265 (
            .O(N__35449),
            .I(N__35446));
    LocalMux I__7264 (
            .O(N__35446),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_9 ));
    CascadeMux I__7263 (
            .O(N__35443),
            .I(N__35434));
    CascadeMux I__7262 (
            .O(N__35442),
            .I(N__35431));
    CascadeMux I__7261 (
            .O(N__35441),
            .I(N__35428));
    InMux I__7260 (
            .O(N__35440),
            .I(N__35421));
    InMux I__7259 (
            .O(N__35439),
            .I(N__35421));
    InMux I__7258 (
            .O(N__35438),
            .I(N__35416));
    InMux I__7257 (
            .O(N__35437),
            .I(N__35413));
    InMux I__7256 (
            .O(N__35434),
            .I(N__35410));
    InMux I__7255 (
            .O(N__35431),
            .I(N__35407));
    InMux I__7254 (
            .O(N__35428),
            .I(N__35402));
    InMux I__7253 (
            .O(N__35427),
            .I(N__35402));
    InMux I__7252 (
            .O(N__35426),
            .I(N__35399));
    LocalMux I__7251 (
            .O(N__35421),
            .I(N__35395));
    InMux I__7250 (
            .O(N__35420),
            .I(N__35390));
    InMux I__7249 (
            .O(N__35419),
            .I(N__35390));
    LocalMux I__7248 (
            .O(N__35416),
            .I(N__35379));
    LocalMux I__7247 (
            .O(N__35413),
            .I(N__35379));
    LocalMux I__7246 (
            .O(N__35410),
            .I(N__35379));
    LocalMux I__7245 (
            .O(N__35407),
            .I(N__35379));
    LocalMux I__7244 (
            .O(N__35402),
            .I(N__35379));
    LocalMux I__7243 (
            .O(N__35399),
            .I(N__35376));
    InMux I__7242 (
            .O(N__35398),
            .I(N__35370));
    Span4Mux_h I__7241 (
            .O(N__35395),
            .I(N__35365));
    LocalMux I__7240 (
            .O(N__35390),
            .I(N__35365));
    Span4Mux_v I__7239 (
            .O(N__35379),
            .I(N__35360));
    Span4Mux_h I__7238 (
            .O(N__35376),
            .I(N__35360));
    InMux I__7237 (
            .O(N__35375),
            .I(N__35357));
    InMux I__7236 (
            .O(N__35374),
            .I(N__35352));
    InMux I__7235 (
            .O(N__35373),
            .I(N__35352));
    LocalMux I__7234 (
            .O(N__35370),
            .I(\u1.DMA_control.readDlw_9 ));
    Odrv4 I__7233 (
            .O(N__35365),
            .I(\u1.DMA_control.readDlw_9 ));
    Odrv4 I__7232 (
            .O(N__35360),
            .I(\u1.DMA_control.readDlw_9 ));
    LocalMux I__7231 (
            .O(N__35357),
            .I(\u1.DMA_control.readDlw_9 ));
    LocalMux I__7230 (
            .O(N__35352),
            .I(\u1.DMA_control.readDlw_9 ));
    InMux I__7229 (
            .O(N__35341),
            .I(N__35332));
    InMux I__7228 (
            .O(N__35340),
            .I(N__35329));
    InMux I__7227 (
            .O(N__35339),
            .I(N__35324));
    InMux I__7226 (
            .O(N__35338),
            .I(N__35324));
    InMux I__7225 (
            .O(N__35337),
            .I(N__35320));
    InMux I__7224 (
            .O(N__35336),
            .I(N__35317));
    CascadeMux I__7223 (
            .O(N__35335),
            .I(N__35314));
    LocalMux I__7222 (
            .O(N__35332),
            .I(N__35307));
    LocalMux I__7221 (
            .O(N__35329),
            .I(N__35304));
    LocalMux I__7220 (
            .O(N__35324),
            .I(N__35301));
    InMux I__7219 (
            .O(N__35323),
            .I(N__35298));
    LocalMux I__7218 (
            .O(N__35320),
            .I(N__35291));
    LocalMux I__7217 (
            .O(N__35317),
            .I(N__35291));
    InMux I__7216 (
            .O(N__35314),
            .I(N__35286));
    InMux I__7215 (
            .O(N__35313),
            .I(N__35286));
    InMux I__7214 (
            .O(N__35312),
            .I(N__35283));
    InMux I__7213 (
            .O(N__35311),
            .I(N__35280));
    InMux I__7212 (
            .O(N__35310),
            .I(N__35277));
    Span4Mux_h I__7211 (
            .O(N__35307),
            .I(N__35272));
    Span4Mux_h I__7210 (
            .O(N__35304),
            .I(N__35272));
    Span4Mux_h I__7209 (
            .O(N__35301),
            .I(N__35269));
    LocalMux I__7208 (
            .O(N__35298),
            .I(N__35266));
    InMux I__7207 (
            .O(N__35297),
            .I(N__35263));
    InMux I__7206 (
            .O(N__35296),
            .I(N__35260));
    Span4Mux_h I__7205 (
            .O(N__35291),
            .I(N__35249));
    LocalMux I__7204 (
            .O(N__35286),
            .I(N__35249));
    LocalMux I__7203 (
            .O(N__35283),
            .I(N__35249));
    LocalMux I__7202 (
            .O(N__35280),
            .I(N__35249));
    LocalMux I__7201 (
            .O(N__35277),
            .I(N__35249));
    Odrv4 I__7200 (
            .O(N__35272),
            .I(\u1.DMA_control.readDfw_9 ));
    Odrv4 I__7199 (
            .O(N__35269),
            .I(\u1.DMA_control.readDfw_9 ));
    Odrv4 I__7198 (
            .O(N__35266),
            .I(\u1.DMA_control.readDfw_9 ));
    LocalMux I__7197 (
            .O(N__35263),
            .I(\u1.DMA_control.readDfw_9 ));
    LocalMux I__7196 (
            .O(N__35260),
            .I(\u1.DMA_control.readDfw_9 ));
    Odrv4 I__7195 (
            .O(N__35249),
            .I(\u1.DMA_control.readDfw_9 ));
    InMux I__7194 (
            .O(N__35236),
            .I(N__35233));
    LocalMux I__7193 (
            .O(N__35233),
            .I(N__35230));
    Odrv4 I__7192 (
            .O(N__35230),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_25 ));
    InMux I__7191 (
            .O(N__35227),
            .I(N__35224));
    LocalMux I__7190 (
            .O(N__35224),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_0 ));
    InMux I__7189 (
            .O(N__35221),
            .I(N__35218));
    LocalMux I__7188 (
            .O(N__35218),
            .I(N__35215));
    Span4Mux_v I__7187 (
            .O(N__35215),
            .I(N__35212));
    Sp12to4 I__7186 (
            .O(N__35212),
            .I(N__35209));
    Odrv12 I__7185 (
            .O(N__35209),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI2R0RZ0Z_24 ));
    InMux I__7184 (
            .O(N__35206),
            .I(N__35203));
    LocalMux I__7183 (
            .O(N__35203),
            .I(N__35200));
    Span4Mux_v I__7182 (
            .O(N__35200),
            .I(N__35197));
    Span4Mux_v I__7181 (
            .O(N__35197),
            .I(N__35194));
    Odrv4 I__7180 (
            .O(N__35194),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI6F9KZ0Z_24 ));
    InMux I__7179 (
            .O(N__35191),
            .I(N__35188));
    LocalMux I__7178 (
            .O(N__35188),
            .I(N__35185));
    Span4Mux_v I__7177 (
            .O(N__35185),
            .I(N__35182));
    Odrv4 I__7176 (
            .O(N__35182),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_24 ));
    CascadeMux I__7175 (
            .O(N__35179),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIA3ITZ0Z_24_cascade_ ));
    InMux I__7174 (
            .O(N__35176),
            .I(N__35173));
    LocalMux I__7173 (
            .O(N__35173),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_24 ));
    InMux I__7172 (
            .O(N__35170),
            .I(N__35167));
    LocalMux I__7171 (
            .O(N__35167),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIQKHM1Z0Z_2 ));
    CascadeMux I__7170 (
            .O(N__35164),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIA2E71Z0Z_24_cascade_ ));
    InMux I__7169 (
            .O(N__35161),
            .I(N__35158));
    LocalMux I__7168 (
            .O(N__35158),
            .I(N__35154));
    InMux I__7167 (
            .O(N__35157),
            .I(N__35151));
    Odrv4 I__7166 (
            .O(N__35154),
            .I(DMA_dev0_Tm_5));
    LocalMux I__7165 (
            .O(N__35151),
            .I(DMA_dev0_Tm_5));
    CascadeMux I__7164 (
            .O(N__35146),
            .I(N__35143));
    InMux I__7163 (
            .O(N__35143),
            .I(N__35139));
    InMux I__7162 (
            .O(N__35142),
            .I(N__35136));
    LocalMux I__7161 (
            .O(N__35139),
            .I(N__35133));
    LocalMux I__7160 (
            .O(N__35136),
            .I(N__35130));
    Span4Mux_v I__7159 (
            .O(N__35133),
            .I(N__35127));
    Span4Mux_h I__7158 (
            .O(N__35130),
            .I(N__35124));
    Odrv4 I__7157 (
            .O(N__35127),
            .I(PIO_cmdport_T4_2));
    Odrv4 I__7156 (
            .O(N__35124),
            .I(PIO_cmdport_T4_2));
    InMux I__7155 (
            .O(N__35119),
            .I(N__35116));
    LocalMux I__7154 (
            .O(N__35116),
            .I(N__35113));
    Span4Mux_v I__7153 (
            .O(N__35113),
            .I(N__35110));
    Span4Mux_h I__7152 (
            .O(N__35110),
            .I(N__35107));
    Odrv4 I__7151 (
            .O(N__35107),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIG7GTZ0Z_18 ));
    InMux I__7150 (
            .O(N__35104),
            .I(N__35101));
    LocalMux I__7149 (
            .O(N__35101),
            .I(N__35098));
    Span4Mux_v I__7148 (
            .O(N__35098),
            .I(N__35095));
    Odrv4 I__7147 (
            .O(N__35095),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_18 ));
    CascadeMux I__7146 (
            .O(N__35092),
            .I(mem_mem_ram6__RNIJ8B71_18_cascade_));
    InMux I__7145 (
            .O(N__35089),
            .I(N__35086));
    LocalMux I__7144 (
            .O(N__35086),
            .I(N__35083));
    Span12Mux_h I__7143 (
            .O(N__35083),
            .I(N__35080));
    Odrv12 I__7142 (
            .O(N__35080),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_18 ));
    InMux I__7141 (
            .O(N__35077),
            .I(N__35074));
    LocalMux I__7140 (
            .O(N__35074),
            .I(N__35071));
    Span4Mux_h I__7139 (
            .O(N__35071),
            .I(N__35068));
    Odrv4 I__7138 (
            .O(N__35068),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_18 ));
    InMux I__7137 (
            .O(N__35065),
            .I(N__35062));
    LocalMux I__7136 (
            .O(N__35062),
            .I(N__35059));
    Span4Mux_v I__7135 (
            .O(N__35059),
            .I(N__35056));
    Odrv4 I__7134 (
            .O(N__35056),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNICJ7KZ0Z_18 ));
    CascadeMux I__7133 (
            .O(N__35053),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI8VUQZ0Z_18_cascade_ ));
    InMux I__7132 (
            .O(N__35050),
            .I(N__35047));
    LocalMux I__7131 (
            .O(N__35047),
            .I(iQ_RNI6TDM1_2));
    InMux I__7130 (
            .O(N__35044),
            .I(N__35040));
    InMux I__7129 (
            .O(N__35043),
            .I(N__35037));
    LocalMux I__7128 (
            .O(N__35040),
            .I(N__35033));
    LocalMux I__7127 (
            .O(N__35037),
            .I(N__35030));
    InMux I__7126 (
            .O(N__35036),
            .I(N__35027));
    Span4Mux_v I__7125 (
            .O(N__35033),
            .I(N__35022));
    Span4Mux_v I__7124 (
            .O(N__35030),
            .I(N__35022));
    LocalMux I__7123 (
            .O(N__35027),
            .I(N__35017));
    Span4Mux_h I__7122 (
            .O(N__35022),
            .I(N__35014));
    InMux I__7121 (
            .O(N__35021),
            .I(N__35011));
    InMux I__7120 (
            .O(N__35020),
            .I(N__35008));
    Span4Mux_v I__7119 (
            .O(N__35017),
            .I(N__35005));
    Span4Mux_h I__7118 (
            .O(N__35014),
            .I(N__35002));
    LocalMux I__7117 (
            .O(N__35011),
            .I(N__34999));
    LocalMux I__7116 (
            .O(N__35008),
            .I(N__34996));
    Sp12to4 I__7115 (
            .O(N__35005),
            .I(N__34989));
    Sp12to4 I__7114 (
            .O(N__35002),
            .I(N__34989));
    Span12Mux_v I__7113 (
            .O(N__34999),
            .I(N__34989));
    Span12Mux_s10_v I__7112 (
            .O(N__34996),
            .I(N__34986));
    Odrv12 I__7111 (
            .O(N__34989),
            .I(wb_dat_i_c_18));
    Odrv12 I__7110 (
            .O(N__34986),
            .I(wb_dat_i_c_18));
    InMux I__7109 (
            .O(N__34981),
            .I(N__34978));
    LocalMux I__7108 (
            .O(N__34978),
            .I(\u0.CtrlRegZ0Z_18 ));
    CascadeMux I__7107 (
            .O(N__34975),
            .I(N__34972));
    InMux I__7106 (
            .O(N__34972),
            .I(N__34968));
    InMux I__7105 (
            .O(N__34971),
            .I(N__34965));
    LocalMux I__7104 (
            .O(N__34968),
            .I(N__34962));
    LocalMux I__7103 (
            .O(N__34965),
            .I(N__34959));
    Span4Mux_v I__7102 (
            .O(N__34962),
            .I(N__34956));
    Odrv12 I__7101 (
            .O(N__34959),
            .I(PIO_dport1_T1_3));
    Odrv4 I__7100 (
            .O(N__34956),
            .I(PIO_dport1_T1_3));
    InMux I__7099 (
            .O(N__34951),
            .I(N__34948));
    LocalMux I__7098 (
            .O(N__34948),
            .I(N__34945));
    Span4Mux_v I__7097 (
            .O(N__34945),
            .I(N__34942));
    Odrv4 I__7096 (
            .O(N__34942),
            .I(\u0.dat_o_0_0_2_3 ));
    InMux I__7095 (
            .O(N__34939),
            .I(N__34936));
    LocalMux I__7094 (
            .O(N__34936),
            .I(\u0.dat_o_0_0_3_3 ));
    CascadeMux I__7093 (
            .O(N__34933),
            .I(\u0.dat_o_0_0_0_3_cascade_ ));
    InMux I__7092 (
            .O(N__34930),
            .I(N__34927));
    LocalMux I__7091 (
            .O(N__34927),
            .I(\u0.dat_o_0_0_1Z0Z_3 ));
    IoInMux I__7090 (
            .O(N__34924),
            .I(N__34921));
    LocalMux I__7089 (
            .O(N__34921),
            .I(N__34918));
    Span12Mux_s6_h I__7088 (
            .O(N__34918),
            .I(N__34915));
    Odrv12 I__7087 (
            .O(N__34915),
            .I(wb_dat_o_c_3));
    InMux I__7086 (
            .O(N__34912),
            .I(N__34905));
    InMux I__7085 (
            .O(N__34911),
            .I(N__34905));
    InMux I__7084 (
            .O(N__34910),
            .I(N__34902));
    LocalMux I__7083 (
            .O(N__34905),
            .I(N__34899));
    LocalMux I__7082 (
            .O(N__34902),
            .I(N__34896));
    Span4Mux_v I__7081 (
            .O(N__34899),
            .I(N__34893));
    Span4Mux_v I__7080 (
            .O(N__34896),
            .I(N__34890));
    Span4Mux_v I__7079 (
            .O(N__34893),
            .I(N__34887));
    Span4Mux_h I__7078 (
            .O(N__34890),
            .I(N__34884));
    Sp12to4 I__7077 (
            .O(N__34887),
            .I(N__34879));
    Sp12to4 I__7076 (
            .O(N__34884),
            .I(N__34879));
    Odrv12 I__7075 (
            .O(N__34879),
            .I(dd_pad_i_c_3));
    InMux I__7074 (
            .O(N__34876),
            .I(N__34873));
    LocalMux I__7073 (
            .O(N__34873),
            .I(PIOq_3));
    InMux I__7072 (
            .O(N__34870),
            .I(N__34867));
    LocalMux I__7071 (
            .O(N__34867),
            .I(N__34864));
    Span4Mux_h I__7070 (
            .O(N__34864),
            .I(N__34861));
    Odrv4 I__7069 (
            .O(N__34861),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_3 ));
    CascadeMux I__7068 (
            .O(N__34858),
            .I(N__34855));
    InMux I__7067 (
            .O(N__34855),
            .I(N__34852));
    LocalMux I__7066 (
            .O(N__34852),
            .I(N__34849));
    Span4Mux_v I__7065 (
            .O(N__34849),
            .I(N__34846));
    Sp12to4 I__7064 (
            .O(N__34846),
            .I(N__34843));
    Odrv12 I__7063 (
            .O(N__34843),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNI43TNZ0Z_3 ));
    InMux I__7062 (
            .O(N__34840),
            .I(N__34837));
    LocalMux I__7061 (
            .O(N__34837),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIHGOD1Z0Z_3 ));
    InMux I__7060 (
            .O(N__34834),
            .I(N__34830));
    InMux I__7059 (
            .O(N__34833),
            .I(N__34827));
    LocalMux I__7058 (
            .O(N__34830),
            .I(DMA_dev0_Tm_3));
    LocalMux I__7057 (
            .O(N__34827),
            .I(DMA_dev0_Tm_3));
    CascadeMux I__7056 (
            .O(N__34822),
            .I(N__34819));
    InMux I__7055 (
            .O(N__34819),
            .I(N__34816));
    LocalMux I__7054 (
            .O(N__34816),
            .I(N__34812));
    InMux I__7053 (
            .O(N__34815),
            .I(N__34809));
    Odrv4 I__7052 (
            .O(N__34812),
            .I(DMA_dev0_Tm_4));
    LocalMux I__7051 (
            .O(N__34809),
            .I(DMA_dev0_Tm_4));
    InMux I__7050 (
            .O(N__34804),
            .I(N__34800));
    InMux I__7049 (
            .O(N__34803),
            .I(N__34797));
    LocalMux I__7048 (
            .O(N__34800),
            .I(N__34792));
    LocalMux I__7047 (
            .O(N__34797),
            .I(N__34792));
    Span4Mux_v I__7046 (
            .O(N__34792),
            .I(N__34789));
    Span4Mux_h I__7045 (
            .O(N__34789),
            .I(N__34784));
    InMux I__7044 (
            .O(N__34788),
            .I(N__34781));
    InMux I__7043 (
            .O(N__34787),
            .I(N__34777));
    Span4Mux_h I__7042 (
            .O(N__34784),
            .I(N__34772));
    LocalMux I__7041 (
            .O(N__34781),
            .I(N__34772));
    InMux I__7040 (
            .O(N__34780),
            .I(N__34769));
    LocalMux I__7039 (
            .O(N__34777),
            .I(N__34766));
    Span4Mux_v I__7038 (
            .O(N__34772),
            .I(N__34761));
    LocalMux I__7037 (
            .O(N__34769),
            .I(N__34761));
    Span12Mux_v I__7036 (
            .O(N__34766),
            .I(N__34758));
    Span4Mux_h I__7035 (
            .O(N__34761),
            .I(N__34755));
    Span12Mux_h I__7034 (
            .O(N__34758),
            .I(N__34752));
    Span4Mux_v I__7033 (
            .O(N__34755),
            .I(N__34749));
    Odrv12 I__7032 (
            .O(N__34752),
            .I(wb_dat_i_c_20));
    Odrv4 I__7031 (
            .O(N__34749),
            .I(wb_dat_i_c_20));
    InMux I__7030 (
            .O(N__34744),
            .I(N__34741));
    LocalMux I__7029 (
            .O(N__34741),
            .I(N__34738));
    Span4Mux_v I__7028 (
            .O(N__34738),
            .I(N__34735));
    Odrv4 I__7027 (
            .O(N__34735),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIS2CMZ0Z_3 ));
    InMux I__7026 (
            .O(N__34732),
            .I(N__34729));
    LocalMux I__7025 (
            .O(N__34729),
            .I(N__34726));
    Span4Mux_h I__7024 (
            .O(N__34726),
            .I(N__34723));
    Span4Mux_h I__7023 (
            .O(N__34723),
            .I(N__34720));
    Span4Mux_v I__7022 (
            .O(N__34720),
            .I(N__34717));
    Odrv4 I__7021 (
            .O(N__34717),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI0J4NZ0Z_3 ));
    CascadeMux I__7020 (
            .O(N__34714),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIE0OK1Z0Z_2_cascade_ ));
    CascadeMux I__7019 (
            .O(N__34711),
            .I(DMAq_3_cascade_));
    InMux I__7018 (
            .O(N__34708),
            .I(N__34705));
    LocalMux I__7017 (
            .O(N__34705),
            .I(N__34700));
    InMux I__7016 (
            .O(N__34704),
            .I(N__34695));
    InMux I__7015 (
            .O(N__34703),
            .I(N__34692));
    Span4Mux_v I__7014 (
            .O(N__34700),
            .I(N__34689));
    InMux I__7013 (
            .O(N__34699),
            .I(N__34684));
    InMux I__7012 (
            .O(N__34698),
            .I(N__34681));
    LocalMux I__7011 (
            .O(N__34695),
            .I(N__34676));
    LocalMux I__7010 (
            .O(N__34692),
            .I(N__34676));
    Span4Mux_h I__7009 (
            .O(N__34689),
            .I(N__34673));
    InMux I__7008 (
            .O(N__34688),
            .I(N__34670));
    InMux I__7007 (
            .O(N__34687),
            .I(N__34667));
    LocalMux I__7006 (
            .O(N__34684),
            .I(N__34663));
    LocalMux I__7005 (
            .O(N__34681),
            .I(N__34658));
    Span4Mux_v I__7004 (
            .O(N__34676),
            .I(N__34658));
    Span4Mux_h I__7003 (
            .O(N__34673),
            .I(N__34653));
    LocalMux I__7002 (
            .O(N__34670),
            .I(N__34653));
    LocalMux I__7001 (
            .O(N__34667),
            .I(N__34650));
    InMux I__7000 (
            .O(N__34666),
            .I(N__34647));
    Sp12to4 I__6999 (
            .O(N__34663),
            .I(N__34643));
    Span4Mux_v I__6998 (
            .O(N__34658),
            .I(N__34640));
    Span4Mux_v I__6997 (
            .O(N__34653),
            .I(N__34637));
    Span4Mux_v I__6996 (
            .O(N__34650),
            .I(N__34632));
    LocalMux I__6995 (
            .O(N__34647),
            .I(N__34632));
    InMux I__6994 (
            .O(N__34646),
            .I(N__34629));
    Span12Mux_v I__6993 (
            .O(N__34643),
            .I(N__34624));
    Sp12to4 I__6992 (
            .O(N__34640),
            .I(N__34624));
    Span4Mux_v I__6991 (
            .O(N__34637),
            .I(N__34621));
    Sp12to4 I__6990 (
            .O(N__34632),
            .I(N__34616));
    LocalMux I__6989 (
            .O(N__34629),
            .I(N__34616));
    Span12Mux_h I__6988 (
            .O(N__34624),
            .I(N__34613));
    Sp12to4 I__6987 (
            .O(N__34621),
            .I(N__34608));
    Span12Mux_v I__6986 (
            .O(N__34616),
            .I(N__34608));
    Span12Mux_h I__6985 (
            .O(N__34613),
            .I(N__34605));
    Span12Mux_h I__6984 (
            .O(N__34608),
            .I(N__34602));
    Odrv12 I__6983 (
            .O(N__34605),
            .I(wb_dat_i_c_13));
    Odrv12 I__6982 (
            .O(N__34602),
            .I(wb_dat_i_c_13));
    CascadeMux I__6981 (
            .O(N__34597),
            .I(N__34594));
    InMux I__6980 (
            .O(N__34594),
            .I(N__34591));
    LocalMux I__6979 (
            .O(N__34591),
            .I(N__34588));
    Span4Mux_v I__6978 (
            .O(N__34588),
            .I(N__34584));
    InMux I__6977 (
            .O(N__34587),
            .I(N__34581));
    Span4Mux_h I__6976 (
            .O(N__34584),
            .I(N__34576));
    LocalMux I__6975 (
            .O(N__34581),
            .I(N__34576));
    Span4Mux_h I__6974 (
            .O(N__34576),
            .I(N__34573));
    Odrv4 I__6973 (
            .O(N__34573),
            .I(PIO_dport0_T2_5));
    InMux I__6972 (
            .O(N__34570),
            .I(N__34565));
    InMux I__6971 (
            .O(N__34569),
            .I(N__34562));
    InMux I__6970 (
            .O(N__34568),
            .I(N__34559));
    LocalMux I__6969 (
            .O(N__34565),
            .I(N__34554));
    LocalMux I__6968 (
            .O(N__34562),
            .I(N__34554));
    LocalMux I__6967 (
            .O(N__34559),
            .I(N__34551));
    Span4Mux_v I__6966 (
            .O(N__34554),
            .I(N__34546));
    Span4Mux_v I__6965 (
            .O(N__34551),
            .I(N__34543));
    InMux I__6964 (
            .O(N__34550),
            .I(N__34538));
    InMux I__6963 (
            .O(N__34549),
            .I(N__34535));
    Span4Mux_v I__6962 (
            .O(N__34546),
            .I(N__34530));
    Span4Mux_h I__6961 (
            .O(N__34543),
            .I(N__34530));
    InMux I__6960 (
            .O(N__34542),
            .I(N__34527));
    InMux I__6959 (
            .O(N__34541),
            .I(N__34524));
    LocalMux I__6958 (
            .O(N__34538),
            .I(N__34519));
    LocalMux I__6957 (
            .O(N__34535),
            .I(N__34516));
    Span4Mux_h I__6956 (
            .O(N__34530),
            .I(N__34513));
    LocalMux I__6955 (
            .O(N__34527),
            .I(N__34508));
    LocalMux I__6954 (
            .O(N__34524),
            .I(N__34508));
    InMux I__6953 (
            .O(N__34523),
            .I(N__34505));
    InMux I__6952 (
            .O(N__34522),
            .I(N__34502));
    Sp12to4 I__6951 (
            .O(N__34519),
            .I(N__34497));
    Sp12to4 I__6950 (
            .O(N__34516),
            .I(N__34497));
    Span4Mux_h I__6949 (
            .O(N__34513),
            .I(N__34492));
    Span4Mux_v I__6948 (
            .O(N__34508),
            .I(N__34492));
    LocalMux I__6947 (
            .O(N__34505),
            .I(N__34489));
    LocalMux I__6946 (
            .O(N__34502),
            .I(N__34486));
    Span12Mux_v I__6945 (
            .O(N__34497),
            .I(N__34483));
    Span4Mux_v I__6944 (
            .O(N__34492),
            .I(N__34480));
    Span12Mux_v I__6943 (
            .O(N__34489),
            .I(N__34477));
    Span4Mux_v I__6942 (
            .O(N__34486),
            .I(N__34474));
    Span12Mux_h I__6941 (
            .O(N__34483),
            .I(N__34471));
    Sp12to4 I__6940 (
            .O(N__34480),
            .I(N__34468));
    Span12Mux_h I__6939 (
            .O(N__34477),
            .I(N__34463));
    Sp12to4 I__6938 (
            .O(N__34474),
            .I(N__34463));
    Span12Mux_h I__6937 (
            .O(N__34471),
            .I(N__34460));
    Span12Mux_h I__6936 (
            .O(N__34468),
            .I(N__34457));
    Span12Mux_h I__6935 (
            .O(N__34463),
            .I(N__34454));
    Odrv12 I__6934 (
            .O(N__34460),
            .I(wb_dat_i_c_15));
    Odrv12 I__6933 (
            .O(N__34457),
            .I(wb_dat_i_c_15));
    Odrv12 I__6932 (
            .O(N__34454),
            .I(wb_dat_i_c_15));
    CascadeMux I__6931 (
            .O(N__34447),
            .I(N__34444));
    InMux I__6930 (
            .O(N__34444),
            .I(N__34441));
    LocalMux I__6929 (
            .O(N__34441),
            .I(N__34437));
    InMux I__6928 (
            .O(N__34440),
            .I(N__34434));
    Span4Mux_h I__6927 (
            .O(N__34437),
            .I(N__34431));
    LocalMux I__6926 (
            .O(N__34434),
            .I(PIO_dport1_T4_3));
    Odrv4 I__6925 (
            .O(N__34431),
            .I(PIO_dport1_T4_3));
    InMux I__6924 (
            .O(N__34426),
            .I(N__34423));
    LocalMux I__6923 (
            .O(N__34423),
            .I(N__34420));
    Span4Mux_v I__6922 (
            .O(N__34420),
            .I(N__34417));
    Span4Mux_h I__6921 (
            .O(N__34417),
            .I(N__34414));
    Odrv4 I__6920 (
            .O(N__34414),
            .I(\u0.dat_o_i_0_0_19 ));
    InMux I__6919 (
            .O(N__34411),
            .I(N__34408));
    LocalMux I__6918 (
            .O(N__34408),
            .I(N__34405));
    Span4Mux_h I__6917 (
            .O(N__34405),
            .I(N__34402));
    Odrv4 I__6916 (
            .O(N__34402),
            .I(\u0.dat_o_0_0_3_4 ));
    InMux I__6915 (
            .O(N__34399),
            .I(N__34395));
    InMux I__6914 (
            .O(N__34398),
            .I(N__34392));
    LocalMux I__6913 (
            .O(N__34395),
            .I(N__34389));
    LocalMux I__6912 (
            .O(N__34392),
            .I(PIO_dport0_T2_7));
    Odrv4 I__6911 (
            .O(N__34389),
            .I(PIO_dport0_T2_7));
    InMux I__6910 (
            .O(N__34384),
            .I(N__34381));
    LocalMux I__6909 (
            .O(N__34381),
            .I(N__34378));
    Span4Mux_v I__6908 (
            .O(N__34378),
            .I(N__34375));
    Span4Mux_h I__6907 (
            .O(N__34375),
            .I(N__34372));
    Odrv4 I__6906 (
            .O(N__34372),
            .I(\u0.N_2033 ));
    InMux I__6905 (
            .O(N__34369),
            .I(N__34365));
    InMux I__6904 (
            .O(N__34368),
            .I(N__34362));
    LocalMux I__6903 (
            .O(N__34365),
            .I(N__34359));
    LocalMux I__6902 (
            .O(N__34362),
            .I(N__34355));
    Span4Mux_v I__6901 (
            .O(N__34359),
            .I(N__34352));
    InMux I__6900 (
            .O(N__34358),
            .I(N__34349));
    Span4Mux_v I__6899 (
            .O(N__34355),
            .I(N__34346));
    Span4Mux_h I__6898 (
            .O(N__34352),
            .I(N__34341));
    LocalMux I__6897 (
            .O(N__34349),
            .I(N__34341));
    Span4Mux_v I__6896 (
            .O(N__34346),
            .I(N__34338));
    Span4Mux_v I__6895 (
            .O(N__34341),
            .I(N__34334));
    Span4Mux_v I__6894 (
            .O(N__34338),
            .I(N__34330));
    InMux I__6893 (
            .O(N__34337),
            .I(N__34327));
    Span4Mux_v I__6892 (
            .O(N__34334),
            .I(N__34324));
    InMux I__6891 (
            .O(N__34333),
            .I(N__34321));
    Span4Mux_h I__6890 (
            .O(N__34330),
            .I(N__34318));
    LocalMux I__6889 (
            .O(N__34327),
            .I(N__34315));
    Span4Mux_h I__6888 (
            .O(N__34324),
            .I(N__34312));
    LocalMux I__6887 (
            .O(N__34321),
            .I(N__34309));
    Sp12to4 I__6886 (
            .O(N__34318),
            .I(N__34304));
    Span12Mux_v I__6885 (
            .O(N__34315),
            .I(N__34304));
    Sp12to4 I__6884 (
            .O(N__34312),
            .I(N__34299));
    Span12Mux_v I__6883 (
            .O(N__34309),
            .I(N__34299));
    Odrv12 I__6882 (
            .O(N__34304),
            .I(wb_dat_i_c_19));
    Odrv12 I__6881 (
            .O(N__34299),
            .I(wb_dat_i_c_19));
    InMux I__6880 (
            .O(N__34294),
            .I(N__34291));
    LocalMux I__6879 (
            .O(N__34291),
            .I(N__34287));
    InMux I__6878 (
            .O(N__34290),
            .I(N__34284));
    Span4Mux_h I__6877 (
            .O(N__34287),
            .I(N__34281));
    LocalMux I__6876 (
            .O(N__34284),
            .I(PIO_dport0_T4_3));
    Odrv4 I__6875 (
            .O(N__34281),
            .I(PIO_dport0_T4_3));
    InMux I__6874 (
            .O(N__34276),
            .I(N__34273));
    LocalMux I__6873 (
            .O(N__34273),
            .I(N__34268));
    InMux I__6872 (
            .O(N__34272),
            .I(N__34265));
    InMux I__6871 (
            .O(N__34271),
            .I(N__34261));
    Span4Mux_v I__6870 (
            .O(N__34268),
            .I(N__34258));
    LocalMux I__6869 (
            .O(N__34265),
            .I(N__34255));
    InMux I__6868 (
            .O(N__34264),
            .I(N__34252));
    LocalMux I__6867 (
            .O(N__34261),
            .I(N__34249));
    Span4Mux_h I__6866 (
            .O(N__34258),
            .I(N__34244));
    Span4Mux_v I__6865 (
            .O(N__34255),
            .I(N__34244));
    LocalMux I__6864 (
            .O(N__34252),
            .I(N__34238));
    Sp12to4 I__6863 (
            .O(N__34249),
            .I(N__34233));
    Span4Mux_v I__6862 (
            .O(N__34244),
            .I(N__34230));
    InMux I__6861 (
            .O(N__34243),
            .I(N__34227));
    InMux I__6860 (
            .O(N__34242),
            .I(N__34224));
    InMux I__6859 (
            .O(N__34241),
            .I(N__34221));
    Sp12to4 I__6858 (
            .O(N__34238),
            .I(N__34218));
    InMux I__6857 (
            .O(N__34237),
            .I(N__34215));
    InMux I__6856 (
            .O(N__34236),
            .I(N__34212));
    Span12Mux_v I__6855 (
            .O(N__34233),
            .I(N__34209));
    Sp12to4 I__6854 (
            .O(N__34230),
            .I(N__34204));
    LocalMux I__6853 (
            .O(N__34227),
            .I(N__34204));
    LocalMux I__6852 (
            .O(N__34224),
            .I(N__34201));
    LocalMux I__6851 (
            .O(N__34221),
            .I(N__34198));
    Span12Mux_v I__6850 (
            .O(N__34218),
            .I(N__34195));
    LocalMux I__6849 (
            .O(N__34215),
            .I(N__34192));
    LocalMux I__6848 (
            .O(N__34212),
            .I(N__34189));
    Span12Mux_v I__6847 (
            .O(N__34209),
            .I(N__34186));
    Span12Mux_h I__6846 (
            .O(N__34204),
            .I(N__34183));
    Span12Mux_v I__6845 (
            .O(N__34201),
            .I(N__34178));
    Sp12to4 I__6844 (
            .O(N__34198),
            .I(N__34178));
    Span12Mux_v I__6843 (
            .O(N__34195),
            .I(N__34175));
    Span12Mux_v I__6842 (
            .O(N__34192),
            .I(N__34170));
    Sp12to4 I__6841 (
            .O(N__34189),
            .I(N__34170));
    Span12Mux_h I__6840 (
            .O(N__34186),
            .I(N__34165));
    Span12Mux_v I__6839 (
            .O(N__34183),
            .I(N__34165));
    Span12Mux_v I__6838 (
            .O(N__34178),
            .I(N__34162));
    Span12Mux_h I__6837 (
            .O(N__34175),
            .I(N__34157));
    Span12Mux_v I__6836 (
            .O(N__34170),
            .I(N__34157));
    Span12Mux_h I__6835 (
            .O(N__34165),
            .I(N__34154));
    Span12Mux_h I__6834 (
            .O(N__34162),
            .I(N__34151));
    Span12Mux_h I__6833 (
            .O(N__34157),
            .I(N__34148));
    Odrv12 I__6832 (
            .O(N__34154),
            .I(wb_dat_i_c_2));
    Odrv12 I__6831 (
            .O(N__34151),
            .I(wb_dat_i_c_2));
    Odrv12 I__6830 (
            .O(N__34148),
            .I(wb_dat_i_c_2));
    CascadeMux I__6829 (
            .O(N__34141),
            .I(N__34138));
    InMux I__6828 (
            .O(N__34138),
            .I(N__34134));
    InMux I__6827 (
            .O(N__34137),
            .I(N__34131));
    LocalMux I__6826 (
            .O(N__34134),
            .I(N__34128));
    LocalMux I__6825 (
            .O(N__34131),
            .I(N__34125));
    Span4Mux_v I__6824 (
            .O(N__34128),
            .I(N__34122));
    Span4Mux_v I__6823 (
            .O(N__34125),
            .I(N__34119));
    Span4Mux_h I__6822 (
            .O(N__34122),
            .I(N__34116));
    Odrv4 I__6821 (
            .O(N__34119),
            .I(PIO_dport1_T1_2));
    Odrv4 I__6820 (
            .O(N__34116),
            .I(PIO_dport1_T1_2));
    InMux I__6819 (
            .O(N__34111),
            .I(N__34108));
    LocalMux I__6818 (
            .O(N__34108),
            .I(N__34105));
    Span4Mux_s3_v I__6817 (
            .O(N__34105),
            .I(N__34102));
    Odrv4 I__6816 (
            .O(N__34102),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_13 ));
    CascadeMux I__6815 (
            .O(N__34099),
            .I(N__34096));
    InMux I__6814 (
            .O(N__34096),
            .I(N__34093));
    LocalMux I__6813 (
            .O(N__34093),
            .I(N__34090));
    Span4Mux_s2_v I__6812 (
            .O(N__34090),
            .I(N__34087));
    Odrv4 I__6811 (
            .O(N__34087),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_13 ));
    CascadeMux I__6810 (
            .O(N__34084),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI297KZ0Z_13_cascade_ ));
    InMux I__6809 (
            .O(N__34081),
            .I(N__34078));
    LocalMux I__6808 (
            .O(N__34078),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNII8DM1Z0Z_2 ));
    InMux I__6807 (
            .O(N__34075),
            .I(N__34072));
    LocalMux I__6806 (
            .O(N__34072),
            .I(DMAq_13));
    InMux I__6805 (
            .O(N__34069),
            .I(N__34066));
    LocalMux I__6804 (
            .O(N__34066),
            .I(N__34063));
    Span4Mux_s1_v I__6803 (
            .O(N__34063),
            .I(N__34060));
    Odrv4 I__6802 (
            .O(N__34060),
            .I(\u0.dat_o_0_0_1Z0Z_13 ));
    InMux I__6801 (
            .O(N__34057),
            .I(N__34054));
    LocalMux I__6800 (
            .O(N__34054),
            .I(N__34051));
    Odrv12 I__6799 (
            .O(N__34051),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_13 ));
    InMux I__6798 (
            .O(N__34048),
            .I(N__34045));
    LocalMux I__6797 (
            .O(N__34045),
            .I(N__34042));
    Span4Mux_v I__6796 (
            .O(N__34042),
            .I(N__34039));
    Odrv4 I__6795 (
            .O(N__34039),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_13 ));
    InMux I__6794 (
            .O(N__34036),
            .I(N__34033));
    LocalMux I__6793 (
            .O(N__34033),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIUKUQZ0Z_13 ));
    InMux I__6792 (
            .O(N__34030),
            .I(N__34027));
    LocalMux I__6791 (
            .O(N__34027),
            .I(N__34022));
    InMux I__6790 (
            .O(N__34026),
            .I(N__34017));
    InMux I__6789 (
            .O(N__34025),
            .I(N__34017));
    Span4Mux_s2_v I__6788 (
            .O(N__34022),
            .I(N__34014));
    LocalMux I__6787 (
            .O(N__34017),
            .I(N__34011));
    Sp12to4 I__6786 (
            .O(N__34014),
            .I(N__34008));
    Span4Mux_v I__6785 (
            .O(N__34011),
            .I(N__34005));
    Span12Mux_h I__6784 (
            .O(N__34008),
            .I(N__34002));
    Span4Mux_v I__6783 (
            .O(N__34005),
            .I(N__33999));
    Span12Mux_v I__6782 (
            .O(N__34002),
            .I(N__33994));
    Sp12to4 I__6781 (
            .O(N__33999),
            .I(N__33994));
    Odrv12 I__6780 (
            .O(N__33994),
            .I(dd_pad_i_c_13));
    InMux I__6779 (
            .O(N__33991),
            .I(N__33988));
    LocalMux I__6778 (
            .O(N__33988),
            .I(PIOq_13));
    CascadeMux I__6777 (
            .O(N__33985),
            .I(N__33982));
    InMux I__6776 (
            .O(N__33982),
            .I(N__33978));
    InMux I__6775 (
            .O(N__33981),
            .I(N__33975));
    LocalMux I__6774 (
            .O(N__33978),
            .I(N__33972));
    LocalMux I__6773 (
            .O(N__33975),
            .I(N__33969));
    Span4Mux_v I__6772 (
            .O(N__33972),
            .I(N__33964));
    Span4Mux_h I__6771 (
            .O(N__33969),
            .I(N__33964));
    Odrv4 I__6770 (
            .O(N__33964),
            .I(PIO_cmdport_T2_1));
    CascadeMux I__6769 (
            .O(N__33961),
            .I(N__33957));
    InMux I__6768 (
            .O(N__33960),
            .I(N__33954));
    InMux I__6767 (
            .O(N__33957),
            .I(N__33951));
    LocalMux I__6766 (
            .O(N__33954),
            .I(N__33948));
    LocalMux I__6765 (
            .O(N__33951),
            .I(N__33945));
    Span4Mux_h I__6764 (
            .O(N__33948),
            .I(N__33942));
    Odrv4 I__6763 (
            .O(N__33945),
            .I(PIO_cmdport_T2_0));
    Odrv4 I__6762 (
            .O(N__33942),
            .I(PIO_cmdport_T2_0));
    InMux I__6761 (
            .O(N__33937),
            .I(N__33933));
    CascadeMux I__6760 (
            .O(N__33936),
            .I(N__33930));
    LocalMux I__6759 (
            .O(N__33933),
            .I(N__33927));
    InMux I__6758 (
            .O(N__33930),
            .I(N__33924));
    Span4Mux_h I__6757 (
            .O(N__33927),
            .I(N__33921));
    LocalMux I__6756 (
            .O(N__33924),
            .I(PIO_dport1_T2_0));
    Odrv4 I__6755 (
            .O(N__33921),
            .I(PIO_dport1_T2_0));
    InMux I__6754 (
            .O(N__33916),
            .I(N__33913));
    LocalMux I__6753 (
            .O(N__33913),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIOEUQZ0Z_10 ));
    CascadeMux I__6752 (
            .O(N__33910),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIS27KZ0Z_10_cascade_ ));
    InMux I__6751 (
            .O(N__33907),
            .I(N__33904));
    LocalMux I__6750 (
            .O(N__33904),
            .I(N__33901));
    Span4Mux_v I__6749 (
            .O(N__33901),
            .I(N__33898));
    Odrv4 I__6748 (
            .O(N__33898),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_10 ));
    InMux I__6747 (
            .O(N__33895),
            .I(N__33892));
    LocalMux I__6746 (
            .O(N__33892),
            .I(N__33889));
    Span4Mux_h I__6745 (
            .O(N__33889),
            .I(N__33886));
    Odrv4 I__6744 (
            .O(N__33886),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_10 ));
    CascadeMux I__6743 (
            .O(N__33883),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI0NFTZ0Z_10_cascade_ ));
    InMux I__6742 (
            .O(N__33880),
            .I(N__33877));
    LocalMux I__6741 (
            .O(N__33877),
            .I(iQ_RNI6SCM1_2));
    CascadeMux I__6740 (
            .O(N__33874),
            .I(mem_mem_ram6__RNIRFA71_10_cascade_));
    InMux I__6739 (
            .O(N__33871),
            .I(N__33868));
    LocalMux I__6738 (
            .O(N__33868),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_10 ));
    CascadeMux I__6737 (
            .O(N__33865),
            .I(N__33856));
    InMux I__6736 (
            .O(N__33864),
            .I(N__33850));
    InMux I__6735 (
            .O(N__33863),
            .I(N__33847));
    InMux I__6734 (
            .O(N__33862),
            .I(N__33842));
    InMux I__6733 (
            .O(N__33861),
            .I(N__33842));
    InMux I__6732 (
            .O(N__33860),
            .I(N__33837));
    InMux I__6731 (
            .O(N__33859),
            .I(N__33837));
    InMux I__6730 (
            .O(N__33856),
            .I(N__33832));
    InMux I__6729 (
            .O(N__33855),
            .I(N__33832));
    InMux I__6728 (
            .O(N__33854),
            .I(N__33825));
    InMux I__6727 (
            .O(N__33853),
            .I(N__33825));
    LocalMux I__6726 (
            .O(N__33850),
            .I(N__33821));
    LocalMux I__6725 (
            .O(N__33847),
            .I(N__33816));
    LocalMux I__6724 (
            .O(N__33842),
            .I(N__33816));
    LocalMux I__6723 (
            .O(N__33837),
            .I(N__33813));
    LocalMux I__6722 (
            .O(N__33832),
            .I(N__33810));
    InMux I__6721 (
            .O(N__33831),
            .I(N__33805));
    InMux I__6720 (
            .O(N__33830),
            .I(N__33805));
    LocalMux I__6719 (
            .O(N__33825),
            .I(N__33802));
    InMux I__6718 (
            .O(N__33824),
            .I(N__33797));
    Span4Mux_v I__6717 (
            .O(N__33821),
            .I(N__33792));
    Span4Mux_v I__6716 (
            .O(N__33816),
            .I(N__33792));
    Span4Mux_v I__6715 (
            .O(N__33813),
            .I(N__33787));
    Span4Mux_h I__6714 (
            .O(N__33810),
            .I(N__33787));
    LocalMux I__6713 (
            .O(N__33805),
            .I(N__33784));
    Span4Mux_h I__6712 (
            .O(N__33802),
            .I(N__33781));
    InMux I__6711 (
            .O(N__33801),
            .I(N__33778));
    InMux I__6710 (
            .O(N__33800),
            .I(N__33775));
    LocalMux I__6709 (
            .O(N__33797),
            .I(\u1.DMA_control.readDlw_10 ));
    Odrv4 I__6708 (
            .O(N__33792),
            .I(\u1.DMA_control.readDlw_10 ));
    Odrv4 I__6707 (
            .O(N__33787),
            .I(\u1.DMA_control.readDlw_10 ));
    Odrv12 I__6706 (
            .O(N__33784),
            .I(\u1.DMA_control.readDlw_10 ));
    Odrv4 I__6705 (
            .O(N__33781),
            .I(\u1.DMA_control.readDlw_10 ));
    LocalMux I__6704 (
            .O(N__33778),
            .I(\u1.DMA_control.readDlw_10 ));
    LocalMux I__6703 (
            .O(N__33775),
            .I(\u1.DMA_control.readDlw_10 ));
    InMux I__6702 (
            .O(N__33760),
            .I(N__33750));
    InMux I__6701 (
            .O(N__33759),
            .I(N__33750));
    InMux I__6700 (
            .O(N__33758),
            .I(N__33745));
    InMux I__6699 (
            .O(N__33757),
            .I(N__33745));
    CascadeMux I__6698 (
            .O(N__33756),
            .I(N__33742));
    CascadeMux I__6697 (
            .O(N__33755),
            .I(N__33738));
    LocalMux I__6696 (
            .O(N__33750),
            .I(N__33730));
    LocalMux I__6695 (
            .O(N__33745),
            .I(N__33730));
    InMux I__6694 (
            .O(N__33742),
            .I(N__33723));
    InMux I__6693 (
            .O(N__33741),
            .I(N__33723));
    InMux I__6692 (
            .O(N__33738),
            .I(N__33718));
    InMux I__6691 (
            .O(N__33737),
            .I(N__33718));
    InMux I__6690 (
            .O(N__33736),
            .I(N__33713));
    InMux I__6689 (
            .O(N__33735),
            .I(N__33713));
    Span4Mux_v I__6688 (
            .O(N__33730),
            .I(N__33709));
    InMux I__6687 (
            .O(N__33729),
            .I(N__33706));
    InMux I__6686 (
            .O(N__33728),
            .I(N__33703));
    LocalMux I__6685 (
            .O(N__33723),
            .I(N__33700));
    LocalMux I__6684 (
            .O(N__33718),
            .I(N__33697));
    LocalMux I__6683 (
            .O(N__33713),
            .I(N__33693));
    InMux I__6682 (
            .O(N__33712),
            .I(N__33690));
    Sp12to4 I__6681 (
            .O(N__33709),
            .I(N__33687));
    LocalMux I__6680 (
            .O(N__33706),
            .I(N__33682));
    LocalMux I__6679 (
            .O(N__33703),
            .I(N__33682));
    Span4Mux_v I__6678 (
            .O(N__33700),
            .I(N__33677));
    Span4Mux_h I__6677 (
            .O(N__33697),
            .I(N__33677));
    InMux I__6676 (
            .O(N__33696),
            .I(N__33674));
    Span4Mux_h I__6675 (
            .O(N__33693),
            .I(N__33669));
    LocalMux I__6674 (
            .O(N__33690),
            .I(N__33669));
    Odrv12 I__6673 (
            .O(N__33687),
            .I(\u1.DMA_control.readDfw_10 ));
    Odrv12 I__6672 (
            .O(N__33682),
            .I(\u1.DMA_control.readDfw_10 ));
    Odrv4 I__6671 (
            .O(N__33677),
            .I(\u1.DMA_control.readDfw_10 ));
    LocalMux I__6670 (
            .O(N__33674),
            .I(\u1.DMA_control.readDfw_10 ));
    Odrv4 I__6669 (
            .O(N__33669),
            .I(\u1.DMA_control.readDfw_10 ));
    InMux I__6668 (
            .O(N__33658),
            .I(N__33655));
    LocalMux I__6667 (
            .O(N__33655),
            .I(N__33652));
    Span4Mux_v I__6666 (
            .O(N__33652),
            .I(N__33649));
    Odrv4 I__6665 (
            .O(N__33649),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_26 ));
    InMux I__6664 (
            .O(N__33646),
            .I(N__33643));
    LocalMux I__6663 (
            .O(N__33643),
            .I(N__33640));
    Span4Mux_s3_v I__6662 (
            .O(N__33640),
            .I(N__33637));
    Sp12to4 I__6661 (
            .O(N__33637),
            .I(N__33634));
    Odrv12 I__6660 (
            .O(N__33634),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_13 ));
    InMux I__6659 (
            .O(N__33631),
            .I(N__33628));
    LocalMux I__6658 (
            .O(N__33628),
            .I(N__33625));
    Span4Mux_v I__6657 (
            .O(N__33625),
            .I(N__33622));
    Odrv4 I__6656 (
            .O(N__33622),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_13 ));
    CascadeMux I__6655 (
            .O(N__33619),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI6TFTZ0Z_13_cascade_ ));
    InMux I__6654 (
            .O(N__33616),
            .I(N__33613));
    LocalMux I__6653 (
            .O(N__33613),
            .I(N__33610));
    Odrv4 I__6652 (
            .O(N__33610),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_13 ));
    CascadeMux I__6651 (
            .O(N__33607),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI4PA71Z0Z_13_cascade_ ));
    InMux I__6650 (
            .O(N__33604),
            .I(N__33601));
    LocalMux I__6649 (
            .O(N__33601),
            .I(N__33595));
    InMux I__6648 (
            .O(N__33600),
            .I(N__33588));
    InMux I__6647 (
            .O(N__33599),
            .I(N__33585));
    InMux I__6646 (
            .O(N__33598),
            .I(N__33582));
    Span4Mux_h I__6645 (
            .O(N__33595),
            .I(N__33579));
    InMux I__6644 (
            .O(N__33594),
            .I(N__33576));
    CascadeMux I__6643 (
            .O(N__33593),
            .I(N__33572));
    InMux I__6642 (
            .O(N__33592),
            .I(N__33566));
    InMux I__6641 (
            .O(N__33591),
            .I(N__33566));
    LocalMux I__6640 (
            .O(N__33588),
            .I(N__33563));
    LocalMux I__6639 (
            .O(N__33585),
            .I(N__33555));
    LocalMux I__6638 (
            .O(N__33582),
            .I(N__33555));
    IoSpan4Mux I__6637 (
            .O(N__33579),
            .I(N__33552));
    LocalMux I__6636 (
            .O(N__33576),
            .I(N__33549));
    InMux I__6635 (
            .O(N__33575),
            .I(N__33546));
    InMux I__6634 (
            .O(N__33572),
            .I(N__33543));
    InMux I__6633 (
            .O(N__33571),
            .I(N__33540));
    LocalMux I__6632 (
            .O(N__33566),
            .I(N__33537));
    Span4Mux_h I__6631 (
            .O(N__33563),
            .I(N__33534));
    InMux I__6630 (
            .O(N__33562),
            .I(N__33531));
    InMux I__6629 (
            .O(N__33561),
            .I(N__33525));
    InMux I__6628 (
            .O(N__33560),
            .I(N__33525));
    Span4Mux_h I__6627 (
            .O(N__33555),
            .I(N__33521));
    Span4Mux_s1_v I__6626 (
            .O(N__33552),
            .I(N__33518));
    Span4Mux_v I__6625 (
            .O(N__33549),
            .I(N__33515));
    LocalMux I__6624 (
            .O(N__33546),
            .I(N__33508));
    LocalMux I__6623 (
            .O(N__33543),
            .I(N__33508));
    LocalMux I__6622 (
            .O(N__33540),
            .I(N__33508));
    Span12Mux_h I__6621 (
            .O(N__33537),
            .I(N__33501));
    Sp12to4 I__6620 (
            .O(N__33534),
            .I(N__33501));
    LocalMux I__6619 (
            .O(N__33531),
            .I(N__33501));
    InMux I__6618 (
            .O(N__33530),
            .I(N__33498));
    LocalMux I__6617 (
            .O(N__33525),
            .I(N__33495));
    InMux I__6616 (
            .O(N__33524),
            .I(N__33492));
    Span4Mux_v I__6615 (
            .O(N__33521),
            .I(N__33489));
    Span4Mux_v I__6614 (
            .O(N__33518),
            .I(N__33482));
    Span4Mux_h I__6613 (
            .O(N__33515),
            .I(N__33482));
    Span4Mux_h I__6612 (
            .O(N__33508),
            .I(N__33482));
    Span12Mux_s4_v I__6611 (
            .O(N__33501),
            .I(N__33477));
    LocalMux I__6610 (
            .O(N__33498),
            .I(N__33477));
    Span4Mux_h I__6609 (
            .O(N__33495),
            .I(N__33474));
    LocalMux I__6608 (
            .O(N__33492),
            .I(\u1.DMA_control.readDlw_13 ));
    Odrv4 I__6607 (
            .O(N__33489),
            .I(\u1.DMA_control.readDlw_13 ));
    Odrv4 I__6606 (
            .O(N__33482),
            .I(\u1.DMA_control.readDlw_13 ));
    Odrv12 I__6605 (
            .O(N__33477),
            .I(\u1.DMA_control.readDlw_13 ));
    Odrv4 I__6604 (
            .O(N__33474),
            .I(\u1.DMA_control.readDlw_13 ));
    CascadeMux I__6603 (
            .O(N__33463),
            .I(N__33451));
    InMux I__6602 (
            .O(N__33462),
            .I(N__33447));
    CascadeMux I__6601 (
            .O(N__33461),
            .I(N__33444));
    CascadeMux I__6600 (
            .O(N__33460),
            .I(N__33441));
    InMux I__6599 (
            .O(N__33459),
            .I(N__33437));
    InMux I__6598 (
            .O(N__33458),
            .I(N__33434));
    InMux I__6597 (
            .O(N__33457),
            .I(N__33431));
    InMux I__6596 (
            .O(N__33456),
            .I(N__33426));
    InMux I__6595 (
            .O(N__33455),
            .I(N__33426));
    InMux I__6594 (
            .O(N__33454),
            .I(N__33421));
    InMux I__6593 (
            .O(N__33451),
            .I(N__33416));
    InMux I__6592 (
            .O(N__33450),
            .I(N__33416));
    LocalMux I__6591 (
            .O(N__33447),
            .I(N__33413));
    InMux I__6590 (
            .O(N__33444),
            .I(N__33410));
    InMux I__6589 (
            .O(N__33441),
            .I(N__33407));
    InMux I__6588 (
            .O(N__33440),
            .I(N__33404));
    LocalMux I__6587 (
            .O(N__33437),
            .I(N__33399));
    LocalMux I__6586 (
            .O(N__33434),
            .I(N__33399));
    LocalMux I__6585 (
            .O(N__33431),
            .I(N__33394));
    LocalMux I__6584 (
            .O(N__33426),
            .I(N__33394));
    InMux I__6583 (
            .O(N__33425),
            .I(N__33391));
    InMux I__6582 (
            .O(N__33424),
            .I(N__33388));
    LocalMux I__6581 (
            .O(N__33421),
            .I(N__33385));
    LocalMux I__6580 (
            .O(N__33416),
            .I(N__33380));
    Span4Mux_v I__6579 (
            .O(N__33413),
            .I(N__33380));
    LocalMux I__6578 (
            .O(N__33410),
            .I(N__33377));
    LocalMux I__6577 (
            .O(N__33407),
            .I(N__33368));
    LocalMux I__6576 (
            .O(N__33404),
            .I(N__33368));
    Span4Mux_h I__6575 (
            .O(N__33399),
            .I(N__33368));
    Span4Mux_v I__6574 (
            .O(N__33394),
            .I(N__33368));
    LocalMux I__6573 (
            .O(N__33391),
            .I(N__33363));
    LocalMux I__6572 (
            .O(N__33388),
            .I(N__33363));
    Span4Mux_h I__6571 (
            .O(N__33385),
            .I(N__33360));
    Span4Mux_h I__6570 (
            .O(N__33380),
            .I(N__33355));
    Span4Mux_v I__6569 (
            .O(N__33377),
            .I(N__33355));
    Span4Mux_v I__6568 (
            .O(N__33368),
            .I(N__33352));
    Odrv12 I__6567 (
            .O(N__33363),
            .I(\u1.DMA_control.readDfw_13 ));
    Odrv4 I__6566 (
            .O(N__33360),
            .I(\u1.DMA_control.readDfw_13 ));
    Odrv4 I__6565 (
            .O(N__33355),
            .I(\u1.DMA_control.readDfw_13 ));
    Odrv4 I__6564 (
            .O(N__33352),
            .I(\u1.DMA_control.readDfw_13 ));
    CascadeMux I__6563 (
            .O(N__33343),
            .I(N__33340));
    InMux I__6562 (
            .O(N__33340),
            .I(N__33337));
    LocalMux I__6561 (
            .O(N__33337),
            .I(N__33334));
    Odrv12 I__6560 (
            .O(N__33334),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_25 ));
    InMux I__6559 (
            .O(N__33331),
            .I(N__33328));
    LocalMux I__6558 (
            .O(N__33328),
            .I(N__33325));
    Span12Mux_s4_v I__6557 (
            .O(N__33325),
            .I(N__33322));
    Odrv12 I__6556 (
            .O(N__33322),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_25 ));
    InMux I__6555 (
            .O(N__33319),
            .I(N__33316));
    LocalMux I__6554 (
            .O(N__33316),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_25 ));
    InMux I__6553 (
            .O(N__33313),
            .I(N__33310));
    LocalMux I__6552 (
            .O(N__33310),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI4T0RZ0Z_25 ));
    CascadeMux I__6551 (
            .O(N__33307),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI8H9KZ0Z_25_cascade_ ));
    InMux I__6550 (
            .O(N__33304),
            .I(N__33301));
    LocalMux I__6549 (
            .O(N__33301),
            .I(N__33298));
    Span4Mux_v I__6548 (
            .O(N__33298),
            .I(N__33295));
    Span4Mux_h I__6547 (
            .O(N__33295),
            .I(N__33292));
    Odrv4 I__6546 (
            .O(N__33292),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_10 ));
    InMux I__6545 (
            .O(N__33289),
            .I(N__33286));
    LocalMux I__6544 (
            .O(N__33286),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_10 ));
    InMux I__6543 (
            .O(N__33283),
            .I(N__33280));
    LocalMux I__6542 (
            .O(N__33280),
            .I(N__33277));
    Odrv4 I__6541 (
            .O(N__33277),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_10 ));
    InMux I__6540 (
            .O(N__33274),
            .I(N__33271));
    LocalMux I__6539 (
            .O(N__33271),
            .I(N__33268));
    Span12Mux_h I__6538 (
            .O(N__33268),
            .I(N__33265));
    Odrv12 I__6537 (
            .O(N__33265),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_10 ));
    CEMux I__6536 (
            .O(N__33262),
            .I(N__33257));
    CEMux I__6535 (
            .O(N__33261),
            .I(N__33253));
    CEMux I__6534 (
            .O(N__33260),
            .I(N__33250));
    LocalMux I__6533 (
            .O(N__33257),
            .I(N__33247));
    CEMux I__6532 (
            .O(N__33256),
            .I(N__33244));
    LocalMux I__6531 (
            .O(N__33253),
            .I(N__33241));
    LocalMux I__6530 (
            .O(N__33250),
            .I(N__33238));
    Span4Mux_h I__6529 (
            .O(N__33247),
            .I(N__33235));
    LocalMux I__6528 (
            .O(N__33244),
            .I(N__33232));
    Span4Mux_h I__6527 (
            .O(N__33241),
            .I(N__33229));
    Span4Mux_h I__6526 (
            .O(N__33238),
            .I(N__33226));
    Odrv4 I__6525 (
            .O(N__33235),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_awe1 ));
    Odrv12 I__6524 (
            .O(N__33232),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_awe1 ));
    Odrv4 I__6523 (
            .O(N__33229),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_awe1 ));
    Odrv4 I__6522 (
            .O(N__33226),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_awe1 ));
    InMux I__6521 (
            .O(N__33217),
            .I(N__33214));
    LocalMux I__6520 (
            .O(N__33214),
            .I(N__33211));
    Span4Mux_h I__6519 (
            .O(N__33211),
            .I(N__33208));
    Odrv4 I__6518 (
            .O(N__33208),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_29 ));
    InMux I__6517 (
            .O(N__33205),
            .I(N__33202));
    LocalMux I__6516 (
            .O(N__33202),
            .I(N__33199));
    Span4Mux_h I__6515 (
            .O(N__33199),
            .I(N__33196));
    Odrv4 I__6514 (
            .O(N__33196),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_29 ));
    InMux I__6513 (
            .O(N__33193),
            .I(N__33190));
    LocalMux I__6512 (
            .O(N__33190),
            .I(N__33187));
    Odrv4 I__6511 (
            .O(N__33187),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_29 ));
    InMux I__6510 (
            .O(N__33184),
            .I(N__33181));
    LocalMux I__6509 (
            .O(N__33181),
            .I(N__33178));
    Span4Mux_v I__6508 (
            .O(N__33178),
            .I(N__33175));
    Span4Mux_h I__6507 (
            .O(N__33175),
            .I(N__33172));
    Odrv4 I__6506 (
            .O(N__33172),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_29 ));
    CascadeMux I__6505 (
            .O(N__33169),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIKDITZ0Z_29_cascade_ ));
    CascadeMux I__6504 (
            .O(N__33166),
            .I(mem_mem_ram6__RNIPHE71_29_cascade_));
    InMux I__6503 (
            .O(N__33163),
            .I(N__33160));
    LocalMux I__6502 (
            .O(N__33160),
            .I(N__33157));
    Span4Mux_v I__6501 (
            .O(N__33157),
            .I(N__33154));
    Odrv4 I__6500 (
            .O(N__33154),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_29 ));
    InMux I__6499 (
            .O(N__33151),
            .I(N__33148));
    LocalMux I__6498 (
            .O(N__33148),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_29 ));
    InMux I__6497 (
            .O(N__33145),
            .I(N__33142));
    LocalMux I__6496 (
            .O(N__33142),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIGP9KZ0Z_29 ));
    CascadeMux I__6495 (
            .O(N__33139),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIC51RZ0Z_29_cascade_ ));
    InMux I__6494 (
            .O(N__33136),
            .I(N__33133));
    LocalMux I__6493 (
            .O(N__33133),
            .I(iQ_RNIE9IM1_2));
    InMux I__6492 (
            .O(N__33130),
            .I(N__33127));
    LocalMux I__6491 (
            .O(N__33127),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_29 ));
    InMux I__6490 (
            .O(N__33124),
            .I(N__33118));
    InMux I__6489 (
            .O(N__33123),
            .I(N__33118));
    LocalMux I__6488 (
            .O(N__33118),
            .I(N__33115));
    Span4Mux_v I__6487 (
            .O(N__33115),
            .I(N__33112));
    Span4Mux_h I__6486 (
            .O(N__33112),
            .I(N__33108));
    InMux I__6485 (
            .O(N__33111),
            .I(N__33105));
    Span4Mux_h I__6484 (
            .O(N__33108),
            .I(N__33102));
    LocalMux I__6483 (
            .O(N__33105),
            .I(N__33099));
    Span4Mux_v I__6482 (
            .O(N__33102),
            .I(N__33096));
    Span4Mux_h I__6481 (
            .O(N__33099),
            .I(N__33093));
    Span4Mux_h I__6480 (
            .O(N__33096),
            .I(N__33088));
    Span4Mux_v I__6479 (
            .O(N__33093),
            .I(N__33088));
    Odrv4 I__6478 (
            .O(N__33088),
            .I(dd_pad_i_c_11));
    InMux I__6477 (
            .O(N__33085),
            .I(N__33082));
    LocalMux I__6476 (
            .O(N__33082),
            .I(N__33079));
    Odrv4 I__6475 (
            .O(N__33079),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_26 ));
    CascadeMux I__6474 (
            .O(N__33076),
            .I(N__33069));
    InMux I__6473 (
            .O(N__33075),
            .I(N__33063));
    InMux I__6472 (
            .O(N__33074),
            .I(N__33063));
    InMux I__6471 (
            .O(N__33073),
            .I(N__33056));
    InMux I__6470 (
            .O(N__33072),
            .I(N__33056));
    InMux I__6469 (
            .O(N__33069),
            .I(N__33049));
    InMux I__6468 (
            .O(N__33068),
            .I(N__33049));
    LocalMux I__6467 (
            .O(N__33063),
            .I(N__33046));
    InMux I__6466 (
            .O(N__33062),
            .I(N__33041));
    InMux I__6465 (
            .O(N__33061),
            .I(N__33041));
    LocalMux I__6464 (
            .O(N__33056),
            .I(N__33036));
    InMux I__6463 (
            .O(N__33055),
            .I(N__33031));
    InMux I__6462 (
            .O(N__33054),
            .I(N__33031));
    LocalMux I__6461 (
            .O(N__33049),
            .I(N__33025));
    Sp12to4 I__6460 (
            .O(N__33046),
            .I(N__33020));
    LocalMux I__6459 (
            .O(N__33041),
            .I(N__33020));
    InMux I__6458 (
            .O(N__33040),
            .I(N__33015));
    InMux I__6457 (
            .O(N__33039),
            .I(N__33015));
    Span4Mux_s3_v I__6456 (
            .O(N__33036),
            .I(N__33010));
    LocalMux I__6455 (
            .O(N__33031),
            .I(N__33010));
    InMux I__6454 (
            .O(N__33030),
            .I(N__33005));
    InMux I__6453 (
            .O(N__33029),
            .I(N__33005));
    InMux I__6452 (
            .O(N__33028),
            .I(N__33002));
    Span4Mux_v I__6451 (
            .O(N__33025),
            .I(N__32999));
    Span12Mux_s7_v I__6450 (
            .O(N__33020),
            .I(N__32994));
    LocalMux I__6449 (
            .O(N__33015),
            .I(N__32994));
    Span4Mux_v I__6448 (
            .O(N__33010),
            .I(N__32989));
    LocalMux I__6447 (
            .O(N__33005),
            .I(N__32989));
    LocalMux I__6446 (
            .O(N__33002),
            .I(\u1.DMA_control.readDlw_14 ));
    Odrv4 I__6445 (
            .O(N__32999),
            .I(\u1.DMA_control.readDlw_14 ));
    Odrv12 I__6444 (
            .O(N__32994),
            .I(\u1.DMA_control.readDlw_14 ));
    Odrv4 I__6443 (
            .O(N__32989),
            .I(\u1.DMA_control.readDlw_14 ));
    CascadeMux I__6442 (
            .O(N__32980),
            .I(N__32974));
    CascadeMux I__6441 (
            .O(N__32979),
            .I(N__32970));
    CascadeMux I__6440 (
            .O(N__32978),
            .I(N__32964));
    CascadeMux I__6439 (
            .O(N__32977),
            .I(N__32960));
    InMux I__6438 (
            .O(N__32974),
            .I(N__32954));
    InMux I__6437 (
            .O(N__32973),
            .I(N__32954));
    InMux I__6436 (
            .O(N__32970),
            .I(N__32949));
    InMux I__6435 (
            .O(N__32969),
            .I(N__32949));
    CascadeMux I__6434 (
            .O(N__32968),
            .I(N__32946));
    CascadeMux I__6433 (
            .O(N__32967),
            .I(N__32941));
    InMux I__6432 (
            .O(N__32964),
            .I(N__32935));
    InMux I__6431 (
            .O(N__32963),
            .I(N__32935));
    InMux I__6430 (
            .O(N__32960),
            .I(N__32930));
    InMux I__6429 (
            .O(N__32959),
            .I(N__32930));
    LocalMux I__6428 (
            .O(N__32954),
            .I(N__32927));
    LocalMux I__6427 (
            .O(N__32949),
            .I(N__32923));
    InMux I__6426 (
            .O(N__32946),
            .I(N__32918));
    InMux I__6425 (
            .O(N__32945),
            .I(N__32918));
    InMux I__6424 (
            .O(N__32944),
            .I(N__32915));
    InMux I__6423 (
            .O(N__32941),
            .I(N__32910));
    InMux I__6422 (
            .O(N__32940),
            .I(N__32910));
    LocalMux I__6421 (
            .O(N__32935),
            .I(N__32903));
    LocalMux I__6420 (
            .O(N__32930),
            .I(N__32903));
    Span4Mux_v I__6419 (
            .O(N__32927),
            .I(N__32903));
    InMux I__6418 (
            .O(N__32926),
            .I(N__32900));
    Span4Mux_v I__6417 (
            .O(N__32923),
            .I(N__32895));
    LocalMux I__6416 (
            .O(N__32918),
            .I(N__32895));
    LocalMux I__6415 (
            .O(N__32915),
            .I(N__32890));
    LocalMux I__6414 (
            .O(N__32910),
            .I(N__32890));
    Span4Mux_h I__6413 (
            .O(N__32903),
            .I(N__32885));
    LocalMux I__6412 (
            .O(N__32900),
            .I(N__32885));
    Span4Mux_h I__6411 (
            .O(N__32895),
            .I(N__32882));
    Span4Mux_v I__6410 (
            .O(N__32890),
            .I(N__32879));
    Span4Mux_v I__6409 (
            .O(N__32885),
            .I(N__32876));
    Span4Mux_v I__6408 (
            .O(N__32882),
            .I(N__32873));
    Odrv4 I__6407 (
            .O(N__32879),
            .I(\u1.DMA_control.readDfw_14 ));
    Odrv4 I__6406 (
            .O(N__32876),
            .I(\u1.DMA_control.readDfw_14 ));
    Odrv4 I__6405 (
            .O(N__32873),
            .I(\u1.DMA_control.readDfw_14 ));
    InMux I__6404 (
            .O(N__32866),
            .I(N__32860));
    InMux I__6403 (
            .O(N__32865),
            .I(N__32860));
    LocalMux I__6402 (
            .O(N__32860),
            .I(N__32857));
    Span4Mux_v I__6401 (
            .O(N__32857),
            .I(N__32854));
    Span4Mux_h I__6400 (
            .O(N__32854),
            .I(N__32851));
    Span4Mux_h I__6399 (
            .O(N__32851),
            .I(N__32847));
    InMux I__6398 (
            .O(N__32850),
            .I(N__32844));
    Span4Mux_h I__6397 (
            .O(N__32847),
            .I(N__32839));
    LocalMux I__6396 (
            .O(N__32844),
            .I(N__32839));
    Span4Mux_v I__6395 (
            .O(N__32839),
            .I(N__32836));
    Span4Mux_v I__6394 (
            .O(N__32836),
            .I(N__32833));
    Odrv4 I__6393 (
            .O(N__32833),
            .I(dd_pad_i_c_14));
    InMux I__6392 (
            .O(N__32830),
            .I(N__32827));
    LocalMux I__6391 (
            .O(N__32827),
            .I(N__32816));
    InMux I__6390 (
            .O(N__32826),
            .I(N__32813));
    InMux I__6389 (
            .O(N__32825),
            .I(N__32810));
    InMux I__6388 (
            .O(N__32824),
            .I(N__32807));
    InMux I__6387 (
            .O(N__32823),
            .I(N__32802));
    InMux I__6386 (
            .O(N__32822),
            .I(N__32799));
    InMux I__6385 (
            .O(N__32821),
            .I(N__32796));
    InMux I__6384 (
            .O(N__32820),
            .I(N__32790));
    InMux I__6383 (
            .O(N__32819),
            .I(N__32790));
    Span4Mux_h I__6382 (
            .O(N__32816),
            .I(N__32786));
    LocalMux I__6381 (
            .O(N__32813),
            .I(N__32779));
    LocalMux I__6380 (
            .O(N__32810),
            .I(N__32779));
    LocalMux I__6379 (
            .O(N__32807),
            .I(N__32779));
    InMux I__6378 (
            .O(N__32806),
            .I(N__32774));
    InMux I__6377 (
            .O(N__32805),
            .I(N__32774));
    LocalMux I__6376 (
            .O(N__32802),
            .I(N__32767));
    LocalMux I__6375 (
            .O(N__32799),
            .I(N__32767));
    LocalMux I__6374 (
            .O(N__32796),
            .I(N__32767));
    CascadeMux I__6373 (
            .O(N__32795),
            .I(N__32764));
    LocalMux I__6372 (
            .O(N__32790),
            .I(N__32759));
    InMux I__6371 (
            .O(N__32789),
            .I(N__32756));
    Span4Mux_h I__6370 (
            .O(N__32786),
            .I(N__32749));
    Span4Mux_h I__6369 (
            .O(N__32779),
            .I(N__32749));
    LocalMux I__6368 (
            .O(N__32774),
            .I(N__32749));
    Span4Mux_h I__6367 (
            .O(N__32767),
            .I(N__32746));
    InMux I__6366 (
            .O(N__32764),
            .I(N__32741));
    InMux I__6365 (
            .O(N__32763),
            .I(N__32741));
    InMux I__6364 (
            .O(N__32762),
            .I(N__32738));
    Span12Mux_s7_v I__6363 (
            .O(N__32759),
            .I(N__32733));
    LocalMux I__6362 (
            .O(N__32756),
            .I(N__32733));
    Span4Mux_v I__6361 (
            .O(N__32749),
            .I(N__32730));
    Span4Mux_v I__6360 (
            .O(N__32746),
            .I(N__32725));
    LocalMux I__6359 (
            .O(N__32741),
            .I(N__32725));
    LocalMux I__6358 (
            .O(N__32738),
            .I(\u1.DMA_control.readDlw_6 ));
    Odrv12 I__6357 (
            .O(N__32733),
            .I(\u1.DMA_control.readDlw_6 ));
    Odrv4 I__6356 (
            .O(N__32730),
            .I(\u1.DMA_control.readDlw_6 ));
    Odrv4 I__6355 (
            .O(N__32725),
            .I(\u1.DMA_control.readDlw_6 ));
    CascadeMux I__6354 (
            .O(N__32716),
            .I(N__32708));
    InMux I__6353 (
            .O(N__32715),
            .I(N__32701));
    InMux I__6352 (
            .O(N__32714),
            .I(N__32701));
    InMux I__6351 (
            .O(N__32713),
            .I(N__32698));
    InMux I__6350 (
            .O(N__32712),
            .I(N__32693));
    InMux I__6349 (
            .O(N__32711),
            .I(N__32693));
    InMux I__6348 (
            .O(N__32708),
            .I(N__32687));
    InMux I__6347 (
            .O(N__32707),
            .I(N__32687));
    InMux I__6346 (
            .O(N__32706),
            .I(N__32684));
    LocalMux I__6345 (
            .O(N__32701),
            .I(N__32676));
    LocalMux I__6344 (
            .O(N__32698),
            .I(N__32676));
    LocalMux I__6343 (
            .O(N__32693),
            .I(N__32673));
    InMux I__6342 (
            .O(N__32692),
            .I(N__32670));
    LocalMux I__6341 (
            .O(N__32687),
            .I(N__32667));
    LocalMux I__6340 (
            .O(N__32684),
            .I(N__32664));
    InMux I__6339 (
            .O(N__32683),
            .I(N__32661));
    InMux I__6338 (
            .O(N__32682),
            .I(N__32658));
    InMux I__6337 (
            .O(N__32681),
            .I(N__32655));
    Span4Mux_h I__6336 (
            .O(N__32676),
            .I(N__32652));
    Span4Mux_h I__6335 (
            .O(N__32673),
            .I(N__32647));
    LocalMux I__6334 (
            .O(N__32670),
            .I(N__32647));
    Span4Mux_v I__6333 (
            .O(N__32667),
            .I(N__32640));
    Span4Mux_h I__6332 (
            .O(N__32664),
            .I(N__32640));
    LocalMux I__6331 (
            .O(N__32661),
            .I(N__32640));
    LocalMux I__6330 (
            .O(N__32658),
            .I(N__32635));
    LocalMux I__6329 (
            .O(N__32655),
            .I(N__32635));
    Span4Mux_v I__6328 (
            .O(N__32652),
            .I(N__32630));
    Span4Mux_v I__6327 (
            .O(N__32647),
            .I(N__32623));
    Span4Mux_h I__6326 (
            .O(N__32640),
            .I(N__32623));
    Span4Mux_v I__6325 (
            .O(N__32635),
            .I(N__32623));
    InMux I__6324 (
            .O(N__32634),
            .I(N__32618));
    InMux I__6323 (
            .O(N__32633),
            .I(N__32618));
    Odrv4 I__6322 (
            .O(N__32630),
            .I(\u1.DMA_control.readDfw_6 ));
    Odrv4 I__6321 (
            .O(N__32623),
            .I(\u1.DMA_control.readDfw_6 ));
    LocalMux I__6320 (
            .O(N__32618),
            .I(\u1.DMA_control.readDfw_6 ));
    InMux I__6319 (
            .O(N__32611),
            .I(N__32602));
    InMux I__6318 (
            .O(N__32610),
            .I(N__32602));
    InMux I__6317 (
            .O(N__32609),
            .I(N__32594));
    InMux I__6316 (
            .O(N__32608),
            .I(N__32591));
    CascadeMux I__6315 (
            .O(N__32607),
            .I(N__32586));
    LocalMux I__6314 (
            .O(N__32602),
            .I(N__32581));
    InMux I__6313 (
            .O(N__32601),
            .I(N__32576));
    InMux I__6312 (
            .O(N__32600),
            .I(N__32576));
    InMux I__6311 (
            .O(N__32599),
            .I(N__32571));
    InMux I__6310 (
            .O(N__32598),
            .I(N__32571));
    InMux I__6309 (
            .O(N__32597),
            .I(N__32568));
    LocalMux I__6308 (
            .O(N__32594),
            .I(N__32563));
    LocalMux I__6307 (
            .O(N__32591),
            .I(N__32563));
    InMux I__6306 (
            .O(N__32590),
            .I(N__32558));
    InMux I__6305 (
            .O(N__32589),
            .I(N__32558));
    InMux I__6304 (
            .O(N__32586),
            .I(N__32553));
    InMux I__6303 (
            .O(N__32585),
            .I(N__32553));
    InMux I__6302 (
            .O(N__32584),
            .I(N__32550));
    Span4Mux_h I__6301 (
            .O(N__32581),
            .I(N__32544));
    LocalMux I__6300 (
            .O(N__32576),
            .I(N__32544));
    LocalMux I__6299 (
            .O(N__32571),
            .I(N__32541));
    LocalMux I__6298 (
            .O(N__32568),
            .I(N__32538));
    Span4Mux_v I__6297 (
            .O(N__32563),
            .I(N__32535));
    LocalMux I__6296 (
            .O(N__32558),
            .I(N__32532));
    LocalMux I__6295 (
            .O(N__32553),
            .I(N__32527));
    LocalMux I__6294 (
            .O(N__32550),
            .I(N__32527));
    InMux I__6293 (
            .O(N__32549),
            .I(N__32524));
    Span4Mux_v I__6292 (
            .O(N__32544),
            .I(N__32521));
    Span4Mux_v I__6291 (
            .O(N__32541),
            .I(N__32516));
    Span4Mux_v I__6290 (
            .O(N__32538),
            .I(N__32516));
    Span4Mux_h I__6289 (
            .O(N__32535),
            .I(N__32511));
    Span4Mux_h I__6288 (
            .O(N__32532),
            .I(N__32511));
    Span4Mux_h I__6287 (
            .O(N__32527),
            .I(N__32508));
    LocalMux I__6286 (
            .O(N__32524),
            .I(\u1.DMA_control.readDlw_15 ));
    Odrv4 I__6285 (
            .O(N__32521),
            .I(\u1.DMA_control.readDlw_15 ));
    Odrv4 I__6284 (
            .O(N__32516),
            .I(\u1.DMA_control.readDlw_15 ));
    Odrv4 I__6283 (
            .O(N__32511),
            .I(\u1.DMA_control.readDlw_15 ));
    Odrv4 I__6282 (
            .O(N__32508),
            .I(\u1.DMA_control.readDlw_15 ));
    CascadeMux I__6281 (
            .O(N__32497),
            .I(N__32493));
    CascadeMux I__6280 (
            .O(N__32496),
            .I(N__32486));
    InMux I__6279 (
            .O(N__32493),
            .I(N__32480));
    InMux I__6278 (
            .O(N__32492),
            .I(N__32480));
    CascadeMux I__6277 (
            .O(N__32491),
            .I(N__32474));
    InMux I__6276 (
            .O(N__32490),
            .I(N__32468));
    InMux I__6275 (
            .O(N__32489),
            .I(N__32468));
    InMux I__6274 (
            .O(N__32486),
            .I(N__32463));
    InMux I__6273 (
            .O(N__32485),
            .I(N__32463));
    LocalMux I__6272 (
            .O(N__32480),
            .I(N__32460));
    InMux I__6271 (
            .O(N__32479),
            .I(N__32457));
    InMux I__6270 (
            .O(N__32478),
            .I(N__32454));
    InMux I__6269 (
            .O(N__32477),
            .I(N__32451));
    InMux I__6268 (
            .O(N__32474),
            .I(N__32446));
    InMux I__6267 (
            .O(N__32473),
            .I(N__32446));
    LocalMux I__6266 (
            .O(N__32468),
            .I(N__32440));
    LocalMux I__6265 (
            .O(N__32463),
            .I(N__32437));
    Span4Mux_h I__6264 (
            .O(N__32460),
            .I(N__32428));
    LocalMux I__6263 (
            .O(N__32457),
            .I(N__32428));
    LocalMux I__6262 (
            .O(N__32454),
            .I(N__32428));
    LocalMux I__6261 (
            .O(N__32451),
            .I(N__32428));
    LocalMux I__6260 (
            .O(N__32446),
            .I(N__32425));
    InMux I__6259 (
            .O(N__32445),
            .I(N__32420));
    InMux I__6258 (
            .O(N__32444),
            .I(N__32420));
    InMux I__6257 (
            .O(N__32443),
            .I(N__32417));
    Span12Mux_h I__6256 (
            .O(N__32440),
            .I(N__32414));
    Span4Mux_v I__6255 (
            .O(N__32437),
            .I(N__32409));
    Span4Mux_v I__6254 (
            .O(N__32428),
            .I(N__32409));
    Span4Mux_h I__6253 (
            .O(N__32425),
            .I(N__32406));
    LocalMux I__6252 (
            .O(N__32420),
            .I(N__32401));
    LocalMux I__6251 (
            .O(N__32417),
            .I(N__32401));
    Odrv12 I__6250 (
            .O(N__32414),
            .I(\u1.DMA_control.readDfw_15 ));
    Odrv4 I__6249 (
            .O(N__32409),
            .I(\u1.DMA_control.readDfw_15 ));
    Odrv4 I__6248 (
            .O(N__32406),
            .I(\u1.DMA_control.readDfw_15 ));
    Odrv12 I__6247 (
            .O(N__32401),
            .I(\u1.DMA_control.readDfw_15 ));
    InMux I__6246 (
            .O(N__32392),
            .I(N__32386));
    InMux I__6245 (
            .O(N__32391),
            .I(N__32386));
    LocalMux I__6244 (
            .O(N__32386),
            .I(N__32383));
    Span4Mux_h I__6243 (
            .O(N__32383),
            .I(N__32379));
    InMux I__6242 (
            .O(N__32382),
            .I(N__32376));
    Span4Mux_h I__6241 (
            .O(N__32379),
            .I(N__32371));
    LocalMux I__6240 (
            .O(N__32376),
            .I(N__32371));
    Span4Mux_v I__6239 (
            .O(N__32371),
            .I(N__32368));
    Span4Mux_v I__6238 (
            .O(N__32368),
            .I(N__32365));
    Span4Mux_v I__6237 (
            .O(N__32365),
            .I(N__32362));
    Sp12to4 I__6236 (
            .O(N__32362),
            .I(N__32359));
    Odrv12 I__6235 (
            .O(N__32359),
            .I(dd_pad_i_c_15));
    InMux I__6234 (
            .O(N__32356),
            .I(N__32352));
    InMux I__6233 (
            .O(N__32355),
            .I(N__32349));
    LocalMux I__6232 (
            .O(N__32352),
            .I(N__32346));
    LocalMux I__6231 (
            .O(N__32349),
            .I(N__32343));
    Span4Mux_v I__6230 (
            .O(N__32346),
            .I(N__32340));
    Span4Mux_v I__6229 (
            .O(N__32343),
            .I(N__32337));
    Span4Mux_h I__6228 (
            .O(N__32340),
            .I(N__32333));
    Span4Mux_h I__6227 (
            .O(N__32337),
            .I(N__32330));
    InMux I__6226 (
            .O(N__32336),
            .I(N__32327));
    Span4Mux_h I__6225 (
            .O(N__32333),
            .I(N__32324));
    Span4Mux_h I__6224 (
            .O(N__32330),
            .I(N__32319));
    LocalMux I__6223 (
            .O(N__32327),
            .I(N__32319));
    Span4Mux_h I__6222 (
            .O(N__32324),
            .I(N__32316));
    Span4Mux_v I__6221 (
            .O(N__32319),
            .I(N__32313));
    Span4Mux_v I__6220 (
            .O(N__32316),
            .I(N__32310));
    Span4Mux_v I__6219 (
            .O(N__32313),
            .I(N__32307));
    Odrv4 I__6218 (
            .O(N__32310),
            .I(dd_pad_i_c_2));
    Odrv4 I__6217 (
            .O(N__32307),
            .I(dd_pad_i_c_2));
    InMux I__6216 (
            .O(N__32302),
            .I(N__32299));
    LocalMux I__6215 (
            .O(N__32299),
            .I(N__32294));
    InMux I__6214 (
            .O(N__32298),
            .I(N__32291));
    InMux I__6213 (
            .O(N__32297),
            .I(N__32288));
    Sp12to4 I__6212 (
            .O(N__32294),
            .I(N__32285));
    LocalMux I__6211 (
            .O(N__32291),
            .I(N__32282));
    LocalMux I__6210 (
            .O(N__32288),
            .I(N__32279));
    Span12Mux_v I__6209 (
            .O(N__32285),
            .I(N__32276));
    Span4Mux_v I__6208 (
            .O(N__32282),
            .I(N__32273));
    Span4Mux_v I__6207 (
            .O(N__32279),
            .I(N__32270));
    Span12Mux_h I__6206 (
            .O(N__32276),
            .I(N__32267));
    Span4Mux_v I__6205 (
            .O(N__32273),
            .I(N__32262));
    Span4Mux_h I__6204 (
            .O(N__32270),
            .I(N__32262));
    Odrv12 I__6203 (
            .O(N__32267),
            .I(dd_pad_i_c_10));
    Odrv4 I__6202 (
            .O(N__32262),
            .I(dd_pad_i_c_10));
    InMux I__6201 (
            .O(N__32257),
            .I(N__32254));
    LocalMux I__6200 (
            .O(N__32254),
            .I(N__32251));
    Span4Mux_v I__6199 (
            .O(N__32251),
            .I(N__32248));
    Odrv4 I__6198 (
            .O(N__32248),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_14 ));
    InMux I__6197 (
            .O(N__32245),
            .I(N__32242));
    LocalMux I__6196 (
            .O(N__32242),
            .I(N__32239));
    Span4Mux_h I__6195 (
            .O(N__32239),
            .I(N__32236));
    Span4Mux_v I__6194 (
            .O(N__32236),
            .I(N__32233));
    Span4Mux_v I__6193 (
            .O(N__32233),
            .I(N__32230));
    Odrv4 I__6192 (
            .O(N__32230),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_14 ));
    InMux I__6191 (
            .O(N__32227),
            .I(N__32224));
    LocalMux I__6190 (
            .O(N__32224),
            .I(N__32221));
    Span4Mux_v I__6189 (
            .O(N__32221),
            .I(N__32218));
    Odrv4 I__6188 (
            .O(N__32218),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI0NUQZ0Z_14 ));
    CascadeMux I__6187 (
            .O(N__32215),
            .I(N__32208));
    InMux I__6186 (
            .O(N__32214),
            .I(N__32201));
    InMux I__6185 (
            .O(N__32213),
            .I(N__32201));
    InMux I__6184 (
            .O(N__32212),
            .I(N__32198));
    CascadeMux I__6183 (
            .O(N__32211),
            .I(N__32195));
    InMux I__6182 (
            .O(N__32208),
            .I(N__32189));
    InMux I__6181 (
            .O(N__32207),
            .I(N__32189));
    InMux I__6180 (
            .O(N__32206),
            .I(N__32186));
    LocalMux I__6179 (
            .O(N__32201),
            .I(N__32179));
    LocalMux I__6178 (
            .O(N__32198),
            .I(N__32179));
    InMux I__6177 (
            .O(N__32195),
            .I(N__32174));
    InMux I__6176 (
            .O(N__32194),
            .I(N__32174));
    LocalMux I__6175 (
            .O(N__32189),
            .I(N__32168));
    LocalMux I__6174 (
            .O(N__32186),
            .I(N__32168));
    InMux I__6173 (
            .O(N__32185),
            .I(N__32165));
    InMux I__6172 (
            .O(N__32184),
            .I(N__32159));
    Span4Mux_v I__6171 (
            .O(N__32179),
            .I(N__32154));
    LocalMux I__6170 (
            .O(N__32174),
            .I(N__32154));
    InMux I__6169 (
            .O(N__32173),
            .I(N__32151));
    Span4Mux_h I__6168 (
            .O(N__32168),
            .I(N__32146));
    LocalMux I__6167 (
            .O(N__32165),
            .I(N__32146));
    InMux I__6166 (
            .O(N__32164),
            .I(N__32141));
    InMux I__6165 (
            .O(N__32163),
            .I(N__32141));
    InMux I__6164 (
            .O(N__32162),
            .I(N__32137));
    LocalMux I__6163 (
            .O(N__32159),
            .I(N__32134));
    Span4Mux_v I__6162 (
            .O(N__32154),
            .I(N__32131));
    LocalMux I__6161 (
            .O(N__32151),
            .I(N__32128));
    Span4Mux_v I__6160 (
            .O(N__32146),
            .I(N__32123));
    LocalMux I__6159 (
            .O(N__32141),
            .I(N__32123));
    InMux I__6158 (
            .O(N__32140),
            .I(N__32120));
    LocalMux I__6157 (
            .O(N__32137),
            .I(\u1.DMA_control.readDlw_12 ));
    Odrv12 I__6156 (
            .O(N__32134),
            .I(\u1.DMA_control.readDlw_12 ));
    Odrv4 I__6155 (
            .O(N__32131),
            .I(\u1.DMA_control.readDlw_12 ));
    Odrv12 I__6154 (
            .O(N__32128),
            .I(\u1.DMA_control.readDlw_12 ));
    Odrv4 I__6153 (
            .O(N__32123),
            .I(\u1.DMA_control.readDlw_12 ));
    LocalMux I__6152 (
            .O(N__32120),
            .I(\u1.DMA_control.readDlw_12 ));
    CascadeMux I__6151 (
            .O(N__32107),
            .I(N__32104));
    InMux I__6150 (
            .O(N__32104),
            .I(N__32097));
    InMux I__6149 (
            .O(N__32103),
            .I(N__32097));
    CascadeMux I__6148 (
            .O(N__32102),
            .I(N__32093));
    LocalMux I__6147 (
            .O(N__32097),
            .I(N__32089));
    InMux I__6146 (
            .O(N__32096),
            .I(N__32084));
    InMux I__6145 (
            .O(N__32093),
            .I(N__32076));
    InMux I__6144 (
            .O(N__32092),
            .I(N__32076));
    Span4Mux_s3_v I__6143 (
            .O(N__32089),
            .I(N__32071));
    InMux I__6142 (
            .O(N__32088),
            .I(N__32066));
    InMux I__6141 (
            .O(N__32087),
            .I(N__32066));
    LocalMux I__6140 (
            .O(N__32084),
            .I(N__32063));
    CascadeMux I__6139 (
            .O(N__32083),
            .I(N__32060));
    InMux I__6138 (
            .O(N__32082),
            .I(N__32056));
    InMux I__6137 (
            .O(N__32081),
            .I(N__32053));
    LocalMux I__6136 (
            .O(N__32076),
            .I(N__32050));
    InMux I__6135 (
            .O(N__32075),
            .I(N__32046));
    InMux I__6134 (
            .O(N__32074),
            .I(N__32043));
    Span4Mux_h I__6133 (
            .O(N__32071),
            .I(N__32040));
    LocalMux I__6132 (
            .O(N__32066),
            .I(N__32035));
    Span4Mux_v I__6131 (
            .O(N__32063),
            .I(N__32035));
    InMux I__6130 (
            .O(N__32060),
            .I(N__32030));
    InMux I__6129 (
            .O(N__32059),
            .I(N__32030));
    LocalMux I__6128 (
            .O(N__32056),
            .I(N__32023));
    LocalMux I__6127 (
            .O(N__32053),
            .I(N__32023));
    Span4Mux_h I__6126 (
            .O(N__32050),
            .I(N__32023));
    InMux I__6125 (
            .O(N__32049),
            .I(N__32020));
    LocalMux I__6124 (
            .O(N__32046),
            .I(N__32017));
    LocalMux I__6123 (
            .O(N__32043),
            .I(N__32014));
    Span4Mux_v I__6122 (
            .O(N__32040),
            .I(N__32011));
    Span4Mux_v I__6121 (
            .O(N__32035),
            .I(N__32008));
    LocalMux I__6120 (
            .O(N__32030),
            .I(N__32003));
    Span4Mux_v I__6119 (
            .O(N__32023),
            .I(N__32003));
    LocalMux I__6118 (
            .O(N__32020),
            .I(\u1.DMA_control.readDfw_12 ));
    Odrv12 I__6117 (
            .O(N__32017),
            .I(\u1.DMA_control.readDfw_12 ));
    Odrv12 I__6116 (
            .O(N__32014),
            .I(\u1.DMA_control.readDfw_12 ));
    Odrv4 I__6115 (
            .O(N__32011),
            .I(\u1.DMA_control.readDfw_12 ));
    Odrv4 I__6114 (
            .O(N__32008),
            .I(\u1.DMA_control.readDfw_12 ));
    Odrv4 I__6113 (
            .O(N__32003),
            .I(\u1.DMA_control.readDfw_12 ));
    InMux I__6112 (
            .O(N__31990),
            .I(N__31987));
    LocalMux I__6111 (
            .O(N__31987),
            .I(N__31984));
    Span4Mux_v I__6110 (
            .O(N__31984),
            .I(N__31981));
    Span4Mux_v I__6109 (
            .O(N__31981),
            .I(N__31978));
    Span4Mux_h I__6108 (
            .O(N__31978),
            .I(N__31975));
    Odrv4 I__6107 (
            .O(N__31975),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_28 ));
    InMux I__6106 (
            .O(N__31972),
            .I(N__31969));
    LocalMux I__6105 (
            .O(N__31969),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_5 ));
    InMux I__6104 (
            .O(N__31966),
            .I(N__31963));
    LocalMux I__6103 (
            .O(N__31963),
            .I(N__31960));
    Span4Mux_v I__6102 (
            .O(N__31960),
            .I(N__31957));
    Span4Mux_v I__6101 (
            .O(N__31957),
            .I(N__31954));
    Odrv4 I__6100 (
            .O(N__31954),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_6 ));
    InMux I__6099 (
            .O(N__31951),
            .I(N__31948));
    LocalMux I__6098 (
            .O(N__31948),
            .I(N__31945));
    Span4Mux_v I__6097 (
            .O(N__31945),
            .I(N__31942));
    Odrv4 I__6096 (
            .O(N__31942),
            .I(\u0.dat_o_0_2_5 ));
    CascadeMux I__6095 (
            .O(N__31939),
            .I(\u0.dat_o_0_1Z0Z_5_cascade_ ));
    InMux I__6094 (
            .O(N__31936),
            .I(N__31933));
    LocalMux I__6093 (
            .O(N__31933),
            .I(\u0.dat_o_0_3_5 ));
    IoInMux I__6092 (
            .O(N__31930),
            .I(N__31927));
    LocalMux I__6091 (
            .O(N__31927),
            .I(N__31924));
    IoSpan4Mux I__6090 (
            .O(N__31924),
            .I(N__31921));
    Sp12to4 I__6089 (
            .O(N__31921),
            .I(N__31918));
    Span12Mux_s9_v I__6088 (
            .O(N__31918),
            .I(N__31915));
    Span12Mux_h I__6087 (
            .O(N__31915),
            .I(N__31912));
    Span12Mux_v I__6086 (
            .O(N__31912),
            .I(N__31909));
    Odrv12 I__6085 (
            .O(N__31909),
            .I(wb_dat_o_c_5));
    CascadeMux I__6084 (
            .O(N__31906),
            .I(N__31903));
    InMux I__6083 (
            .O(N__31903),
            .I(N__31900));
    LocalMux I__6082 (
            .O(N__31900),
            .I(N__31896));
    InMux I__6081 (
            .O(N__31899),
            .I(N__31893));
    Span4Mux_h I__6080 (
            .O(N__31896),
            .I(N__31890));
    LocalMux I__6079 (
            .O(N__31893),
            .I(N__31887));
    Sp12to4 I__6078 (
            .O(N__31890),
            .I(N__31884));
    Span4Mux_h I__6077 (
            .O(N__31887),
            .I(N__31881));
    Odrv12 I__6076 (
            .O(N__31884),
            .I(PIO_dport1_T1_5));
    Odrv4 I__6075 (
            .O(N__31881),
            .I(PIO_dport1_T1_5));
    InMux I__6074 (
            .O(N__31876),
            .I(N__31873));
    LocalMux I__6073 (
            .O(N__31873),
            .I(\u0.dat_o_0_0_5 ));
    InMux I__6072 (
            .O(N__31870),
            .I(N__31867));
    LocalMux I__6071 (
            .O(N__31867),
            .I(N__31864));
    Span4Mux_v I__6070 (
            .O(N__31864),
            .I(N__31859));
    InMux I__6069 (
            .O(N__31863),
            .I(N__31854));
    InMux I__6068 (
            .O(N__31862),
            .I(N__31854));
    Span4Mux_h I__6067 (
            .O(N__31859),
            .I(N__31849));
    LocalMux I__6066 (
            .O(N__31854),
            .I(N__31849));
    Sp12to4 I__6065 (
            .O(N__31849),
            .I(N__31846));
    Span12Mux_v I__6064 (
            .O(N__31846),
            .I(N__31843));
    Odrv12 I__6063 (
            .O(N__31843),
            .I(dd_pad_i_c_5));
    InMux I__6062 (
            .O(N__31840),
            .I(N__31837));
    LocalMux I__6061 (
            .O(N__31837),
            .I(PIOq_5));
    InMux I__6060 (
            .O(N__31834),
            .I(N__31831));
    LocalMux I__6059 (
            .O(N__31831),
            .I(N__31828));
    Span12Mux_s7_h I__6058 (
            .O(N__31828),
            .I(N__31825));
    Odrv12 I__6057 (
            .O(N__31825),
            .I(\u1.DMA_control.Tm_3 ));
    InMux I__6056 (
            .O(N__31822),
            .I(N__31819));
    LocalMux I__6055 (
            .O(N__31819),
            .I(N__31816));
    Span12Mux_s6_h I__6054 (
            .O(N__31816),
            .I(N__31813));
    Odrv12 I__6053 (
            .O(N__31813),
            .I(\u1.DMA_control.Tm_4 ));
    InMux I__6052 (
            .O(N__31810),
            .I(N__31807));
    LocalMux I__6051 (
            .O(N__31807),
            .I(N__31804));
    Sp12to4 I__6050 (
            .O(N__31804),
            .I(N__31801));
    Span12Mux_s5_h I__6049 (
            .O(N__31801),
            .I(N__31798));
    Odrv12 I__6048 (
            .O(N__31798),
            .I(\u1.DMA_control.Tm_5 ));
    InMux I__6047 (
            .O(N__31795),
            .I(N__31792));
    LocalMux I__6046 (
            .O(N__31792),
            .I(N__31789));
    Sp12to4 I__6045 (
            .O(N__31789),
            .I(N__31786));
    Span12Mux_s4_h I__6044 (
            .O(N__31786),
            .I(N__31783));
    Odrv12 I__6043 (
            .O(N__31783),
            .I(\u1.DMA_control.Tm_6 ));
    InMux I__6042 (
            .O(N__31780),
            .I(N__31777));
    LocalMux I__6041 (
            .O(N__31777),
            .I(N__31774));
    Span4Mux_v I__6040 (
            .O(N__31774),
            .I(N__31771));
    Odrv4 I__6039 (
            .O(N__31771),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_5 ));
    InMux I__6038 (
            .O(N__31768),
            .I(N__31765));
    LocalMux I__6037 (
            .O(N__31765),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI07CMZ0Z_5 ));
    InMux I__6036 (
            .O(N__31762),
            .I(N__31758));
    CascadeMux I__6035 (
            .O(N__31761),
            .I(N__31755));
    LocalMux I__6034 (
            .O(N__31758),
            .I(N__31752));
    InMux I__6033 (
            .O(N__31755),
            .I(N__31749));
    Span4Mux_h I__6032 (
            .O(N__31752),
            .I(N__31746));
    LocalMux I__6031 (
            .O(N__31749),
            .I(N__31743));
    Span4Mux_v I__6030 (
            .O(N__31746),
            .I(N__31740));
    Odrv12 I__6029 (
            .O(N__31743),
            .I(DMA_dev1_Tm_1));
    Odrv4 I__6028 (
            .O(N__31740),
            .I(DMA_dev1_Tm_1));
    InMux I__6027 (
            .O(N__31735),
            .I(N__31732));
    LocalMux I__6026 (
            .O(N__31732),
            .I(N__31728));
    InMux I__6025 (
            .O(N__31731),
            .I(N__31725));
    Span4Mux_h I__6024 (
            .O(N__31728),
            .I(N__31720));
    LocalMux I__6023 (
            .O(N__31725),
            .I(N__31720));
    Span4Mux_v I__6022 (
            .O(N__31720),
            .I(N__31717));
    Odrv4 I__6021 (
            .O(N__31717),
            .I(PIO_dport0_T1_1));
    CascadeMux I__6020 (
            .O(N__31714),
            .I(N__31711));
    InMux I__6019 (
            .O(N__31711),
            .I(N__31708));
    LocalMux I__6018 (
            .O(N__31708),
            .I(N__31705));
    Span4Mux_h I__6017 (
            .O(N__31705),
            .I(N__31702));
    Span4Mux_h I__6016 (
            .O(N__31702),
            .I(N__31698));
    InMux I__6015 (
            .O(N__31701),
            .I(N__31695));
    Span4Mux_v I__6014 (
            .O(N__31698),
            .I(N__31690));
    LocalMux I__6013 (
            .O(N__31695),
            .I(N__31690));
    Span4Mux_h I__6012 (
            .O(N__31690),
            .I(N__31687));
    Odrv4 I__6011 (
            .O(N__31687),
            .I(PIO_dport0_T1_2));
    InMux I__6010 (
            .O(N__31684),
            .I(N__31680));
    InMux I__6009 (
            .O(N__31683),
            .I(N__31677));
    LocalMux I__6008 (
            .O(N__31680),
            .I(N__31674));
    LocalMux I__6007 (
            .O(N__31677),
            .I(N__31671));
    Span12Mux_s6_h I__6006 (
            .O(N__31674),
            .I(N__31668));
    Odrv12 I__6005 (
            .O(N__31671),
            .I(DMA_dev1_Tm_2));
    Odrv12 I__6004 (
            .O(N__31668),
            .I(DMA_dev1_Tm_2));
    InMux I__6003 (
            .O(N__31663),
            .I(N__31660));
    LocalMux I__6002 (
            .O(N__31660),
            .I(N__31657));
    Span4Mux_v I__6001 (
            .O(N__31657),
            .I(N__31654));
    Odrv4 I__6000 (
            .O(N__31654),
            .I(\u0.dat_o_0_0_3_2 ));
    InMux I__5999 (
            .O(N__31651),
            .I(N__31648));
    LocalMux I__5998 (
            .O(N__31648),
            .I(N__31644));
    InMux I__5997 (
            .O(N__31647),
            .I(N__31641));
    Span4Mux_v I__5996 (
            .O(N__31644),
            .I(N__31638));
    LocalMux I__5995 (
            .O(N__31641),
            .I(N__31635));
    Odrv4 I__5994 (
            .O(N__31638),
            .I(PIO_dport0_T1_3));
    Odrv12 I__5993 (
            .O(N__31635),
            .I(PIO_dport0_T1_3));
    InMux I__5992 (
            .O(N__31630),
            .I(N__31627));
    LocalMux I__5991 (
            .O(N__31627),
            .I(N__31624));
    Span4Mux_h I__5990 (
            .O(N__31624),
            .I(N__31621));
    Span4Mux_h I__5989 (
            .O(N__31621),
            .I(N__31618));
    Odrv4 I__5988 (
            .O(N__31618),
            .I(\u1.DMA_control.Td_6 ));
    InMux I__5987 (
            .O(N__31615),
            .I(N__31612));
    LocalMux I__5986 (
            .O(N__31612),
            .I(N__31609));
    Span4Mux_h I__5985 (
            .O(N__31609),
            .I(N__31606));
    Odrv4 I__5984 (
            .O(N__31606),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNI87TNZ0Z_5 ));
    InMux I__5983 (
            .O(N__31603),
            .I(N__31600));
    LocalMux I__5982 (
            .O(N__31600),
            .I(N__31597));
    Span4Mux_v I__5981 (
            .O(N__31597),
            .I(N__31594));
    Odrv4 I__5980 (
            .O(N__31594),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_5 ));
    InMux I__5979 (
            .O(N__31591),
            .I(N__31588));
    LocalMux I__5978 (
            .O(N__31588),
            .I(N__31585));
    Span4Mux_v I__5977 (
            .O(N__31585),
            .I(N__31582));
    Span4Mux_v I__5976 (
            .O(N__31582),
            .I(N__31579));
    Sp12to4 I__5975 (
            .O(N__31579),
            .I(N__31576));
    Odrv12 I__5974 (
            .O(N__31576),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI4N4NZ0Z_5 ));
    InMux I__5973 (
            .O(N__31573),
            .I(N__31570));
    LocalMux I__5972 (
            .O(N__31570),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNINMOD1Z0Z_5 ));
    CascadeMux I__5971 (
            .O(N__31567),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIM8OK1Z0Z_2_cascade_ ));
    CascadeMux I__5970 (
            .O(N__31564),
            .I(DMAq_5_cascade_));
    InMux I__5969 (
            .O(N__31561),
            .I(N__31557));
    InMux I__5968 (
            .O(N__31560),
            .I(N__31554));
    LocalMux I__5967 (
            .O(N__31557),
            .I(N__31551));
    LocalMux I__5966 (
            .O(N__31554),
            .I(N__31548));
    Span4Mux_h I__5965 (
            .O(N__31551),
            .I(N__31545));
    Span4Mux_v I__5964 (
            .O(N__31548),
            .I(N__31540));
    Span4Mux_h I__5963 (
            .O(N__31545),
            .I(N__31540));
    Odrv4 I__5962 (
            .O(N__31540),
            .I(DMA_dev1_Td_4));
    InMux I__5961 (
            .O(N__31537),
            .I(N__31534));
    LocalMux I__5960 (
            .O(N__31534),
            .I(N__31530));
    InMux I__5959 (
            .O(N__31533),
            .I(N__31527));
    Span4Mux_v I__5958 (
            .O(N__31530),
            .I(N__31524));
    LocalMux I__5957 (
            .O(N__31527),
            .I(N__31521));
    Span4Mux_v I__5956 (
            .O(N__31524),
            .I(N__31516));
    Span4Mux_h I__5955 (
            .O(N__31521),
            .I(N__31516));
    Span4Mux_h I__5954 (
            .O(N__31516),
            .I(N__31513));
    Span4Mux_v I__5953 (
            .O(N__31513),
            .I(N__31510));
    Odrv4 I__5952 (
            .O(N__31510),
            .I(DMA_dev1_Td_5));
    InMux I__5951 (
            .O(N__31507),
            .I(N__31503));
    InMux I__5950 (
            .O(N__31506),
            .I(N__31500));
    LocalMux I__5949 (
            .O(N__31503),
            .I(N__31497));
    LocalMux I__5948 (
            .O(N__31500),
            .I(N__31494));
    Span4Mux_h I__5947 (
            .O(N__31497),
            .I(N__31491));
    Span4Mux_v I__5946 (
            .O(N__31494),
            .I(N__31488));
    Odrv4 I__5945 (
            .O(N__31491),
            .I(PIO_dport1_T2_5));
    Odrv4 I__5944 (
            .O(N__31488),
            .I(PIO_dport1_T2_5));
    InMux I__5943 (
            .O(N__31483),
            .I(N__31479));
    InMux I__5942 (
            .O(N__31482),
            .I(N__31476));
    LocalMux I__5941 (
            .O(N__31479),
            .I(N__31473));
    LocalMux I__5940 (
            .O(N__31476),
            .I(N__31470));
    Span4Mux_h I__5939 (
            .O(N__31473),
            .I(N__31467));
    Odrv4 I__5938 (
            .O(N__31470),
            .I(PIO_dport1_T2_7));
    Odrv4 I__5937 (
            .O(N__31467),
            .I(PIO_dport1_T2_7));
    InMux I__5936 (
            .O(N__31462),
            .I(N__31459));
    LocalMux I__5935 (
            .O(N__31459),
            .I(N__31456));
    Span4Mux_h I__5934 (
            .O(N__31456),
            .I(N__31453));
    Span4Mux_h I__5933 (
            .O(N__31453),
            .I(N__31450));
    Odrv4 I__5932 (
            .O(N__31450),
            .I(\u0.dat_o_0_0_3_8 ));
    InMux I__5931 (
            .O(N__31447),
            .I(N__31444));
    LocalMux I__5930 (
            .O(N__31444),
            .I(N__31439));
    InMux I__5929 (
            .O(N__31443),
            .I(N__31436));
    InMux I__5928 (
            .O(N__31442),
            .I(N__31433));
    Span4Mux_h I__5927 (
            .O(N__31439),
            .I(N__31430));
    LocalMux I__5926 (
            .O(N__31436),
            .I(N__31426));
    LocalMux I__5925 (
            .O(N__31433),
            .I(N__31422));
    Span4Mux_h I__5924 (
            .O(N__31430),
            .I(N__31419));
    InMux I__5923 (
            .O(N__31429),
            .I(N__31416));
    Span4Mux_v I__5922 (
            .O(N__31426),
            .I(N__31413));
    InMux I__5921 (
            .O(N__31425),
            .I(N__31410));
    Span4Mux_v I__5920 (
            .O(N__31422),
            .I(N__31407));
    Odrv4 I__5919 (
            .O(N__31419),
            .I(DMATxFull));
    LocalMux I__5918 (
            .O(N__31416),
            .I(DMATxFull));
    Odrv4 I__5917 (
            .O(N__31413),
            .I(DMATxFull));
    LocalMux I__5916 (
            .O(N__31410),
            .I(DMATxFull));
    Odrv4 I__5915 (
            .O(N__31407),
            .I(DMATxFull));
    CascadeMux I__5914 (
            .O(N__31396),
            .I(N__31392));
    InMux I__5913 (
            .O(N__31395),
            .I(N__31389));
    InMux I__5912 (
            .O(N__31392),
            .I(N__31386));
    LocalMux I__5911 (
            .O(N__31389),
            .I(N__31383));
    LocalMux I__5910 (
            .O(N__31386),
            .I(N__31380));
    Odrv4 I__5909 (
            .O(N__31383),
            .I(PIO_dport1_T2_1));
    Odrv4 I__5908 (
            .O(N__31380),
            .I(PIO_dport1_T2_1));
    CascadeMux I__5907 (
            .O(N__31375),
            .I(N__31372));
    InMux I__5906 (
            .O(N__31372),
            .I(N__31369));
    LocalMux I__5905 (
            .O(N__31369),
            .I(N__31366));
    Span4Mux_v I__5904 (
            .O(N__31366),
            .I(N__31362));
    CascadeMux I__5903 (
            .O(N__31365),
            .I(N__31359));
    Span4Mux_h I__5902 (
            .O(N__31362),
            .I(N__31356));
    InMux I__5901 (
            .O(N__31359),
            .I(N__31353));
    Odrv4 I__5900 (
            .O(N__31356),
            .I(DMA_dev1_Td_7));
    LocalMux I__5899 (
            .O(N__31353),
            .I(DMA_dev1_Td_7));
    InMux I__5898 (
            .O(N__31348),
            .I(N__31345));
    LocalMux I__5897 (
            .O(N__31345),
            .I(N__31342));
    Span4Mux_h I__5896 (
            .O(N__31342),
            .I(N__31339));
    Span4Mux_v I__5895 (
            .O(N__31339),
            .I(N__31336));
    Odrv4 I__5894 (
            .O(N__31336),
            .I(\u0.dat_o_0_0_0_15 ));
    InMux I__5893 (
            .O(N__31333),
            .I(N__31330));
    LocalMux I__5892 (
            .O(N__31330),
            .I(N__31327));
    Span4Mux_v I__5891 (
            .O(N__31327),
            .I(N__31323));
    InMux I__5890 (
            .O(N__31326),
            .I(N__31320));
    Span4Mux_h I__5889 (
            .O(N__31323),
            .I(N__31317));
    LocalMux I__5888 (
            .O(N__31320),
            .I(N__31314));
    Span4Mux_h I__5887 (
            .O(N__31317),
            .I(N__31311));
    Odrv12 I__5886 (
            .O(N__31314),
            .I(DMA_dev1_Td_0));
    Odrv4 I__5885 (
            .O(N__31311),
            .I(DMA_dev1_Td_0));
    InMux I__5884 (
            .O(N__31306),
            .I(N__31303));
    LocalMux I__5883 (
            .O(N__31303),
            .I(N__31299));
    InMux I__5882 (
            .O(N__31302),
            .I(N__31296));
    Span4Mux_h I__5881 (
            .O(N__31299),
            .I(N__31293));
    LocalMux I__5880 (
            .O(N__31296),
            .I(DMA_dev1_Td_1));
    Odrv4 I__5879 (
            .O(N__31293),
            .I(DMA_dev1_Td_1));
    InMux I__5878 (
            .O(N__31288),
            .I(N__31284));
    InMux I__5877 (
            .O(N__31287),
            .I(N__31281));
    LocalMux I__5876 (
            .O(N__31284),
            .I(N__31278));
    LocalMux I__5875 (
            .O(N__31281),
            .I(N__31275));
    Span4Mux_v I__5874 (
            .O(N__31278),
            .I(N__31272));
    Span4Mux_v I__5873 (
            .O(N__31275),
            .I(N__31269));
    Span4Mux_h I__5872 (
            .O(N__31272),
            .I(N__31266));
    Odrv4 I__5871 (
            .O(N__31269),
            .I(DMA_dev1_Td_3));
    Odrv4 I__5870 (
            .O(N__31266),
            .I(DMA_dev1_Td_3));
    InMux I__5869 (
            .O(N__31261),
            .I(N__31258));
    LocalMux I__5868 (
            .O(N__31258),
            .I(N__31255));
    Odrv4 I__5867 (
            .O(N__31255),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_6 ));
    InMux I__5866 (
            .O(N__31252),
            .I(N__31249));
    LocalMux I__5865 (
            .O(N__31249),
            .I(N__31246));
    Span4Mux_s2_v I__5864 (
            .O(N__31246),
            .I(N__31243));
    Odrv4 I__5863 (
            .O(N__31243),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_6 ));
    CascadeMux I__5862 (
            .O(N__31240),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI6P4NZ0Z_6_cascade_ ));
    InMux I__5861 (
            .O(N__31237),
            .I(N__31234));
    LocalMux I__5860 (
            .O(N__31234),
            .I(N__31231));
    Span12Mux_s11_h I__5859 (
            .O(N__31231),
            .I(N__31228));
    Odrv12 I__5858 (
            .O(N__31228),
            .I(iQ_RNIQCOK1_2));
    InMux I__5857 (
            .O(N__31225),
            .I(N__31222));
    LocalMux I__5856 (
            .O(N__31222),
            .I(N__31219));
    Odrv12 I__5855 (
            .O(N__31219),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_6 ));
    InMux I__5854 (
            .O(N__31216),
            .I(N__31213));
    LocalMux I__5853 (
            .O(N__31213),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI29CMZ0Z_6 ));
    InMux I__5852 (
            .O(N__31210),
            .I(N__31207));
    LocalMux I__5851 (
            .O(N__31207),
            .I(N__31203));
    CascadeMux I__5850 (
            .O(N__31206),
            .I(N__31200));
    Span4Mux_v I__5849 (
            .O(N__31203),
            .I(N__31197));
    InMux I__5848 (
            .O(N__31200),
            .I(N__31194));
    Sp12to4 I__5847 (
            .O(N__31197),
            .I(N__31191));
    LocalMux I__5846 (
            .O(N__31194),
            .I(N__31188));
    Span12Mux_h I__5845 (
            .O(N__31191),
            .I(N__31185));
    Odrv4 I__5844 (
            .O(N__31188),
            .I(DMA_dev0_Tm_2));
    Odrv12 I__5843 (
            .O(N__31185),
            .I(DMA_dev0_Tm_2));
    InMux I__5842 (
            .O(N__31180),
            .I(N__31177));
    LocalMux I__5841 (
            .O(N__31177),
            .I(N__31173));
    InMux I__5840 (
            .O(N__31176),
            .I(N__31170));
    Span4Mux_v I__5839 (
            .O(N__31173),
            .I(N__31167));
    LocalMux I__5838 (
            .O(N__31170),
            .I(N__31164));
    Span4Mux_v I__5837 (
            .O(N__31167),
            .I(N__31161));
    Span4Mux_h I__5836 (
            .O(N__31164),
            .I(N__31158));
    Odrv4 I__5835 (
            .O(N__31161),
            .I(PIO_cmdport_T1_5));
    Odrv4 I__5834 (
            .O(N__31158),
            .I(PIO_cmdport_T1_5));
    InMux I__5833 (
            .O(N__31153),
            .I(N__31150));
    LocalMux I__5832 (
            .O(N__31150),
            .I(N__31147));
    Span12Mux_s8_h I__5831 (
            .O(N__31147),
            .I(N__31144));
    Odrv12 I__5830 (
            .O(N__31144),
            .I(\u0.dat_o_0_0_0_8 ));
    InMux I__5829 (
            .O(N__31141),
            .I(N__31138));
    LocalMux I__5828 (
            .O(N__31138),
            .I(N__31135));
    Span4Mux_s2_v I__5827 (
            .O(N__31135),
            .I(N__31132));
    Span4Mux_v I__5826 (
            .O(N__31132),
            .I(N__31129));
    Odrv4 I__5825 (
            .O(N__31129),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_28 ));
    CascadeMux I__5824 (
            .O(N__31126),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIA31RZ0Z_28_cascade_ ));
    InMux I__5823 (
            .O(N__31123),
            .I(N__31120));
    LocalMux I__5822 (
            .O(N__31120),
            .I(N__31117));
    Span4Mux_h I__5821 (
            .O(N__31117),
            .I(N__31114));
    Odrv4 I__5820 (
            .O(N__31114),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_28 ));
    InMux I__5819 (
            .O(N__31111),
            .I(N__31108));
    LocalMux I__5818 (
            .O(N__31108),
            .I(N__31105));
    Span4Mux_v I__5817 (
            .O(N__31105),
            .I(N__31102));
    Odrv4 I__5816 (
            .O(N__31102),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_28 ));
    CascadeMux I__5815 (
            .O(N__31099),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_N_1197_cascade_ ));
    CascadeMux I__5814 (
            .O(N__31096),
            .I(u1_DMA_control_gen_DMAbuf_Rxbuf_mem_N_1229_cascade_));
    InMux I__5813 (
            .O(N__31093),
            .I(N__31090));
    LocalMux I__5812 (
            .O(N__31090),
            .I(u1_DMA_control_gen_DMAbuf_Rxbuf_mem_N_1165));
    InMux I__5811 (
            .O(N__31087),
            .I(N__31084));
    LocalMux I__5810 (
            .O(N__31084),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_28 ));
    InMux I__5809 (
            .O(N__31081),
            .I(N__31078));
    LocalMux I__5808 (
            .O(N__31078),
            .I(N__31075));
    Span4Mux_s2_v I__5807 (
            .O(N__31075),
            .I(N__31072));
    Odrv4 I__5806 (
            .O(N__31072),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_28 ));
    InMux I__5805 (
            .O(N__31069),
            .I(N__31066));
    LocalMux I__5804 (
            .O(N__31066),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIEN9KZ0Z_28 ));
    InMux I__5803 (
            .O(N__31063),
            .I(N__31060));
    LocalMux I__5802 (
            .O(N__31060),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_28 ));
    InMux I__5801 (
            .O(N__31057),
            .I(N__31054));
    LocalMux I__5800 (
            .O(N__31054),
            .I(N__31051));
    Span12Mux_v I__5799 (
            .O(N__31051),
            .I(N__31048));
    Odrv12 I__5798 (
            .O(N__31048),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_12 ));
    InMux I__5797 (
            .O(N__31045),
            .I(N__31042));
    LocalMux I__5796 (
            .O(N__31042),
            .I(N__31039));
    Span4Mux_v I__5795 (
            .O(N__31039),
            .I(N__31036));
    Odrv4 I__5794 (
            .O(N__31036),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_20 ));
    InMux I__5793 (
            .O(N__31033),
            .I(N__31030));
    LocalMux I__5792 (
            .O(N__31030),
            .I(N__31027));
    Span4Mux_v I__5791 (
            .O(N__31027),
            .I(N__31024));
    Span4Mux_v I__5790 (
            .O(N__31024),
            .I(N__31021));
    Odrv4 I__5789 (
            .O(N__31021),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIU69KZ0Z_20 ));
    InMux I__5788 (
            .O(N__31018),
            .I(N__31014));
    InMux I__5787 (
            .O(N__31017),
            .I(N__31011));
    LocalMux I__5786 (
            .O(N__31014),
            .I(N__30996));
    LocalMux I__5785 (
            .O(N__31011),
            .I(N__30996));
    InMux I__5784 (
            .O(N__31010),
            .I(N__30993));
    InMux I__5783 (
            .O(N__31009),
            .I(N__30990));
    InMux I__5782 (
            .O(N__31008),
            .I(N__30985));
    InMux I__5781 (
            .O(N__31007),
            .I(N__30985));
    InMux I__5780 (
            .O(N__31006),
            .I(N__30980));
    InMux I__5779 (
            .O(N__31005),
            .I(N__30980));
    InMux I__5778 (
            .O(N__31004),
            .I(N__30976));
    InMux I__5777 (
            .O(N__31003),
            .I(N__30973));
    InMux I__5776 (
            .O(N__31002),
            .I(N__30968));
    InMux I__5775 (
            .O(N__31001),
            .I(N__30968));
    Span4Mux_v I__5774 (
            .O(N__30996),
            .I(N__30959));
    LocalMux I__5773 (
            .O(N__30993),
            .I(N__30959));
    LocalMux I__5772 (
            .O(N__30990),
            .I(N__30959));
    LocalMux I__5771 (
            .O(N__30985),
            .I(N__30959));
    LocalMux I__5770 (
            .O(N__30980),
            .I(N__30956));
    InMux I__5769 (
            .O(N__30979),
            .I(N__30951));
    LocalMux I__5768 (
            .O(N__30976),
            .I(N__30946));
    LocalMux I__5767 (
            .O(N__30973),
            .I(N__30946));
    LocalMux I__5766 (
            .O(N__30968),
            .I(N__30943));
    Span4Mux_v I__5765 (
            .O(N__30959),
            .I(N__30938));
    Span4Mux_h I__5764 (
            .O(N__30956),
            .I(N__30938));
    InMux I__5763 (
            .O(N__30955),
            .I(N__30933));
    InMux I__5762 (
            .O(N__30954),
            .I(N__30933));
    LocalMux I__5761 (
            .O(N__30951),
            .I(\u1.DMA_control.readDlw_4 ));
    Odrv12 I__5760 (
            .O(N__30946),
            .I(\u1.DMA_control.readDlw_4 ));
    Odrv4 I__5759 (
            .O(N__30943),
            .I(\u1.DMA_control.readDlw_4 ));
    Odrv4 I__5758 (
            .O(N__30938),
            .I(\u1.DMA_control.readDlw_4 ));
    LocalMux I__5757 (
            .O(N__30933),
            .I(\u1.DMA_control.readDlw_4 ));
    InMux I__5756 (
            .O(N__30922),
            .I(N__30918));
    InMux I__5755 (
            .O(N__30921),
            .I(N__30915));
    LocalMux I__5754 (
            .O(N__30918),
            .I(N__30906));
    LocalMux I__5753 (
            .O(N__30915),
            .I(N__30906));
    InMux I__5752 (
            .O(N__30914),
            .I(N__30901));
    InMux I__5751 (
            .O(N__30913),
            .I(N__30901));
    InMux I__5750 (
            .O(N__30912),
            .I(N__30896));
    InMux I__5749 (
            .O(N__30911),
            .I(N__30893));
    Span4Mux_v I__5748 (
            .O(N__30906),
            .I(N__30884));
    LocalMux I__5747 (
            .O(N__30901),
            .I(N__30884));
    InMux I__5746 (
            .O(N__30900),
            .I(N__30879));
    InMux I__5745 (
            .O(N__30899),
            .I(N__30879));
    LocalMux I__5744 (
            .O(N__30896),
            .I(N__30874));
    LocalMux I__5743 (
            .O(N__30893),
            .I(N__30874));
    InMux I__5742 (
            .O(N__30892),
            .I(N__30869));
    InMux I__5741 (
            .O(N__30891),
            .I(N__30869));
    InMux I__5740 (
            .O(N__30890),
            .I(N__30866));
    InMux I__5739 (
            .O(N__30889),
            .I(N__30863));
    Span4Mux_v I__5738 (
            .O(N__30884),
            .I(N__30858));
    LocalMux I__5737 (
            .O(N__30879),
            .I(N__30855));
    Span4Mux_h I__5736 (
            .O(N__30874),
            .I(N__30852));
    LocalMux I__5735 (
            .O(N__30869),
            .I(N__30849));
    LocalMux I__5734 (
            .O(N__30866),
            .I(N__30844));
    LocalMux I__5733 (
            .O(N__30863),
            .I(N__30844));
    InMux I__5732 (
            .O(N__30862),
            .I(N__30841));
    InMux I__5731 (
            .O(N__30861),
            .I(N__30838));
    Odrv4 I__5730 (
            .O(N__30858),
            .I(\u1.DMA_control.readDfw_4 ));
    Odrv12 I__5729 (
            .O(N__30855),
            .I(\u1.DMA_control.readDfw_4 ));
    Odrv4 I__5728 (
            .O(N__30852),
            .I(\u1.DMA_control.readDfw_4 ));
    Odrv4 I__5727 (
            .O(N__30849),
            .I(\u1.DMA_control.readDfw_4 ));
    Odrv4 I__5726 (
            .O(N__30844),
            .I(\u1.DMA_control.readDfw_4 ));
    LocalMux I__5725 (
            .O(N__30841),
            .I(\u1.DMA_control.readDfw_4 ));
    LocalMux I__5724 (
            .O(N__30838),
            .I(\u1.DMA_control.readDfw_4 ));
    InMux I__5723 (
            .O(N__30823),
            .I(N__30820));
    LocalMux I__5722 (
            .O(N__30820),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_20 ));
    CEMux I__5721 (
            .O(N__30817),
            .I(N__30814));
    LocalMux I__5720 (
            .O(N__30814),
            .I(N__30809));
    CEMux I__5719 (
            .O(N__30813),
            .I(N__30803));
    CEMux I__5718 (
            .O(N__30812),
            .I(N__30800));
    Span4Mux_v I__5717 (
            .O(N__30809),
            .I(N__30797));
    CEMux I__5716 (
            .O(N__30808),
            .I(N__30794));
    CEMux I__5715 (
            .O(N__30807),
            .I(N__30791));
    CEMux I__5714 (
            .O(N__30806),
            .I(N__30788));
    LocalMux I__5713 (
            .O(N__30803),
            .I(N__30784));
    LocalMux I__5712 (
            .O(N__30800),
            .I(N__30781));
    Span4Mux_h I__5711 (
            .O(N__30797),
            .I(N__30776));
    LocalMux I__5710 (
            .O(N__30794),
            .I(N__30776));
    LocalMux I__5709 (
            .O(N__30791),
            .I(N__30773));
    LocalMux I__5708 (
            .O(N__30788),
            .I(N__30770));
    CEMux I__5707 (
            .O(N__30787),
            .I(N__30767));
    Span4Mux_h I__5706 (
            .O(N__30784),
            .I(N__30761));
    Span4Mux_s3_v I__5705 (
            .O(N__30781),
            .I(N__30761));
    Span4Mux_v I__5704 (
            .O(N__30776),
            .I(N__30758));
    Span4Mux_v I__5703 (
            .O(N__30773),
            .I(N__30755));
    Span4Mux_h I__5702 (
            .O(N__30770),
            .I(N__30750));
    LocalMux I__5701 (
            .O(N__30767),
            .I(N__30750));
    CEMux I__5700 (
            .O(N__30766),
            .I(N__30747));
    Span4Mux_h I__5699 (
            .O(N__30761),
            .I(N__30744));
    Span4Mux_h I__5698 (
            .O(N__30758),
            .I(N__30739));
    Span4Mux_h I__5697 (
            .O(N__30755),
            .I(N__30739));
    Span4Mux_h I__5696 (
            .O(N__30750),
            .I(N__30736));
    LocalMux I__5695 (
            .O(N__30747),
            .I(N__30733));
    Odrv4 I__5694 (
            .O(N__30744),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_awe2 ));
    Odrv4 I__5693 (
            .O(N__30739),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_awe2 ));
    Odrv4 I__5692 (
            .O(N__30736),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_awe2 ));
    Odrv12 I__5691 (
            .O(N__30733),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_awe2 ));
    InMux I__5690 (
            .O(N__30724),
            .I(N__30721));
    LocalMux I__5689 (
            .O(N__30721),
            .I(N__30718));
    Odrv12 I__5688 (
            .O(N__30718),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_7 ));
    InMux I__5687 (
            .O(N__30715),
            .I(N__30712));
    LocalMux I__5686 (
            .O(N__30712),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_7 ));
    InMux I__5685 (
            .O(N__30709),
            .I(N__30706));
    LocalMux I__5684 (
            .O(N__30706),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_26 ));
    InMux I__5683 (
            .O(N__30703),
            .I(N__30700));
    LocalMux I__5682 (
            .O(N__30700),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_26 ));
    InMux I__5681 (
            .O(N__30697),
            .I(N__30694));
    LocalMux I__5680 (
            .O(N__30694),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_26 ));
    InMux I__5679 (
            .O(N__30691),
            .I(N__30688));
    LocalMux I__5678 (
            .O(N__30688),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIAJ9KZ0Z_26 ));
    CascadeMux I__5677 (
            .O(N__30685),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI6V0RZ0Z_26_cascade_ ));
    InMux I__5676 (
            .O(N__30682),
            .I(N__30679));
    LocalMux I__5675 (
            .O(N__30679),
            .I(N__30676));
    Odrv4 I__5674 (
            .O(N__30676),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI2THM1Z0Z_2 ));
    CascadeMux I__5673 (
            .O(N__30673),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIE7ITZ0Z_26_cascade_ ));
    CascadeMux I__5672 (
            .O(N__30670),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIG8E71Z0Z_26_cascade_ ));
    InMux I__5671 (
            .O(N__30667),
            .I(N__30664));
    LocalMux I__5670 (
            .O(N__30664),
            .I(N__30661));
    Span4Mux_v I__5669 (
            .O(N__30661),
            .I(N__30658));
    Sp12to4 I__5668 (
            .O(N__30658),
            .I(N__30655));
    Odrv12 I__5667 (
            .O(N__30655),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_23 ));
    InMux I__5666 (
            .O(N__30652),
            .I(N__30649));
    LocalMux I__5665 (
            .O(N__30649),
            .I(N__30646));
    Span4Mux_v I__5664 (
            .O(N__30646),
            .I(N__30643));
    Odrv4 I__5663 (
            .O(N__30643),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_23 ));
    InMux I__5662 (
            .O(N__30640),
            .I(N__30637));
    LocalMux I__5661 (
            .O(N__30637),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_9 ));
    InMux I__5660 (
            .O(N__30634),
            .I(N__30631));
    LocalMux I__5659 (
            .O(N__30631),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_9 ));
    InMux I__5658 (
            .O(N__30628),
            .I(N__30625));
    LocalMux I__5657 (
            .O(N__30625),
            .I(N__30622));
    Span4Mux_v I__5656 (
            .O(N__30622),
            .I(N__30619));
    Odrv4 I__5655 (
            .O(N__30619),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_11 ));
    InMux I__5654 (
            .O(N__30616),
            .I(N__30613));
    LocalMux I__5653 (
            .O(N__30613),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_11 ));
    InMux I__5652 (
            .O(N__30610),
            .I(N__30607));
    LocalMux I__5651 (
            .O(N__30607),
            .I(N__30604));
    Odrv12 I__5650 (
            .O(N__30604),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_14 ));
    CascadeMux I__5649 (
            .O(N__30601),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI4B7KZ0Z_14_cascade_ ));
    InMux I__5648 (
            .O(N__30598),
            .I(N__30595));
    LocalMux I__5647 (
            .O(N__30595),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_14 ));
    InMux I__5646 (
            .O(N__30592),
            .I(N__30589));
    LocalMux I__5645 (
            .O(N__30589),
            .I(N__30586));
    Span4Mux_v I__5644 (
            .O(N__30586),
            .I(N__30583));
    Odrv4 I__5643 (
            .O(N__30583),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_30 ));
    InMux I__5642 (
            .O(N__30580),
            .I(N__30577));
    LocalMux I__5641 (
            .O(N__30577),
            .I(N__30574));
    Odrv4 I__5640 (
            .O(N__30574),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_26 ));
    InMux I__5639 (
            .O(N__30571),
            .I(N__30568));
    LocalMux I__5638 (
            .O(N__30568),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_26 ));
    CascadeMux I__5637 (
            .O(N__30565),
            .I(N__30562));
    InMux I__5636 (
            .O(N__30562),
            .I(N__30559));
    LocalMux I__5635 (
            .O(N__30559),
            .I(N__30556));
    Span4Mux_v I__5634 (
            .O(N__30556),
            .I(N__30553));
    Span4Mux_s3_v I__5633 (
            .O(N__30553),
            .I(N__30550));
    Odrv4 I__5632 (
            .O(N__30550),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_17 ));
    InMux I__5631 (
            .O(N__30547),
            .I(N__30544));
    LocalMux I__5630 (
            .O(N__30544),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_17 ));
    InMux I__5629 (
            .O(N__30541),
            .I(N__30538));
    LocalMux I__5628 (
            .O(N__30538),
            .I(N__30535));
    Span4Mux_h I__5627 (
            .O(N__30535),
            .I(N__30532));
    Span4Mux_v I__5626 (
            .O(N__30532),
            .I(N__30529));
    Odrv4 I__5625 (
            .O(N__30529),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_1 ));
    InMux I__5624 (
            .O(N__30526),
            .I(N__30523));
    LocalMux I__5623 (
            .O(N__30523),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_1 ));
    InMux I__5622 (
            .O(N__30520),
            .I(N__30517));
    LocalMux I__5621 (
            .O(N__30517),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_18 ));
    InMux I__5620 (
            .O(N__30514),
            .I(N__30511));
    LocalMux I__5619 (
            .O(N__30511),
            .I(N__30508));
    Span4Mux_v I__5618 (
            .O(N__30508),
            .I(N__30505));
    Sp12to4 I__5617 (
            .O(N__30505),
            .I(N__30502));
    Odrv12 I__5616 (
            .O(N__30502),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_18 ));
    CascadeMux I__5615 (
            .O(N__30499),
            .I(N__30495));
    CascadeMux I__5614 (
            .O(N__30498),
            .I(N__30488));
    InMux I__5613 (
            .O(N__30495),
            .I(N__30481));
    InMux I__5612 (
            .O(N__30494),
            .I(N__30481));
    InMux I__5611 (
            .O(N__30493),
            .I(N__30474));
    InMux I__5610 (
            .O(N__30492),
            .I(N__30474));
    InMux I__5609 (
            .O(N__30491),
            .I(N__30469));
    InMux I__5608 (
            .O(N__30488),
            .I(N__30464));
    InMux I__5607 (
            .O(N__30487),
            .I(N__30464));
    InMux I__5606 (
            .O(N__30486),
            .I(N__30461));
    LocalMux I__5605 (
            .O(N__30481),
            .I(N__30457));
    InMux I__5604 (
            .O(N__30480),
            .I(N__30454));
    InMux I__5603 (
            .O(N__30479),
            .I(N__30451));
    LocalMux I__5602 (
            .O(N__30474),
            .I(N__30448));
    InMux I__5601 (
            .O(N__30473),
            .I(N__30445));
    InMux I__5600 (
            .O(N__30472),
            .I(N__30442));
    LocalMux I__5599 (
            .O(N__30469),
            .I(N__30439));
    LocalMux I__5598 (
            .O(N__30464),
            .I(N__30434));
    LocalMux I__5597 (
            .O(N__30461),
            .I(N__30434));
    InMux I__5596 (
            .O(N__30460),
            .I(N__30429));
    Span4Mux_v I__5595 (
            .O(N__30457),
            .I(N__30426));
    LocalMux I__5594 (
            .O(N__30454),
            .I(N__30423));
    LocalMux I__5593 (
            .O(N__30451),
            .I(N__30420));
    Span4Mux_v I__5592 (
            .O(N__30448),
            .I(N__30417));
    LocalMux I__5591 (
            .O(N__30445),
            .I(N__30412));
    LocalMux I__5590 (
            .O(N__30442),
            .I(N__30412));
    Span4Mux_h I__5589 (
            .O(N__30439),
            .I(N__30407));
    Span4Mux_v I__5588 (
            .O(N__30434),
            .I(N__30407));
    InMux I__5587 (
            .O(N__30433),
            .I(N__30404));
    InMux I__5586 (
            .O(N__30432),
            .I(N__30401));
    LocalMux I__5585 (
            .O(N__30429),
            .I(N__30398));
    Span4Mux_h I__5584 (
            .O(N__30426),
            .I(N__30393));
    Span4Mux_v I__5583 (
            .O(N__30423),
            .I(N__30393));
    Span4Mux_h I__5582 (
            .O(N__30420),
            .I(N__30390));
    Sp12to4 I__5581 (
            .O(N__30417),
            .I(N__30381));
    Span12Mux_s5_v I__5580 (
            .O(N__30412),
            .I(N__30381));
    Sp12to4 I__5579 (
            .O(N__30407),
            .I(N__30381));
    LocalMux I__5578 (
            .O(N__30404),
            .I(N__30381));
    LocalMux I__5577 (
            .O(N__30401),
            .I(N__30378));
    Odrv12 I__5576 (
            .O(N__30398),
            .I(\u1.DMA_control.readDlw_2 ));
    Odrv4 I__5575 (
            .O(N__30393),
            .I(\u1.DMA_control.readDlw_2 ));
    Odrv4 I__5574 (
            .O(N__30390),
            .I(\u1.DMA_control.readDlw_2 ));
    Odrv12 I__5573 (
            .O(N__30381),
            .I(\u1.DMA_control.readDlw_2 ));
    Odrv4 I__5572 (
            .O(N__30378),
            .I(\u1.DMA_control.readDlw_2 ));
    CascadeMux I__5571 (
            .O(N__30367),
            .I(N__30364));
    InMux I__5570 (
            .O(N__30364),
            .I(N__30353));
    InMux I__5569 (
            .O(N__30363),
            .I(N__30353));
    InMux I__5568 (
            .O(N__30362),
            .I(N__30348));
    InMux I__5567 (
            .O(N__30361),
            .I(N__30348));
    InMux I__5566 (
            .O(N__30360),
            .I(N__30343));
    InMux I__5565 (
            .O(N__30359),
            .I(N__30343));
    InMux I__5564 (
            .O(N__30358),
            .I(N__30340));
    LocalMux I__5563 (
            .O(N__30353),
            .I(N__30332));
    LocalMux I__5562 (
            .O(N__30348),
            .I(N__30327));
    LocalMux I__5561 (
            .O(N__30343),
            .I(N__30327));
    LocalMux I__5560 (
            .O(N__30340),
            .I(N__30324));
    InMux I__5559 (
            .O(N__30339),
            .I(N__30321));
    InMux I__5558 (
            .O(N__30338),
            .I(N__30318));
    InMux I__5557 (
            .O(N__30337),
            .I(N__30315));
    InMux I__5556 (
            .O(N__30336),
            .I(N__30310));
    InMux I__5555 (
            .O(N__30335),
            .I(N__30310));
    Span4Mux_v I__5554 (
            .O(N__30332),
            .I(N__30306));
    Span4Mux_v I__5553 (
            .O(N__30327),
            .I(N__30299));
    Span4Mux_h I__5552 (
            .O(N__30324),
            .I(N__30299));
    LocalMux I__5551 (
            .O(N__30321),
            .I(N__30299));
    LocalMux I__5550 (
            .O(N__30318),
            .I(N__30296));
    LocalMux I__5549 (
            .O(N__30315),
            .I(N__30293));
    LocalMux I__5548 (
            .O(N__30310),
            .I(N__30290));
    InMux I__5547 (
            .O(N__30309),
            .I(N__30287));
    Span4Mux_h I__5546 (
            .O(N__30306),
            .I(N__30283));
    Span4Mux_h I__5545 (
            .O(N__30299),
            .I(N__30280));
    Span4Mux_h I__5544 (
            .O(N__30296),
            .I(N__30275));
    Span4Mux_v I__5543 (
            .O(N__30293),
            .I(N__30275));
    Span4Mux_v I__5542 (
            .O(N__30290),
            .I(N__30272));
    LocalMux I__5541 (
            .O(N__30287),
            .I(N__30269));
    InMux I__5540 (
            .O(N__30286),
            .I(N__30266));
    Span4Mux_h I__5539 (
            .O(N__30283),
            .I(N__30263));
    Span4Mux_h I__5538 (
            .O(N__30280),
            .I(N__30260));
    Span4Mux_v I__5537 (
            .O(N__30275),
            .I(N__30253));
    Span4Mux_h I__5536 (
            .O(N__30272),
            .I(N__30253));
    Span4Mux_s2_v I__5535 (
            .O(N__30269),
            .I(N__30253));
    LocalMux I__5534 (
            .O(N__30266),
            .I(N__30250));
    Odrv4 I__5533 (
            .O(N__30263),
            .I(\u1.DMA_control.readDfw_2 ));
    Odrv4 I__5532 (
            .O(N__30260),
            .I(\u1.DMA_control.readDfw_2 ));
    Odrv4 I__5531 (
            .O(N__30253),
            .I(\u1.DMA_control.readDfw_2 ));
    Odrv12 I__5530 (
            .O(N__30250),
            .I(\u1.DMA_control.readDfw_2 ));
    InMux I__5529 (
            .O(N__30241),
            .I(N__30238));
    LocalMux I__5528 (
            .O(N__30238),
            .I(N__30235));
    Span4Mux_h I__5527 (
            .O(N__30235),
            .I(N__30232));
    Odrv4 I__5526 (
            .O(N__30232),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_1 ));
    InMux I__5525 (
            .O(N__30229),
            .I(N__30226));
    LocalMux I__5524 (
            .O(N__30226),
            .I(N__30223));
    Odrv4 I__5523 (
            .O(N__30223),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_1 ));
    InMux I__5522 (
            .O(N__30220),
            .I(N__30217));
    LocalMux I__5521 (
            .O(N__30217),
            .I(N__30214));
    Span4Mux_v I__5520 (
            .O(N__30214),
            .I(N__30211));
    Span4Mux_h I__5519 (
            .O(N__30211),
            .I(N__30208));
    Odrv4 I__5518 (
            .O(N__30208),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_2 ));
    InMux I__5517 (
            .O(N__30205),
            .I(N__30202));
    LocalMux I__5516 (
            .O(N__30202),
            .I(N__30199));
    Odrv12 I__5515 (
            .O(N__30199),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_2 ));
    InMux I__5514 (
            .O(N__30196),
            .I(N__30193));
    LocalMux I__5513 (
            .O(N__30193),
            .I(N__30190));
    Odrv4 I__5512 (
            .O(N__30190),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNI21TNZ0Z_2 ));
    InMux I__5511 (
            .O(N__30187),
            .I(N__30184));
    LocalMux I__5510 (
            .O(N__30184),
            .I(N__30181));
    Span4Mux_h I__5509 (
            .O(N__30181),
            .I(N__30178));
    Odrv4 I__5508 (
            .O(N__30178),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_3 ));
    InMux I__5507 (
            .O(N__30175),
            .I(N__30172));
    LocalMux I__5506 (
            .O(N__30172),
            .I(N__30169));
    Span12Mux_v I__5505 (
            .O(N__30169),
            .I(N__30166));
    Odrv12 I__5504 (
            .O(N__30166),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_3 ));
    InMux I__5503 (
            .O(N__30163),
            .I(N__30160));
    LocalMux I__5502 (
            .O(N__30160),
            .I(N__30157));
    Span4Mux_v I__5501 (
            .O(N__30157),
            .I(N__30154));
    Span4Mux_v I__5500 (
            .O(N__30154),
            .I(N__30151));
    Sp12to4 I__5499 (
            .O(N__30151),
            .I(N__30148));
    Odrv12 I__5498 (
            .O(N__30148),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_4 ));
    InMux I__5497 (
            .O(N__30145),
            .I(N__30142));
    LocalMux I__5496 (
            .O(N__30142),
            .I(N__30139));
    Odrv12 I__5495 (
            .O(N__30139),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_4 ));
    InMux I__5494 (
            .O(N__30136),
            .I(N__30133));
    LocalMux I__5493 (
            .O(N__30133),
            .I(N__30130));
    Odrv4 I__5492 (
            .O(N__30130),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNI65TNZ0Z_4 ));
    InMux I__5491 (
            .O(N__30127),
            .I(N__30124));
    LocalMux I__5490 (
            .O(N__30124),
            .I(N__30121));
    Span12Mux_h I__5489 (
            .O(N__30121),
            .I(N__30118));
    Odrv12 I__5488 (
            .O(N__30118),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_5 ));
    InMux I__5487 (
            .O(N__30115),
            .I(N__30112));
    LocalMux I__5486 (
            .O(N__30112),
            .I(N__30109));
    Span4Mux_h I__5485 (
            .O(N__30109),
            .I(N__30106));
    Sp12to4 I__5484 (
            .O(N__30106),
            .I(N__30103));
    Odrv12 I__5483 (
            .O(N__30103),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_5 ));
    InMux I__5482 (
            .O(N__30100),
            .I(N__30097));
    LocalMux I__5481 (
            .O(N__30097),
            .I(N__30094));
    Span4Mux_h I__5480 (
            .O(N__30094),
            .I(N__30091));
    Odrv4 I__5479 (
            .O(N__30091),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_7 ));
    InMux I__5478 (
            .O(N__30088),
            .I(N__30085));
    LocalMux I__5477 (
            .O(N__30085),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_7 ));
    InMux I__5476 (
            .O(N__30082),
            .I(N__30079));
    LocalMux I__5475 (
            .O(N__30079),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_4 ));
    InMux I__5474 (
            .O(N__30076),
            .I(N__30073));
    LocalMux I__5473 (
            .O(N__30073),
            .I(N__30070));
    Span4Mux_v I__5472 (
            .O(N__30070),
            .I(N__30067));
    Span4Mux_v I__5471 (
            .O(N__30067),
            .I(N__30064));
    Odrv4 I__5470 (
            .O(N__30064),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_12 ));
    InMux I__5469 (
            .O(N__30061),
            .I(N__30058));
    LocalMux I__5468 (
            .O(N__30058),
            .I(N__30055));
    Odrv4 I__5467 (
            .O(N__30055),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_12 ));
    CascadeMux I__5466 (
            .O(N__30052),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI4RFTZ0Z_12_cascade_ ));
    InMux I__5465 (
            .O(N__30049),
            .I(N__30046));
    LocalMux I__5464 (
            .O(N__30046),
            .I(N__30043));
    Odrv4 I__5463 (
            .O(N__30043),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI1MA71Z0Z_12 ));
    InMux I__5462 (
            .O(N__30040),
            .I(N__30037));
    LocalMux I__5461 (
            .O(N__30037),
            .I(N__30034));
    Odrv4 I__5460 (
            .O(N__30034),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_20 ));
    InMux I__5459 (
            .O(N__30031),
            .I(N__30028));
    LocalMux I__5458 (
            .O(N__30028),
            .I(N__30025));
    Span4Mux_h I__5457 (
            .O(N__30025),
            .I(N__30022));
    Odrv4 I__5456 (
            .O(N__30022),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_12 ));
    InMux I__5455 (
            .O(N__30019),
            .I(N__30016));
    LocalMux I__5454 (
            .O(N__30016),
            .I(N__30013));
    Span4Mux_v I__5453 (
            .O(N__30013),
            .I(N__30010));
    Span4Mux_v I__5452 (
            .O(N__30010),
            .I(N__30007));
    Odrv4 I__5451 (
            .O(N__30007),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_12 ));
    CascadeMux I__5450 (
            .O(N__30004),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI077KZ0Z_12_cascade_ ));
    InMux I__5449 (
            .O(N__30001),
            .I(N__29998));
    LocalMux I__5448 (
            .O(N__29998),
            .I(N__29995));
    Odrv12 I__5447 (
            .O(N__29995),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNISIUQZ0Z_12 ));
    InMux I__5446 (
            .O(N__29992),
            .I(N__29989));
    LocalMux I__5445 (
            .O(N__29989),
            .I(N__29986));
    Odrv4 I__5444 (
            .O(N__29986),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIE4DM1Z0Z_2 ));
    InMux I__5443 (
            .O(N__29983),
            .I(N__29980));
    LocalMux I__5442 (
            .O(N__29980),
            .I(N__29977));
    Span4Mux_v I__5441 (
            .O(N__29977),
            .I(N__29974));
    Odrv4 I__5440 (
            .O(N__29974),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_14 ));
    InMux I__5439 (
            .O(N__29971),
            .I(N__29968));
    LocalMux I__5438 (
            .O(N__29968),
            .I(N__29965));
    Span4Mux_v I__5437 (
            .O(N__29965),
            .I(N__29962));
    Odrv4 I__5436 (
            .O(N__29962),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI8VFTZ0Z_14 ));
    InMux I__5435 (
            .O(N__29959),
            .I(N__29956));
    LocalMux I__5434 (
            .O(N__29956),
            .I(N__29953));
    Span4Mux_h I__5433 (
            .O(N__29953),
            .I(N__29950));
    Odrv4 I__5432 (
            .O(N__29950),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_2 ));
    InMux I__5431 (
            .O(N__29947),
            .I(N__29944));
    LocalMux I__5430 (
            .O(N__29944),
            .I(N__29941));
    Odrv4 I__5429 (
            .O(N__29941),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIUG4NZ0Z_2 ));
    InMux I__5428 (
            .O(N__29938),
            .I(N__29935));
    LocalMux I__5427 (
            .O(N__29935),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_2 ));
    CascadeMux I__5426 (
            .O(N__29932),
            .I(DMAq_12_cascade_));
    InMux I__5425 (
            .O(N__29929),
            .I(N__29926));
    LocalMux I__5424 (
            .O(N__29926),
            .I(N__29923));
    Span4Mux_v I__5423 (
            .O(N__29923),
            .I(N__29920));
    Span4Mux_h I__5422 (
            .O(N__29920),
            .I(N__29917));
    Span4Mux_h I__5421 (
            .O(N__29917),
            .I(N__29914));
    Odrv4 I__5420 (
            .O(N__29914),
            .I(PIOq_12));
    InMux I__5419 (
            .O(N__29911),
            .I(N__29908));
    LocalMux I__5418 (
            .O(N__29908),
            .I(\u0.dat_o_0_0_1Z0Z_12 ));
    CascadeMux I__5417 (
            .O(N__29905),
            .I(\u0.dat_o_0_0_1Z0Z_4_cascade_ ));
    InMux I__5416 (
            .O(N__29902),
            .I(N__29899));
    LocalMux I__5415 (
            .O(N__29899),
            .I(N__29896));
    Odrv4 I__5414 (
            .O(N__29896),
            .I(\u0.dat_o_0_0_2_4 ));
    IoInMux I__5413 (
            .O(N__29893),
            .I(N__29890));
    LocalMux I__5412 (
            .O(N__29890),
            .I(N__29887));
    IoSpan4Mux I__5411 (
            .O(N__29887),
            .I(N__29884));
    Span4Mux_s3_h I__5410 (
            .O(N__29884),
            .I(N__29881));
    Sp12to4 I__5409 (
            .O(N__29881),
            .I(N__29878));
    Span12Mux_h I__5408 (
            .O(N__29878),
            .I(N__29875));
    Odrv12 I__5407 (
            .O(N__29875),
            .I(wb_dat_o_c_4));
    CascadeMux I__5406 (
            .O(N__29872),
            .I(N__29869));
    InMux I__5405 (
            .O(N__29869),
            .I(N__29865));
    InMux I__5404 (
            .O(N__29868),
            .I(N__29862));
    LocalMux I__5403 (
            .O(N__29865),
            .I(N__29859));
    LocalMux I__5402 (
            .O(N__29862),
            .I(N__29856));
    Span4Mux_h I__5401 (
            .O(N__29859),
            .I(N__29853));
    Odrv12 I__5400 (
            .O(N__29856),
            .I(PIO_dport1_T1_4));
    Odrv4 I__5399 (
            .O(N__29853),
            .I(PIO_dport1_T1_4));
    InMux I__5398 (
            .O(N__29848),
            .I(N__29845));
    LocalMux I__5397 (
            .O(N__29845),
            .I(N__29842));
    Odrv12 I__5396 (
            .O(N__29842),
            .I(\u0.dat_o_0_0_0_4 ));
    InMux I__5395 (
            .O(N__29839),
            .I(N__29836));
    LocalMux I__5394 (
            .O(N__29836),
            .I(N__29833));
    Span4Mux_v I__5393 (
            .O(N__29833),
            .I(N__29830));
    Span4Mux_v I__5392 (
            .O(N__29830),
            .I(N__29827));
    Odrv4 I__5391 (
            .O(N__29827),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI2L4NZ0Z_4 ));
    CascadeMux I__5390 (
            .O(N__29824),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNII4OK1Z0Z_2_cascade_ ));
    InMux I__5389 (
            .O(N__29821),
            .I(N__29818));
    LocalMux I__5388 (
            .O(N__29818),
            .I(DMAq_4));
    InMux I__5387 (
            .O(N__29815),
            .I(N__29812));
    LocalMux I__5386 (
            .O(N__29812),
            .I(N__29807));
    InMux I__5385 (
            .O(N__29811),
            .I(N__29802));
    InMux I__5384 (
            .O(N__29810),
            .I(N__29802));
    Span4Mux_v I__5383 (
            .O(N__29807),
            .I(N__29799));
    LocalMux I__5382 (
            .O(N__29802),
            .I(N__29796));
    Span4Mux_v I__5381 (
            .O(N__29799),
            .I(N__29793));
    Span4Mux_v I__5380 (
            .O(N__29796),
            .I(N__29790));
    Span4Mux_h I__5379 (
            .O(N__29793),
            .I(N__29785));
    Span4Mux_v I__5378 (
            .O(N__29790),
            .I(N__29785));
    Sp12to4 I__5377 (
            .O(N__29785),
            .I(N__29782));
    Odrv12 I__5376 (
            .O(N__29782),
            .I(dd_pad_i_c_4));
    InMux I__5375 (
            .O(N__29779),
            .I(N__29776));
    LocalMux I__5374 (
            .O(N__29776),
            .I(N__29773));
    Odrv12 I__5373 (
            .O(N__29773),
            .I(PIOq_4));
    InMux I__5372 (
            .O(N__29770),
            .I(N__29767));
    LocalMux I__5371 (
            .O(N__29767),
            .I(N__29764));
    Odrv4 I__5370 (
            .O(N__29764),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_4 ));
    InMux I__5369 (
            .O(N__29761),
            .I(N__29758));
    LocalMux I__5368 (
            .O(N__29758),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIKJOD1Z0Z_4 ));
    InMux I__5367 (
            .O(N__29755),
            .I(N__29752));
    LocalMux I__5366 (
            .O(N__29752),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_4 ));
    InMux I__5365 (
            .O(N__29749),
            .I(N__29746));
    LocalMux I__5364 (
            .O(N__29746),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIU4CMZ0Z_4 ));
    InMux I__5363 (
            .O(N__29743),
            .I(N__29740));
    LocalMux I__5362 (
            .O(N__29740),
            .I(N__29737));
    Span4Mux_v I__5361 (
            .O(N__29737),
            .I(N__29734));
    Span4Mux_v I__5360 (
            .O(N__29734),
            .I(N__29731));
    Odrv4 I__5359 (
            .O(N__29731),
            .I(\u0.dat_o_0_0_3_12 ));
    CascadeMux I__5358 (
            .O(N__29728),
            .I(\u0.dat_o_0_0_2_12_cascade_ ));
    IoInMux I__5357 (
            .O(N__29725),
            .I(N__29722));
    LocalMux I__5356 (
            .O(N__29722),
            .I(N__29719));
    IoSpan4Mux I__5355 (
            .O(N__29719),
            .I(N__29716));
    Span4Mux_s1_v I__5354 (
            .O(N__29716),
            .I(N__29713));
    Span4Mux_h I__5353 (
            .O(N__29713),
            .I(N__29710));
    Sp12to4 I__5352 (
            .O(N__29710),
            .I(N__29707));
    Span12Mux_h I__5351 (
            .O(N__29707),
            .I(N__29704));
    Odrv12 I__5350 (
            .O(N__29704),
            .I(wb_dat_o_c_12));
    InMux I__5349 (
            .O(N__29701),
            .I(N__29698));
    LocalMux I__5348 (
            .O(N__29698),
            .I(\u0.CtrlRegZ0Z_12 ));
    CascadeMux I__5347 (
            .O(N__29695),
            .I(N__29692));
    InMux I__5346 (
            .O(N__29692),
            .I(N__29689));
    LocalMux I__5345 (
            .O(N__29689),
            .I(N__29686));
    Span4Mux_v I__5344 (
            .O(N__29686),
            .I(N__29683));
    Span4Mux_h I__5343 (
            .O(N__29683),
            .I(N__29679));
    InMux I__5342 (
            .O(N__29682),
            .I(N__29676));
    Odrv4 I__5341 (
            .O(N__29679),
            .I(DMA_dev0_Td_4));
    LocalMux I__5340 (
            .O(N__29676),
            .I(DMA_dev0_Td_4));
    InMux I__5339 (
            .O(N__29671),
            .I(N__29668));
    LocalMux I__5338 (
            .O(N__29668),
            .I(N__29665));
    Odrv12 I__5337 (
            .O(N__29665),
            .I(\u0.dat_o_0_0_0_12 ));
    InMux I__5336 (
            .O(N__29662),
            .I(N__29659));
    LocalMux I__5335 (
            .O(N__29659),
            .I(N__29656));
    Span4Mux_s3_h I__5334 (
            .O(N__29656),
            .I(N__29653));
    Span4Mux_h I__5333 (
            .O(N__29653),
            .I(N__29650));
    Span4Mux_h I__5332 (
            .O(N__29650),
            .I(N__29647));
    Odrv4 I__5331 (
            .O(N__29647),
            .I(\u1.PIO_control.PIO_access_control.TeocZ0Z_0 ));
    InMux I__5330 (
            .O(N__29644),
            .I(N__29641));
    LocalMux I__5329 (
            .O(N__29641),
            .I(N__29638));
    Span4Mux_v I__5328 (
            .O(N__29638),
            .I(N__29635));
    Span4Mux_h I__5327 (
            .O(N__29635),
            .I(N__29631));
    InMux I__5326 (
            .O(N__29634),
            .I(N__29628));
    Span4Mux_h I__5325 (
            .O(N__29631),
            .I(N__29623));
    LocalMux I__5324 (
            .O(N__29628),
            .I(N__29623));
    Odrv4 I__5323 (
            .O(N__29623),
            .I(PIO_cmdport_T2_5));
    InMux I__5322 (
            .O(N__29620),
            .I(N__29616));
    InMux I__5321 (
            .O(N__29619),
            .I(N__29613));
    LocalMux I__5320 (
            .O(N__29616),
            .I(N__29610));
    LocalMux I__5319 (
            .O(N__29613),
            .I(N__29607));
    Span4Mux_h I__5318 (
            .O(N__29610),
            .I(N__29604));
    Odrv12 I__5317 (
            .O(N__29607),
            .I(PIO_cmdport_T2_7));
    Odrv4 I__5316 (
            .O(N__29604),
            .I(PIO_cmdport_T2_7));
    InMux I__5315 (
            .O(N__29599),
            .I(N__29596));
    LocalMux I__5314 (
            .O(N__29596),
            .I(N__29592));
    InMux I__5313 (
            .O(N__29595),
            .I(N__29589));
    Span4Mux_v I__5312 (
            .O(N__29592),
            .I(N__29584));
    LocalMux I__5311 (
            .O(N__29589),
            .I(N__29584));
    Odrv4 I__5310 (
            .O(N__29584),
            .I(PIO_cmdport_T4_3));
    InMux I__5309 (
            .O(N__29581),
            .I(N__29577));
    InMux I__5308 (
            .O(N__29580),
            .I(N__29574));
    LocalMux I__5307 (
            .O(N__29577),
            .I(N__29571));
    LocalMux I__5306 (
            .O(N__29574),
            .I(N__29568));
    Odrv4 I__5305 (
            .O(N__29571),
            .I(PIO_cmdport_T4_4));
    Odrv4 I__5304 (
            .O(N__29568),
            .I(PIO_cmdport_T4_4));
    InMux I__5303 (
            .O(N__29563),
            .I(N__29559));
    CascadeMux I__5302 (
            .O(N__29562),
            .I(N__29556));
    LocalMux I__5301 (
            .O(N__29559),
            .I(N__29553));
    InMux I__5300 (
            .O(N__29556),
            .I(N__29550));
    Odrv4 I__5299 (
            .O(N__29553),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.QiZ0Z_7 ));
    LocalMux I__5298 (
            .O(N__29550),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.QiZ0Z_7 ));
    InMux I__5297 (
            .O(N__29545),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_cry_6 ));
    InMux I__5296 (
            .O(N__29542),
            .I(N__29539));
    LocalMux I__5295 (
            .O(N__29539),
            .I(N__29536));
    Odrv4 I__5294 (
            .O(N__29536),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_s_7 ));
    InMux I__5293 (
            .O(N__29533),
            .I(N__29530));
    LocalMux I__5292 (
            .O(N__29530),
            .I(\u1.PIO_control.PIO_access_control.iteoc_1_iv_i_i_0_1 ));
    InMux I__5291 (
            .O(N__29527),
            .I(N__29524));
    LocalMux I__5290 (
            .O(N__29524),
            .I(N__29521));
    Span4Mux_s3_h I__5289 (
            .O(N__29521),
            .I(N__29518));
    Span4Mux_h I__5288 (
            .O(N__29518),
            .I(N__29515));
    Span4Mux_h I__5287 (
            .O(N__29515),
            .I(N__29512));
    Odrv4 I__5286 (
            .O(N__29512),
            .I(\u1.PIO_control.PIO_access_control.TeocZ0Z_1 ));
    CascadeMux I__5285 (
            .O(N__29509),
            .I(\u1.PIO_control.PIO_access_control.it4_1_iv_0_0_1_cascade_ ));
    InMux I__5284 (
            .O(N__29506),
            .I(N__29503));
    LocalMux I__5283 (
            .O(N__29503),
            .I(N__29500));
    Span4Mux_h I__5282 (
            .O(N__29500),
            .I(N__29497));
    Span4Mux_h I__5281 (
            .O(N__29497),
            .I(N__29494));
    Span4Mux_h I__5280 (
            .O(N__29494),
            .I(N__29491));
    Odrv4 I__5279 (
            .O(N__29491),
            .I(\u1.PIO_control.PIO_access_control.T4Z0Z_1 ));
    InMux I__5278 (
            .O(N__29488),
            .I(N__29485));
    LocalMux I__5277 (
            .O(N__29485),
            .I(\u1.PIO_control.PIO_access_control.iteoc_1_iv_i_i_0_3 ));
    InMux I__5276 (
            .O(N__29482),
            .I(N__29479));
    LocalMux I__5275 (
            .O(N__29479),
            .I(N__29476));
    Span4Mux_v I__5274 (
            .O(N__29476),
            .I(N__29473));
    Span4Mux_h I__5273 (
            .O(N__29473),
            .I(N__29470));
    Span4Mux_h I__5272 (
            .O(N__29470),
            .I(N__29467));
    Odrv4 I__5271 (
            .O(N__29467),
            .I(\u1.PIO_control.PIO_access_control.TeocZ0Z_3 ));
    CascadeMux I__5270 (
            .O(N__29464),
            .I(N__29453));
    CascadeMux I__5269 (
            .O(N__29463),
            .I(N__29442));
    InMux I__5268 (
            .O(N__29462),
            .I(N__29429));
    InMux I__5267 (
            .O(N__29461),
            .I(N__29429));
    InMux I__5266 (
            .O(N__29460),
            .I(N__29429));
    InMux I__5265 (
            .O(N__29459),
            .I(N__29420));
    InMux I__5264 (
            .O(N__29458),
            .I(N__29420));
    InMux I__5263 (
            .O(N__29457),
            .I(N__29420));
    InMux I__5262 (
            .O(N__29456),
            .I(N__29420));
    InMux I__5261 (
            .O(N__29453),
            .I(N__29415));
    InMux I__5260 (
            .O(N__29452),
            .I(N__29415));
    InMux I__5259 (
            .O(N__29451),
            .I(N__29412));
    CascadeMux I__5258 (
            .O(N__29450),
            .I(N__29407));
    CascadeMux I__5257 (
            .O(N__29449),
            .I(N__29403));
    CascadeMux I__5256 (
            .O(N__29448),
            .I(N__29399));
    CascadeMux I__5255 (
            .O(N__29447),
            .I(N__29396));
    CascadeMux I__5254 (
            .O(N__29446),
            .I(N__29393));
    CascadeMux I__5253 (
            .O(N__29445),
            .I(N__29390));
    InMux I__5252 (
            .O(N__29442),
            .I(N__29381));
    InMux I__5251 (
            .O(N__29441),
            .I(N__29381));
    InMux I__5250 (
            .O(N__29440),
            .I(N__29381));
    CascadeMux I__5249 (
            .O(N__29439),
            .I(N__29377));
    CascadeMux I__5248 (
            .O(N__29438),
            .I(N__29373));
    CascadeMux I__5247 (
            .O(N__29437),
            .I(N__29370));
    CascadeMux I__5246 (
            .O(N__29436),
            .I(N__29367));
    LocalMux I__5245 (
            .O(N__29429),
            .I(N__29362));
    LocalMux I__5244 (
            .O(N__29420),
            .I(N__29359));
    LocalMux I__5243 (
            .O(N__29415),
            .I(N__29356));
    LocalMux I__5242 (
            .O(N__29412),
            .I(N__29353));
    InMux I__5241 (
            .O(N__29411),
            .I(N__29340));
    InMux I__5240 (
            .O(N__29410),
            .I(N__29340));
    InMux I__5239 (
            .O(N__29407),
            .I(N__29340));
    InMux I__5238 (
            .O(N__29406),
            .I(N__29340));
    InMux I__5237 (
            .O(N__29403),
            .I(N__29340));
    InMux I__5236 (
            .O(N__29402),
            .I(N__29340));
    InMux I__5235 (
            .O(N__29399),
            .I(N__29329));
    InMux I__5234 (
            .O(N__29396),
            .I(N__29329));
    InMux I__5233 (
            .O(N__29393),
            .I(N__29329));
    InMux I__5232 (
            .O(N__29390),
            .I(N__29329));
    InMux I__5231 (
            .O(N__29389),
            .I(N__29329));
    InMux I__5230 (
            .O(N__29388),
            .I(N__29326));
    LocalMux I__5229 (
            .O(N__29381),
            .I(N__29323));
    InMux I__5228 (
            .O(N__29380),
            .I(N__29316));
    InMux I__5227 (
            .O(N__29377),
            .I(N__29316));
    InMux I__5226 (
            .O(N__29376),
            .I(N__29316));
    InMux I__5225 (
            .O(N__29373),
            .I(N__29307));
    InMux I__5224 (
            .O(N__29370),
            .I(N__29307));
    InMux I__5223 (
            .O(N__29367),
            .I(N__29307));
    InMux I__5222 (
            .O(N__29366),
            .I(N__29307));
    InMux I__5221 (
            .O(N__29365),
            .I(N__29304));
    Odrv4 I__5220 (
            .O(N__29362),
            .I(\u1.PIO_control.PIO_access_control.N_1319 ));
    Odrv4 I__5219 (
            .O(N__29359),
            .I(\u1.PIO_control.PIO_access_control.N_1319 ));
    Odrv4 I__5218 (
            .O(N__29356),
            .I(\u1.PIO_control.PIO_access_control.N_1319 ));
    Odrv12 I__5217 (
            .O(N__29353),
            .I(\u1.PIO_control.PIO_access_control.N_1319 ));
    LocalMux I__5216 (
            .O(N__29340),
            .I(\u1.PIO_control.PIO_access_control.N_1319 ));
    LocalMux I__5215 (
            .O(N__29329),
            .I(\u1.PIO_control.PIO_access_control.N_1319 ));
    LocalMux I__5214 (
            .O(N__29326),
            .I(\u1.PIO_control.PIO_access_control.N_1319 ));
    Odrv4 I__5213 (
            .O(N__29323),
            .I(\u1.PIO_control.PIO_access_control.N_1319 ));
    LocalMux I__5212 (
            .O(N__29316),
            .I(\u1.PIO_control.PIO_access_control.N_1319 ));
    LocalMux I__5211 (
            .O(N__29307),
            .I(\u1.PIO_control.PIO_access_control.N_1319 ));
    LocalMux I__5210 (
            .O(N__29304),
            .I(\u1.PIO_control.PIO_access_control.N_1319 ));
    InMux I__5209 (
            .O(N__29281),
            .I(N__29271));
    InMux I__5208 (
            .O(N__29280),
            .I(N__29271));
    InMux I__5207 (
            .O(N__29279),
            .I(N__29258));
    InMux I__5206 (
            .O(N__29278),
            .I(N__29258));
    InMux I__5205 (
            .O(N__29277),
            .I(N__29258));
    InMux I__5204 (
            .O(N__29276),
            .I(N__29258));
    LocalMux I__5203 (
            .O(N__29271),
            .I(N__29249));
    InMux I__5202 (
            .O(N__29270),
            .I(N__29234));
    InMux I__5201 (
            .O(N__29269),
            .I(N__29234));
    InMux I__5200 (
            .O(N__29268),
            .I(N__29234));
    InMux I__5199 (
            .O(N__29267),
            .I(N__29234));
    LocalMux I__5198 (
            .O(N__29258),
            .I(N__29231));
    InMux I__5197 (
            .O(N__29257),
            .I(N__29228));
    InMux I__5196 (
            .O(N__29256),
            .I(N__29225));
    InMux I__5195 (
            .O(N__29255),
            .I(N__29216));
    InMux I__5194 (
            .O(N__29254),
            .I(N__29216));
    InMux I__5193 (
            .O(N__29253),
            .I(N__29216));
    InMux I__5192 (
            .O(N__29252),
            .I(N__29216));
    Span4Mux_h I__5191 (
            .O(N__29249),
            .I(N__29203));
    InMux I__5190 (
            .O(N__29248),
            .I(N__29194));
    InMux I__5189 (
            .O(N__29247),
            .I(N__29194));
    InMux I__5188 (
            .O(N__29246),
            .I(N__29194));
    InMux I__5187 (
            .O(N__29245),
            .I(N__29194));
    InMux I__5186 (
            .O(N__29244),
            .I(N__29189));
    InMux I__5185 (
            .O(N__29243),
            .I(N__29189));
    LocalMux I__5184 (
            .O(N__29234),
            .I(N__29186));
    Span4Mux_h I__5183 (
            .O(N__29231),
            .I(N__29181));
    LocalMux I__5182 (
            .O(N__29228),
            .I(N__29181));
    LocalMux I__5181 (
            .O(N__29225),
            .I(N__29176));
    LocalMux I__5180 (
            .O(N__29216),
            .I(N__29176));
    InMux I__5179 (
            .O(N__29215),
            .I(N__29167));
    InMux I__5178 (
            .O(N__29214),
            .I(N__29167));
    InMux I__5177 (
            .O(N__29213),
            .I(N__29167));
    InMux I__5176 (
            .O(N__29212),
            .I(N__29167));
    InMux I__5175 (
            .O(N__29211),
            .I(N__29154));
    InMux I__5174 (
            .O(N__29210),
            .I(N__29154));
    InMux I__5173 (
            .O(N__29209),
            .I(N__29154));
    InMux I__5172 (
            .O(N__29208),
            .I(N__29154));
    InMux I__5171 (
            .O(N__29207),
            .I(N__29154));
    InMux I__5170 (
            .O(N__29206),
            .I(N__29154));
    Odrv4 I__5169 (
            .O(N__29203),
            .I(\u1.PIO_control.PIO_access_control.N_2112 ));
    LocalMux I__5168 (
            .O(N__29194),
            .I(\u1.PIO_control.PIO_access_control.N_2112 ));
    LocalMux I__5167 (
            .O(N__29189),
            .I(\u1.PIO_control.PIO_access_control.N_2112 ));
    Odrv4 I__5166 (
            .O(N__29186),
            .I(\u1.PIO_control.PIO_access_control.N_2112 ));
    Odrv4 I__5165 (
            .O(N__29181),
            .I(\u1.PIO_control.PIO_access_control.N_2112 ));
    Odrv12 I__5164 (
            .O(N__29176),
            .I(\u1.PIO_control.PIO_access_control.N_2112 ));
    LocalMux I__5163 (
            .O(N__29167),
            .I(\u1.PIO_control.PIO_access_control.N_2112 ));
    LocalMux I__5162 (
            .O(N__29154),
            .I(\u1.PIO_control.PIO_access_control.N_2112 ));
    CascadeMux I__5161 (
            .O(N__29137),
            .I(\u1.PIO_control.PIO_access_control.iteoc_1_iv_i_i_0_4_cascade_ ));
    InMux I__5160 (
            .O(N__29134),
            .I(N__29131));
    LocalMux I__5159 (
            .O(N__29131),
            .I(N__29128));
    Span12Mux_v I__5158 (
            .O(N__29128),
            .I(N__29125));
    Odrv12 I__5157 (
            .O(N__29125),
            .I(\u1.PIO_control.PIO_access_control.TeocZ0Z_4 ));
    InMux I__5156 (
            .O(N__29122),
            .I(N__29119));
    LocalMux I__5155 (
            .O(N__29119),
            .I(\u1.PIO_control.PIO_access_control.it4_1_iv_i_i_0_6 ));
    InMux I__5154 (
            .O(N__29116),
            .I(N__29113));
    LocalMux I__5153 (
            .O(N__29113),
            .I(N__29110));
    Span4Mux_s3_h I__5152 (
            .O(N__29110),
            .I(N__29107));
    Span4Mux_h I__5151 (
            .O(N__29107),
            .I(N__29104));
    Span4Mux_h I__5150 (
            .O(N__29104),
            .I(N__29101));
    Odrv4 I__5149 (
            .O(N__29101),
            .I(\u1.PIO_control.PIO_access_control.T4Z0Z_6 ));
    InMux I__5148 (
            .O(N__29098),
            .I(N__29085));
    InMux I__5147 (
            .O(N__29097),
            .I(N__29085));
    InMux I__5146 (
            .O(N__29096),
            .I(N__29072));
    InMux I__5145 (
            .O(N__29095),
            .I(N__29072));
    InMux I__5144 (
            .O(N__29094),
            .I(N__29072));
    InMux I__5143 (
            .O(N__29093),
            .I(N__29072));
    InMux I__5142 (
            .O(N__29092),
            .I(N__29072));
    InMux I__5141 (
            .O(N__29091),
            .I(N__29072));
    InMux I__5140 (
            .O(N__29090),
            .I(N__29063));
    LocalMux I__5139 (
            .O(N__29085),
            .I(N__29056));
    LocalMux I__5138 (
            .O(N__29072),
            .I(N__29056));
    InMux I__5137 (
            .O(N__29071),
            .I(N__29051));
    InMux I__5136 (
            .O(N__29070),
            .I(N__29051));
    InMux I__5135 (
            .O(N__29069),
            .I(N__29042));
    InMux I__5134 (
            .O(N__29068),
            .I(N__29042));
    InMux I__5133 (
            .O(N__29067),
            .I(N__29042));
    InMux I__5132 (
            .O(N__29066),
            .I(N__29042));
    LocalMux I__5131 (
            .O(N__29063),
            .I(N__29024));
    InMux I__5130 (
            .O(N__29062),
            .I(N__29019));
    InMux I__5129 (
            .O(N__29061),
            .I(N__29019));
    Span4Mux_v I__5128 (
            .O(N__29056),
            .I(N__29016));
    LocalMux I__5127 (
            .O(N__29051),
            .I(N__29011));
    LocalMux I__5126 (
            .O(N__29042),
            .I(N__29011));
    InMux I__5125 (
            .O(N__29041),
            .I(N__29002));
    InMux I__5124 (
            .O(N__29040),
            .I(N__29002));
    InMux I__5123 (
            .O(N__29039),
            .I(N__29002));
    InMux I__5122 (
            .O(N__29038),
            .I(N__29002));
    InMux I__5121 (
            .O(N__29037),
            .I(N__28993));
    InMux I__5120 (
            .O(N__29036),
            .I(N__28993));
    InMux I__5119 (
            .O(N__29035),
            .I(N__28993));
    InMux I__5118 (
            .O(N__29034),
            .I(N__28993));
    InMux I__5117 (
            .O(N__29033),
            .I(N__28986));
    InMux I__5116 (
            .O(N__29032),
            .I(N__28986));
    InMux I__5115 (
            .O(N__29031),
            .I(N__28986));
    InMux I__5114 (
            .O(N__29030),
            .I(N__28977));
    InMux I__5113 (
            .O(N__29029),
            .I(N__28977));
    InMux I__5112 (
            .O(N__29028),
            .I(N__28977));
    InMux I__5111 (
            .O(N__29027),
            .I(N__28977));
    Odrv4 I__5110 (
            .O(N__29024),
            .I(\u1.PIO_control.PIO_access_control.N_2110 ));
    LocalMux I__5109 (
            .O(N__29019),
            .I(\u1.PIO_control.PIO_access_control.N_2110 ));
    Odrv4 I__5108 (
            .O(N__29016),
            .I(\u1.PIO_control.PIO_access_control.N_2110 ));
    Odrv4 I__5107 (
            .O(N__29011),
            .I(\u1.PIO_control.PIO_access_control.N_2110 ));
    LocalMux I__5106 (
            .O(N__29002),
            .I(\u1.PIO_control.PIO_access_control.N_2110 ));
    LocalMux I__5105 (
            .O(N__28993),
            .I(\u1.PIO_control.PIO_access_control.N_2110 ));
    LocalMux I__5104 (
            .O(N__28986),
            .I(\u1.PIO_control.PIO_access_control.N_2110 ));
    LocalMux I__5103 (
            .O(N__28977),
            .I(\u1.PIO_control.PIO_access_control.N_2110 ));
    InMux I__5102 (
            .O(N__28960),
            .I(N__28957));
    LocalMux I__5101 (
            .O(N__28957),
            .I(\u1.PIO_control.PIO_access_control.iteoc_1_iv_i_i_0_0 ));
    CascadeMux I__5100 (
            .O(N__28954),
            .I(N__28951));
    InMux I__5099 (
            .O(N__28951),
            .I(N__28948));
    LocalMux I__5098 (
            .O(N__28948),
            .I(N__28945));
    Span4Mux_h I__5097 (
            .O(N__28945),
            .I(N__28939));
    InMux I__5096 (
            .O(N__28944),
            .I(N__28934));
    InMux I__5095 (
            .O(N__28943),
            .I(N__28934));
    InMux I__5094 (
            .O(N__28942),
            .I(N__28931));
    Span4Mux_h I__5093 (
            .O(N__28939),
            .I(N__28924));
    LocalMux I__5092 (
            .O(N__28934),
            .I(N__28924));
    LocalMux I__5091 (
            .O(N__28931),
            .I(N__28924));
    Odrv4 I__5090 (
            .O(N__28924),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.QiZ0Z_0 ));
    InMux I__5089 (
            .O(N__28921),
            .I(N__28917));
    InMux I__5088 (
            .O(N__28920),
            .I(N__28914));
    LocalMux I__5087 (
            .O(N__28917),
            .I(N__28908));
    LocalMux I__5086 (
            .O(N__28914),
            .I(N__28908));
    InMux I__5085 (
            .O(N__28913),
            .I(N__28905));
    Odrv12 I__5084 (
            .O(N__28908),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.QiZ0Z_1 ));
    LocalMux I__5083 (
            .O(N__28905),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.QiZ0Z_1 ));
    InMux I__5082 (
            .O(N__28900),
            .I(N__28897));
    LocalMux I__5081 (
            .O(N__28897),
            .I(N__28894));
    Span4Mux_h I__5080 (
            .O(N__28894),
            .I(N__28891));
    Odrv4 I__5079 (
            .O(N__28891),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_s_1 ));
    InMux I__5078 (
            .O(N__28888),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_cry_0 ));
    InMux I__5077 (
            .O(N__28885),
            .I(N__28881));
    InMux I__5076 (
            .O(N__28884),
            .I(N__28878));
    LocalMux I__5075 (
            .O(N__28881),
            .I(N__28873));
    LocalMux I__5074 (
            .O(N__28878),
            .I(N__28873));
    Odrv12 I__5073 (
            .O(N__28873),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.QiZ0Z_2 ));
    InMux I__5072 (
            .O(N__28870),
            .I(N__28867));
    LocalMux I__5071 (
            .O(N__28867),
            .I(N__28864));
    Odrv12 I__5070 (
            .O(N__28864),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_s_2 ));
    InMux I__5069 (
            .O(N__28861),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_cry_1 ));
    InMux I__5068 (
            .O(N__28858),
            .I(N__28854));
    InMux I__5067 (
            .O(N__28857),
            .I(N__28851));
    LocalMux I__5066 (
            .O(N__28854),
            .I(N__28847));
    LocalMux I__5065 (
            .O(N__28851),
            .I(N__28844));
    InMux I__5064 (
            .O(N__28850),
            .I(N__28841));
    Odrv4 I__5063 (
            .O(N__28847),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.QiZ0Z_3 ));
    Odrv12 I__5062 (
            .O(N__28844),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.QiZ0Z_3 ));
    LocalMux I__5061 (
            .O(N__28841),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.QiZ0Z_3 ));
    InMux I__5060 (
            .O(N__28834),
            .I(N__28831));
    LocalMux I__5059 (
            .O(N__28831),
            .I(N__28828));
    Odrv12 I__5058 (
            .O(N__28828),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_s_3 ));
    InMux I__5057 (
            .O(N__28825),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_cry_2 ));
    InMux I__5056 (
            .O(N__28822),
            .I(N__28818));
    InMux I__5055 (
            .O(N__28821),
            .I(N__28815));
    LocalMux I__5054 (
            .O(N__28818),
            .I(N__28811));
    LocalMux I__5053 (
            .O(N__28815),
            .I(N__28808));
    InMux I__5052 (
            .O(N__28814),
            .I(N__28805));
    Odrv4 I__5051 (
            .O(N__28811),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.QiZ0Z_4 ));
    Odrv12 I__5050 (
            .O(N__28808),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.QiZ0Z_4 ));
    LocalMux I__5049 (
            .O(N__28805),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.QiZ0Z_4 ));
    CascadeMux I__5048 (
            .O(N__28798),
            .I(N__28795));
    InMux I__5047 (
            .O(N__28795),
            .I(N__28792));
    LocalMux I__5046 (
            .O(N__28792),
            .I(N__28789));
    Odrv4 I__5045 (
            .O(N__28789),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_s_4 ));
    InMux I__5044 (
            .O(N__28786),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_cry_3 ));
    InMux I__5043 (
            .O(N__28783),
            .I(N__28779));
    InMux I__5042 (
            .O(N__28782),
            .I(N__28776));
    LocalMux I__5041 (
            .O(N__28779),
            .I(N__28771));
    LocalMux I__5040 (
            .O(N__28776),
            .I(N__28771));
    Span4Mux_h I__5039 (
            .O(N__28771),
            .I(N__28768));
    Odrv4 I__5038 (
            .O(N__28768),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.QiZ0Z_5 ));
    CascadeMux I__5037 (
            .O(N__28765),
            .I(N__28762));
    InMux I__5036 (
            .O(N__28762),
            .I(N__28759));
    LocalMux I__5035 (
            .O(N__28759),
            .I(N__28756));
    Span4Mux_h I__5034 (
            .O(N__28756),
            .I(N__28753));
    Odrv4 I__5033 (
            .O(N__28753),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_s_5 ));
    InMux I__5032 (
            .O(N__28750),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_cry_4 ));
    InMux I__5031 (
            .O(N__28747),
            .I(N__28744));
    LocalMux I__5030 (
            .O(N__28744),
            .I(N__28740));
    InMux I__5029 (
            .O(N__28743),
            .I(N__28737));
    Odrv4 I__5028 (
            .O(N__28740),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.QiZ0Z_6 ));
    LocalMux I__5027 (
            .O(N__28737),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.QiZ0Z_6 ));
    CascadeMux I__5026 (
            .O(N__28732),
            .I(N__28724));
    CascadeMux I__5025 (
            .O(N__28731),
            .I(N__28721));
    CascadeMux I__5024 (
            .O(N__28730),
            .I(N__28718));
    CascadeMux I__5023 (
            .O(N__28729),
            .I(N__28715));
    CascadeMux I__5022 (
            .O(N__28728),
            .I(N__28712));
    CascadeMux I__5021 (
            .O(N__28727),
            .I(N__28709));
    InMux I__5020 (
            .O(N__28724),
            .I(N__28692));
    InMux I__5019 (
            .O(N__28721),
            .I(N__28692));
    InMux I__5018 (
            .O(N__28718),
            .I(N__28692));
    InMux I__5017 (
            .O(N__28715),
            .I(N__28685));
    InMux I__5016 (
            .O(N__28712),
            .I(N__28685));
    InMux I__5015 (
            .O(N__28709),
            .I(N__28685));
    InMux I__5014 (
            .O(N__28708),
            .I(N__28679));
    InMux I__5013 (
            .O(N__28707),
            .I(N__28674));
    InMux I__5012 (
            .O(N__28706),
            .I(N__28674));
    CascadeMux I__5011 (
            .O(N__28705),
            .I(N__28671));
    CascadeMux I__5010 (
            .O(N__28704),
            .I(N__28668));
    CascadeMux I__5009 (
            .O(N__28703),
            .I(N__28665));
    InMux I__5008 (
            .O(N__28702),
            .I(N__28662));
    CascadeMux I__5007 (
            .O(N__28701),
            .I(N__28659));
    CascadeMux I__5006 (
            .O(N__28700),
            .I(N__28656));
    CascadeMux I__5005 (
            .O(N__28699),
            .I(N__28653));
    LocalMux I__5004 (
            .O(N__28692),
            .I(N__28642));
    LocalMux I__5003 (
            .O(N__28685),
            .I(N__28642));
    CascadeMux I__5002 (
            .O(N__28684),
            .I(N__28638));
    CascadeMux I__5001 (
            .O(N__28683),
            .I(N__28634));
    CascadeMux I__5000 (
            .O(N__28682),
            .I(N__28630));
    LocalMux I__4999 (
            .O(N__28679),
            .I(N__28627));
    LocalMux I__4998 (
            .O(N__28674),
            .I(N__28624));
    InMux I__4997 (
            .O(N__28671),
            .I(N__28617));
    InMux I__4996 (
            .O(N__28668),
            .I(N__28617));
    InMux I__4995 (
            .O(N__28665),
            .I(N__28617));
    LocalMux I__4994 (
            .O(N__28662),
            .I(N__28614));
    InMux I__4993 (
            .O(N__28659),
            .I(N__28607));
    InMux I__4992 (
            .O(N__28656),
            .I(N__28607));
    InMux I__4991 (
            .O(N__28653),
            .I(N__28607));
    CascadeMux I__4990 (
            .O(N__28652),
            .I(N__28604));
    CascadeMux I__4989 (
            .O(N__28651),
            .I(N__28601));
    CascadeMux I__4988 (
            .O(N__28650),
            .I(N__28598));
    CascadeMux I__4987 (
            .O(N__28649),
            .I(N__28595));
    CascadeMux I__4986 (
            .O(N__28648),
            .I(N__28592));
    CascadeMux I__4985 (
            .O(N__28647),
            .I(N__28589));
    Span4Mux_v I__4984 (
            .O(N__28642),
            .I(N__28586));
    InMux I__4983 (
            .O(N__28641),
            .I(N__28562));
    InMux I__4982 (
            .O(N__28638),
            .I(N__28562));
    InMux I__4981 (
            .O(N__28637),
            .I(N__28562));
    InMux I__4980 (
            .O(N__28634),
            .I(N__28562));
    InMux I__4979 (
            .O(N__28633),
            .I(N__28562));
    InMux I__4978 (
            .O(N__28630),
            .I(N__28562));
    Span4Mux_v I__4977 (
            .O(N__28627),
            .I(N__28557));
    Span4Mux_v I__4976 (
            .O(N__28624),
            .I(N__28557));
    LocalMux I__4975 (
            .O(N__28617),
            .I(N__28554));
    Span4Mux_v I__4974 (
            .O(N__28614),
            .I(N__28549));
    LocalMux I__4973 (
            .O(N__28607),
            .I(N__28549));
    InMux I__4972 (
            .O(N__28604),
            .I(N__28542));
    InMux I__4971 (
            .O(N__28601),
            .I(N__28542));
    InMux I__4970 (
            .O(N__28598),
            .I(N__28542));
    InMux I__4969 (
            .O(N__28595),
            .I(N__28535));
    InMux I__4968 (
            .O(N__28592),
            .I(N__28535));
    InMux I__4967 (
            .O(N__28589),
            .I(N__28535));
    Span4Mux_h I__4966 (
            .O(N__28586),
            .I(N__28532));
    InMux I__4965 (
            .O(N__28585),
            .I(N__28527));
    InMux I__4964 (
            .O(N__28584),
            .I(N__28527));
    InMux I__4963 (
            .O(N__28583),
            .I(N__28524));
    CascadeMux I__4962 (
            .O(N__28582),
            .I(N__28520));
    CascadeMux I__4961 (
            .O(N__28581),
            .I(N__28516));
    CascadeMux I__4960 (
            .O(N__28580),
            .I(N__28512));
    CascadeMux I__4959 (
            .O(N__28579),
            .I(N__28504));
    CascadeMux I__4958 (
            .O(N__28578),
            .I(N__28501));
    CascadeMux I__4957 (
            .O(N__28577),
            .I(N__28497));
    CascadeMux I__4956 (
            .O(N__28576),
            .I(N__28494));
    CascadeMux I__4955 (
            .O(N__28575),
            .I(N__28491));
    LocalMux I__4954 (
            .O(N__28562),
            .I(N__28488));
    Span4Mux_h I__4953 (
            .O(N__28557),
            .I(N__28477));
    Span4Mux_h I__4952 (
            .O(N__28554),
            .I(N__28477));
    Span4Mux_h I__4951 (
            .O(N__28549),
            .I(N__28477));
    LocalMux I__4950 (
            .O(N__28542),
            .I(N__28477));
    LocalMux I__4949 (
            .O(N__28535),
            .I(N__28477));
    Span4Mux_h I__4948 (
            .O(N__28532),
            .I(N__28470));
    LocalMux I__4947 (
            .O(N__28527),
            .I(N__28470));
    LocalMux I__4946 (
            .O(N__28524),
            .I(N__28470));
    InMux I__4945 (
            .O(N__28523),
            .I(N__28457));
    InMux I__4944 (
            .O(N__28520),
            .I(N__28457));
    InMux I__4943 (
            .O(N__28519),
            .I(N__28457));
    InMux I__4942 (
            .O(N__28516),
            .I(N__28457));
    InMux I__4941 (
            .O(N__28515),
            .I(N__28457));
    InMux I__4940 (
            .O(N__28512),
            .I(N__28457));
    CascadeMux I__4939 (
            .O(N__28511),
            .I(N__28454));
    CascadeMux I__4938 (
            .O(N__28510),
            .I(N__28451));
    CascadeMux I__4937 (
            .O(N__28509),
            .I(N__28448));
    CascadeMux I__4936 (
            .O(N__28508),
            .I(N__28444));
    CascadeMux I__4935 (
            .O(N__28507),
            .I(N__28441));
    InMux I__4934 (
            .O(N__28504),
            .I(N__28432));
    InMux I__4933 (
            .O(N__28501),
            .I(N__28432));
    InMux I__4932 (
            .O(N__28500),
            .I(N__28432));
    InMux I__4931 (
            .O(N__28497),
            .I(N__28432));
    InMux I__4930 (
            .O(N__28494),
            .I(N__28427));
    InMux I__4929 (
            .O(N__28491),
            .I(N__28427));
    Span4Mux_v I__4928 (
            .O(N__28488),
            .I(N__28418));
    Span4Mux_h I__4927 (
            .O(N__28477),
            .I(N__28418));
    Span4Mux_v I__4926 (
            .O(N__28470),
            .I(N__28415));
    LocalMux I__4925 (
            .O(N__28457),
            .I(N__28412));
    InMux I__4924 (
            .O(N__28454),
            .I(N__28407));
    InMux I__4923 (
            .O(N__28451),
            .I(N__28407));
    InMux I__4922 (
            .O(N__28448),
            .I(N__28398));
    InMux I__4921 (
            .O(N__28447),
            .I(N__28398));
    InMux I__4920 (
            .O(N__28444),
            .I(N__28398));
    InMux I__4919 (
            .O(N__28441),
            .I(N__28398));
    LocalMux I__4918 (
            .O(N__28432),
            .I(N__28393));
    LocalMux I__4917 (
            .O(N__28427),
            .I(N__28393));
    InMux I__4916 (
            .O(N__28426),
            .I(N__28390));
    InMux I__4915 (
            .O(N__28425),
            .I(N__28383));
    InMux I__4914 (
            .O(N__28424),
            .I(N__28383));
    InMux I__4913 (
            .O(N__28423),
            .I(N__28383));
    Odrv4 I__4912 (
            .O(N__28418),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__4911 (
            .O(N__28415),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__4910 (
            .O(N__28412),
            .I(CONSTANT_ONE_NET));
    LocalMux I__4909 (
            .O(N__28407),
            .I(CONSTANT_ONE_NET));
    LocalMux I__4908 (
            .O(N__28398),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__4907 (
            .O(N__28393),
            .I(CONSTANT_ONE_NET));
    LocalMux I__4906 (
            .O(N__28390),
            .I(CONSTANT_ONE_NET));
    LocalMux I__4905 (
            .O(N__28383),
            .I(CONSTANT_ONE_NET));
    InMux I__4904 (
            .O(N__28366),
            .I(N__28363));
    LocalMux I__4903 (
            .O(N__28363),
            .I(N__28360));
    Odrv12 I__4902 (
            .O(N__28360),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_s_6 ));
    InMux I__4901 (
            .O(N__28357),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_cry_5 ));
    CascadeMux I__4900 (
            .O(N__28354),
            .I(N__28351));
    InMux I__4899 (
            .O(N__28351),
            .I(N__28348));
    LocalMux I__4898 (
            .O(N__28348),
            .I(N__28345));
    Span4Mux_v I__4897 (
            .O(N__28345),
            .I(N__28341));
    InMux I__4896 (
            .O(N__28344),
            .I(N__28338));
    Odrv4 I__4895 (
            .O(N__28341),
            .I(PIO_dport0_T2_4));
    LocalMux I__4894 (
            .O(N__28338),
            .I(PIO_dport0_T2_4));
    CascadeMux I__4893 (
            .O(N__28333),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI4VJTZ0Z_30_cascade_ ));
    InMux I__4892 (
            .O(N__28330),
            .I(N__28327));
    LocalMux I__4891 (
            .O(N__28327),
            .I(N__28324));
    Odrv12 I__4890 (
            .O(N__28324),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_30 ));
    InMux I__4889 (
            .O(N__28321),
            .I(N__28318));
    LocalMux I__4888 (
            .O(N__28318),
            .I(N__28315));
    Span4Mux_h I__4887 (
            .O(N__28315),
            .I(N__28312));
    Odrv4 I__4886 (
            .O(N__28312),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_30 ));
    InMux I__4885 (
            .O(N__28309),
            .I(N__28306));
    LocalMux I__4884 (
            .O(N__28306),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNISM2RZ0Z_30 ));
    CascadeMux I__4883 (
            .O(N__28303),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI0BBKZ0Z_30_cascade_ ));
    InMux I__4882 (
            .O(N__28300),
            .I(N__28297));
    LocalMux I__4881 (
            .O(N__28297),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_30 ));
    CEMux I__4880 (
            .O(N__28294),
            .I(N__28286));
    CEMux I__4879 (
            .O(N__28293),
            .I(N__28283));
    CEMux I__4878 (
            .O(N__28292),
            .I(N__28280));
    CEMux I__4877 (
            .O(N__28291),
            .I(N__28277));
    CEMux I__4876 (
            .O(N__28290),
            .I(N__28274));
    CEMux I__4875 (
            .O(N__28289),
            .I(N__28271));
    LocalMux I__4874 (
            .O(N__28286),
            .I(N__28264));
    LocalMux I__4873 (
            .O(N__28283),
            .I(N__28264));
    LocalMux I__4872 (
            .O(N__28280),
            .I(N__28264));
    LocalMux I__4871 (
            .O(N__28277),
            .I(N__28261));
    LocalMux I__4870 (
            .O(N__28274),
            .I(N__28257));
    LocalMux I__4869 (
            .O(N__28271),
            .I(N__28254));
    Span4Mux_v I__4868 (
            .O(N__28264),
            .I(N__28251));
    Span4Mux_h I__4867 (
            .O(N__28261),
            .I(N__28248));
    CEMux I__4866 (
            .O(N__28260),
            .I(N__28245));
    Span4Mux_v I__4865 (
            .O(N__28257),
            .I(N__28240));
    Span4Mux_h I__4864 (
            .O(N__28254),
            .I(N__28240));
    Span4Mux_h I__4863 (
            .O(N__28251),
            .I(N__28233));
    Span4Mux_v I__4862 (
            .O(N__28248),
            .I(N__28233));
    LocalMux I__4861 (
            .O(N__28245),
            .I(N__28233));
    Span4Mux_h I__4860 (
            .O(N__28240),
            .I(N__28230));
    Sp12to4 I__4859 (
            .O(N__28233),
            .I(N__28227));
    Odrv4 I__4858 (
            .O(N__28230),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_awe5 ));
    Odrv12 I__4857 (
            .O(N__28227),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_awe5 ));
    InMux I__4856 (
            .O(N__28222),
            .I(N__28219));
    LocalMux I__4855 (
            .O(N__28219),
            .I(N__28216));
    Odrv12 I__4854 (
            .O(N__28216),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_4 ));
    InMux I__4853 (
            .O(N__28213),
            .I(N__28210));
    LocalMux I__4852 (
            .O(N__28210),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_0 ));
    InMux I__4851 (
            .O(N__28207),
            .I(N__28204));
    LocalMux I__4850 (
            .O(N__28204),
            .I(N__28201));
    Odrv12 I__4849 (
            .O(N__28201),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_30 ));
    InMux I__4848 (
            .O(N__28198),
            .I(N__28195));
    LocalMux I__4847 (
            .O(N__28195),
            .I(N__28192));
    Span4Mux_v I__4846 (
            .O(N__28192),
            .I(N__28189));
    Odrv4 I__4845 (
            .O(N__28189),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_30 ));
    InMux I__4844 (
            .O(N__28186),
            .I(N__28183));
    LocalMux I__4843 (
            .O(N__28183),
            .I(N__28180));
    Span4Mux_v I__4842 (
            .O(N__28180),
            .I(N__28177));
    Odrv4 I__4841 (
            .O(N__28177),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_30 ));
    InMux I__4840 (
            .O(N__28174),
            .I(N__28171));
    LocalMux I__4839 (
            .O(N__28171),
            .I(N__28168));
    Span4Mux_h I__4838 (
            .O(N__28168),
            .I(N__28165));
    Odrv4 I__4837 (
            .O(N__28165),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_15 ));
    InMux I__4836 (
            .O(N__28162),
            .I(N__28159));
    LocalMux I__4835 (
            .O(N__28159),
            .I(N__28156));
    Span4Mux_s3_v I__4834 (
            .O(N__28156),
            .I(N__28153));
    Span4Mux_h I__4833 (
            .O(N__28153),
            .I(N__28150));
    Odrv4 I__4832 (
            .O(N__28150),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_31 ));
    CEMux I__4831 (
            .O(N__28147),
            .I(N__28142));
    CEMux I__4830 (
            .O(N__28146),
            .I(N__28139));
    CEMux I__4829 (
            .O(N__28145),
            .I(N__28134));
    LocalMux I__4828 (
            .O(N__28142),
            .I(N__28129));
    LocalMux I__4827 (
            .O(N__28139),
            .I(N__28129));
    CEMux I__4826 (
            .O(N__28138),
            .I(N__28126));
    CEMux I__4825 (
            .O(N__28137),
            .I(N__28123));
    LocalMux I__4824 (
            .O(N__28134),
            .I(N__28120));
    Span4Mux_s3_v I__4823 (
            .O(N__28129),
            .I(N__28115));
    LocalMux I__4822 (
            .O(N__28126),
            .I(N__28115));
    LocalMux I__4821 (
            .O(N__28123),
            .I(N__28112));
    Span4Mux_h I__4820 (
            .O(N__28120),
            .I(N__28107));
    Span4Mux_v I__4819 (
            .O(N__28115),
            .I(N__28107));
    Span4Mux_v I__4818 (
            .O(N__28112),
            .I(N__28104));
    Span4Mux_h I__4817 (
            .O(N__28107),
            .I(N__28101));
    Span4Mux_h I__4816 (
            .O(N__28104),
            .I(N__28098));
    Odrv4 I__4815 (
            .O(N__28101),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_awe3 ));
    Odrv4 I__4814 (
            .O(N__28098),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_awe3 ));
    InMux I__4813 (
            .O(N__28093),
            .I(N__28090));
    LocalMux I__4812 (
            .O(N__28090),
            .I(N__28087));
    Span4Mux_h I__4811 (
            .O(N__28087),
            .I(N__28084));
    Odrv4 I__4810 (
            .O(N__28084),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_19 ));
    InMux I__4809 (
            .O(N__28081),
            .I(N__28078));
    LocalMux I__4808 (
            .O(N__28078),
            .I(N__28075));
    Odrv12 I__4807 (
            .O(N__28075),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_20 ));
    InMux I__4806 (
            .O(N__28072),
            .I(N__28069));
    LocalMux I__4805 (
            .O(N__28069),
            .I(N__28066));
    Odrv12 I__4804 (
            .O(N__28066),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_20 ));
    InMux I__4803 (
            .O(N__28063),
            .I(N__28060));
    LocalMux I__4802 (
            .O(N__28060),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_15 ));
    CascadeMux I__4801 (
            .O(N__28057),
            .I(N__28054));
    InMux I__4800 (
            .O(N__28054),
            .I(N__28051));
    LocalMux I__4799 (
            .O(N__28051),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_8 ));
    InMux I__4798 (
            .O(N__28048),
            .I(N__28045));
    LocalMux I__4797 (
            .O(N__28045),
            .I(N__28042));
    Odrv12 I__4796 (
            .O(N__28042),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_2 ));
    InMux I__4795 (
            .O(N__28039),
            .I(N__28036));
    LocalMux I__4794 (
            .O(N__28036),
            .I(N__28033));
    Span4Mux_h I__4793 (
            .O(N__28033),
            .I(N__28030));
    Sp12to4 I__4792 (
            .O(N__28030),
            .I(N__28027));
    Odrv12 I__4791 (
            .O(N__28027),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI2PUQZ0Z_15 ));
    InMux I__4790 (
            .O(N__28024),
            .I(N__28021));
    LocalMux I__4789 (
            .O(N__28021),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_15 ));
    InMux I__4788 (
            .O(N__28018),
            .I(N__28015));
    LocalMux I__4787 (
            .O(N__28015),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_31 ));
    InMux I__4786 (
            .O(N__28012),
            .I(N__28009));
    LocalMux I__4785 (
            .O(N__28009),
            .I(N__28006));
    Odrv4 I__4784 (
            .O(N__28006),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_31 ));
    InMux I__4783 (
            .O(N__28003),
            .I(N__28000));
    LocalMux I__4782 (
            .O(N__28000),
            .I(N__27997));
    Span12Mux_s10_h I__4781 (
            .O(N__27997),
            .I(N__27994));
    Odrv12 I__4780 (
            .O(N__27994),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIUO2RZ0Z_31 ));
    InMux I__4779 (
            .O(N__27991),
            .I(N__27988));
    LocalMux I__4778 (
            .O(N__27988),
            .I(N__27985));
    Odrv4 I__4777 (
            .O(N__27985),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_24 ));
    InMux I__4776 (
            .O(N__27982),
            .I(N__27979));
    LocalMux I__4775 (
            .O(N__27979),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_24 ));
    InMux I__4774 (
            .O(N__27976),
            .I(N__27973));
    LocalMux I__4773 (
            .O(N__27973),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_8 ));
    InMux I__4772 (
            .O(N__27970),
            .I(N__27967));
    LocalMux I__4771 (
            .O(N__27967),
            .I(N__27964));
    Span4Mux_h I__4770 (
            .O(N__27964),
            .I(N__27961));
    Span4Mux_h I__4769 (
            .O(N__27961),
            .I(N__27958));
    Odrv4 I__4768 (
            .O(N__27958),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.N_1386_i ));
    InMux I__4767 (
            .O(N__27955),
            .I(N__27952));
    LocalMux I__4766 (
            .O(N__27952),
            .I(N__27949));
    Span4Mux_v I__4765 (
            .O(N__27949),
            .I(N__27946));
    Odrv4 I__4764 (
            .O(N__27946),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI2RHTZ0Z_20 ));
    InMux I__4763 (
            .O(N__27943),
            .I(N__27940));
    LocalMux I__4762 (
            .O(N__27940),
            .I(iQ_RNIA4HM1_2));
    CascadeMux I__4761 (
            .O(N__27937),
            .I(mem_mem_ram6__RNIULD71_20_cascade_));
    InMux I__4760 (
            .O(N__27934),
            .I(N__27931));
    LocalMux I__4759 (
            .O(N__27931),
            .I(N__27928));
    Odrv4 I__4758 (
            .O(N__27928),
            .I(\u0.N_1559 ));
    CascadeMux I__4757 (
            .O(N__27925),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIEDOD1Z0Z_2_cascade_ ));
    CascadeMux I__4756 (
            .O(N__27922),
            .I(DMAq_2_cascade_));
    InMux I__4755 (
            .O(N__27919),
            .I(N__27916));
    LocalMux I__4754 (
            .O(N__27916),
            .I(N__27913));
    Sp12to4 I__4753 (
            .O(N__27913),
            .I(N__27910));
    Odrv12 I__4752 (
            .O(N__27910),
            .I(\u0.dat_o_0_0_0_2 ));
    CascadeMux I__4751 (
            .O(N__27907),
            .I(\u0.dat_o_0_0_1Z0Z_2_cascade_ ));
    InMux I__4750 (
            .O(N__27904),
            .I(N__27901));
    LocalMux I__4749 (
            .O(N__27901),
            .I(N__27898));
    Odrv12 I__4748 (
            .O(N__27898),
            .I(\u0.dat_o_0_0_2_2 ));
    IoInMux I__4747 (
            .O(N__27895),
            .I(N__27892));
    LocalMux I__4746 (
            .O(N__27892),
            .I(N__27889));
    Span12Mux_s4_h I__4745 (
            .O(N__27889),
            .I(N__27886));
    Span12Mux_h I__4744 (
            .O(N__27886),
            .I(N__27883));
    Odrv12 I__4743 (
            .O(N__27883),
            .I(wb_dat_o_c_2));
    InMux I__4742 (
            .O(N__27880),
            .I(N__27877));
    LocalMux I__4741 (
            .O(N__27877),
            .I(PIOq_2));
    InMux I__4740 (
            .O(N__27874),
            .I(N__27871));
    LocalMux I__4739 (
            .O(N__27871),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIQ0CMZ0Z_2 ));
    InMux I__4738 (
            .O(N__27868),
            .I(N__27865));
    LocalMux I__4737 (
            .O(N__27865),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIASNK1Z0Z_2 ));
    CascadeMux I__4736 (
            .O(N__27862),
            .I(N__27859));
    InMux I__4735 (
            .O(N__27859),
            .I(N__27856));
    LocalMux I__4734 (
            .O(N__27856),
            .I(N__27852));
    InMux I__4733 (
            .O(N__27855),
            .I(N__27849));
    Span4Mux_h I__4732 (
            .O(N__27852),
            .I(N__27846));
    LocalMux I__4731 (
            .O(N__27849),
            .I(N__27843));
    Span4Mux_v I__4730 (
            .O(N__27846),
            .I(N__27838));
    Span4Mux_h I__4729 (
            .O(N__27843),
            .I(N__27838));
    Odrv4 I__4728 (
            .O(N__27838),
            .I(PIO_cmdport_T1_2));
    InMux I__4727 (
            .O(N__27835),
            .I(N__27832));
    LocalMux I__4726 (
            .O(N__27832),
            .I(N__27828));
    InMux I__4725 (
            .O(N__27831),
            .I(N__27825));
    Span4Mux_v I__4724 (
            .O(N__27828),
            .I(N__27822));
    LocalMux I__4723 (
            .O(N__27825),
            .I(N__27819));
    Odrv4 I__4722 (
            .O(N__27822),
            .I(PIO_dport0_IORDYen));
    Odrv12 I__4721 (
            .O(N__27819),
            .I(PIO_dport0_IORDYen));
    CascadeMux I__4720 (
            .O(N__27814),
            .I(N__27811));
    InMux I__4719 (
            .O(N__27811),
            .I(N__27808));
    LocalMux I__4718 (
            .O(N__27808),
            .I(N__27804));
    InMux I__4717 (
            .O(N__27807),
            .I(N__27801));
    Odrv12 I__4716 (
            .O(N__27804),
            .I(PIO_cmdport_T1_3));
    LocalMux I__4715 (
            .O(N__27801),
            .I(PIO_cmdport_T1_3));
    InMux I__4714 (
            .O(N__27796),
            .I(N__27793));
    LocalMux I__4713 (
            .O(N__27793),
            .I(N__27789));
    InMux I__4712 (
            .O(N__27792),
            .I(N__27786));
    Span4Mux_h I__4711 (
            .O(N__27789),
            .I(N__27783));
    LocalMux I__4710 (
            .O(N__27786),
            .I(N__27780));
    Sp12to4 I__4709 (
            .O(N__27783),
            .I(N__27775));
    Sp12to4 I__4708 (
            .O(N__27780),
            .I(N__27775));
    Odrv12 I__4707 (
            .O(N__27775),
            .I(PIO_dport1_IORDYen));
    InMux I__4706 (
            .O(N__27772),
            .I(N__27768));
    CascadeMux I__4705 (
            .O(N__27771),
            .I(N__27765));
    LocalMux I__4704 (
            .O(N__27768),
            .I(N__27762));
    InMux I__4703 (
            .O(N__27765),
            .I(N__27759));
    Span4Mux_v I__4702 (
            .O(N__27762),
            .I(N__27756));
    LocalMux I__4701 (
            .O(N__27759),
            .I(N__27753));
    Span4Mux_v I__4700 (
            .O(N__27756),
            .I(N__27750));
    Odrv12 I__4699 (
            .O(N__27753),
            .I(PIO_cmdport_T1_4));
    Odrv4 I__4698 (
            .O(N__27750),
            .I(PIO_cmdport_T1_4));
    CascadeMux I__4697 (
            .O(N__27745),
            .I(N__27739));
    InMux I__4696 (
            .O(N__27744),
            .I(N__27733));
    InMux I__4695 (
            .O(N__27743),
            .I(N__27733));
    InMux I__4694 (
            .O(N__27742),
            .I(N__27730));
    InMux I__4693 (
            .O(N__27739),
            .I(N__27727));
    InMux I__4692 (
            .O(N__27738),
            .I(N__27724));
    LocalMux I__4691 (
            .O(N__27733),
            .I(N__27719));
    LocalMux I__4690 (
            .O(N__27730),
            .I(N__27719));
    LocalMux I__4689 (
            .O(N__27727),
            .I(N__27716));
    LocalMux I__4688 (
            .O(N__27724),
            .I(N__27713));
    Span4Mux_v I__4687 (
            .O(N__27719),
            .I(N__27708));
    Span4Mux_v I__4686 (
            .O(N__27716),
            .I(N__27708));
    Span4Mux_v I__4685 (
            .O(N__27713),
            .I(N__27705));
    Span4Mux_h I__4684 (
            .O(N__27708),
            .I(N__27702));
    Odrv4 I__4683 (
            .O(N__27705),
            .I(IDEctrl_ppen));
    Odrv4 I__4682 (
            .O(N__27702),
            .I(IDEctrl_ppen));
    CascadeMux I__4681 (
            .O(N__27697),
            .I(N__27694));
    InMux I__4680 (
            .O(N__27694),
            .I(N__27691));
    LocalMux I__4679 (
            .O(N__27691),
            .I(N__27687));
    InMux I__4678 (
            .O(N__27690),
            .I(N__27684));
    Span4Mux_v I__4677 (
            .O(N__27687),
            .I(N__27678));
    LocalMux I__4676 (
            .O(N__27684),
            .I(N__27678));
    InMux I__4675 (
            .O(N__27683),
            .I(N__27675));
    Span4Mux_h I__4674 (
            .O(N__27678),
            .I(N__27672));
    LocalMux I__4673 (
            .O(N__27675),
            .I(N__27669));
    Span4Mux_v I__4672 (
            .O(N__27672),
            .I(N__27666));
    Span4Mux_h I__4671 (
            .O(N__27669),
            .I(N__27663));
    Odrv4 I__4670 (
            .O(N__27666),
            .I(IDEctrl_FATR0));
    Odrv4 I__4669 (
            .O(N__27663),
            .I(IDEctrl_FATR0));
    InMux I__4668 (
            .O(N__27658),
            .I(N__27655));
    LocalMux I__4667 (
            .O(N__27655),
            .I(N__27652));
    Span4Mux_v I__4666 (
            .O(N__27652),
            .I(N__27648));
    InMux I__4665 (
            .O(N__27651),
            .I(N__27645));
    Span4Mux_v I__4664 (
            .O(N__27648),
            .I(N__27642));
    LocalMux I__4663 (
            .O(N__27645),
            .I(N__27639));
    Odrv4 I__4662 (
            .O(N__27642),
            .I(PIO_cmdport_T1_1));
    Odrv12 I__4661 (
            .O(N__27639),
            .I(PIO_cmdport_T1_1));
    InMux I__4660 (
            .O(N__27634),
            .I(N__27631));
    LocalMux I__4659 (
            .O(N__27631),
            .I(N__27628));
    Span4Mux_h I__4658 (
            .O(N__27628),
            .I(N__27625));
    Span4Mux_h I__4657 (
            .O(N__27625),
            .I(N__27622));
    Odrv4 I__4656 (
            .O(N__27622),
            .I(\u0.CtrlRegZ0Z_20 ));
    CascadeMux I__4655 (
            .O(N__27619),
            .I(\u0.dat_o_0_a2_i_2_20_cascade_ ));
    IoInMux I__4654 (
            .O(N__27616),
            .I(N__27613));
    LocalMux I__4653 (
            .O(N__27613),
            .I(N__27610));
    IoSpan4Mux I__4652 (
            .O(N__27610),
            .I(N__27607));
    Span4Mux_s3_h I__4651 (
            .O(N__27607),
            .I(N__27604));
    Span4Mux_h I__4650 (
            .O(N__27604),
            .I(N__27601));
    Span4Mux_h I__4649 (
            .O(N__27601),
            .I(N__27598));
    Span4Mux_h I__4648 (
            .O(N__27598),
            .I(N__27595));
    Span4Mux_h I__4647 (
            .O(N__27595),
            .I(N__27592));
    Odrv4 I__4646 (
            .O(N__27592),
            .I(N_211_i));
    CascadeMux I__4645 (
            .O(N__27589),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIQI0RZ0Z_20_cascade_ ));
    CascadeMux I__4644 (
            .O(N__27586),
            .I(\u1.PIO_control.PIO_access_control.it4_1_iv_i_i_0_7_cascade_ ));
    InMux I__4643 (
            .O(N__27583),
            .I(N__27580));
    LocalMux I__4642 (
            .O(N__27580),
            .I(N__27577));
    Span4Mux_v I__4641 (
            .O(N__27577),
            .I(N__27574));
    Span4Mux_h I__4640 (
            .O(N__27574),
            .I(N__27571));
    Odrv4 I__4639 (
            .O(N__27571),
            .I(\u1.PIO_control.PIO_access_control.T4Z0Z_7 ));
    CascadeMux I__4638 (
            .O(N__27568),
            .I(\u1.PIO_control.PIO_access_control.iteoc_1_iv_i_i_0_5_cascade_ ));
    InMux I__4637 (
            .O(N__27565),
            .I(N__27562));
    LocalMux I__4636 (
            .O(N__27562),
            .I(N__27559));
    Span4Mux_v I__4635 (
            .O(N__27559),
            .I(N__27556));
    Span4Mux_h I__4634 (
            .O(N__27556),
            .I(N__27553));
    Odrv4 I__4633 (
            .O(N__27553),
            .I(\u1.PIO_control.PIO_access_control.TeocZ0Z_5 ));
    InMux I__4632 (
            .O(N__27550),
            .I(N__27547));
    LocalMux I__4631 (
            .O(N__27547),
            .I(\u1.PIO_control.PIO_access_control.iteoc_1_iv_i_i_0_2 ));
    InMux I__4630 (
            .O(N__27544),
            .I(N__27541));
    LocalMux I__4629 (
            .O(N__27541),
            .I(N__27538));
    Span4Mux_h I__4628 (
            .O(N__27538),
            .I(N__27535));
    Span4Mux_h I__4627 (
            .O(N__27535),
            .I(N__27532));
    Odrv4 I__4626 (
            .O(N__27532),
            .I(\u1.DMA_control.Teoc_3 ));
    CascadeMux I__4625 (
            .O(N__27529),
            .I(\u1.PIO_control.PIO_access_control.it2_1_iv_0_0_5_cascade_ ));
    InMux I__4624 (
            .O(N__27526),
            .I(N__27523));
    LocalMux I__4623 (
            .O(N__27523),
            .I(N__27520));
    Odrv12 I__4622 (
            .O(N__27520),
            .I(\u1.PIO_control.PIO_access_control.T2Z0Z_5 ));
    CascadeMux I__4621 (
            .O(N__27517),
            .I(\u1.PIO_control.PIO_access_control.it2_1_iv_i_i_0_6_cascade_ ));
    CascadeMux I__4620 (
            .O(N__27514),
            .I(N__27511));
    InMux I__4619 (
            .O(N__27511),
            .I(N__27508));
    LocalMux I__4618 (
            .O(N__27508),
            .I(\u1.PIO_control.PIO_access_control.T2Z0Z_6 ));
    CascadeMux I__4617 (
            .O(N__27505),
            .I(\u1.PIO_control.PIO_access_control.it2_1_iv_i_i_0_7_cascade_ ));
    InMux I__4616 (
            .O(N__27502),
            .I(N__27499));
    LocalMux I__4615 (
            .O(N__27499),
            .I(\u1.PIO_control.PIO_access_control.T2Z0Z_7 ));
    CascadeMux I__4614 (
            .O(N__27496),
            .I(\u1.PIO_control.PIO_access_control.it4_1_iv_0_0_0_cascade_ ));
    InMux I__4613 (
            .O(N__27493),
            .I(N__27490));
    LocalMux I__4612 (
            .O(N__27490),
            .I(N__27487));
    Sp12to4 I__4611 (
            .O(N__27487),
            .I(N__27484));
    Odrv12 I__4610 (
            .O(N__27484),
            .I(\u1.PIO_control.PIO_access_control.T4Z0Z_0 ));
    InMux I__4609 (
            .O(N__27481),
            .I(N__27478));
    LocalMux I__4608 (
            .O(N__27478),
            .I(N__27475));
    Span4Mux_s3_h I__4607 (
            .O(N__27475),
            .I(N__27472));
    Span4Mux_h I__4606 (
            .O(N__27472),
            .I(N__27469));
    Span4Mux_h I__4605 (
            .O(N__27469),
            .I(N__27466));
    Odrv4 I__4604 (
            .O(N__27466),
            .I(\u1.PIO_control.PIO_access_control.TeocZ0Z_2 ));
    CascadeMux I__4603 (
            .O(N__27463),
            .I(\u1.PIO_control.PIO_access_control.it2_1_iv_0_0_0_cascade_ ));
    InMux I__4602 (
            .O(N__27460),
            .I(N__27457));
    LocalMux I__4601 (
            .O(N__27457),
            .I(\u1.PIO_control.PIO_access_control.T2Z0Z_0 ));
    CascadeMux I__4600 (
            .O(N__27454),
            .I(\u1.PIO_control.PIO_access_control.it2_1_iv_i_i_0_1_cascade_ ));
    CascadeMux I__4599 (
            .O(N__27451),
            .I(N__27448));
    InMux I__4598 (
            .O(N__27448),
            .I(N__27445));
    LocalMux I__4597 (
            .O(N__27445),
            .I(\u1.PIO_control.PIO_access_control.T2Z0Z_1 ));
    CascadeMux I__4596 (
            .O(N__27442),
            .I(\u1.PIO_control.PIO_access_control.it2_1_iv_0_0_2_cascade_ ));
    InMux I__4595 (
            .O(N__27439),
            .I(N__27436));
    LocalMux I__4594 (
            .O(N__27436),
            .I(N__27433));
    Odrv12 I__4593 (
            .O(N__27433),
            .I(\u1.PIO_control.PIO_access_control.T2Z0Z_2 ));
    CascadeMux I__4592 (
            .O(N__27430),
            .I(\u1.PIO_control.PIO_access_control.it2_1_iv_i_i_0_3_cascade_ ));
    InMux I__4591 (
            .O(N__27427),
            .I(N__27424));
    LocalMux I__4590 (
            .O(N__27424),
            .I(N__27420));
    InMux I__4589 (
            .O(N__27423),
            .I(N__27417));
    Span4Mux_v I__4588 (
            .O(N__27420),
            .I(N__27414));
    LocalMux I__4587 (
            .O(N__27417),
            .I(N__27411));
    Span4Mux_v I__4586 (
            .O(N__27414),
            .I(N__27408));
    Span12Mux_h I__4585 (
            .O(N__27411),
            .I(N__27405));
    Span4Mux_v I__4584 (
            .O(N__27408),
            .I(N__27402));
    Span12Mux_v I__4583 (
            .O(N__27405),
            .I(N__27399));
    Odrv4 I__4582 (
            .O(N__27402),
            .I(PIO_dport0_T2_3));
    Odrv12 I__4581 (
            .O(N__27399),
            .I(PIO_dport0_T2_3));
    InMux I__4580 (
            .O(N__27394),
            .I(N__27391));
    LocalMux I__4579 (
            .O(N__27391),
            .I(\u1.PIO_control.PIO_access_control.T2Z0Z_3 ));
    InMux I__4578 (
            .O(N__27388),
            .I(N__27385));
    LocalMux I__4577 (
            .O(N__27385),
            .I(\u1.PIO_control.PIO_access_control.it2_1_iv_0_0_4 ));
    InMux I__4576 (
            .O(N__27382),
            .I(N__27379));
    LocalMux I__4575 (
            .O(N__27379),
            .I(\u1.PIO_control.PIO_access_control.it1_1_iv_i_i_0_7 ));
    CascadeMux I__4574 (
            .O(N__27376),
            .I(\u1.PIO_control.PIO_access_control.it1_1_iv_i_i_0_6_cascade_ ));
    InMux I__4573 (
            .O(N__27373),
            .I(N__27370));
    LocalMux I__4572 (
            .O(N__27370),
            .I(N__27367));
    Odrv12 I__4571 (
            .O(N__27367),
            .I(\u1.PIO_control.PIO_access_control.T1Z0Z_6 ));
    InMux I__4570 (
            .O(N__27364),
            .I(N__27360));
    InMux I__4569 (
            .O(N__27363),
            .I(N__27357));
    LocalMux I__4568 (
            .O(N__27360),
            .I(PIO_dport1_T2_4));
    LocalMux I__4567 (
            .O(N__27357),
            .I(PIO_dport1_T2_4));
    InMux I__4566 (
            .O(N__27352),
            .I(N__27349));
    LocalMux I__4565 (
            .O(N__27349),
            .I(N__27346));
    Odrv4 I__4564 (
            .O(N__27346),
            .I(\u1.PIO_control.PIO_access_control.T2Z0Z_4 ));
    InMux I__4563 (
            .O(N__27343),
            .I(N__27340));
    LocalMux I__4562 (
            .O(N__27340),
            .I(N__27337));
    Span4Mux_h I__4561 (
            .O(N__27337),
            .I(N__27334));
    Odrv4 I__4560 (
            .O(N__27334),
            .I(\u1.PIO_control.PIO_access_control.T1Z0Z_7 ));
    InMux I__4559 (
            .O(N__27331),
            .I(N__27328));
    LocalMux I__4558 (
            .O(N__27328),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_24 ));
    InMux I__4557 (
            .O(N__27325),
            .I(N__27322));
    LocalMux I__4556 (
            .O(N__27322),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_8 ));
    InMux I__4555 (
            .O(N__27319),
            .I(N__27316));
    LocalMux I__4554 (
            .O(N__27316),
            .I(N__27313));
    Odrv4 I__4553 (
            .O(N__27313),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_8 ));
    InMux I__4552 (
            .O(N__27310),
            .I(N__27307));
    LocalMux I__4551 (
            .O(N__27307),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_16 ));
    InMux I__4550 (
            .O(N__27304),
            .I(N__27301));
    LocalMux I__4549 (
            .O(N__27301),
            .I(N__27298));
    Odrv4 I__4548 (
            .O(N__27298),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_16 ));
    InMux I__4547 (
            .O(N__27295),
            .I(N__27292));
    LocalMux I__4546 (
            .O(N__27292),
            .I(N__27289));
    Odrv4 I__4545 (
            .O(N__27289),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_0 ));
    InMux I__4544 (
            .O(N__27286),
            .I(N__27283));
    LocalMux I__4543 (
            .O(N__27283),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_24 ));
    InMux I__4542 (
            .O(N__27280),
            .I(N__27277));
    LocalMux I__4541 (
            .O(N__27277),
            .I(N__27274));
    Span4Mux_h I__4540 (
            .O(N__27274),
            .I(N__27271));
    Span4Mux_v I__4539 (
            .O(N__27271),
            .I(N__27268));
    Odrv4 I__4538 (
            .O(N__27268),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_19 ));
    InMux I__4537 (
            .O(N__27265),
            .I(N__27262));
    LocalMux I__4536 (
            .O(N__27262),
            .I(N__27259));
    Odrv4 I__4535 (
            .O(N__27259),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_22 ));
    InMux I__4534 (
            .O(N__27256),
            .I(N__27253));
    LocalMux I__4533 (
            .O(N__27253),
            .I(N__27250));
    Span4Mux_v I__4532 (
            .O(N__27250),
            .I(N__27247));
    Odrv4 I__4531 (
            .O(N__27247),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_21 ));
    InMux I__4530 (
            .O(N__27244),
            .I(N__27241));
    LocalMux I__4529 (
            .O(N__27241),
            .I(N__27238));
    Odrv4 I__4528 (
            .O(N__27238),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_19 ));
    InMux I__4527 (
            .O(N__27235),
            .I(N__27232));
    LocalMux I__4526 (
            .O(N__27232),
            .I(N__27229));
    Span4Mux_v I__4525 (
            .O(N__27229),
            .I(N__27226));
    Odrv4 I__4524 (
            .O(N__27226),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_17 ));
    InMux I__4523 (
            .O(N__27223),
            .I(N__27220));
    LocalMux I__4522 (
            .O(N__27220),
            .I(N__27217));
    Span4Mux_h I__4521 (
            .O(N__27217),
            .I(N__27214));
    Odrv4 I__4520 (
            .O(N__27214),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_3 ));
    InMux I__4519 (
            .O(N__27211),
            .I(N__27208));
    LocalMux I__4518 (
            .O(N__27208),
            .I(N__27205));
    Span4Mux_v I__4517 (
            .O(N__27205),
            .I(N__27202));
    Odrv4 I__4516 (
            .O(N__27202),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_19 ));
    InMux I__4515 (
            .O(N__27199),
            .I(N__27196));
    LocalMux I__4514 (
            .O(N__27196),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_15 ));
    InMux I__4513 (
            .O(N__27193),
            .I(N__27190));
    LocalMux I__4512 (
            .O(N__27190),
            .I(N__27187));
    Span4Mux_v I__4511 (
            .O(N__27187),
            .I(N__27184));
    Odrv4 I__4510 (
            .O(N__27184),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_31 ));
    InMux I__4509 (
            .O(N__27181),
            .I(N__27178));
    LocalMux I__4508 (
            .O(N__27178),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_17 ));
    InMux I__4507 (
            .O(N__27175),
            .I(N__27172));
    LocalMux I__4506 (
            .O(N__27172),
            .I(N__27169));
    Odrv4 I__4505 (
            .O(N__27169),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_2 ));
    InMux I__4504 (
            .O(N__27166),
            .I(N__27163));
    LocalMux I__4503 (
            .O(N__27163),
            .I(N__27160));
    Odrv4 I__4502 (
            .O(N__27160),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_12 ));
    InMux I__4501 (
            .O(N__27157),
            .I(N__27154));
    LocalMux I__4500 (
            .O(N__27154),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_3 ));
    InMux I__4499 (
            .O(N__27151),
            .I(N__27148));
    LocalMux I__4498 (
            .O(N__27148),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_19 ));
    InMux I__4497 (
            .O(N__27145),
            .I(N__27142));
    LocalMux I__4496 (
            .O(N__27142),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_12 ));
    InMux I__4495 (
            .O(N__27139),
            .I(N__27136));
    LocalMux I__4494 (
            .O(N__27136),
            .I(N__27133));
    Odrv4 I__4493 (
            .O(N__27133),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_14 ));
    CascadeMux I__4492 (
            .O(N__27130),
            .I(N__27127));
    InMux I__4491 (
            .O(N__27127),
            .I(N__27124));
    LocalMux I__4490 (
            .O(N__27124),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_14 ));
    InMux I__4489 (
            .O(N__27121),
            .I(N__27118));
    LocalMux I__4488 (
            .O(N__27118),
            .I(N__27115));
    Span4Mux_v I__4487 (
            .O(N__27115),
            .I(N__27112));
    Odrv4 I__4486 (
            .O(N__27112),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_15 ));
    InMux I__4485 (
            .O(N__27109),
            .I(N__27106));
    LocalMux I__4484 (
            .O(N__27106),
            .I(N__27103));
    Span4Mux_h I__4483 (
            .O(N__27103),
            .I(N__27100));
    Odrv4 I__4482 (
            .O(N__27100),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIA1GTZ0Z_15 ));
    InMux I__4481 (
            .O(N__27097),
            .I(N__27094));
    LocalMux I__4480 (
            .O(N__27094),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_15 ));
    InMux I__4479 (
            .O(N__27091),
            .I(N__27088));
    LocalMux I__4478 (
            .O(N__27088),
            .I(N__27085));
    Span4Mux_v I__4477 (
            .O(N__27085),
            .I(N__27082));
    Odrv4 I__4476 (
            .O(N__27082),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_31 ));
    CascadeMux I__4475 (
            .O(N__27079),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI61KTZ0Z_31_cascade_ ));
    InMux I__4474 (
            .O(N__27076),
            .I(N__27073));
    LocalMux I__4473 (
            .O(N__27073),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_31 ));
    InMux I__4472 (
            .O(N__27070),
            .I(N__27067));
    LocalMux I__4471 (
            .O(N__27067),
            .I(N__27064));
    Span4Mux_v I__4470 (
            .O(N__27064),
            .I(N__27061));
    Odrv4 I__4469 (
            .O(N__27061),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI2DBKZ0Z_31 ));
    InMux I__4468 (
            .O(N__27058),
            .I(N__27055));
    LocalMux I__4467 (
            .O(N__27055),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI4VG71Z0Z_31 ));
    CascadeMux I__4466 (
            .O(N__27052),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIIGLM1Z0Z_2_cascade_ ));
    InMux I__4465 (
            .O(N__27049),
            .I(N__27046));
    LocalMux I__4464 (
            .O(N__27046),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_2 ));
    InMux I__4463 (
            .O(N__27043),
            .I(N__27040));
    LocalMux I__4462 (
            .O(N__27040),
            .I(N__27037));
    Span12Mux_h I__4461 (
            .O(N__27037),
            .I(N__27034));
    Odrv12 I__4460 (
            .O(N__27034),
            .I(\u1.DMAd_0 ));
    IoInMux I__4459 (
            .O(N__27031),
            .I(N__27028));
    LocalMux I__4458 (
            .O(N__27028),
            .I(N__27025));
    IoSpan4Mux I__4457 (
            .O(N__27025),
            .I(N__27022));
    Span4Mux_s2_v I__4456 (
            .O(N__27022),
            .I(N__27019));
    Sp12to4 I__4455 (
            .O(N__27019),
            .I(N__27016));
    Span12Mux_h I__4454 (
            .O(N__27016),
            .I(N__27013));
    Odrv12 I__4453 (
            .O(N__27013),
            .I(dd_pad_o_c_0));
    InMux I__4452 (
            .O(N__27010),
            .I(N__27007));
    LocalMux I__4451 (
            .O(N__27007),
            .I(N__27003));
    InMux I__4450 (
            .O(N__27006),
            .I(N__27000));
    Odrv4 I__4449 (
            .O(N__27003),
            .I(\u1.PIO_control.pong_a_3 ));
    LocalMux I__4448 (
            .O(N__27000),
            .I(\u1.PIO_control.pong_a_3 ));
    InMux I__4447 (
            .O(N__26995),
            .I(N__26992));
    LocalMux I__4446 (
            .O(N__26992),
            .I(N__26987));
    InMux I__4445 (
            .O(N__26991),
            .I(N__26982));
    InMux I__4444 (
            .O(N__26990),
            .I(N__26982));
    Odrv4 I__4443 (
            .O(N__26987),
            .I(\u1.PIO_control.ping_a_3 ));
    LocalMux I__4442 (
            .O(N__26982),
            .I(\u1.PIO_control.ping_a_3 ));
    CascadeMux I__4441 (
            .O(N__26977),
            .I(\u1.N_1425_cascade_ ));
    IoInMux I__4440 (
            .O(N__26974),
            .I(N__26971));
    LocalMux I__4439 (
            .O(N__26971),
            .I(N__26968));
    Span4Mux_s0_v I__4438 (
            .O(N__26968),
            .I(N__26965));
    Sp12to4 I__4437 (
            .O(N__26965),
            .I(N__26962));
    Span12Mux_h I__4436 (
            .O(N__26962),
            .I(N__26959));
    Odrv12 I__4435 (
            .O(N__26959),
            .I(cs0n_pad_o_c));
    InMux I__4434 (
            .O(N__26956),
            .I(N__26953));
    LocalMux I__4433 (
            .O(N__26953),
            .I(N__26950));
    Span4Mux_v I__4432 (
            .O(N__26950),
            .I(N__26947));
    Odrv4 I__4431 (
            .O(N__26947),
            .I(\u1.PIO_control.pong_d_0 ));
    InMux I__4430 (
            .O(N__26944),
            .I(N__26941));
    LocalMux I__4429 (
            .O(N__26941),
            .I(N__26938));
    Odrv4 I__4428 (
            .O(N__26938),
            .I(\u1.PIO_control.ping_d_0 ));
    InMux I__4427 (
            .O(N__26935),
            .I(N__26932));
    LocalMux I__4426 (
            .O(N__26932),
            .I(\u1.N_1426 ));
    InMux I__4425 (
            .O(N__26929),
            .I(N__26922));
    CascadeMux I__4424 (
            .O(N__26928),
            .I(N__26914));
    CascadeMux I__4423 (
            .O(N__26927),
            .I(N__26911));
    CascadeMux I__4422 (
            .O(N__26926),
            .I(N__26908));
    CascadeMux I__4421 (
            .O(N__26925),
            .I(N__26905));
    LocalMux I__4420 (
            .O(N__26922),
            .I(N__26900));
    InMux I__4419 (
            .O(N__26921),
            .I(N__26897));
    InMux I__4418 (
            .O(N__26920),
            .I(N__26879));
    InMux I__4417 (
            .O(N__26919),
            .I(N__26879));
    InMux I__4416 (
            .O(N__26918),
            .I(N__26879));
    InMux I__4415 (
            .O(N__26917),
            .I(N__26879));
    InMux I__4414 (
            .O(N__26914),
            .I(N__26867));
    InMux I__4413 (
            .O(N__26911),
            .I(N__26867));
    InMux I__4412 (
            .O(N__26908),
            .I(N__26867));
    InMux I__4411 (
            .O(N__26905),
            .I(N__26867));
    InMux I__4410 (
            .O(N__26904),
            .I(N__26862));
    InMux I__4409 (
            .O(N__26903),
            .I(N__26862));
    Span4Mux_h I__4408 (
            .O(N__26900),
            .I(N__26857));
    LocalMux I__4407 (
            .O(N__26897),
            .I(N__26857));
    InMux I__4406 (
            .O(N__26896),
            .I(N__26850));
    InMux I__4405 (
            .O(N__26895),
            .I(N__26841));
    InMux I__4404 (
            .O(N__26894),
            .I(N__26841));
    InMux I__4403 (
            .O(N__26893),
            .I(N__26841));
    InMux I__4402 (
            .O(N__26892),
            .I(N__26841));
    InMux I__4401 (
            .O(N__26891),
            .I(N__26832));
    InMux I__4400 (
            .O(N__26890),
            .I(N__26832));
    InMux I__4399 (
            .O(N__26889),
            .I(N__26832));
    InMux I__4398 (
            .O(N__26888),
            .I(N__26832));
    LocalMux I__4397 (
            .O(N__26879),
            .I(N__26829));
    InMux I__4396 (
            .O(N__26878),
            .I(N__26822));
    InMux I__4395 (
            .O(N__26877),
            .I(N__26822));
    InMux I__4394 (
            .O(N__26876),
            .I(N__26822));
    LocalMux I__4393 (
            .O(N__26867),
            .I(N__26819));
    LocalMux I__4392 (
            .O(N__26862),
            .I(N__26814));
    Span4Mux_v I__4391 (
            .O(N__26857),
            .I(N__26814));
    InMux I__4390 (
            .O(N__26856),
            .I(N__26805));
    InMux I__4389 (
            .O(N__26855),
            .I(N__26805));
    InMux I__4388 (
            .O(N__26854),
            .I(N__26805));
    InMux I__4387 (
            .O(N__26853),
            .I(N__26805));
    LocalMux I__4386 (
            .O(N__26850),
            .I(N__26802));
    LocalMux I__4385 (
            .O(N__26841),
            .I(N__26795));
    LocalMux I__4384 (
            .O(N__26832),
            .I(N__26795));
    Sp12to4 I__4383 (
            .O(N__26829),
            .I(N__26795));
    LocalMux I__4382 (
            .O(N__26822),
            .I(N__26785));
    Span12Mux_s9_h I__4381 (
            .O(N__26819),
            .I(N__26785));
    Sp12to4 I__4380 (
            .O(N__26814),
            .I(N__26776));
    LocalMux I__4379 (
            .O(N__26805),
            .I(N__26776));
    Span12Mux_s4_h I__4378 (
            .O(N__26802),
            .I(N__26776));
    Span12Mux_v I__4377 (
            .O(N__26795),
            .I(N__26776));
    InMux I__4376 (
            .O(N__26794),
            .I(N__26769));
    InMux I__4375 (
            .O(N__26793),
            .I(N__26769));
    InMux I__4374 (
            .O(N__26792),
            .I(N__26769));
    InMux I__4373 (
            .O(N__26791),
            .I(N__26764));
    InMux I__4372 (
            .O(N__26790),
            .I(N__26764));
    Odrv12 I__4371 (
            .O(N__26785),
            .I(\u1.rpp ));
    Odrv12 I__4370 (
            .O(N__26776),
            .I(\u1.rpp ));
    LocalMux I__4369 (
            .O(N__26769),
            .I(\u1.rpp ));
    LocalMux I__4368 (
            .O(N__26764),
            .I(\u1.rpp ));
    CascadeMux I__4367 (
            .O(N__26755),
            .I(N__26752));
    InMux I__4366 (
            .O(N__26752),
            .I(N__26749));
    LocalMux I__4365 (
            .O(N__26749),
            .I(N__26746));
    Odrv4 I__4364 (
            .O(N__26746),
            .I(\u1.PIO_control.ping_d_1 ));
    InMux I__4363 (
            .O(N__26743),
            .I(N__26740));
    LocalMux I__4362 (
            .O(N__26740),
            .I(N__26737));
    Span4Mux_h I__4361 (
            .O(N__26737),
            .I(N__26734));
    Odrv4 I__4360 (
            .O(N__26734),
            .I(\u1.PIO_control.pong_d_1 ));
    CascadeMux I__4359 (
            .O(N__26731),
            .I(\u1.N_1427_cascade_ ));
    InMux I__4358 (
            .O(N__26728),
            .I(N__26725));
    LocalMux I__4357 (
            .O(N__26725),
            .I(N__26722));
    Span4Mux_h I__4356 (
            .O(N__26722),
            .I(N__26719));
    Span4Mux_v I__4355 (
            .O(N__26719),
            .I(N__26716));
    Odrv4 I__4354 (
            .O(N__26716),
            .I(\u1.DMAd_1 ));
    IoInMux I__4353 (
            .O(N__26713),
            .I(N__26710));
    LocalMux I__4352 (
            .O(N__26710),
            .I(N__26707));
    Span12Mux_s10_v I__4351 (
            .O(N__26707),
            .I(N__26704));
    Odrv12 I__4350 (
            .O(N__26704),
            .I(dd_pad_o_c_1));
    InMux I__4349 (
            .O(N__26701),
            .I(N__26698));
    LocalMux I__4348 (
            .O(N__26698),
            .I(\u1.N_1425 ));
    IoInMux I__4347 (
            .O(N__26695),
            .I(N__26692));
    LocalMux I__4346 (
            .O(N__26692),
            .I(N__26689));
    Span12Mux_s10_v I__4345 (
            .O(N__26689),
            .I(N__26686));
    Odrv12 I__4344 (
            .O(N__26686),
            .I(cs1n_pad_o_c));
    InMux I__4343 (
            .O(N__26683),
            .I(N__26680));
    LocalMux I__4342 (
            .O(N__26680),
            .I(N__26674));
    InMux I__4341 (
            .O(N__26679),
            .I(N__26671));
    InMux I__4340 (
            .O(N__26678),
            .I(N__26668));
    InMux I__4339 (
            .O(N__26677),
            .I(N__26665));
    Odrv4 I__4338 (
            .O(N__26674),
            .I(\u1.PIO_control.N_1315 ));
    LocalMux I__4337 (
            .O(N__26671),
            .I(\u1.PIO_control.N_1315 ));
    LocalMux I__4336 (
            .O(N__26668),
            .I(\u1.PIO_control.N_1315 ));
    LocalMux I__4335 (
            .O(N__26665),
            .I(\u1.PIO_control.N_1315 ));
    CascadeMux I__4334 (
            .O(N__26656),
            .I(\u1.PIO_control.PIO_access_control.N_2112_cascade_ ));
    InMux I__4333 (
            .O(N__26653),
            .I(N__26650));
    LocalMux I__4332 (
            .O(N__26650),
            .I(N__26647));
    Odrv12 I__4331 (
            .O(N__26647),
            .I(\u1.PIO_control.PIO_access_control.iteoc_1_iv_i_i_0_7 ));
    CascadeMux I__4330 (
            .O(N__26644),
            .I(\u1.PIO_control.PIO_access_control.it4_1_iv_i_i_0_2_cascade_ ));
    InMux I__4329 (
            .O(N__26641),
            .I(N__26638));
    LocalMux I__4328 (
            .O(N__26638),
            .I(N__26635));
    Span4Mux_h I__4327 (
            .O(N__26635),
            .I(N__26632));
    Span4Mux_h I__4326 (
            .O(N__26632),
            .I(N__26629));
    Odrv4 I__4325 (
            .O(N__26629),
            .I(\u1.PIO_control.PIO_access_control.T4Z0Z_2 ));
    CascadeMux I__4324 (
            .O(N__26626),
            .I(\u1.PIO_control.PIO_access_control.it4_1_iv_i_i_0_3_cascade_ ));
    InMux I__4323 (
            .O(N__26623),
            .I(N__26620));
    LocalMux I__4322 (
            .O(N__26620),
            .I(N__26617));
    Span12Mux_v I__4321 (
            .O(N__26617),
            .I(N__26614));
    Odrv12 I__4320 (
            .O(N__26614),
            .I(\u1.PIO_control.PIO_access_control.T4Z0Z_3 ));
    CascadeMux I__4319 (
            .O(N__26611),
            .I(\u1.PIO_control.PIO_access_control.it4_1_iv_0_0_4_cascade_ ));
    InMux I__4318 (
            .O(N__26608),
            .I(N__26605));
    LocalMux I__4317 (
            .O(N__26605),
            .I(N__26602));
    Span4Mux_h I__4316 (
            .O(N__26602),
            .I(N__26599));
    Span4Mux_h I__4315 (
            .O(N__26599),
            .I(N__26596));
    Odrv4 I__4314 (
            .O(N__26596),
            .I(\u1.PIO_control.PIO_access_control.T4Z0Z_4 ));
    CascadeMux I__4313 (
            .O(N__26593),
            .I(\u1.PIO_control.PIO_access_control.it4_1_iv_i_i_0_5_cascade_ ));
    InMux I__4312 (
            .O(N__26590),
            .I(N__26587));
    LocalMux I__4311 (
            .O(N__26587),
            .I(N__26584));
    Span4Mux_h I__4310 (
            .O(N__26584),
            .I(N__26581));
    Span4Mux_h I__4309 (
            .O(N__26581),
            .I(N__26578));
    Odrv4 I__4308 (
            .O(N__26578),
            .I(\u1.PIO_control.PIO_access_control.T4Z0Z_5 ));
    InMux I__4307 (
            .O(N__26575),
            .I(N__26571));
    InMux I__4306 (
            .O(N__26574),
            .I(N__26568));
    LocalMux I__4305 (
            .O(N__26571),
            .I(\u1.PIO_control.pong_a_1 ));
    LocalMux I__4304 (
            .O(N__26568),
            .I(\u1.PIO_control.pong_a_1 ));
    CascadeMux I__4303 (
            .O(N__26563),
            .I(\u1.PIO_control.PIO_access_control.it4_1_iv_i_i_o2_0_x0Z0Z_2_cascade_ ));
    InMux I__4302 (
            .O(N__26560),
            .I(N__26557));
    LocalMux I__4301 (
            .O(N__26557),
            .I(\u1.PIO_control.PIO_access_control.it4_1_iv_i_i_o2_0_x1Z0Z_2 ));
    CascadeMux I__4300 (
            .O(N__26554),
            .I(\u1.PIO_control.PIO_access_control.it4_1_iv_i_i_o2_0_2_cascade_ ));
    CascadeMux I__4299 (
            .O(N__26551),
            .I(\u1.PIO_control.PIO_access_control.it4_1_iv_i_i_o3_x0Z0Z_2_cascade_ ));
    CascadeMux I__4298 (
            .O(N__26548),
            .I(\u1.PIO_control.PIO_access_control.iiordyen_1_iv_i_i_0_cascade_ ));
    InMux I__4297 (
            .O(N__26545),
            .I(N__26542));
    LocalMux I__4296 (
            .O(N__26542),
            .I(N__26539));
    Span4Mux_h I__4295 (
            .O(N__26539),
            .I(N__26536));
    Span4Mux_h I__4294 (
            .O(N__26536),
            .I(N__26533));
    Odrv4 I__4293 (
            .O(N__26533),
            .I(\u1.PIO_control.PIO_access_control.IORDYenZ0 ));
    CascadeMux I__4292 (
            .O(N__26530),
            .I(\u1.PIO_control.PIO_access_control.it1_1_iv_i_i_0_1_cascade_ ));
    InMux I__4291 (
            .O(N__26527),
            .I(N__26524));
    LocalMux I__4290 (
            .O(N__26524),
            .I(N__26521));
    Span4Mux_v I__4289 (
            .O(N__26521),
            .I(N__26518));
    Span4Mux_h I__4288 (
            .O(N__26518),
            .I(N__26515));
    Odrv4 I__4287 (
            .O(N__26515),
            .I(\u1.PIO_control.PIO_access_control.T1Z0Z_1 ));
    InMux I__4286 (
            .O(N__26512),
            .I(N__26509));
    LocalMux I__4285 (
            .O(N__26509),
            .I(N__26506));
    Span4Mux_v I__4284 (
            .O(N__26506),
            .I(N__26503));
    Sp12to4 I__4283 (
            .O(N__26503),
            .I(N__26500));
    Span12Mux_s8_h I__4282 (
            .O(N__26500),
            .I(N__26497));
    Odrv12 I__4281 (
            .O(N__26497),
            .I(\u1.DMA_control.Td_1 ));
    InMux I__4280 (
            .O(N__26494),
            .I(N__26490));
    InMux I__4279 (
            .O(N__26493),
            .I(N__26487));
    LocalMux I__4278 (
            .O(N__26490),
            .I(\u1.PIO_control.PIO_access_control.it4_1_iv_i_i_o2_0_2 ));
    LocalMux I__4277 (
            .O(N__26487),
            .I(\u1.PIO_control.PIO_access_control.it4_1_iv_i_i_o2_0_2 ));
    CascadeMux I__4276 (
            .O(N__26482),
            .I(\u1.PIO_control.PIO_access_control.N_2110_cascade_ ));
    InMux I__4275 (
            .O(N__26479),
            .I(N__26476));
    LocalMux I__4274 (
            .O(N__26476),
            .I(\u1.PIO_control.PIO_access_control.it1_1_iv_i_i_0_5 ));
    InMux I__4273 (
            .O(N__26473),
            .I(N__26455));
    InMux I__4272 (
            .O(N__26472),
            .I(N__26455));
    InMux I__4271 (
            .O(N__26471),
            .I(N__26455));
    InMux I__4270 (
            .O(N__26470),
            .I(N__26455));
    InMux I__4269 (
            .O(N__26469),
            .I(N__26455));
    InMux I__4268 (
            .O(N__26468),
            .I(N__26455));
    LocalMux I__4267 (
            .O(N__26455),
            .I(N__26452));
    Span4Mux_h I__4266 (
            .O(N__26452),
            .I(N__26447));
    InMux I__4265 (
            .O(N__26451),
            .I(N__26442));
    InMux I__4264 (
            .O(N__26450),
            .I(N__26442));
    Odrv4 I__4263 (
            .O(N__26447),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_1_sqmuxa_i ));
    LocalMux I__4262 (
            .O(N__26442),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_1_sqmuxa_i ));
    CEMux I__4261 (
            .O(N__26437),
            .I(N__26434));
    LocalMux I__4260 (
            .O(N__26434),
            .I(N__26431));
    Span4Mux_h I__4259 (
            .O(N__26431),
            .I(N__26428));
    Span4Mux_h I__4258 (
            .O(N__26428),
            .I(N__26424));
    CEMux I__4257 (
            .O(N__26427),
            .I(N__26421));
    Odrv4 I__4256 (
            .O(N__26424),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qie_0_iZ0 ));
    LocalMux I__4255 (
            .O(N__26421),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qie_0_iZ0 ));
    InMux I__4254 (
            .O(N__26416),
            .I(N__26412));
    InMux I__4253 (
            .O(N__26415),
            .I(N__26409));
    LocalMux I__4252 (
            .O(N__26412),
            .I(\u1.pong_a_0 ));
    LocalMux I__4251 (
            .O(N__26409),
            .I(\u1.pong_a_0 ));
    CascadeMux I__4250 (
            .O(N__26404),
            .I(N__26400));
    InMux I__4249 (
            .O(N__26403),
            .I(N__26396));
    InMux I__4248 (
            .O(N__26400),
            .I(N__26391));
    InMux I__4247 (
            .O(N__26399),
            .I(N__26391));
    LocalMux I__4246 (
            .O(N__26396),
            .I(\u1.ping_a_0 ));
    LocalMux I__4245 (
            .O(N__26391),
            .I(\u1.ping_a_0 ));
    IoInMux I__4244 (
            .O(N__26386),
            .I(N__26383));
    LocalMux I__4243 (
            .O(N__26383),
            .I(N__26380));
    IoSpan4Mux I__4242 (
            .O(N__26380),
            .I(N__26377));
    Span4Mux_s3_h I__4241 (
            .O(N__26377),
            .I(N__26374));
    Sp12to4 I__4240 (
            .O(N__26374),
            .I(N__26371));
    Span12Mux_h I__4239 (
            .O(N__26371),
            .I(N__26368));
    Odrv12 I__4238 (
            .O(N__26368),
            .I(da_pad_o_c_0));
    InMux I__4237 (
            .O(N__26365),
            .I(N__26361));
    InMux I__4236 (
            .O(N__26364),
            .I(N__26357));
    LocalMux I__4235 (
            .O(N__26361),
            .I(N__26354));
    InMux I__4234 (
            .O(N__26360),
            .I(N__26351));
    LocalMux I__4233 (
            .O(N__26357),
            .I(N__26348));
    Span4Mux_h I__4232 (
            .O(N__26354),
            .I(N__26345));
    LocalMux I__4231 (
            .O(N__26351),
            .I(N__26341));
    Span4Mux_v I__4230 (
            .O(N__26348),
            .I(N__26336));
    Span4Mux_h I__4229 (
            .O(N__26345),
            .I(N__26336));
    InMux I__4228 (
            .O(N__26344),
            .I(N__26333));
    Odrv12 I__4227 (
            .O(N__26341),
            .I(\u1.PIO_control.N_1450 ));
    Odrv4 I__4226 (
            .O(N__26336),
            .I(\u1.PIO_control.N_1450 ));
    LocalMux I__4225 (
            .O(N__26333),
            .I(\u1.PIO_control.N_1450 ));
    CascadeMux I__4224 (
            .O(N__26326),
            .I(N__26323));
    InMux I__4223 (
            .O(N__26323),
            .I(N__26320));
    LocalMux I__4222 (
            .O(N__26320),
            .I(N__26317));
    Span4Mux_h I__4221 (
            .O(N__26317),
            .I(N__26314));
    Span4Mux_h I__4220 (
            .O(N__26314),
            .I(N__26311));
    Odrv4 I__4219 (
            .O(N__26311),
            .I(\u1.PIO_control.rpp_2_i_0 ));
    InMux I__4218 (
            .O(N__26308),
            .I(N__26304));
    InMux I__4217 (
            .O(N__26307),
            .I(N__26301));
    LocalMux I__4216 (
            .O(N__26304),
            .I(N__26298));
    LocalMux I__4215 (
            .O(N__26301),
            .I(N__26292));
    Span4Mux_h I__4214 (
            .O(N__26298),
            .I(N__26289));
    InMux I__4213 (
            .O(N__26297),
            .I(N__26282));
    InMux I__4212 (
            .O(N__26296),
            .I(N__26282));
    InMux I__4211 (
            .O(N__26295),
            .I(N__26282));
    Odrv12 I__4210 (
            .O(N__26292),
            .I(\u1.PIOdone_i ));
    Odrv4 I__4209 (
            .O(N__26289),
            .I(\u1.PIOdone_i ));
    LocalMux I__4208 (
            .O(N__26282),
            .I(\u1.PIOdone_i ));
    InMux I__4207 (
            .O(N__26275),
            .I(N__26268));
    InMux I__4206 (
            .O(N__26274),
            .I(N__26268));
    InMux I__4205 (
            .O(N__26273),
            .I(N__26265));
    LocalMux I__4204 (
            .O(N__26268),
            .I(N__26262));
    LocalMux I__4203 (
            .O(N__26265),
            .I(\u1.PIO_control.ping_a_1 ));
    Odrv4 I__4202 (
            .O(N__26262),
            .I(\u1.PIO_control.ping_a_1 ));
    CascadeMux I__4201 (
            .O(N__26257),
            .I(N__26254));
    InMux I__4200 (
            .O(N__26254),
            .I(N__26249));
    InMux I__4199 (
            .O(N__26253),
            .I(N__26246));
    InMux I__4198 (
            .O(N__26252),
            .I(N__26243));
    LocalMux I__4197 (
            .O(N__26249),
            .I(N__26240));
    LocalMux I__4196 (
            .O(N__26246),
            .I(\u1.pong_a_2 ));
    LocalMux I__4195 (
            .O(N__26243),
            .I(\u1.pong_a_2 ));
    Odrv12 I__4194 (
            .O(N__26240),
            .I(\u1.pong_a_2 ));
    InMux I__4193 (
            .O(N__26233),
            .I(N__26227));
    InMux I__4192 (
            .O(N__26232),
            .I(N__26227));
    LocalMux I__4191 (
            .O(N__26227),
            .I(N__26223));
    CascadeMux I__4190 (
            .O(N__26226),
            .I(N__26220));
    Span4Mux_h I__4189 (
            .O(N__26223),
            .I(N__26216));
    InMux I__4188 (
            .O(N__26220),
            .I(N__26211));
    InMux I__4187 (
            .O(N__26219),
            .I(N__26211));
    Odrv4 I__4186 (
            .O(N__26216),
            .I(\u1.ping_a_2 ));
    LocalMux I__4185 (
            .O(N__26211),
            .I(\u1.ping_a_2 ));
    CascadeMux I__4184 (
            .O(N__26206),
            .I(\u1.PIO_control.PIO_access_control.iteoc_1_iv_0_0_6_cascade_ ));
    InMux I__4183 (
            .O(N__26203),
            .I(N__26200));
    LocalMux I__4182 (
            .O(N__26200),
            .I(N__26197));
    Span4Mux_s3_h I__4181 (
            .O(N__26197),
            .I(N__26194));
    Span4Mux_h I__4180 (
            .O(N__26194),
            .I(N__26191));
    Odrv4 I__4179 (
            .O(N__26191),
            .I(\u1.PIO_control.PIO_access_control.TeocZ0Z_6 ));
    InMux I__4178 (
            .O(N__26188),
            .I(N__26185));
    LocalMux I__4177 (
            .O(N__26185),
            .I(N__26182));
    Span4Mux_h I__4176 (
            .O(N__26182),
            .I(N__26179));
    Odrv4 I__4175 (
            .O(N__26179),
            .I(\u1.PIO_control.PIO_access_control.T1Z0Z_5 ));
    InMux I__4174 (
            .O(N__26176),
            .I(N__26173));
    LocalMux I__4173 (
            .O(N__26173),
            .I(N__26170));
    Sp12to4 I__4172 (
            .O(N__26170),
            .I(N__26167));
    Odrv12 I__4171 (
            .O(N__26167),
            .I(\u1.PIO_control.PIO_access_control.TeocZ0Z_7 ));
    CascadeMux I__4170 (
            .O(N__26164),
            .I(\u1.PIO_control.PIO_access_control.it1_1_iv_i_i_0_3_cascade_ ));
    InMux I__4169 (
            .O(N__26161),
            .I(N__26158));
    LocalMux I__4168 (
            .O(N__26158),
            .I(N__26155));
    Span4Mux_h I__4167 (
            .O(N__26155),
            .I(N__26152));
    Odrv4 I__4166 (
            .O(N__26152),
            .I(\u1.PIO_control.PIO_access_control.T1Z0Z_3 ));
    InMux I__4165 (
            .O(N__26149),
            .I(N__26146));
    LocalMux I__4164 (
            .O(N__26146),
            .I(\u1.PIO_control.PIO_access_control.it1_1_iv_0_0_2 ));
    InMux I__4163 (
            .O(N__26143),
            .I(N__26140));
    LocalMux I__4162 (
            .O(N__26140),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_s_0 ));
    InMux I__4161 (
            .O(N__26137),
            .I(N__26134));
    LocalMux I__4160 (
            .O(N__26134),
            .I(N__26131));
    Span12Mux_s2_v I__4159 (
            .O(N__26131),
            .I(N__26128));
    Odrv12 I__4158 (
            .O(N__26128),
            .I(\u0.dat_o_0_0_3_13 ));
    CascadeMux I__4157 (
            .O(N__26125),
            .I(N__26122));
    InMux I__4156 (
            .O(N__26122),
            .I(N__26119));
    LocalMux I__4155 (
            .O(N__26119),
            .I(N__26116));
    Odrv12 I__4154 (
            .O(N__26116),
            .I(\u0.dat_o_0_0_0_13 ));
    InMux I__4153 (
            .O(N__26113),
            .I(N__26110));
    LocalMux I__4152 (
            .O(N__26110),
            .I(N__26107));
    Span4Mux_s3_v I__4151 (
            .O(N__26107),
            .I(N__26104));
    Sp12to4 I__4150 (
            .O(N__26104),
            .I(N__26101));
    Span12Mux_h I__4149 (
            .O(N__26101),
            .I(N__26098));
    Odrv12 I__4148 (
            .O(N__26098),
            .I(\u0.dat_o_0_0_2_13 ));
    IoInMux I__4147 (
            .O(N__26095),
            .I(N__26092));
    LocalMux I__4146 (
            .O(N__26092),
            .I(N__26089));
    Span4Mux_s0_v I__4145 (
            .O(N__26089),
            .I(N__26086));
    Span4Mux_h I__4144 (
            .O(N__26086),
            .I(N__26083));
    Odrv4 I__4143 (
            .O(N__26083),
            .I(wb_dat_o_c_13));
    InMux I__4142 (
            .O(N__26080),
            .I(N__26075));
    InMux I__4141 (
            .O(N__26079),
            .I(N__26070));
    InMux I__4140 (
            .O(N__26078),
            .I(N__26070));
    LocalMux I__4139 (
            .O(N__26075),
            .I(N__26065));
    LocalMux I__4138 (
            .O(N__26070),
            .I(N__26062));
    InMux I__4137 (
            .O(N__26069),
            .I(N__26057));
    InMux I__4136 (
            .O(N__26068),
            .I(N__26057));
    Span4Mux_h I__4135 (
            .O(N__26065),
            .I(N__26053));
    Span4Mux_h I__4134 (
            .O(N__26062),
            .I(N__26048));
    LocalMux I__4133 (
            .O(N__26057),
            .I(N__26048));
    InMux I__4132 (
            .O(N__26056),
            .I(N__26045));
    Odrv4 I__4131 (
            .O(N__26053),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.Qi_0_0 ));
    Odrv4 I__4130 (
            .O(N__26048),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.Qi_0_0 ));
    LocalMux I__4129 (
            .O(N__26045),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.Qi_0_0 ));
    InMux I__4128 (
            .O(N__26038),
            .I(N__26035));
    LocalMux I__4127 (
            .O(N__26035),
            .I(N__26032));
    Span4Mux_v I__4126 (
            .O(N__26032),
            .I(N__26029));
    Odrv4 I__4125 (
            .O(N__26029),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_s_0 ));
    CascadeMux I__4124 (
            .O(N__26026),
            .I(N__26023));
    InMux I__4123 (
            .O(N__26023),
            .I(N__26020));
    LocalMux I__4122 (
            .O(N__26020),
            .I(N__26017));
    Span4Mux_h I__4121 (
            .O(N__26017),
            .I(N__26014));
    Span4Mux_v I__4120 (
            .O(N__26014),
            .I(N__26011));
    Span4Mux_h I__4119 (
            .O(N__26011),
            .I(N__26008));
    Odrv4 I__4118 (
            .O(N__26008),
            .I(\u0.int_3_i_0_0 ));
    InMux I__4117 (
            .O(N__26005),
            .I(N__26002));
    LocalMux I__4116 (
            .O(N__26002),
            .I(N__25999));
    Span4Mux_v I__4115 (
            .O(N__25999),
            .I(N__25995));
    CascadeMux I__4114 (
            .O(N__25998),
            .I(N__25992));
    Span4Mux_h I__4113 (
            .O(N__25995),
            .I(N__25989));
    InMux I__4112 (
            .O(N__25992),
            .I(N__25986));
    Odrv4 I__4111 (
            .O(N__25989),
            .I(PIO_dport1_T1_0));
    LocalMux I__4110 (
            .O(N__25986),
            .I(PIO_dport1_T1_0));
    InMux I__4109 (
            .O(N__25981),
            .I(N__25978));
    LocalMux I__4108 (
            .O(N__25978),
            .I(\u1.PIO_control.PIO_access_control.it1_1_iv_i_i_0_0 ));
    InMux I__4107 (
            .O(N__25975),
            .I(N__25972));
    LocalMux I__4106 (
            .O(N__25972),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_22 ));
    InMux I__4105 (
            .O(N__25969),
            .I(N__25966));
    LocalMux I__4104 (
            .O(N__25966),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_31 ));
    InMux I__4103 (
            .O(N__25963),
            .I(N__25960));
    LocalMux I__4102 (
            .O(N__25960),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_15 ));
    InMux I__4101 (
            .O(N__25957),
            .I(N__25954));
    LocalMux I__4100 (
            .O(N__25954),
            .I(N__25951));
    Span4Mux_v I__4099 (
            .O(N__25951),
            .I(N__25948));
    Span4Mux_v I__4098 (
            .O(N__25948),
            .I(N__25945));
    Odrv4 I__4097 (
            .O(N__25945),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI6D7KZ0Z_15 ));
    InMux I__4096 (
            .O(N__25942),
            .I(N__25939));
    LocalMux I__4095 (
            .O(N__25939),
            .I(N__25936));
    Odrv12 I__4094 (
            .O(N__25936),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_4 ));
    InMux I__4093 (
            .O(N__25933),
            .I(N__25930));
    LocalMux I__4092 (
            .O(N__25930),
            .I(N__25927));
    Odrv4 I__4091 (
            .O(N__25927),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_5 ));
    InMux I__4090 (
            .O(N__25924),
            .I(N__25921));
    LocalMux I__4089 (
            .O(N__25921),
            .I(N__25918));
    Span4Mux_h I__4088 (
            .O(N__25918),
            .I(N__25915));
    Odrv4 I__4087 (
            .O(N__25915),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_6 ));
    InMux I__4086 (
            .O(N__25912),
            .I(N__25909));
    LocalMux I__4085 (
            .O(N__25909),
            .I(N__25906));
    Span4Mux_v I__4084 (
            .O(N__25906),
            .I(N__25903));
    Odrv4 I__4083 (
            .O(N__25903),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_22 ));
    InMux I__4082 (
            .O(N__25900),
            .I(N__25897));
    LocalMux I__4081 (
            .O(N__25897),
            .I(N__25894));
    Odrv4 I__4080 (
            .O(N__25894),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_21 ));
    InMux I__4079 (
            .O(N__25891),
            .I(N__25888));
    LocalMux I__4078 (
            .O(N__25888),
            .I(N__25885));
    Odrv12 I__4077 (
            .O(N__25885),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_3 ));
    InMux I__4076 (
            .O(N__25882),
            .I(N__25878));
    InMux I__4075 (
            .O(N__25881),
            .I(N__25875));
    LocalMux I__4074 (
            .O(N__25878),
            .I(N__25872));
    LocalMux I__4073 (
            .O(N__25875),
            .I(N__25869));
    Span12Mux_h I__4072 (
            .O(N__25872),
            .I(N__25866));
    Odrv4 I__4071 (
            .O(N__25869),
            .I(\u1.DMA_control.TxbufQ_18 ));
    Odrv12 I__4070 (
            .O(N__25866),
            .I(\u1.DMA_control.TxbufQ_18 ));
    CascadeMux I__4069 (
            .O(N__25861),
            .I(N__25858));
    InMux I__4068 (
            .O(N__25858),
            .I(N__25855));
    LocalMux I__4067 (
            .O(N__25855),
            .I(N__25852));
    Span4Mux_h I__4066 (
            .O(N__25852),
            .I(N__25849));
    Odrv4 I__4065 (
            .O(N__25849),
            .I(\u1.DMA_control.writeDlw_2 ));
    InMux I__4064 (
            .O(N__25846),
            .I(N__25842));
    InMux I__4063 (
            .O(N__25845),
            .I(N__25839));
    LocalMux I__4062 (
            .O(N__25842),
            .I(N__25836));
    LocalMux I__4061 (
            .O(N__25839),
            .I(N__25833));
    Span4Mux_h I__4060 (
            .O(N__25836),
            .I(N__25830));
    Span12Mux_h I__4059 (
            .O(N__25833),
            .I(N__25827));
    Odrv4 I__4058 (
            .O(N__25830),
            .I(\u1.DMA_control.TxbufQ_10 ));
    Odrv12 I__4057 (
            .O(N__25827),
            .I(\u1.DMA_control.TxbufQ_10 ));
    CascadeMux I__4056 (
            .O(N__25822),
            .I(\u1.DMA_control.writeDfw_6_i_0_2_cascade_ ));
    InMux I__4055 (
            .O(N__25819),
            .I(N__25816));
    LocalMux I__4054 (
            .O(N__25816),
            .I(N__25813));
    Span4Mux_h I__4053 (
            .O(N__25813),
            .I(N__25810));
    Span4Mux_h I__4052 (
            .O(N__25810),
            .I(N__25807));
    Odrv4 I__4051 (
            .O(N__25807),
            .I(\u1.DMAd_2 ));
    InMux I__4050 (
            .O(N__25804),
            .I(N__25800));
    InMux I__4049 (
            .O(N__25803),
            .I(N__25797));
    LocalMux I__4048 (
            .O(N__25800),
            .I(N__25794));
    LocalMux I__4047 (
            .O(N__25797),
            .I(N__25791));
    Span4Mux_h I__4046 (
            .O(N__25794),
            .I(N__25788));
    Odrv4 I__4045 (
            .O(N__25791),
            .I(\u1.DMA_control.TxbufQ_19 ));
    Odrv4 I__4044 (
            .O(N__25788),
            .I(\u1.DMA_control.TxbufQ_19 ));
    CascadeMux I__4043 (
            .O(N__25783),
            .I(N__25780));
    InMux I__4042 (
            .O(N__25780),
            .I(N__25777));
    LocalMux I__4041 (
            .O(N__25777),
            .I(N__25774));
    Span4Mux_v I__4040 (
            .O(N__25774),
            .I(N__25771));
    Odrv4 I__4039 (
            .O(N__25771),
            .I(\u1.DMA_control.writeDlw_3 ));
    InMux I__4038 (
            .O(N__25768),
            .I(N__25765));
    LocalMux I__4037 (
            .O(N__25765),
            .I(N__25762));
    Sp12to4 I__4036 (
            .O(N__25762),
            .I(N__25758));
    InMux I__4035 (
            .O(N__25761),
            .I(N__25755));
    Odrv12 I__4034 (
            .O(N__25758),
            .I(\u1.DMA_control.TxbufQ_11 ));
    LocalMux I__4033 (
            .O(N__25755),
            .I(\u1.DMA_control.TxbufQ_11 ));
    CascadeMux I__4032 (
            .O(N__25750),
            .I(\u1.DMA_control.writeDfw_6_i_0_3_cascade_ ));
    InMux I__4031 (
            .O(N__25747),
            .I(N__25744));
    LocalMux I__4030 (
            .O(N__25744),
            .I(N__25741));
    Span4Mux_v I__4029 (
            .O(N__25741),
            .I(N__25738));
    Span4Mux_h I__4028 (
            .O(N__25738),
            .I(N__25735));
    Odrv4 I__4027 (
            .O(N__25735),
            .I(\u1.DMAd_3 ));
    InMux I__4026 (
            .O(N__25732),
            .I(N__25729));
    LocalMux I__4025 (
            .O(N__25729),
            .I(N__25725));
    InMux I__4024 (
            .O(N__25728),
            .I(N__25722));
    Span4Mux_h I__4023 (
            .O(N__25725),
            .I(N__25719));
    LocalMux I__4022 (
            .O(N__25722),
            .I(N__25716));
    Span4Mux_h I__4021 (
            .O(N__25719),
            .I(N__25713));
    Odrv4 I__4020 (
            .O(N__25716),
            .I(\u1.DMA_control.TxbufQ_20 ));
    Odrv4 I__4019 (
            .O(N__25713),
            .I(\u1.DMA_control.TxbufQ_20 ));
    CascadeMux I__4018 (
            .O(N__25708),
            .I(N__25705));
    InMux I__4017 (
            .O(N__25705),
            .I(N__25702));
    LocalMux I__4016 (
            .O(N__25702),
            .I(N__25699));
    Span4Mux_v I__4015 (
            .O(N__25699),
            .I(N__25696));
    Odrv4 I__4014 (
            .O(N__25696),
            .I(\u1.DMA_control.writeDlw_4 ));
    InMux I__4013 (
            .O(N__25693),
            .I(N__25690));
    LocalMux I__4012 (
            .O(N__25690),
            .I(\u1.DMA_control.writeDfw_6_i_0_4 ));
    InMux I__4011 (
            .O(N__25687),
            .I(N__25684));
    LocalMux I__4010 (
            .O(N__25684),
            .I(N__25681));
    Span4Mux_h I__4009 (
            .O(N__25681),
            .I(N__25678));
    Odrv4 I__4008 (
            .O(N__25678),
            .I(\u1.DMA_control.writeDlw_15 ));
    InMux I__4007 (
            .O(N__25675),
            .I(N__25671));
    InMux I__4006 (
            .O(N__25674),
            .I(N__25668));
    LocalMux I__4005 (
            .O(N__25671),
            .I(N__25665));
    LocalMux I__4004 (
            .O(N__25668),
            .I(N__25662));
    Span12Mux_s8_v I__4003 (
            .O(N__25665),
            .I(N__25659));
    Odrv4 I__4002 (
            .O(N__25662),
            .I(\u1.DMA_control.TxbufQ_31 ));
    Odrv12 I__4001 (
            .O(N__25659),
            .I(\u1.DMA_control.TxbufQ_31 ));
    InMux I__4000 (
            .O(N__25654),
            .I(N__25651));
    LocalMux I__3999 (
            .O(N__25651),
            .I(N__25648));
    Span4Mux_h I__3998 (
            .O(N__25648),
            .I(N__25644));
    InMux I__3997 (
            .O(N__25647),
            .I(N__25641));
    Span4Mux_h I__3996 (
            .O(N__25644),
            .I(N__25638));
    LocalMux I__3995 (
            .O(N__25641),
            .I(N__25635));
    Odrv4 I__3994 (
            .O(N__25638),
            .I(\u1.DMA_control.TxbufQ_7 ));
    Odrv4 I__3993 (
            .O(N__25635),
            .I(\u1.DMA_control.TxbufQ_7 ));
    CascadeMux I__3992 (
            .O(N__25630),
            .I(N__25626));
    CascadeMux I__3991 (
            .O(N__25629),
            .I(N__25615));
    InMux I__3990 (
            .O(N__25626),
            .I(N__25604));
    InMux I__3989 (
            .O(N__25625),
            .I(N__25597));
    InMux I__3988 (
            .O(N__25624),
            .I(N__25597));
    InMux I__3987 (
            .O(N__25623),
            .I(N__25597));
    CascadeMux I__3986 (
            .O(N__25622),
            .I(N__25594));
    InMux I__3985 (
            .O(N__25621),
            .I(N__25589));
    InMux I__3984 (
            .O(N__25620),
            .I(N__25589));
    CascadeMux I__3983 (
            .O(N__25619),
            .I(N__25586));
    InMux I__3982 (
            .O(N__25618),
            .I(N__25574));
    InMux I__3981 (
            .O(N__25615),
            .I(N__25574));
    InMux I__3980 (
            .O(N__25614),
            .I(N__25574));
    InMux I__3979 (
            .O(N__25613),
            .I(N__25574));
    InMux I__3978 (
            .O(N__25612),
            .I(N__25574));
    CascadeMux I__3977 (
            .O(N__25611),
            .I(N__25564));
    CascadeMux I__3976 (
            .O(N__25610),
            .I(N__25558));
    CascadeMux I__3975 (
            .O(N__25609),
            .I(N__25555));
    CascadeMux I__3974 (
            .O(N__25608),
            .I(N__25552));
    CEMux I__3973 (
            .O(N__25607),
            .I(N__25546));
    LocalMux I__3972 (
            .O(N__25604),
            .I(N__25543));
    LocalMux I__3971 (
            .O(N__25597),
            .I(N__25540));
    InMux I__3970 (
            .O(N__25594),
            .I(N__25537));
    LocalMux I__3969 (
            .O(N__25589),
            .I(N__25534));
    InMux I__3968 (
            .O(N__25586),
            .I(N__25531));
    CascadeMux I__3967 (
            .O(N__25585),
            .I(N__25524));
    LocalMux I__3966 (
            .O(N__25574),
            .I(N__25521));
    InMux I__3965 (
            .O(N__25573),
            .I(N__25506));
    InMux I__3964 (
            .O(N__25572),
            .I(N__25506));
    InMux I__3963 (
            .O(N__25571),
            .I(N__25506));
    InMux I__3962 (
            .O(N__25570),
            .I(N__25506));
    InMux I__3961 (
            .O(N__25569),
            .I(N__25506));
    InMux I__3960 (
            .O(N__25568),
            .I(N__25506));
    InMux I__3959 (
            .O(N__25567),
            .I(N__25506));
    InMux I__3958 (
            .O(N__25564),
            .I(N__25489));
    InMux I__3957 (
            .O(N__25563),
            .I(N__25489));
    InMux I__3956 (
            .O(N__25562),
            .I(N__25489));
    InMux I__3955 (
            .O(N__25561),
            .I(N__25489));
    InMux I__3954 (
            .O(N__25558),
            .I(N__25489));
    InMux I__3953 (
            .O(N__25555),
            .I(N__25489));
    InMux I__3952 (
            .O(N__25552),
            .I(N__25489));
    InMux I__3951 (
            .O(N__25551),
            .I(N__25489));
    InMux I__3950 (
            .O(N__25550),
            .I(N__25486));
    CEMux I__3949 (
            .O(N__25549),
            .I(N__25483));
    LocalMux I__3948 (
            .O(N__25546),
            .I(N__25480));
    Span4Mux_h I__3947 (
            .O(N__25543),
            .I(N__25477));
    Span4Mux_h I__3946 (
            .O(N__25540),
            .I(N__25472));
    LocalMux I__3945 (
            .O(N__25537),
            .I(N__25472));
    Span4Mux_v I__3944 (
            .O(N__25534),
            .I(N__25467));
    LocalMux I__3943 (
            .O(N__25531),
            .I(N__25467));
    InMux I__3942 (
            .O(N__25530),
            .I(N__25462));
    InMux I__3941 (
            .O(N__25529),
            .I(N__25462));
    InMux I__3940 (
            .O(N__25528),
            .I(N__25455));
    InMux I__3939 (
            .O(N__25527),
            .I(N__25455));
    InMux I__3938 (
            .O(N__25524),
            .I(N__25455));
    Span4Mux_v I__3937 (
            .O(N__25521),
            .I(N__25452));
    LocalMux I__3936 (
            .O(N__25506),
            .I(N__25445));
    LocalMux I__3935 (
            .O(N__25489),
            .I(N__25445));
    LocalMux I__3934 (
            .O(N__25486),
            .I(N__25445));
    LocalMux I__3933 (
            .O(N__25483),
            .I(N__25442));
    Span4Mux_h I__3932 (
            .O(N__25480),
            .I(N__25439));
    Span4Mux_v I__3931 (
            .O(N__25477),
            .I(N__25432));
    Span4Mux_v I__3930 (
            .O(N__25472),
            .I(N__25432));
    Span4Mux_v I__3929 (
            .O(N__25467),
            .I(N__25432));
    LocalMux I__3928 (
            .O(N__25462),
            .I(N__25423));
    LocalMux I__3927 (
            .O(N__25455),
            .I(N__25423));
    Span4Mux_h I__3926 (
            .O(N__25452),
            .I(N__25423));
    Span4Mux_v I__3925 (
            .O(N__25445),
            .I(N__25423));
    Odrv12 I__3924 (
            .O(N__25442),
            .I(\u1.DMA_control.TxRdZ0 ));
    Odrv4 I__3923 (
            .O(N__25439),
            .I(\u1.DMA_control.TxRdZ0 ));
    Odrv4 I__3922 (
            .O(N__25432),
            .I(\u1.DMA_control.TxRdZ0 ));
    Odrv4 I__3921 (
            .O(N__25423),
            .I(\u1.DMA_control.TxRdZ0 ));
    CascadeMux I__3920 (
            .O(N__25414),
            .I(\u1.DMA_control.writeDfw_6_i_m3_i_0_15_cascade_ ));
    InMux I__3919 (
            .O(N__25411),
            .I(N__25408));
    LocalMux I__3918 (
            .O(N__25408),
            .I(N__25405));
    Span4Mux_h I__3917 (
            .O(N__25405),
            .I(N__25402));
    Span4Mux_h I__3916 (
            .O(N__25402),
            .I(N__25399));
    Odrv4 I__3915 (
            .O(N__25399),
            .I(\u1.DMAd_15 ));
    CEMux I__3914 (
            .O(N__25396),
            .I(N__25392));
    CEMux I__3913 (
            .O(N__25395),
            .I(N__25388));
    LocalMux I__3912 (
            .O(N__25392),
            .I(N__25385));
    CEMux I__3911 (
            .O(N__25391),
            .I(N__25382));
    LocalMux I__3910 (
            .O(N__25388),
            .I(N__25378));
    Span4Mux_h I__3909 (
            .O(N__25385),
            .I(N__25373));
    LocalMux I__3908 (
            .O(N__25382),
            .I(N__25373));
    CEMux I__3907 (
            .O(N__25381),
            .I(N__25370));
    Span4Mux_v I__3906 (
            .O(N__25378),
            .I(N__25367));
    Sp12to4 I__3905 (
            .O(N__25373),
            .I(N__25364));
    LocalMux I__3904 (
            .O(N__25370),
            .I(N__25361));
    Odrv4 I__3903 (
            .O(N__25367),
            .I(\u1.DMA_control.N_53 ));
    Odrv12 I__3902 (
            .O(N__25364),
            .I(\u1.DMA_control.N_53 ));
    Odrv4 I__3901 (
            .O(N__25361),
            .I(\u1.DMA_control.N_53 ));
    InMux I__3900 (
            .O(N__25354),
            .I(N__25351));
    LocalMux I__3899 (
            .O(N__25351),
            .I(N__25348));
    Odrv4 I__3898 (
            .O(N__25348),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_20 ));
    InMux I__3897 (
            .O(N__25345),
            .I(N__25342));
    LocalMux I__3896 (
            .O(N__25342),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_20 ));
    InMux I__3895 (
            .O(N__25339),
            .I(N__25336));
    LocalMux I__3894 (
            .O(N__25336),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_21 ));
    InMux I__3893 (
            .O(N__25333),
            .I(N__25330));
    LocalMux I__3892 (
            .O(N__25330),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_22 ));
    CascadeMux I__3891 (
            .O(N__25327),
            .I(N__25324));
    InMux I__3890 (
            .O(N__25324),
            .I(N__25321));
    LocalMux I__3889 (
            .O(N__25321),
            .I(N__25318));
    Span4Mux_h I__3888 (
            .O(N__25318),
            .I(N__25314));
    InMux I__3887 (
            .O(N__25317),
            .I(N__25311));
    Odrv4 I__3886 (
            .O(N__25314),
            .I(\u1.DMA_control.TxbufQ_12 ));
    LocalMux I__3885 (
            .O(N__25311),
            .I(\u1.DMA_control.TxbufQ_12 ));
    InMux I__3884 (
            .O(N__25306),
            .I(N__25303));
    LocalMux I__3883 (
            .O(N__25303),
            .I(N__25300));
    Span4Mux_h I__3882 (
            .O(N__25300),
            .I(N__25297));
    Odrv4 I__3881 (
            .O(N__25297),
            .I(\u1.DMAd_4 ));
    InMux I__3880 (
            .O(N__25294),
            .I(N__25291));
    LocalMux I__3879 (
            .O(N__25291),
            .I(N__25288));
    Span4Mux_v I__3878 (
            .O(N__25288),
            .I(N__25285));
    Span4Mux_h I__3877 (
            .O(N__25285),
            .I(N__25282));
    Span4Mux_h I__3876 (
            .O(N__25282),
            .I(N__25279));
    Odrv4 I__3875 (
            .O(N__25279),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNII9GTZ0Z_19 ));
    InMux I__3874 (
            .O(N__25276),
            .I(N__25273));
    LocalMux I__3873 (
            .O(N__25273),
            .I(mem_mem_ram6__RNIMBB71_19));
    InMux I__3872 (
            .O(N__25270),
            .I(N__25267));
    LocalMux I__3871 (
            .O(N__25267),
            .I(\u0.CtrlRegZ0Z_19 ));
    CascadeMux I__3870 (
            .O(N__25264),
            .I(\u0.dat_o_i_0_2_19_cascade_ ));
    InMux I__3869 (
            .O(N__25261),
            .I(N__25258));
    LocalMux I__3868 (
            .O(N__25258),
            .I(\u0.N_1724 ));
    IoInMux I__3867 (
            .O(N__25255),
            .I(N__25252));
    LocalMux I__3866 (
            .O(N__25252),
            .I(N__25249));
    IoSpan4Mux I__3865 (
            .O(N__25249),
            .I(N__25246));
    Span4Mux_s2_h I__3864 (
            .O(N__25246),
            .I(N__25243));
    Sp12to4 I__3863 (
            .O(N__25243),
            .I(N__25240));
    Span12Mux_s11_h I__3862 (
            .O(N__25240),
            .I(N__25237));
    Span12Mux_h I__3861 (
            .O(N__25237),
            .I(N__25234));
    Odrv12 I__3860 (
            .O(N__25234),
            .I(N_327_i));
    InMux I__3859 (
            .O(N__25231),
            .I(N__25225));
    InMux I__3858 (
            .O(N__25230),
            .I(N__25225));
    LocalMux I__3857 (
            .O(N__25225),
            .I(N__25222));
    Span4Mux_v I__3856 (
            .O(N__25222),
            .I(N__25218));
    InMux I__3855 (
            .O(N__25221),
            .I(N__25215));
    Span4Mux_h I__3854 (
            .O(N__25218),
            .I(N__25212));
    LocalMux I__3853 (
            .O(N__25215),
            .I(N__25209));
    Span4Mux_h I__3852 (
            .O(N__25212),
            .I(N__25204));
    Span4Mux_v I__3851 (
            .O(N__25209),
            .I(N__25204));
    Span4Mux_v I__3850 (
            .O(N__25204),
            .I(N__25201));
    Odrv4 I__3849 (
            .O(N__25201),
            .I(dd_pad_i_c_12));
    InMux I__3848 (
            .O(N__25198),
            .I(N__25195));
    LocalMux I__3847 (
            .O(N__25195),
            .I(N__25192));
    Span4Mux_v I__3846 (
            .O(N__25192),
            .I(N__25189));
    Odrv4 I__3845 (
            .O(N__25189),
            .I(\u0.dat_o_0_0_3_15 ));
    CascadeMux I__3844 (
            .O(N__25186),
            .I(\u0.dat_o_0_0_5_15_cascade_ ));
    IoInMux I__3843 (
            .O(N__25183),
            .I(N__25180));
    LocalMux I__3842 (
            .O(N__25180),
            .I(N__25177));
    IoSpan4Mux I__3841 (
            .O(N__25177),
            .I(N__25174));
    Span4Mux_s2_h I__3840 (
            .O(N__25174),
            .I(N__25171));
    Sp12to4 I__3839 (
            .O(N__25171),
            .I(N__25168));
    Span12Mux_s11_h I__3838 (
            .O(N__25168),
            .I(N__25165));
    Span12Mux_h I__3837 (
            .O(N__25165),
            .I(N__25162));
    Odrv12 I__3836 (
            .O(N__25162),
            .I(wb_dat_o_c_15));
    CascadeMux I__3835 (
            .O(N__25159),
            .I(mem_mem_ram6__RNIAVA71_15_cascade_));
    InMux I__3834 (
            .O(N__25156),
            .I(N__25153));
    LocalMux I__3833 (
            .O(N__25153),
            .I(\u0.N_2029 ));
    InMux I__3832 (
            .O(N__25150),
            .I(N__25147));
    LocalMux I__3831 (
            .O(N__25147),
            .I(iQ_RNIQGDM1_2));
    InMux I__3830 (
            .O(N__25144),
            .I(N__25141));
    LocalMux I__3829 (
            .O(N__25141),
            .I(PIOq_15));
    InMux I__3828 (
            .O(N__25138),
            .I(N__25135));
    LocalMux I__3827 (
            .O(N__25135),
            .I(N__25132));
    Span4Mux_h I__3826 (
            .O(N__25132),
            .I(N__25129));
    Span4Mux_v I__3825 (
            .O(N__25129),
            .I(N__25126));
    Odrv4 I__3824 (
            .O(N__25126),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIEL7KZ0Z_19 ));
    CascadeMux I__3823 (
            .O(N__25123),
            .I(iQ_RNIA1EM1_2_cascade_));
    InMux I__3822 (
            .O(N__25120),
            .I(N__25117));
    LocalMux I__3821 (
            .O(N__25117),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIA1VQZ0Z_19 ));
    InMux I__3820 (
            .O(N__25114),
            .I(N__25111));
    LocalMux I__3819 (
            .O(N__25111),
            .I(N__25108));
    Span4Mux_h I__3818 (
            .O(N__25108),
            .I(N__25105));
    Odrv4 I__3817 (
            .O(N__25105),
            .I(\u1.PIO_control.ping_d_10 ));
    InMux I__3816 (
            .O(N__25102),
            .I(N__25099));
    LocalMux I__3815 (
            .O(N__25099),
            .I(N__25096));
    Span4Mux_v I__3814 (
            .O(N__25096),
            .I(N__25093));
    Span4Mux_v I__3813 (
            .O(N__25093),
            .I(N__25090));
    Odrv4 I__3812 (
            .O(N__25090),
            .I(\u1.PIO_control.ping_d_11 ));
    CEMux I__3811 (
            .O(N__25087),
            .I(N__25082));
    CEMux I__3810 (
            .O(N__25086),
            .I(N__25079));
    CEMux I__3809 (
            .O(N__25085),
            .I(N__25076));
    LocalMux I__3808 (
            .O(N__25082),
            .I(N__25073));
    LocalMux I__3807 (
            .O(N__25079),
            .I(N__25070));
    LocalMux I__3806 (
            .O(N__25076),
            .I(N__25067));
    Span4Mux_h I__3805 (
            .O(N__25073),
            .I(N__25064));
    Span4Mux_h I__3804 (
            .O(N__25070),
            .I(N__25061));
    Odrv12 I__3803 (
            .O(N__25067),
            .I(\u1.PIO_control.ping_we_0_sqmuxa ));
    Odrv4 I__3802 (
            .O(N__25064),
            .I(\u1.PIO_control.ping_we_0_sqmuxa ));
    Odrv4 I__3801 (
            .O(N__25061),
            .I(\u1.PIO_control.ping_we_0_sqmuxa ));
    CascadeMux I__3800 (
            .O(N__25054),
            .I(N__25051));
    InMux I__3799 (
            .O(N__25051),
            .I(N__25048));
    LocalMux I__3798 (
            .O(N__25048),
            .I(N__25044));
    InMux I__3797 (
            .O(N__25047),
            .I(N__25041));
    Span4Mux_v I__3796 (
            .O(N__25044),
            .I(N__25038));
    LocalMux I__3795 (
            .O(N__25041),
            .I(N__25035));
    Odrv4 I__3794 (
            .O(N__25038),
            .I(DMA_dev0_Td_5));
    Odrv12 I__3793 (
            .O(N__25035),
            .I(DMA_dev0_Td_5));
    InMux I__3792 (
            .O(N__25030),
            .I(N__25027));
    LocalMux I__3791 (
            .O(N__25027),
            .I(N__25023));
    InMux I__3790 (
            .O(N__25026),
            .I(N__25020));
    Span4Mux_h I__3789 (
            .O(N__25023),
            .I(N__25015));
    LocalMux I__3788 (
            .O(N__25020),
            .I(N__25015));
    Odrv4 I__3787 (
            .O(N__25015),
            .I(\u1.N_1423 ));
    CascadeMux I__3786 (
            .O(N__25012),
            .I(N__25009));
    InMux I__3785 (
            .O(N__25009),
            .I(N__25006));
    LocalMux I__3784 (
            .O(N__25006),
            .I(N__25003));
    Span4Mux_h I__3783 (
            .O(N__25003),
            .I(N__25000));
    Odrv4 I__3782 (
            .O(N__25000),
            .I(\u1.PIO_control.un3_idone_0_a2_0 ));
    InMux I__3781 (
            .O(N__24997),
            .I(N__24994));
    LocalMux I__3780 (
            .O(N__24994),
            .I(N__24991));
    Span4Mux_v I__3779 (
            .O(N__24991),
            .I(N__24988));
    Span4Mux_h I__3778 (
            .O(N__24988),
            .I(N__24984));
    InMux I__3777 (
            .O(N__24987),
            .I(N__24981));
    Odrv4 I__3776 (
            .O(N__24984),
            .I(\u1.N_1429 ));
    LocalMux I__3775 (
            .O(N__24981),
            .I(\u1.N_1429 ));
    CascadeMux I__3774 (
            .O(N__24976),
            .I(\u1.PIO_control.SelDev_e_1_cascade_ ));
    CascadeMux I__3773 (
            .O(N__24973),
            .I(N__24968));
    CascadeMux I__3772 (
            .O(N__24972),
            .I(N__24965));
    InMux I__3771 (
            .O(N__24971),
            .I(N__24961));
    InMux I__3770 (
            .O(N__24968),
            .I(N__24954));
    InMux I__3769 (
            .O(N__24965),
            .I(N__24954));
    InMux I__3768 (
            .O(N__24964),
            .I(N__24954));
    LocalMux I__3767 (
            .O(N__24961),
            .I(N__24950));
    LocalMux I__3766 (
            .O(N__24954),
            .I(N__24947));
    InMux I__3765 (
            .O(N__24953),
            .I(N__24944));
    Span4Mux_h I__3764 (
            .O(N__24950),
            .I(N__24939));
    Span4Mux_h I__3763 (
            .O(N__24947),
            .I(N__24939));
    LocalMux I__3762 (
            .O(N__24944),
            .I(N__24936));
    Odrv4 I__3761 (
            .O(N__24939),
            .I(DMActrl_DMAen));
    Odrv4 I__3760 (
            .O(N__24936),
            .I(DMActrl_DMAen));
    CascadeMux I__3759 (
            .O(N__24931),
            .I(\u0.dat_o_0_0_2_15_cascade_ ));
    InMux I__3758 (
            .O(N__24928),
            .I(N__24925));
    LocalMux I__3757 (
            .O(N__24925),
            .I(N__24921));
    InMux I__3756 (
            .O(N__24924),
            .I(N__24918));
    Span4Mux_v I__3755 (
            .O(N__24921),
            .I(N__24913));
    LocalMux I__3754 (
            .O(N__24918),
            .I(N__24913));
    Span4Mux_h I__3753 (
            .O(N__24913),
            .I(N__24910));
    Span4Mux_h I__3752 (
            .O(N__24910),
            .I(N__24907));
    Odrv4 I__3751 (
            .O(N__24907),
            .I(DMA_dev0_Td_7));
    CascadeMux I__3750 (
            .O(N__24904),
            .I(\u1.PIO_control.pong_a_RNI914A1_0_cascade_ ));
    InMux I__3749 (
            .O(N__24901),
            .I(N__24898));
    LocalMux I__3748 (
            .O(N__24898),
            .I(\u1.PIO_control.ping_a_RNIQNVQ_0 ));
    CEMux I__3747 (
            .O(N__24895),
            .I(N__24891));
    CEMux I__3746 (
            .O(N__24894),
            .I(N__24888));
    LocalMux I__3745 (
            .O(N__24891),
            .I(N__24885));
    LocalMux I__3744 (
            .O(N__24888),
            .I(N__24879));
    Span4Mux_h I__3743 (
            .O(N__24885),
            .I(N__24876));
    CEMux I__3742 (
            .O(N__24884),
            .I(N__24873));
    CEMux I__3741 (
            .O(N__24883),
            .I(N__24870));
    CEMux I__3740 (
            .O(N__24882),
            .I(N__24867));
    Span4Mux_h I__3739 (
            .O(N__24879),
            .I(N__24864));
    Span4Mux_h I__3738 (
            .O(N__24876),
            .I(N__24859));
    LocalMux I__3737 (
            .O(N__24873),
            .I(N__24859));
    LocalMux I__3736 (
            .O(N__24870),
            .I(N__24856));
    LocalMux I__3735 (
            .O(N__24867),
            .I(N__24853));
    Span4Mux_v I__3734 (
            .O(N__24864),
            .I(N__24848));
    Span4Mux_h I__3733 (
            .O(N__24859),
            .I(N__24848));
    Span4Mux_v I__3732 (
            .O(N__24856),
            .I(N__24845));
    Span4Mux_h I__3731 (
            .O(N__24853),
            .I(N__24842));
    Odrv4 I__3730 (
            .O(N__24848),
            .I(\u1.PIO_control.pong_we_1_sqmuxa ));
    Odrv4 I__3729 (
            .O(N__24845),
            .I(\u1.PIO_control.pong_we_1_sqmuxa ));
    Odrv4 I__3728 (
            .O(N__24842),
            .I(\u1.PIO_control.pong_we_1_sqmuxa ));
    InMux I__3727 (
            .O(N__24835),
            .I(N__24832));
    LocalMux I__3726 (
            .O(N__24832),
            .I(N__24829));
    Span4Mux_h I__3725 (
            .O(N__24829),
            .I(N__24819));
    InMux I__3724 (
            .O(N__24828),
            .I(N__24806));
    InMux I__3723 (
            .O(N__24827),
            .I(N__24806));
    InMux I__3722 (
            .O(N__24826),
            .I(N__24806));
    InMux I__3721 (
            .O(N__24825),
            .I(N__24806));
    InMux I__3720 (
            .O(N__24824),
            .I(N__24806));
    InMux I__3719 (
            .O(N__24823),
            .I(N__24806));
    InMux I__3718 (
            .O(N__24822),
            .I(N__24803));
    Odrv4 I__3717 (
            .O(N__24819),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.N_1073 ));
    LocalMux I__3716 (
            .O(N__24806),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.N_1073 ));
    LocalMux I__3715 (
            .O(N__24803),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.N_1073 ));
    InMux I__3714 (
            .O(N__24796),
            .I(N__24793));
    LocalMux I__3713 (
            .O(N__24793),
            .I(N__24790));
    Span4Mux_h I__3712 (
            .O(N__24790),
            .I(N__24787));
    Odrv4 I__3711 (
            .O(N__24787),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_s_7 ));
    CascadeMux I__3710 (
            .O(N__24784),
            .I(N__24780));
    InMux I__3709 (
            .O(N__24783),
            .I(N__24777));
    InMux I__3708 (
            .O(N__24780),
            .I(N__24774));
    LocalMux I__3707 (
            .O(N__24777),
            .I(N__24771));
    LocalMux I__3706 (
            .O(N__24774),
            .I(N__24768));
    Span4Mux_v I__3705 (
            .O(N__24771),
            .I(N__24763));
    Span4Mux_h I__3704 (
            .O(N__24768),
            .I(N__24763));
    Odrv4 I__3703 (
            .O(N__24763),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.QiZ0Z_7 ));
    CEMux I__3702 (
            .O(N__24760),
            .I(N__24756));
    CEMux I__3701 (
            .O(N__24759),
            .I(N__24753));
    LocalMux I__3700 (
            .O(N__24756),
            .I(N__24749));
    LocalMux I__3699 (
            .O(N__24753),
            .I(N__24746));
    CEMux I__3698 (
            .O(N__24752),
            .I(N__24743));
    Span4Mux_h I__3697 (
            .O(N__24749),
            .I(N__24740));
    Span4Mux_v I__3696 (
            .O(N__24746),
            .I(N__24735));
    LocalMux I__3695 (
            .O(N__24743),
            .I(N__24735));
    Span4Mux_h I__3694 (
            .O(N__24740),
            .I(N__24732));
    Span4Mux_v I__3693 (
            .O(N__24735),
            .I(N__24729));
    Odrv4 I__3692 (
            .O(N__24732),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.N_1071 ));
    Odrv4 I__3691 (
            .O(N__24729),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.N_1071 ));
    InMux I__3690 (
            .O(N__24724),
            .I(N__24720));
    CascadeMux I__3689 (
            .O(N__24723),
            .I(N__24717));
    LocalMux I__3688 (
            .O(N__24720),
            .I(N__24712));
    InMux I__3687 (
            .O(N__24717),
            .I(N__24709));
    InMux I__3686 (
            .O(N__24716),
            .I(N__24706));
    InMux I__3685 (
            .O(N__24715),
            .I(N__24703));
    Span12Mux_s4_h I__3684 (
            .O(N__24712),
            .I(N__24698));
    LocalMux I__3683 (
            .O(N__24709),
            .I(N__24698));
    LocalMux I__3682 (
            .O(N__24706),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.rciZ0 ));
    LocalMux I__3681 (
            .O(N__24703),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.rciZ0 ));
    Odrv12 I__3680 (
            .O(N__24698),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.rciZ0 ));
    CascadeMux I__3679 (
            .O(N__24691),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNI9LFIZ0Z_1_cascade_ ));
    InMux I__3678 (
            .O(N__24688),
            .I(N__24685));
    LocalMux I__3677 (
            .O(N__24685),
            .I(N__24682));
    Span4Mux_h I__3676 (
            .O(N__24682),
            .I(N__24679));
    Odrv4 I__3675 (
            .O(N__24679),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.Qi_RNI7F9K_0 ));
    InMux I__3674 (
            .O(N__24676),
            .I(N__24673));
    LocalMux I__3673 (
            .O(N__24673),
            .I(N__24670));
    Span4Mux_v I__3672 (
            .O(N__24670),
            .I(N__24666));
    InMux I__3671 (
            .O(N__24669),
            .I(N__24663));
    Span4Mux_h I__3670 (
            .O(N__24666),
            .I(N__24660));
    LocalMux I__3669 (
            .O(N__24663),
            .I(N__24657));
    Odrv4 I__3668 (
            .O(N__24660),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.val_c8_0_4_0 ));
    Odrv12 I__3667 (
            .O(N__24657),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.val_c8_0_4_0 ));
    InMux I__3666 (
            .O(N__24652),
            .I(N__24649));
    LocalMux I__3665 (
            .O(N__24649),
            .I(\u1.PIO_control.PIO_access_control.it1_1_iv_0_0_4 ));
    InMux I__3664 (
            .O(N__24646),
            .I(N__24643));
    LocalMux I__3663 (
            .O(N__24643),
            .I(N__24640));
    Odrv12 I__3662 (
            .O(N__24640),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_18 ));
    InMux I__3661 (
            .O(N__24637),
            .I(N__24634));
    LocalMux I__3660 (
            .O(N__24634),
            .I(N__24631));
    Span4Mux_v I__3659 (
            .O(N__24631),
            .I(N__24628));
    Span4Mux_h I__3658 (
            .O(N__24628),
            .I(N__24625));
    Span4Mux_h I__3657 (
            .O(N__24625),
            .I(N__24622));
    Span4Mux_v I__3656 (
            .O(N__24622),
            .I(N__24619));
    Odrv4 I__3655 (
            .O(N__24619),
            .I(\u1.DMA_control.Tm_1 ));
    InMux I__3654 (
            .O(N__24616),
            .I(N__24613));
    LocalMux I__3653 (
            .O(N__24613),
            .I(N__24610));
    Odrv12 I__3652 (
            .O(N__24610),
            .I(\u1.PIO_control.PIO_access_control.T1Z0Z_0 ));
    InMux I__3651 (
            .O(N__24607),
            .I(N__24604));
    LocalMux I__3650 (
            .O(N__24604),
            .I(N__24600));
    CascadeMux I__3649 (
            .O(N__24603),
            .I(N__24596));
    Span4Mux_v I__3648 (
            .O(N__24600),
            .I(N__24593));
    InMux I__3647 (
            .O(N__24599),
            .I(N__24590));
    InMux I__3646 (
            .O(N__24596),
            .I(N__24584));
    Span4Mux_h I__3645 (
            .O(N__24593),
            .I(N__24579));
    LocalMux I__3644 (
            .O(N__24590),
            .I(N__24579));
    InMux I__3643 (
            .O(N__24589),
            .I(N__24572));
    InMux I__3642 (
            .O(N__24588),
            .I(N__24572));
    InMux I__3641 (
            .O(N__24587),
            .I(N__24572));
    LocalMux I__3640 (
            .O(N__24584),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.hT2doneZ0 ));
    Odrv4 I__3639 (
            .O(N__24579),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.hT2doneZ0 ));
    LocalMux I__3638 (
            .O(N__24572),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.hT2doneZ0 ));
    InMux I__3637 (
            .O(N__24565),
            .I(N__24562));
    LocalMux I__3636 (
            .O(N__24562),
            .I(N__24557));
    CascadeMux I__3635 (
            .O(N__24561),
            .I(N__24554));
    InMux I__3634 (
            .O(N__24560),
            .I(N__24551));
    Span4Mux_h I__3633 (
            .O(N__24557),
            .I(N__24548));
    InMux I__3632 (
            .O(N__24554),
            .I(N__24543));
    LocalMux I__3631 (
            .O(N__24551),
            .I(N__24540));
    Span4Mux_h I__3630 (
            .O(N__24548),
            .I(N__24537));
    InMux I__3629 (
            .O(N__24547),
            .I(N__24534));
    InMux I__3628 (
            .O(N__24546),
            .I(N__24531));
    LocalMux I__3627 (
            .O(N__24543),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.val_c8 ));
    Odrv12 I__3626 (
            .O(N__24540),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.val_c8 ));
    Odrv4 I__3625 (
            .O(N__24537),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.val_c8 ));
    LocalMux I__3624 (
            .O(N__24534),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.val_c8 ));
    LocalMux I__3623 (
            .O(N__24531),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.val_c8 ));
    InMux I__3622 (
            .O(N__24520),
            .I(N__24517));
    LocalMux I__3621 (
            .O(N__24517),
            .I(N__24512));
    InMux I__3620 (
            .O(N__24516),
            .I(N__24506));
    InMux I__3619 (
            .O(N__24515),
            .I(N__24506));
    Span4Mux_h I__3618 (
            .O(N__24512),
            .I(N__24499));
    InMux I__3617 (
            .O(N__24511),
            .I(N__24496));
    LocalMux I__3616 (
            .O(N__24506),
            .I(N__24493));
    InMux I__3615 (
            .O(N__24505),
            .I(N__24484));
    InMux I__3614 (
            .O(N__24504),
            .I(N__24484));
    InMux I__3613 (
            .O(N__24503),
            .I(N__24484));
    InMux I__3612 (
            .O(N__24502),
            .I(N__24484));
    Odrv4 I__3611 (
            .O(N__24499),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.iordy_done_0 ));
    LocalMux I__3610 (
            .O(N__24496),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.iordy_done_0 ));
    Odrv12 I__3609 (
            .O(N__24493),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.iordy_done_0 ));
    LocalMux I__3608 (
            .O(N__24484),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.iordy_done_0 ));
    InMux I__3607 (
            .O(N__24475),
            .I(N__24472));
    LocalMux I__3606 (
            .O(N__24472),
            .I(N__24469));
    Odrv12 I__3605 (
            .O(N__24469),
            .I(\u1.PIO_control.PIO_access_control.T1Z0Z_2 ));
    InMux I__3604 (
            .O(N__24466),
            .I(N__24463));
    LocalMux I__3603 (
            .O(N__24463),
            .I(N__24460));
    Span4Mux_h I__3602 (
            .O(N__24460),
            .I(N__24457));
    Odrv4 I__3601 (
            .O(N__24457),
            .I(\u1.PIO_control.PIO_access_control.T1Z0Z_4 ));
    InMux I__3600 (
            .O(N__24454),
            .I(N__24451));
    LocalMux I__3599 (
            .O(N__24451),
            .I(N__24448));
    Span4Mux_h I__3598 (
            .O(N__24448),
            .I(N__24442));
    InMux I__3597 (
            .O(N__24447),
            .I(N__24439));
    InMux I__3596 (
            .O(N__24446),
            .I(N__24436));
    CascadeMux I__3595 (
            .O(N__24445),
            .I(N__24433));
    Span4Mux_v I__3594 (
            .O(N__24442),
            .I(N__24430));
    LocalMux I__3593 (
            .O(N__24439),
            .I(N__24427));
    LocalMux I__3592 (
            .O(N__24436),
            .I(N__24424));
    InMux I__3591 (
            .O(N__24433),
            .I(N__24421));
    Span4Mux_h I__3590 (
            .O(N__24430),
            .I(N__24418));
    Span4Mux_v I__3589 (
            .O(N__24427),
            .I(N__24413));
    Span4Mux_h I__3588 (
            .O(N__24424),
            .I(N__24413));
    LocalMux I__3587 (
            .O(N__24421),
            .I(\u1.c_stateZ0Z_0 ));
    Odrv4 I__3586 (
            .O(N__24418),
            .I(\u1.c_stateZ0Z_0 ));
    Odrv4 I__3585 (
            .O(N__24413),
            .I(\u1.c_stateZ0Z_0 ));
    InMux I__3584 (
            .O(N__24406),
            .I(N__24400));
    InMux I__3583 (
            .O(N__24405),
            .I(N__24397));
    InMux I__3582 (
            .O(N__24404),
            .I(N__24394));
    InMux I__3581 (
            .O(N__24403),
            .I(N__24391));
    LocalMux I__3580 (
            .O(N__24400),
            .I(N__24388));
    LocalMux I__3579 (
            .O(N__24397),
            .I(N__24385));
    LocalMux I__3578 (
            .O(N__24394),
            .I(N__24382));
    LocalMux I__3577 (
            .O(N__24391),
            .I(N__24379));
    Span4Mux_s3_h I__3576 (
            .O(N__24388),
            .I(N__24376));
    Span4Mux_v I__3575 (
            .O(N__24385),
            .I(N__24371));
    Span4Mux_h I__3574 (
            .O(N__24382),
            .I(N__24371));
    Odrv12 I__3573 (
            .O(N__24379),
            .I(\u1.c_stateZ0Z_1 ));
    Odrv4 I__3572 (
            .O(N__24376),
            .I(\u1.c_stateZ0Z_1 ));
    Odrv4 I__3571 (
            .O(N__24371),
            .I(\u1.c_stateZ0Z_1 ));
    CascadeMux I__3570 (
            .O(N__24364),
            .I(N__24361));
    InMux I__3569 (
            .O(N__24361),
            .I(N__24358));
    LocalMux I__3568 (
            .O(N__24358),
            .I(N__24355));
    Odrv12 I__3567 (
            .O(N__24355),
            .I(\u1.c_state_ns_i_i_i_a2_1_1 ));
    InMux I__3566 (
            .O(N__24352),
            .I(N__24349));
    LocalMux I__3565 (
            .O(N__24349),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_3 ));
    InMux I__3564 (
            .O(N__24346),
            .I(N__24343));
    LocalMux I__3563 (
            .O(N__24343),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_19 ));
    InMux I__3562 (
            .O(N__24340),
            .I(N__24337));
    LocalMux I__3561 (
            .O(N__24337),
            .I(N__24334));
    Odrv12 I__3560 (
            .O(N__24334),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNIA9TNZ0Z_6 ));
    CascadeMux I__3559 (
            .O(N__24331),
            .I(mem_mem_ram6__RNIQPOD1_6_cascade_));
    InMux I__3558 (
            .O(N__24328),
            .I(N__24325));
    LocalMux I__3557 (
            .O(N__24325),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_6 ));
    CascadeMux I__3556 (
            .O(N__24322),
            .I(N__24317));
    InMux I__3555 (
            .O(N__24321),
            .I(N__24310));
    InMux I__3554 (
            .O(N__24320),
            .I(N__24310));
    InMux I__3553 (
            .O(N__24317),
            .I(N__24310));
    LocalMux I__3552 (
            .O(N__24310),
            .I(N__24297));
    InMux I__3551 (
            .O(N__24309),
            .I(N__24284));
    InMux I__3550 (
            .O(N__24308),
            .I(N__24284));
    InMux I__3549 (
            .O(N__24307),
            .I(N__24284));
    InMux I__3548 (
            .O(N__24306),
            .I(N__24284));
    InMux I__3547 (
            .O(N__24305),
            .I(N__24284));
    InMux I__3546 (
            .O(N__24304),
            .I(N__24284));
    InMux I__3545 (
            .O(N__24303),
            .I(N__24275));
    InMux I__3544 (
            .O(N__24302),
            .I(N__24275));
    InMux I__3543 (
            .O(N__24301),
            .I(N__24275));
    InMux I__3542 (
            .O(N__24300),
            .I(N__24275));
    Span4Mux_v I__3541 (
            .O(N__24297),
            .I(N__24272));
    LocalMux I__3540 (
            .O(N__24284),
            .I(N__24269));
    LocalMux I__3539 (
            .O(N__24275),
            .I(\u1.DMA_control.wr_ptr_0 ));
    Odrv4 I__3538 (
            .O(N__24272),
            .I(\u1.DMA_control.wr_ptr_0 ));
    Odrv4 I__3537 (
            .O(N__24269),
            .I(\u1.DMA_control.wr_ptr_0 ));
    CascadeMux I__3536 (
            .O(N__24262),
            .I(N__24253));
    CascadeMux I__3535 (
            .O(N__24261),
            .I(N__24248));
    CascadeMux I__3534 (
            .O(N__24260),
            .I(N__24244));
    CascadeMux I__3533 (
            .O(N__24259),
            .I(N__24240));
    CascadeMux I__3532 (
            .O(N__24258),
            .I(N__24236));
    CascadeMux I__3531 (
            .O(N__24257),
            .I(N__24233));
    InMux I__3530 (
            .O(N__24256),
            .I(N__24222));
    InMux I__3529 (
            .O(N__24253),
            .I(N__24222));
    InMux I__3528 (
            .O(N__24252),
            .I(N__24222));
    InMux I__3527 (
            .O(N__24251),
            .I(N__24222));
    InMux I__3526 (
            .O(N__24248),
            .I(N__24222));
    InMux I__3525 (
            .O(N__24247),
            .I(N__24209));
    InMux I__3524 (
            .O(N__24244),
            .I(N__24209));
    InMux I__3523 (
            .O(N__24243),
            .I(N__24209));
    InMux I__3522 (
            .O(N__24240),
            .I(N__24209));
    InMux I__3521 (
            .O(N__24239),
            .I(N__24209));
    InMux I__3520 (
            .O(N__24236),
            .I(N__24209));
    InMux I__3519 (
            .O(N__24233),
            .I(N__24206));
    LocalMux I__3518 (
            .O(N__24222),
            .I(N__24203));
    LocalMux I__3517 (
            .O(N__24209),
            .I(N__24200));
    LocalMux I__3516 (
            .O(N__24206),
            .I(N__24197));
    Span4Mux_v I__3515 (
            .O(N__24203),
            .I(N__24192));
    Span4Mux_v I__3514 (
            .O(N__24200),
            .I(N__24192));
    Span4Mux_h I__3513 (
            .O(N__24197),
            .I(N__24187));
    Span4Mux_h I__3512 (
            .O(N__24192),
            .I(N__24187));
    Odrv4 I__3511 (
            .O(N__24187),
            .I(\u1.DMA_control.RxWrZ0 ));
    CascadeMux I__3510 (
            .O(N__24184),
            .I(N__24178));
    CascadeMux I__3509 (
            .O(N__24183),
            .I(N__24175));
    CascadeMux I__3508 (
            .O(N__24182),
            .I(N__24170));
    InMux I__3507 (
            .O(N__24181),
            .I(N__24165));
    InMux I__3506 (
            .O(N__24178),
            .I(N__24152));
    InMux I__3505 (
            .O(N__24175),
            .I(N__24152));
    InMux I__3504 (
            .O(N__24174),
            .I(N__24152));
    InMux I__3503 (
            .O(N__24173),
            .I(N__24152));
    InMux I__3502 (
            .O(N__24170),
            .I(N__24152));
    InMux I__3501 (
            .O(N__24169),
            .I(N__24152));
    CascadeMux I__3500 (
            .O(N__24168),
            .I(N__24149));
    LocalMux I__3499 (
            .O(N__24165),
            .I(N__24141));
    LocalMux I__3498 (
            .O(N__24152),
            .I(N__24141));
    InMux I__3497 (
            .O(N__24149),
            .I(N__24132));
    InMux I__3496 (
            .O(N__24148),
            .I(N__24132));
    InMux I__3495 (
            .O(N__24147),
            .I(N__24132));
    InMux I__3494 (
            .O(N__24146),
            .I(N__24132));
    Odrv12 I__3493 (
            .O(N__24141),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.wr_ptr_1 ));
    LocalMux I__3492 (
            .O(N__24132),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.wr_ptr_1 ));
    InMux I__3491 (
            .O(N__24127),
            .I(N__24109));
    InMux I__3490 (
            .O(N__24126),
            .I(N__24109));
    InMux I__3489 (
            .O(N__24125),
            .I(N__24109));
    InMux I__3488 (
            .O(N__24124),
            .I(N__24109));
    InMux I__3487 (
            .O(N__24123),
            .I(N__24109));
    InMux I__3486 (
            .O(N__24122),
            .I(N__24109));
    LocalMux I__3485 (
            .O(N__24109),
            .I(N__24103));
    InMux I__3484 (
            .O(N__24108),
            .I(N__24100));
    InMux I__3483 (
            .O(N__24107),
            .I(N__24095));
    InMux I__3482 (
            .O(N__24106),
            .I(N__24095));
    Odrv4 I__3481 (
            .O(N__24103),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.wr_ptr_2 ));
    LocalMux I__3480 (
            .O(N__24100),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.wr_ptr_2 ));
    LocalMux I__3479 (
            .O(N__24095),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.wr_ptr_2 ));
    InMux I__3478 (
            .O(N__24088),
            .I(N__24085));
    LocalMux I__3477 (
            .O(N__24085),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_21 ));
    InMux I__3476 (
            .O(N__24082),
            .I(N__24079));
    LocalMux I__3475 (
            .O(N__24079),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_5 ));
    CascadeMux I__3474 (
            .O(N__24076),
            .I(\u1.DMA_control.gen_DMAbuf_Txbuf.N_1602_cascade_ ));
    IoInMux I__3473 (
            .O(N__24073),
            .I(N__24070));
    LocalMux I__3472 (
            .O(N__24070),
            .I(N__24067));
    Span4Mux_s3_h I__3471 (
            .O(N__24067),
            .I(N__24064));
    Span4Mux_v I__3470 (
            .O(N__24064),
            .I(N__24061));
    Span4Mux_v I__3469 (
            .O(N__24061),
            .I(N__24058));
    Odrv4 I__3468 (
            .O(N__24058),
            .I(\u1.DMA_control.gen_DMAbuf_Txbuf.N_319 ));
    InMux I__3467 (
            .O(N__24055),
            .I(N__24052));
    LocalMux I__3466 (
            .O(N__24052),
            .I(N__24049));
    Span4Mux_h I__3465 (
            .O(N__24049),
            .I(N__24046));
    Odrv4 I__3464 (
            .O(N__24046),
            .I(\u1.DMA_control.writeDlw_13 ));
    InMux I__3463 (
            .O(N__24043),
            .I(N__24040));
    LocalMux I__3462 (
            .O(N__24040),
            .I(N__24036));
    InMux I__3461 (
            .O(N__24039),
            .I(N__24033));
    Span4Mux_h I__3460 (
            .O(N__24036),
            .I(N__24030));
    LocalMux I__3459 (
            .O(N__24033),
            .I(\u1.DMA_control.TxbufQ_29 ));
    Odrv4 I__3458 (
            .O(N__24030),
            .I(\u1.DMA_control.TxbufQ_29 ));
    InMux I__3457 (
            .O(N__24025),
            .I(N__24022));
    LocalMux I__3456 (
            .O(N__24022),
            .I(\u1.DMA_control.writeDfw_6_i_m2_i_0_13 ));
    InMux I__3455 (
            .O(N__24019),
            .I(N__24016));
    LocalMux I__3454 (
            .O(N__24016),
            .I(N__24013));
    Span4Mux_v I__3453 (
            .O(N__24013),
            .I(N__24010));
    Odrv4 I__3452 (
            .O(N__24010),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_6 ));
    InMux I__3451 (
            .O(N__24007),
            .I(N__24003));
    InMux I__3450 (
            .O(N__24006),
            .I(N__24000));
    LocalMux I__3449 (
            .O(N__24003),
            .I(N__23997));
    LocalMux I__3448 (
            .O(N__24000),
            .I(N__23994));
    Span4Mux_h I__3447 (
            .O(N__23997),
            .I(N__23991));
    Odrv4 I__3446 (
            .O(N__23994),
            .I(\u1.DMA_control.TxbufQ_26 ));
    Odrv4 I__3445 (
            .O(N__23991),
            .I(\u1.DMA_control.TxbufQ_26 ));
    InMux I__3444 (
            .O(N__23986),
            .I(N__23983));
    LocalMux I__3443 (
            .O(N__23983),
            .I(N__23980));
    Odrv4 I__3442 (
            .O(N__23980),
            .I(\u1.DMA_control.writeDlw_10 ));
    InMux I__3441 (
            .O(N__23977),
            .I(N__23974));
    LocalMux I__3440 (
            .O(N__23974),
            .I(\u1.DMA_control.writeDfw_6_i_0_10 ));
    InMux I__3439 (
            .O(N__23971),
            .I(N__23968));
    LocalMux I__3438 (
            .O(N__23968),
            .I(N__23965));
    Span4Mux_h I__3437 (
            .O(N__23965),
            .I(N__23962));
    Span4Mux_v I__3436 (
            .O(N__23962),
            .I(N__23959));
    Odrv4 I__3435 (
            .O(N__23959),
            .I(\u1.DMA_control.Td_5 ));
    InMux I__3434 (
            .O(N__23956),
            .I(N__23952));
    InMux I__3433 (
            .O(N__23955),
            .I(N__23949));
    LocalMux I__3432 (
            .O(N__23952),
            .I(N__23944));
    LocalMux I__3431 (
            .O(N__23949),
            .I(N__23944));
    Span4Mux_h I__3430 (
            .O(N__23944),
            .I(N__23941));
    Odrv4 I__3429 (
            .O(N__23941),
            .I(\u1.DMA_control.TxbufQ_25 ));
    CascadeMux I__3428 (
            .O(N__23938),
            .I(N__23935));
    InMux I__3427 (
            .O(N__23935),
            .I(N__23932));
    LocalMux I__3426 (
            .O(N__23932),
            .I(N__23929));
    Odrv4 I__3425 (
            .O(N__23929),
            .I(\u1.DMA_control.writeDlw_9 ));
    InMux I__3424 (
            .O(N__23926),
            .I(N__23923));
    LocalMux I__3423 (
            .O(N__23923),
            .I(N__23919));
    InMux I__3422 (
            .O(N__23922),
            .I(N__23916));
    Span4Mux_h I__3421 (
            .O(N__23919),
            .I(N__23913));
    LocalMux I__3420 (
            .O(N__23916),
            .I(N__23910));
    Span4Mux_h I__3419 (
            .O(N__23913),
            .I(N__23907));
    Span4Mux_v I__3418 (
            .O(N__23910),
            .I(N__23904));
    Odrv4 I__3417 (
            .O(N__23907),
            .I(\u1.DMA_control.TxbufQ_1 ));
    Odrv4 I__3416 (
            .O(N__23904),
            .I(\u1.DMA_control.TxbufQ_1 ));
    CascadeMux I__3415 (
            .O(N__23899),
            .I(\u1.DMA_control.writeDfw_6_i_0_9_cascade_ ));
    InMux I__3414 (
            .O(N__23896),
            .I(N__23893));
    LocalMux I__3413 (
            .O(N__23893),
            .I(N__23890));
    Span4Mux_s3_h I__3412 (
            .O(N__23890),
            .I(N__23887));
    Span4Mux_h I__3411 (
            .O(N__23887),
            .I(N__23884));
    Odrv4 I__3410 (
            .O(N__23884),
            .I(\u1.DMAd_9 ));
    CascadeMux I__3409 (
            .O(N__23881),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.N_1385_i_cascade_ ));
    InMux I__3408 (
            .O(N__23878),
            .I(N__23841));
    InMux I__3407 (
            .O(N__23877),
            .I(N__23841));
    InMux I__3406 (
            .O(N__23876),
            .I(N__23841));
    InMux I__3405 (
            .O(N__23875),
            .I(N__23841));
    InMux I__3404 (
            .O(N__23874),
            .I(N__23841));
    InMux I__3403 (
            .O(N__23873),
            .I(N__23841));
    InMux I__3402 (
            .O(N__23872),
            .I(N__23841));
    InMux I__3401 (
            .O(N__23871),
            .I(N__23841));
    InMux I__3400 (
            .O(N__23870),
            .I(N__23813));
    InMux I__3399 (
            .O(N__23869),
            .I(N__23813));
    InMux I__3398 (
            .O(N__23868),
            .I(N__23813));
    InMux I__3397 (
            .O(N__23867),
            .I(N__23813));
    InMux I__3396 (
            .O(N__23866),
            .I(N__23813));
    InMux I__3395 (
            .O(N__23865),
            .I(N__23796));
    InMux I__3394 (
            .O(N__23864),
            .I(N__23796));
    InMux I__3393 (
            .O(N__23863),
            .I(N__23796));
    InMux I__3392 (
            .O(N__23862),
            .I(N__23796));
    InMux I__3391 (
            .O(N__23861),
            .I(N__23796));
    InMux I__3390 (
            .O(N__23860),
            .I(N__23796));
    InMux I__3389 (
            .O(N__23859),
            .I(N__23796));
    InMux I__3388 (
            .O(N__23858),
            .I(N__23796));
    LocalMux I__3387 (
            .O(N__23841),
            .I(N__23793));
    InMux I__3386 (
            .O(N__23840),
            .I(N__23776));
    InMux I__3385 (
            .O(N__23839),
            .I(N__23776));
    InMux I__3384 (
            .O(N__23838),
            .I(N__23776));
    InMux I__3383 (
            .O(N__23837),
            .I(N__23776));
    InMux I__3382 (
            .O(N__23836),
            .I(N__23776));
    InMux I__3381 (
            .O(N__23835),
            .I(N__23776));
    InMux I__3380 (
            .O(N__23834),
            .I(N__23776));
    InMux I__3379 (
            .O(N__23833),
            .I(N__23776));
    InMux I__3378 (
            .O(N__23832),
            .I(N__23759));
    InMux I__3377 (
            .O(N__23831),
            .I(N__23759));
    InMux I__3376 (
            .O(N__23830),
            .I(N__23759));
    InMux I__3375 (
            .O(N__23829),
            .I(N__23759));
    InMux I__3374 (
            .O(N__23828),
            .I(N__23759));
    InMux I__3373 (
            .O(N__23827),
            .I(N__23759));
    InMux I__3372 (
            .O(N__23826),
            .I(N__23759));
    InMux I__3371 (
            .O(N__23825),
            .I(N__23759));
    InMux I__3370 (
            .O(N__23824),
            .I(N__23756));
    LocalMux I__3369 (
            .O(N__23813),
            .I(N__23749));
    LocalMux I__3368 (
            .O(N__23796),
            .I(N__23746));
    Span4Mux_v I__3367 (
            .O(N__23793),
            .I(N__23739));
    LocalMux I__3366 (
            .O(N__23776),
            .I(N__23739));
    LocalMux I__3365 (
            .O(N__23759),
            .I(N__23739));
    LocalMux I__3364 (
            .O(N__23756),
            .I(N__23736));
    InMux I__3363 (
            .O(N__23755),
            .I(N__23727));
    InMux I__3362 (
            .O(N__23754),
            .I(N__23727));
    InMux I__3361 (
            .O(N__23753),
            .I(N__23727));
    InMux I__3360 (
            .O(N__23752),
            .I(N__23727));
    Odrv12 I__3359 (
            .O(N__23749),
            .I(\u1.DMA_control.N_1326 ));
    Odrv12 I__3358 (
            .O(N__23746),
            .I(\u1.DMA_control.N_1326 ));
    Odrv4 I__3357 (
            .O(N__23739),
            .I(\u1.DMA_control.N_1326 ));
    Odrv4 I__3356 (
            .O(N__23736),
            .I(\u1.DMA_control.N_1326 ));
    LocalMux I__3355 (
            .O(N__23727),
            .I(\u1.DMA_control.N_1326 ));
    InMux I__3354 (
            .O(N__23716),
            .I(N__23706));
    InMux I__3353 (
            .O(N__23715),
            .I(N__23706));
    InMux I__3352 (
            .O(N__23714),
            .I(N__23706));
    CascadeMux I__3351 (
            .O(N__23713),
            .I(N__23703));
    LocalMux I__3350 (
            .O(N__23706),
            .I(N__23700));
    InMux I__3349 (
            .O(N__23703),
            .I(N__23697));
    Span4Mux_v I__3348 (
            .O(N__23700),
            .I(N__23694));
    LocalMux I__3347 (
            .O(N__23697),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.iQ_fast_2 ));
    Odrv4 I__3346 (
            .O(N__23694),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.iQ_fast_2 ));
    InMux I__3345 (
            .O(N__23689),
            .I(N__23686));
    LocalMux I__3344 (
            .O(N__23686),
            .I(N__23683));
    Odrv12 I__3343 (
            .O(N__23683),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_18 ));
    InMux I__3342 (
            .O(N__23680),
            .I(N__23677));
    LocalMux I__3341 (
            .O(N__23677),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_19 ));
    InMux I__3340 (
            .O(N__23674),
            .I(N__23671));
    LocalMux I__3339 (
            .O(N__23671),
            .I(N__23668));
    Span4Mux_v I__3338 (
            .O(N__23668),
            .I(N__23665));
    Odrv4 I__3337 (
            .O(N__23665),
            .I(\u1.DMA_control.gen_DMAbuf_Txbuf.N_1602 ));
    InMux I__3336 (
            .O(N__23662),
            .I(N__23643));
    InMux I__3335 (
            .O(N__23661),
            .I(N__23643));
    InMux I__3334 (
            .O(N__23660),
            .I(N__23643));
    InMux I__3333 (
            .O(N__23659),
            .I(N__23638));
    InMux I__3332 (
            .O(N__23658),
            .I(N__23638));
    InMux I__3331 (
            .O(N__23657),
            .I(N__23635));
    InMux I__3330 (
            .O(N__23656),
            .I(N__23632));
    InMux I__3329 (
            .O(N__23655),
            .I(N__23629));
    InMux I__3328 (
            .O(N__23654),
            .I(N__23626));
    InMux I__3327 (
            .O(N__23653),
            .I(N__23619));
    InMux I__3326 (
            .O(N__23652),
            .I(N__23619));
    InMux I__3325 (
            .O(N__23651),
            .I(N__23619));
    InMux I__3324 (
            .O(N__23650),
            .I(N__23616));
    LocalMux I__3323 (
            .O(N__23643),
            .I(N__23611));
    LocalMux I__3322 (
            .O(N__23638),
            .I(N__23611));
    LocalMux I__3321 (
            .O(N__23635),
            .I(N__23608));
    LocalMux I__3320 (
            .O(N__23632),
            .I(N__23603));
    LocalMux I__3319 (
            .O(N__23629),
            .I(N__23603));
    LocalMux I__3318 (
            .O(N__23626),
            .I(N__23598));
    LocalMux I__3317 (
            .O(N__23619),
            .I(N__23598));
    LocalMux I__3316 (
            .O(N__23616),
            .I(N__23595));
    Span4Mux_v I__3315 (
            .O(N__23611),
            .I(N__23592));
    Span4Mux_v I__3314 (
            .O(N__23608),
            .I(N__23585));
    Span4Mux_v I__3313 (
            .O(N__23603),
            .I(N__23585));
    Span4Mux_h I__3312 (
            .O(N__23598),
            .I(N__23585));
    Odrv12 I__3311 (
            .O(N__23595),
            .I(DMActrl_dir));
    Odrv4 I__3310 (
            .O(N__23592),
            .I(DMActrl_dir));
    Odrv4 I__3309 (
            .O(N__23585),
            .I(DMActrl_dir));
    CascadeMux I__3308 (
            .O(N__23578),
            .I(N__23575));
    InMux I__3307 (
            .O(N__23575),
            .I(N__23569));
    InMux I__3306 (
            .O(N__23574),
            .I(N__23569));
    LocalMux I__3305 (
            .O(N__23569),
            .I(DMA_dev1_Tm_0));
    IoInMux I__3304 (
            .O(N__23566),
            .I(N__23563));
    LocalMux I__3303 (
            .O(N__23563),
            .I(N__23560));
    IoSpan4Mux I__3302 (
            .O(N__23560),
            .I(N__23557));
    Span4Mux_s2_v I__3301 (
            .O(N__23557),
            .I(N__23554));
    Span4Mux_v I__3300 (
            .O(N__23554),
            .I(N__23551));
    Span4Mux_v I__3299 (
            .O(N__23551),
            .I(N__23548));
    Odrv4 I__3298 (
            .O(N__23548),
            .I(da_pad_o_c_1));
    IoInMux I__3297 (
            .O(N__23545),
            .I(N__23542));
    LocalMux I__3296 (
            .O(N__23542),
            .I(N__23539));
    Span4Mux_s2_v I__3295 (
            .O(N__23539),
            .I(N__23536));
    Span4Mux_v I__3294 (
            .O(N__23536),
            .I(N__23533));
    Span4Mux_v I__3293 (
            .O(N__23533),
            .I(N__23530));
    Odrv4 I__3292 (
            .O(N__23530),
            .I(resetn_pad_o_c));
    InMux I__3291 (
            .O(N__23527),
            .I(N__23521));
    CascadeMux I__3290 (
            .O(N__23526),
            .I(N__23518));
    CascadeMux I__3289 (
            .O(N__23525),
            .I(N__23515));
    InMux I__3288 (
            .O(N__23524),
            .I(N__23507));
    LocalMux I__3287 (
            .O(N__23521),
            .I(N__23504));
    InMux I__3286 (
            .O(N__23518),
            .I(N__23501));
    InMux I__3285 (
            .O(N__23515),
            .I(N__23492));
    InMux I__3284 (
            .O(N__23514),
            .I(N__23492));
    InMux I__3283 (
            .O(N__23513),
            .I(N__23492));
    InMux I__3282 (
            .O(N__23512),
            .I(N__23492));
    InMux I__3281 (
            .O(N__23511),
            .I(N__23487));
    InMux I__3280 (
            .O(N__23510),
            .I(N__23487));
    LocalMux I__3279 (
            .O(N__23507),
            .I(N__23484));
    Span4Mux_h I__3278 (
            .O(N__23504),
            .I(N__23477));
    LocalMux I__3277 (
            .O(N__23501),
            .I(N__23477));
    LocalMux I__3276 (
            .O(N__23492),
            .I(N__23477));
    LocalMux I__3275 (
            .O(N__23487),
            .I(u1_PIO_control_gen_pingpong_ping_valid));
    Odrv12 I__3274 (
            .O(N__23484),
            .I(u1_PIO_control_gen_pingpong_ping_valid));
    Odrv4 I__3273 (
            .O(N__23477),
            .I(u1_PIO_control_gen_pingpong_ping_valid));
    InMux I__3272 (
            .O(N__23470),
            .I(N__23464));
    InMux I__3271 (
            .O(N__23469),
            .I(N__23464));
    LocalMux I__3270 (
            .O(N__23464),
            .I(N__23461));
    Span4Mux_h I__3269 (
            .O(N__23461),
            .I(N__23458));
    Odrv4 I__3268 (
            .O(N__23458),
            .I(\u1.PIO_control.dping_valid ));
    CascadeMux I__3267 (
            .O(N__23455),
            .I(N__23451));
    CascadeMux I__3266 (
            .O(N__23454),
            .I(N__23447));
    InMux I__3265 (
            .O(N__23451),
            .I(N__23440));
    InMux I__3264 (
            .O(N__23450),
            .I(N__23440));
    InMux I__3263 (
            .O(N__23447),
            .I(N__23440));
    LocalMux I__3262 (
            .O(N__23440),
            .I(N__23436));
    InMux I__3261 (
            .O(N__23439),
            .I(N__23433));
    Span4Mux_h I__3260 (
            .O(N__23436),
            .I(N__23430));
    LocalMux I__3259 (
            .O(N__23433),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.iQ_fast_3 ));
    Odrv4 I__3258 (
            .O(N__23430),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.iQ_fast_3 ));
    InMux I__3257 (
            .O(N__23425),
            .I(N__23421));
    InMux I__3256 (
            .O(N__23424),
            .I(N__23418));
    LocalMux I__3255 (
            .O(N__23421),
            .I(N__23415));
    LocalMux I__3254 (
            .O(N__23418),
            .I(N__23412));
    Odrv12 I__3253 (
            .O(N__23415),
            .I(DMA_dev0_Td_0));
    Odrv4 I__3252 (
            .O(N__23412),
            .I(DMA_dev0_Td_0));
    CascadeMux I__3251 (
            .O(N__23407),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.un1_ena_i_0_o3_sx_cascade_ ));
    InMux I__3250 (
            .O(N__23404),
            .I(N__23401));
    LocalMux I__3249 (
            .O(N__23401),
            .I(N__23398));
    Span4Mux_v I__3248 (
            .O(N__23398),
            .I(N__23395));
    Odrv4 I__3247 (
            .O(N__23395),
            .I(N_1364));
    InMux I__3246 (
            .O(N__23392),
            .I(N__23389));
    LocalMux I__3245 (
            .O(N__23389),
            .I(PIOq_10));
    CascadeMux I__3244 (
            .O(N__23386),
            .I(N_1364_cascade_));
    CascadeMux I__3243 (
            .O(N__23383),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.un1_ena_i_0_o3_0_cascade_ ));
    InMux I__3242 (
            .O(N__23380),
            .I(N__23377));
    LocalMux I__3241 (
            .O(N__23377),
            .I(N__23374));
    Span4Mux_v I__3240 (
            .O(N__23374),
            .I(N__23371));
    Odrv4 I__3239 (
            .O(N__23371),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.un1_ena_i_0_a2_sx ));
    CascadeMux I__3238 (
            .O(N__23368),
            .I(N__23363));
    CascadeMux I__3237 (
            .O(N__23367),
            .I(N__23359));
    InMux I__3236 (
            .O(N__23366),
            .I(N__23350));
    InMux I__3235 (
            .O(N__23363),
            .I(N__23350));
    InMux I__3234 (
            .O(N__23362),
            .I(N__23350));
    InMux I__3233 (
            .O(N__23359),
            .I(N__23350));
    LocalMux I__3232 (
            .O(N__23350),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.N_2092 ));
    InMux I__3231 (
            .O(N__23347),
            .I(N__23343));
    InMux I__3230 (
            .O(N__23346),
            .I(N__23340));
    LocalMux I__3229 (
            .O(N__23343),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.drd_ptr_2 ));
    LocalMux I__3228 (
            .O(N__23340),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.drd_ptr_2 ));
    InMux I__3227 (
            .O(N__23335),
            .I(N__23332));
    LocalMux I__3226 (
            .O(N__23332),
            .I(N__23329));
    Span4Mux_h I__3225 (
            .O(N__23329),
            .I(N__23325));
    InMux I__3224 (
            .O(N__23328),
            .I(N__23322));
    Odrv4 I__3223 (
            .O(N__23325),
            .I(\u1.DMA_control.N_1346 ));
    LocalMux I__3222 (
            .O(N__23322),
            .I(\u1.DMA_control.N_1346 ));
    CascadeMux I__3221 (
            .O(N__23317),
            .I(N__23314));
    InMux I__3220 (
            .O(N__23314),
            .I(N__23311));
    LocalMux I__3219 (
            .O(N__23311),
            .I(N__23308));
    Span4Mux_h I__3218 (
            .O(N__23308),
            .I(N__23304));
    InMux I__3217 (
            .O(N__23307),
            .I(N__23301));
    Odrv4 I__3216 (
            .O(N__23304),
            .I(\u1.DMA_control.gen_DMAbuf_Txbuf.N_1341 ));
    LocalMux I__3215 (
            .O(N__23301),
            .I(\u1.DMA_control.gen_DMAbuf_Txbuf.N_1341 ));
    InMux I__3214 (
            .O(N__23296),
            .I(N__23293));
    LocalMux I__3213 (
            .O(N__23293),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_s_6 ));
    InMux I__3212 (
            .O(N__23290),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_cry_5 ));
    InMux I__3211 (
            .O(N__23287),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_cry_6 ));
    InMux I__3210 (
            .O(N__23284),
            .I(N__23281));
    LocalMux I__3209 (
            .O(N__23281),
            .I(N__23277));
    InMux I__3208 (
            .O(N__23280),
            .I(N__23274));
    Span4Mux_h I__3207 (
            .O(N__23277),
            .I(N__23271));
    LocalMux I__3206 (
            .O(N__23274),
            .I(N__23268));
    Span4Mux_v I__3205 (
            .O(N__23271),
            .I(N__23265));
    Span4Mux_h I__3204 (
            .O(N__23268),
            .I(N__23262));
    Odrv4 I__3203 (
            .O(N__23265),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.N_1371 ));
    Odrv4 I__3202 (
            .O(N__23262),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.N_1371 ));
    CascadeMux I__3201 (
            .O(N__23257),
            .I(N__23253));
    InMux I__3200 (
            .O(N__23256),
            .I(N__23248));
    InMux I__3199 (
            .O(N__23253),
            .I(N__23245));
    InMux I__3198 (
            .O(N__23252),
            .I(N__23242));
    CascadeMux I__3197 (
            .O(N__23251),
            .I(N__23239));
    LocalMux I__3196 (
            .O(N__23248),
            .I(N__23234));
    LocalMux I__3195 (
            .O(N__23245),
            .I(N__23231));
    LocalMux I__3194 (
            .O(N__23242),
            .I(N__23228));
    InMux I__3193 (
            .O(N__23239),
            .I(N__23223));
    InMux I__3192 (
            .O(N__23238),
            .I(N__23223));
    InMux I__3191 (
            .O(N__23237),
            .I(N__23220));
    Span4Mux_v I__3190 (
            .O(N__23234),
            .I(N__23211));
    Span4Mux_v I__3189 (
            .O(N__23231),
            .I(N__23211));
    Span4Mux_v I__3188 (
            .O(N__23228),
            .I(N__23211));
    LocalMux I__3187 (
            .O(N__23223),
            .I(N__23211));
    LocalMux I__3186 (
            .O(N__23220),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.rci_0 ));
    Odrv4 I__3185 (
            .O(N__23211),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.rci_0 ));
    InMux I__3184 (
            .O(N__23206),
            .I(N__23200));
    InMux I__3183 (
            .O(N__23205),
            .I(N__23200));
    LocalMux I__3182 (
            .O(N__23200),
            .I(N__23196));
    InMux I__3181 (
            .O(N__23199),
            .I(N__23193));
    Odrv4 I__3180 (
            .O(N__23196),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.T1done_i ));
    LocalMux I__3179 (
            .O(N__23193),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.T1done_i ));
    CascadeMux I__3178 (
            .O(N__23188),
            .I(N__23185));
    InMux I__3177 (
            .O(N__23185),
            .I(N__23182));
    LocalMux I__3176 (
            .O(N__23182),
            .I(N__23179));
    Span4Mux_h I__3175 (
            .O(N__23179),
            .I(N__23176));
    Odrv4 I__3174 (
            .O(N__23176),
            .I(\u1.PIO_control.dsel_3_0_a2_0 ));
    InMux I__3173 (
            .O(N__23173),
            .I(N__23170));
    LocalMux I__3172 (
            .O(N__23170),
            .I(N__23167));
    Span4Mux_v I__3171 (
            .O(N__23167),
            .I(N__23163));
    InMux I__3170 (
            .O(N__23166),
            .I(N__23160));
    Odrv4 I__3169 (
            .O(N__23163),
            .I(\u1.PIO_control.N_2409 ));
    LocalMux I__3168 (
            .O(N__23160),
            .I(\u1.PIO_control.N_2409 ));
    CascadeMux I__3167 (
            .O(N__23155),
            .I(N__23152));
    InMux I__3166 (
            .O(N__23152),
            .I(N__23146));
    InMux I__3165 (
            .O(N__23151),
            .I(N__23146));
    LocalMux I__3164 (
            .O(N__23146),
            .I(N__23142));
    InMux I__3163 (
            .O(N__23145),
            .I(N__23139));
    Span4Mux_h I__3162 (
            .O(N__23142),
            .I(N__23136));
    LocalMux I__3161 (
            .O(N__23139),
            .I(\u1.PIO_control.dsel ));
    Odrv4 I__3160 (
            .O(N__23136),
            .I(\u1.PIO_control.dsel ));
    InMux I__3159 (
            .O(N__23131),
            .I(N__23127));
    InMux I__3158 (
            .O(N__23130),
            .I(N__23124));
    LocalMux I__3157 (
            .O(N__23127),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.QiZ0Z_1 ));
    LocalMux I__3156 (
            .O(N__23124),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.QiZ0Z_1 ));
    InMux I__3155 (
            .O(N__23119),
            .I(N__23116));
    LocalMux I__3154 (
            .O(N__23116),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_s_1 ));
    InMux I__3153 (
            .O(N__23113),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_cry_0 ));
    InMux I__3152 (
            .O(N__23110),
            .I(N__23106));
    InMux I__3151 (
            .O(N__23109),
            .I(N__23103));
    LocalMux I__3150 (
            .O(N__23106),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.QiZ0Z_2 ));
    LocalMux I__3149 (
            .O(N__23103),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.QiZ0Z_2 ));
    InMux I__3148 (
            .O(N__23098),
            .I(N__23095));
    LocalMux I__3147 (
            .O(N__23095),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_s_2 ));
    InMux I__3146 (
            .O(N__23092),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_cry_1 ));
    InMux I__3145 (
            .O(N__23089),
            .I(N__23085));
    InMux I__3144 (
            .O(N__23088),
            .I(N__23082));
    LocalMux I__3143 (
            .O(N__23085),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.QiZ0Z_3 ));
    LocalMux I__3142 (
            .O(N__23082),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.QiZ0Z_3 ));
    InMux I__3141 (
            .O(N__23077),
            .I(N__23074));
    LocalMux I__3140 (
            .O(N__23074),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_s_3 ));
    InMux I__3139 (
            .O(N__23071),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_cry_2 ));
    InMux I__3138 (
            .O(N__23068),
            .I(N__23064));
    InMux I__3137 (
            .O(N__23067),
            .I(N__23061));
    LocalMux I__3136 (
            .O(N__23064),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.QiZ0Z_4 ));
    LocalMux I__3135 (
            .O(N__23061),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.QiZ0Z_4 ));
    InMux I__3134 (
            .O(N__23056),
            .I(N__23053));
    LocalMux I__3133 (
            .O(N__23053),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_s_4 ));
    InMux I__3132 (
            .O(N__23050),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_cry_3 ));
    InMux I__3131 (
            .O(N__23047),
            .I(N__23043));
    InMux I__3130 (
            .O(N__23046),
            .I(N__23040));
    LocalMux I__3129 (
            .O(N__23043),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.QiZ0Z_5 ));
    LocalMux I__3128 (
            .O(N__23040),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.QiZ0Z_5 ));
    InMux I__3127 (
            .O(N__23035),
            .I(N__23032));
    LocalMux I__3126 (
            .O(N__23032),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_s_5 ));
    InMux I__3125 (
            .O(N__23029),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_cry_4 ));
    InMux I__3124 (
            .O(N__23026),
            .I(N__23022));
    InMux I__3123 (
            .O(N__23025),
            .I(N__23019));
    LocalMux I__3122 (
            .O(N__23022),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.QiZ0Z_6 ));
    LocalMux I__3121 (
            .O(N__23019),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.QiZ0Z_6 ));
    InMux I__3120 (
            .O(N__23014),
            .I(N__23011));
    LocalMux I__3119 (
            .O(N__23011),
            .I(N__23008));
    Span12Mux_s8_v I__3118 (
            .O(N__23008),
            .I(N__23005));
    Odrv12 I__3117 (
            .O(N__23005),
            .I(\u1.PIO_control.pong_d_12 ));
    InMux I__3116 (
            .O(N__23002),
            .I(N__22999));
    LocalMux I__3115 (
            .O(N__22999),
            .I(N__22996));
    Odrv4 I__3114 (
            .O(N__22996),
            .I(\u1.PIO_control.ping_d_12 ));
    InMux I__3113 (
            .O(N__22993),
            .I(N__22990));
    LocalMux I__3112 (
            .O(N__22990),
            .I(N__22987));
    Span12Mux_s6_v I__3111 (
            .O(N__22987),
            .I(N__22984));
    Odrv12 I__3110 (
            .O(N__22984),
            .I(\u1.PIO_control.pong_d_14 ));
    InMux I__3109 (
            .O(N__22981),
            .I(N__22978));
    LocalMux I__3108 (
            .O(N__22978),
            .I(N__22975));
    Odrv4 I__3107 (
            .O(N__22975),
            .I(\u1.PIO_control.ping_d_14 ));
    InMux I__3106 (
            .O(N__22972),
            .I(N__22969));
    LocalMux I__3105 (
            .O(N__22969),
            .I(N__22966));
    Span12Mux_s7_v I__3104 (
            .O(N__22966),
            .I(N__22963));
    Odrv12 I__3103 (
            .O(N__22963),
            .I(\u1.PIO_control.pong_d_13 ));
    InMux I__3102 (
            .O(N__22960),
            .I(N__22957));
    LocalMux I__3101 (
            .O(N__22957),
            .I(N__22954));
    Odrv4 I__3100 (
            .O(N__22954),
            .I(\u1.PIO_control.ping_d_13 ));
    InMux I__3099 (
            .O(N__22951),
            .I(N__22948));
    LocalMux I__3098 (
            .O(N__22948),
            .I(N__22945));
    Odrv4 I__3097 (
            .O(N__22945),
            .I(\u1.N_1446 ));
    InMux I__3096 (
            .O(N__22942),
            .I(N__22939));
    LocalMux I__3095 (
            .O(N__22939),
            .I(N__22936));
    Odrv4 I__3094 (
            .O(N__22936),
            .I(\u1.DMAd_12 ));
    InMux I__3093 (
            .O(N__22933),
            .I(N__22930));
    LocalMux I__3092 (
            .O(N__22930),
            .I(\u1.N_1447 ));
    IoInMux I__3091 (
            .O(N__22927),
            .I(N__22924));
    LocalMux I__3090 (
            .O(N__22924),
            .I(N__22921));
    Span4Mux_s3_v I__3089 (
            .O(N__22921),
            .I(N__22918));
    Odrv4 I__3088 (
            .O(N__22918),
            .I(dd_pad_o_c_12));
    InMux I__3087 (
            .O(N__22915),
            .I(N__22912));
    LocalMux I__3086 (
            .O(N__22912),
            .I(\u1.N_1445 ));
    InMux I__3085 (
            .O(N__22909),
            .I(N__22906));
    LocalMux I__3084 (
            .O(N__22906),
            .I(N__22903));
    Odrv4 I__3083 (
            .O(N__22903),
            .I(\u1.DMAd_14 ));
    IoInMux I__3082 (
            .O(N__22900),
            .I(N__22897));
    LocalMux I__3081 (
            .O(N__22897),
            .I(N__22894));
    Span4Mux_s3_v I__3080 (
            .O(N__22894),
            .I(N__22891));
    Odrv4 I__3079 (
            .O(N__22891),
            .I(dd_pad_o_c_14));
    InMux I__3078 (
            .O(N__22888),
            .I(N__22885));
    LocalMux I__3077 (
            .O(N__22885),
            .I(N__22882));
    Odrv4 I__3076 (
            .O(N__22882),
            .I(\u1.DMAd_8 ));
    InMux I__3075 (
            .O(N__22879),
            .I(N__22876));
    LocalMux I__3074 (
            .O(N__22876),
            .I(\u1.N_1433 ));
    IoInMux I__3073 (
            .O(N__22873),
            .I(N__22870));
    LocalMux I__3072 (
            .O(N__22870),
            .I(N__22867));
    Span4Mux_s3_v I__3071 (
            .O(N__22867),
            .I(N__22864));
    Odrv4 I__3070 (
            .O(N__22864),
            .I(dd_pad_o_c_8));
    InMux I__3069 (
            .O(N__22861),
            .I(N__22858));
    LocalMux I__3068 (
            .O(N__22858),
            .I(N__22855));
    Odrv4 I__3067 (
            .O(N__22855),
            .I(\u1.DMAd_7 ));
    InMux I__3066 (
            .O(N__22852),
            .I(N__22849));
    LocalMux I__3065 (
            .O(N__22849),
            .I(\u1.N_1432 ));
    IoInMux I__3064 (
            .O(N__22846),
            .I(N__22843));
    LocalMux I__3063 (
            .O(N__22843),
            .I(N__22840));
    Odrv12 I__3062 (
            .O(N__22840),
            .I(dd_pad_o_c_7));
    InMux I__3061 (
            .O(N__22837),
            .I(N__22834));
    LocalMux I__3060 (
            .O(N__22834),
            .I(N__22831));
    Span4Mux_v I__3059 (
            .O(N__22831),
            .I(N__22828));
    Span4Mux_v I__3058 (
            .O(N__22828),
            .I(N__22825));
    Odrv4 I__3057 (
            .O(N__22825),
            .I(\u0.N_1384 ));
    InMux I__3056 (
            .O(N__22822),
            .I(N__22819));
    LocalMux I__3055 (
            .O(N__22819),
            .I(N__22815));
    InMux I__3054 (
            .O(N__22818),
            .I(N__22812));
    Sp12to4 I__3053 (
            .O(N__22815),
            .I(N__22809));
    LocalMux I__3052 (
            .O(N__22812),
            .I(N__22806));
    Span12Mux_v I__3051 (
            .O(N__22809),
            .I(N__22803));
    Span4Mux_v I__3050 (
            .O(N__22806),
            .I(N__22800));
    Odrv12 I__3049 (
            .O(N__22803),
            .I(wb_sel_i_c_1));
    Odrv4 I__3048 (
            .O(N__22800),
            .I(wb_sel_i_c_1));
    CascadeMux I__3047 (
            .O(N__22795),
            .I(N__22792));
    InMux I__3046 (
            .O(N__22792),
            .I(N__22789));
    LocalMux I__3045 (
            .O(N__22789),
            .I(N__22786));
    Span12Mux_h I__3044 (
            .O(N__22786),
            .I(N__22783));
    Odrv12 I__3043 (
            .O(N__22783),
            .I(\u0.un1_piosel ));
    InMux I__3042 (
            .O(N__22780),
            .I(N__22777));
    LocalMux I__3041 (
            .O(N__22777),
            .I(N__22774));
    Span4Mux_v I__3040 (
            .O(N__22774),
            .I(N__22771));
    Span4Mux_h I__3039 (
            .O(N__22771),
            .I(N__22767));
    InMux I__3038 (
            .O(N__22770),
            .I(N__22764));
    Span4Mux_v I__3037 (
            .O(N__22767),
            .I(N__22759));
    LocalMux I__3036 (
            .O(N__22764),
            .I(N__22759));
    Span4Mux_v I__3035 (
            .O(N__22759),
            .I(N__22756));
    Odrv4 I__3034 (
            .O(N__22756),
            .I(wb_sel_i_c_0));
    IoInMux I__3033 (
            .O(N__22753),
            .I(N__22750));
    LocalMux I__3032 (
            .O(N__22750),
            .I(N__22747));
    IoSpan4Mux I__3031 (
            .O(N__22747),
            .I(N__22744));
    Span4Mux_s2_v I__3030 (
            .O(N__22744),
            .I(N__22741));
    Span4Mux_v I__3029 (
            .O(N__22741),
            .I(N__22738));
    Sp12to4 I__3028 (
            .O(N__22738),
            .I(N__22735));
    Span12Mux_v I__3027 (
            .O(N__22735),
            .I(N__22732));
    Span12Mux_h I__3026 (
            .O(N__22732),
            .I(N__22729));
    Odrv12 I__3025 (
            .O(N__22729),
            .I(N_284_i));
    InMux I__3024 (
            .O(N__22726),
            .I(N__22723));
    LocalMux I__3023 (
            .O(N__22723),
            .I(N__22720));
    Span4Mux_h I__3022 (
            .O(N__22720),
            .I(N__22716));
    InMux I__3021 (
            .O(N__22719),
            .I(N__22713));
    Odrv4 I__3020 (
            .O(N__22716),
            .I(\u1.DMA_control.TxbufQ_14 ));
    LocalMux I__3019 (
            .O(N__22713),
            .I(\u1.DMA_control.TxbufQ_14 ));
    CascadeMux I__3018 (
            .O(N__22708),
            .I(\u1.DMA_control.writeDfw_6_i_0_6_cascade_ ));
    InMux I__3017 (
            .O(N__22705),
            .I(N__22702));
    LocalMux I__3016 (
            .O(N__22702),
            .I(N__22699));
    Odrv4 I__3015 (
            .O(N__22699),
            .I(\u1.DMAd_6 ));
    InMux I__3014 (
            .O(N__22696),
            .I(N__22693));
    LocalMux I__3013 (
            .O(N__22693),
            .I(N__22690));
    Odrv4 I__3012 (
            .O(N__22690),
            .I(\u1.DMA_control.writeDlw_7 ));
    CascadeMux I__3011 (
            .O(N__22687),
            .I(N__22683));
    InMux I__3010 (
            .O(N__22686),
            .I(N__22680));
    InMux I__3009 (
            .O(N__22683),
            .I(N__22677));
    LocalMux I__3008 (
            .O(N__22680),
            .I(N__22674));
    LocalMux I__3007 (
            .O(N__22677),
            .I(N__22671));
    Span4Mux_v I__3006 (
            .O(N__22674),
            .I(N__22668));
    Odrv12 I__3005 (
            .O(N__22671),
            .I(\u1.DMA_control.TxbufQ_23 ));
    Odrv4 I__3004 (
            .O(N__22668),
            .I(\u1.DMA_control.TxbufQ_23 ));
    InMux I__3003 (
            .O(N__22663),
            .I(N__22660));
    LocalMux I__3002 (
            .O(N__22660),
            .I(N__22657));
    Span4Mux_h I__3001 (
            .O(N__22657),
            .I(N__22654));
    Span4Mux_h I__3000 (
            .O(N__22654),
            .I(N__22650));
    InMux I__2999 (
            .O(N__22653),
            .I(N__22647));
    Odrv4 I__2998 (
            .O(N__22650),
            .I(\u1.DMA_control.TxbufQ_15 ));
    LocalMux I__2997 (
            .O(N__22647),
            .I(\u1.DMA_control.TxbufQ_15 ));
    CascadeMux I__2996 (
            .O(N__22642),
            .I(\u1.DMA_control.writeDfw_6_i_0_7_cascade_ ));
    InMux I__2995 (
            .O(N__22639),
            .I(N__22636));
    LocalMux I__2994 (
            .O(N__22636),
            .I(N__22633));
    Odrv12 I__2993 (
            .O(N__22633),
            .I(\u1.DMA_control.writeDlw_8 ));
    InMux I__2992 (
            .O(N__22630),
            .I(N__22626));
    InMux I__2991 (
            .O(N__22629),
            .I(N__22623));
    LocalMux I__2990 (
            .O(N__22626),
            .I(N__22620));
    LocalMux I__2989 (
            .O(N__22623),
            .I(N__22617));
    Span4Mux_v I__2988 (
            .O(N__22620),
            .I(N__22614));
    Odrv12 I__2987 (
            .O(N__22617),
            .I(\u1.DMA_control.TxbufQ_24 ));
    Odrv4 I__2986 (
            .O(N__22614),
            .I(\u1.DMA_control.TxbufQ_24 ));
    InMux I__2985 (
            .O(N__22609),
            .I(N__22605));
    InMux I__2984 (
            .O(N__22608),
            .I(N__22602));
    LocalMux I__2983 (
            .O(N__22605),
            .I(N__22599));
    LocalMux I__2982 (
            .O(N__22602),
            .I(N__22594));
    Span4Mux_h I__2981 (
            .O(N__22599),
            .I(N__22594));
    Sp12to4 I__2980 (
            .O(N__22594),
            .I(N__22591));
    Span12Mux_s3_h I__2979 (
            .O(N__22591),
            .I(N__22588));
    Odrv12 I__2978 (
            .O(N__22588),
            .I(\u1.DMA_control.TxbufQ_0 ));
    CascadeMux I__2977 (
            .O(N__22585),
            .I(\u1.DMA_control.writeDfw_6_i_0_8_cascade_ ));
    InMux I__2976 (
            .O(N__22582),
            .I(N__22579));
    LocalMux I__2975 (
            .O(N__22579),
            .I(N__22576));
    Sp12to4 I__2974 (
            .O(N__22576),
            .I(N__22572));
    InMux I__2973 (
            .O(N__22575),
            .I(N__22569));
    Span12Mux_s6_v I__2972 (
            .O(N__22572),
            .I(N__22566));
    LocalMux I__2971 (
            .O(N__22569),
            .I(N__22563));
    Odrv12 I__2970 (
            .O(N__22566),
            .I(\u1.DMA_control.TxbufQ_13 ));
    Odrv4 I__2969 (
            .O(N__22563),
            .I(\u1.DMA_control.TxbufQ_13 ));
    InMux I__2968 (
            .O(N__22558),
            .I(N__22555));
    LocalMux I__2967 (
            .O(N__22555),
            .I(\u1.DMA_control.writeDfw_6_i_0_5 ));
    InMux I__2966 (
            .O(N__22552),
            .I(N__22549));
    LocalMux I__2965 (
            .O(N__22549),
            .I(N__22546));
    Odrv4 I__2964 (
            .O(N__22546),
            .I(\u1.DMAd_5 ));
    InMux I__2963 (
            .O(N__22543),
            .I(N__22540));
    LocalMux I__2962 (
            .O(N__22540),
            .I(N__22537));
    Span12Mux_s9_v I__2961 (
            .O(N__22537),
            .I(N__22534));
    Odrv12 I__2960 (
            .O(N__22534),
            .I(\u1.PIO_control.pong_d_11 ));
    InMux I__2959 (
            .O(N__22531),
            .I(N__22528));
    LocalMux I__2958 (
            .O(N__22528),
            .I(N__22525));
    Odrv4 I__2957 (
            .O(N__22525),
            .I(\u1.DMAd_11 ));
    CascadeMux I__2956 (
            .O(N__22522),
            .I(\u1.N_1448_cascade_ ));
    IoInMux I__2955 (
            .O(N__22519),
            .I(N__22516));
    LocalMux I__2954 (
            .O(N__22516),
            .I(N__22513));
    Span4Mux_s1_v I__2953 (
            .O(N__22513),
            .I(N__22510));
    Span4Mux_h I__2952 (
            .O(N__22510),
            .I(N__22507));
    Odrv4 I__2951 (
            .O(N__22507),
            .I(dd_pad_o_c_11));
    InMux I__2950 (
            .O(N__22504),
            .I(N__22501));
    LocalMux I__2949 (
            .O(N__22501),
            .I(N__22498));
    Span4Mux_v I__2948 (
            .O(N__22498),
            .I(N__22495));
    Span4Mux_h I__2947 (
            .O(N__22495),
            .I(N__22490));
    InMux I__2946 (
            .O(N__22494),
            .I(N__22487));
    InMux I__2945 (
            .O(N__22493),
            .I(N__22484));
    Odrv4 I__2944 (
            .O(N__22490),
            .I(\u1.DMA_control.dstrb ));
    LocalMux I__2943 (
            .O(N__22487),
            .I(\u1.DMA_control.dstrb ));
    LocalMux I__2942 (
            .O(N__22484),
            .I(\u1.DMA_control.dstrb ));
    InMux I__2941 (
            .O(N__22477),
            .I(N__22474));
    LocalMux I__2940 (
            .O(N__22474),
            .I(\u1.DMA_control.writeDfw_6_i_0_1 ));
    InMux I__2939 (
            .O(N__22471),
            .I(N__22467));
    CascadeMux I__2938 (
            .O(N__22470),
            .I(N__22464));
    LocalMux I__2937 (
            .O(N__22467),
            .I(N__22461));
    InMux I__2936 (
            .O(N__22464),
            .I(N__22458));
    Odrv4 I__2935 (
            .O(N__22461),
            .I(\u1.DMA_control.TxbufQ_9 ));
    LocalMux I__2934 (
            .O(N__22458),
            .I(\u1.DMA_control.TxbufQ_9 ));
    CascadeMux I__2933 (
            .O(N__22453),
            .I(N__22450));
    InMux I__2932 (
            .O(N__22450),
            .I(N__22447));
    LocalMux I__2931 (
            .O(N__22447),
            .I(N__22443));
    InMux I__2930 (
            .O(N__22446),
            .I(N__22440));
    Span4Mux_h I__2929 (
            .O(N__22443),
            .I(N__22437));
    LocalMux I__2928 (
            .O(N__22440),
            .I(N__22434));
    Odrv4 I__2927 (
            .O(N__22437),
            .I(\u1.DMA_control.TxbufQ_2 ));
    Odrv12 I__2926 (
            .O(N__22434),
            .I(\u1.DMA_control.TxbufQ_2 ));
    InMux I__2925 (
            .O(N__22429),
            .I(N__22426));
    LocalMux I__2924 (
            .O(N__22426),
            .I(N__22423));
    Odrv4 I__2923 (
            .O(N__22423),
            .I(\u1.DMAd_10 ));
    InMux I__2922 (
            .O(N__22420),
            .I(N__22417));
    LocalMux I__2921 (
            .O(N__22417),
            .I(\u1.DMA_control.writeDfw_6_i_0_11 ));
    CascadeMux I__2920 (
            .O(N__22414),
            .I(N__22411));
    InMux I__2919 (
            .O(N__22411),
            .I(N__22407));
    InMux I__2918 (
            .O(N__22410),
            .I(N__22404));
    LocalMux I__2917 (
            .O(N__22407),
            .I(N__22401));
    LocalMux I__2916 (
            .O(N__22404),
            .I(N__22398));
    Span4Mux_h I__2915 (
            .O(N__22401),
            .I(N__22395));
    Span4Mux_v I__2914 (
            .O(N__22398),
            .I(N__22392));
    Odrv4 I__2913 (
            .O(N__22395),
            .I(\u1.DMA_control.TxbufQ_3 ));
    Odrv4 I__2912 (
            .O(N__22392),
            .I(\u1.DMA_control.TxbufQ_3 ));
    CascadeMux I__2911 (
            .O(N__22387),
            .I(N__22384));
    InMux I__2910 (
            .O(N__22384),
            .I(N__22381));
    LocalMux I__2909 (
            .O(N__22381),
            .I(N__22377));
    InMux I__2908 (
            .O(N__22380),
            .I(N__22374));
    Span4Mux_h I__2907 (
            .O(N__22377),
            .I(N__22371));
    LocalMux I__2906 (
            .O(N__22374),
            .I(N__22368));
    Odrv4 I__2905 (
            .O(N__22371),
            .I(\u1.DMA_control.TxbufQ_4 ));
    Odrv12 I__2904 (
            .O(N__22368),
            .I(\u1.DMA_control.TxbufQ_4 ));
    InMux I__2903 (
            .O(N__22363),
            .I(N__22360));
    LocalMux I__2902 (
            .O(N__22360),
            .I(\u1.DMA_control.writeDfw_6_i_0_12 ));
    CascadeMux I__2901 (
            .O(N__22357),
            .I(N__22354));
    InMux I__2900 (
            .O(N__22354),
            .I(N__22351));
    LocalMux I__2899 (
            .O(N__22351),
            .I(N__22347));
    InMux I__2898 (
            .O(N__22350),
            .I(N__22344));
    Span4Mux_v I__2897 (
            .O(N__22347),
            .I(N__22339));
    LocalMux I__2896 (
            .O(N__22344),
            .I(N__22339));
    Odrv4 I__2895 (
            .O(N__22339),
            .I(\u1.DMA_control.TxbufQ_5 ));
    InMux I__2894 (
            .O(N__22336),
            .I(N__22333));
    LocalMux I__2893 (
            .O(N__22333),
            .I(N__22330));
    Span4Mux_v I__2892 (
            .O(N__22330),
            .I(N__22327));
    Odrv4 I__2891 (
            .O(N__22327),
            .I(\u1.DMAd_13 ));
    CascadeMux I__2890 (
            .O(N__22324),
            .I(N__22321));
    InMux I__2889 (
            .O(N__22321),
            .I(N__22317));
    InMux I__2888 (
            .O(N__22320),
            .I(N__22314));
    LocalMux I__2887 (
            .O(N__22317),
            .I(N__22311));
    LocalMux I__2886 (
            .O(N__22314),
            .I(N__22308));
    Span4Mux_h I__2885 (
            .O(N__22311),
            .I(N__22305));
    Span4Mux_h I__2884 (
            .O(N__22308),
            .I(N__22302));
    Odrv4 I__2883 (
            .O(N__22305),
            .I(\u1.DMA_control.TxbufQ_6 ));
    Odrv4 I__2882 (
            .O(N__22302),
            .I(\u1.DMA_control.TxbufQ_6 ));
    InMux I__2881 (
            .O(N__22297),
            .I(N__22294));
    LocalMux I__2880 (
            .O(N__22294),
            .I(\u1.DMA_control.writeDfw_6_i_m3_i_0_14 ));
    CascadeMux I__2879 (
            .O(N__22291),
            .I(N__22288));
    InMux I__2878 (
            .O(N__22288),
            .I(N__22284));
    InMux I__2877 (
            .O(N__22287),
            .I(N__22281));
    LocalMux I__2876 (
            .O(N__22284),
            .I(N__22276));
    LocalMux I__2875 (
            .O(N__22281),
            .I(N__22276));
    Span4Mux_v I__2874 (
            .O(N__22276),
            .I(N__22273));
    Odrv4 I__2873 (
            .O(N__22273),
            .I(\u1.DMA_control.TxbufQ_21 ));
    CascadeMux I__2872 (
            .O(N__22270),
            .I(N__22267));
    InMux I__2871 (
            .O(N__22267),
            .I(N__22264));
    LocalMux I__2870 (
            .O(N__22264),
            .I(N__22261));
    Odrv4 I__2869 (
            .O(N__22261),
            .I(\u1.DMA_control.writeDlw_5 ));
    InMux I__2868 (
            .O(N__22258),
            .I(N__22255));
    LocalMux I__2867 (
            .O(N__22255),
            .I(N__22252));
    Span4Mux_v I__2866 (
            .O(N__22252),
            .I(N__22249));
    Odrv4 I__2865 (
            .O(N__22249),
            .I(\u1.DMA_control.writeDlw_6 ));
    InMux I__2864 (
            .O(N__22246),
            .I(N__22243));
    LocalMux I__2863 (
            .O(N__22243),
            .I(N__22239));
    InMux I__2862 (
            .O(N__22242),
            .I(N__22236));
    Span4Mux_h I__2861 (
            .O(N__22239),
            .I(N__22233));
    LocalMux I__2860 (
            .O(N__22236),
            .I(\u1.DMA_control.TxbufQ_22 ));
    Odrv4 I__2859 (
            .O(N__22233),
            .I(\u1.DMA_control.TxbufQ_22 ));
    InMux I__2858 (
            .O(N__22228),
            .I(N__22225));
    LocalMux I__2857 (
            .O(N__22225),
            .I(N__22222));
    Span4Mux_h I__2856 (
            .O(N__22222),
            .I(N__22213));
    InMux I__2855 (
            .O(N__22221),
            .I(N__22200));
    InMux I__2854 (
            .O(N__22220),
            .I(N__22200));
    InMux I__2853 (
            .O(N__22219),
            .I(N__22200));
    InMux I__2852 (
            .O(N__22218),
            .I(N__22200));
    InMux I__2851 (
            .O(N__22217),
            .I(N__22200));
    InMux I__2850 (
            .O(N__22216),
            .I(N__22200));
    Odrv4 I__2849 (
            .O(N__22213),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.N_2413_iZ0 ));
    LocalMux I__2848 (
            .O(N__22200),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.N_2413_iZ0 ));
    InMux I__2847 (
            .O(N__22195),
            .I(N__22192));
    LocalMux I__2846 (
            .O(N__22192),
            .I(N__22189));
    Span4Mux_h I__2845 (
            .O(N__22189),
            .I(N__22186));
    Odrv4 I__2844 (
            .O(N__22186),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_s_7 ));
    InMux I__2843 (
            .O(N__22183),
            .I(N__22180));
    LocalMux I__2842 (
            .O(N__22180),
            .I(N__22176));
    InMux I__2841 (
            .O(N__22179),
            .I(N__22173));
    Span4Mux_v I__2840 (
            .O(N__22176),
            .I(N__22168));
    LocalMux I__2839 (
            .O(N__22173),
            .I(N__22168));
    Span4Mux_h I__2838 (
            .O(N__22168),
            .I(N__22165));
    Odrv4 I__2837 (
            .O(N__22165),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.QiZ0Z_7 ));
    CEMux I__2836 (
            .O(N__22162),
            .I(N__22159));
    LocalMux I__2835 (
            .O(N__22159),
            .I(N__22155));
    CEMux I__2834 (
            .O(N__22158),
            .I(N__22152));
    Span4Mux_v I__2833 (
            .O(N__22155),
            .I(N__22149));
    LocalMux I__2832 (
            .O(N__22152),
            .I(N__22146));
    Sp12to4 I__2831 (
            .O(N__22149),
            .I(N__22143));
    Span4Mux_s3_h I__2830 (
            .O(N__22146),
            .I(N__22140));
    Odrv12 I__2829 (
            .O(N__22143),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qie_0_iZ0 ));
    Odrv4 I__2828 (
            .O(N__22140),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qie_0_iZ0 ));
    InMux I__2827 (
            .O(N__22135),
            .I(N__22131));
    InMux I__2826 (
            .O(N__22134),
            .I(N__22128));
    LocalMux I__2825 (
            .O(N__22131),
            .I(\u1.DMA_control.TxbufQ_16 ));
    LocalMux I__2824 (
            .O(N__22128),
            .I(\u1.DMA_control.TxbufQ_16 ));
    InMux I__2823 (
            .O(N__22123),
            .I(N__22120));
    LocalMux I__2822 (
            .O(N__22120),
            .I(N__22117));
    Odrv4 I__2821 (
            .O(N__22117),
            .I(\u1.DMA_control.writeDlw_0 ));
    InMux I__2820 (
            .O(N__22114),
            .I(N__22110));
    InMux I__2819 (
            .O(N__22113),
            .I(N__22107));
    LocalMux I__2818 (
            .O(N__22110),
            .I(\u1.DMA_control.TxbufQ_17 ));
    LocalMux I__2817 (
            .O(N__22107),
            .I(\u1.DMA_control.TxbufQ_17 ));
    CascadeMux I__2816 (
            .O(N__22102),
            .I(N__22099));
    InMux I__2815 (
            .O(N__22099),
            .I(N__22096));
    LocalMux I__2814 (
            .O(N__22096),
            .I(N__22093));
    Odrv4 I__2813 (
            .O(N__22093),
            .I(\u1.DMA_control.writeDlw_1 ));
    InMux I__2812 (
            .O(N__22090),
            .I(N__22087));
    LocalMux I__2811 (
            .O(N__22087),
            .I(N__22083));
    InMux I__2810 (
            .O(N__22086),
            .I(N__22080));
    Odrv4 I__2809 (
            .O(N__22083),
            .I(\u1.DMA_control.TxbufQ_27 ));
    LocalMux I__2808 (
            .O(N__22080),
            .I(\u1.DMA_control.TxbufQ_27 ));
    CascadeMux I__2807 (
            .O(N__22075),
            .I(N__22072));
    InMux I__2806 (
            .O(N__22072),
            .I(N__22069));
    LocalMux I__2805 (
            .O(N__22069),
            .I(N__22066));
    Odrv4 I__2804 (
            .O(N__22066),
            .I(\u1.DMA_control.writeDlw_11 ));
    InMux I__2803 (
            .O(N__22063),
            .I(N__22059));
    InMux I__2802 (
            .O(N__22062),
            .I(N__22056));
    LocalMux I__2801 (
            .O(N__22059),
            .I(N__22053));
    LocalMux I__2800 (
            .O(N__22056),
            .I(\u1.DMA_control.TxbufQ_28 ));
    Odrv4 I__2799 (
            .O(N__22053),
            .I(\u1.DMA_control.TxbufQ_28 ));
    CascadeMux I__2798 (
            .O(N__22048),
            .I(N__22045));
    InMux I__2797 (
            .O(N__22045),
            .I(N__22042));
    LocalMux I__2796 (
            .O(N__22042),
            .I(N__22039));
    Odrv4 I__2795 (
            .O(N__22039),
            .I(\u1.DMA_control.writeDlw_12 ));
    InMux I__2794 (
            .O(N__22036),
            .I(N__22032));
    InMux I__2793 (
            .O(N__22035),
            .I(N__22029));
    LocalMux I__2792 (
            .O(N__22032),
            .I(N__22026));
    LocalMux I__2791 (
            .O(N__22029),
            .I(N__22023));
    Span4Mux_h I__2790 (
            .O(N__22026),
            .I(N__22020));
    Odrv4 I__2789 (
            .O(N__22023),
            .I(\u1.DMA_control.TxbufQ_30 ));
    Odrv4 I__2788 (
            .O(N__22020),
            .I(\u1.DMA_control.TxbufQ_30 ));
    CascadeMux I__2787 (
            .O(N__22015),
            .I(N__22012));
    InMux I__2786 (
            .O(N__22012),
            .I(N__22009));
    LocalMux I__2785 (
            .O(N__22009),
            .I(N__22006));
    Span4Mux_h I__2784 (
            .O(N__22006),
            .I(N__22003));
    Odrv4 I__2783 (
            .O(N__22003),
            .I(\u1.DMA_control.writeDlw_14 ));
    InMux I__2782 (
            .O(N__22000),
            .I(N__21997));
    LocalMux I__2781 (
            .O(N__21997),
            .I(\u1.DMA_control.writeDfw_6_i_0_0 ));
    CascadeMux I__2780 (
            .O(N__21994),
            .I(N__21991));
    InMux I__2779 (
            .O(N__21991),
            .I(N__21988));
    LocalMux I__2778 (
            .O(N__21988),
            .I(N__21984));
    InMux I__2777 (
            .O(N__21987),
            .I(N__21981));
    Span4Mux_h I__2776 (
            .O(N__21984),
            .I(N__21978));
    LocalMux I__2775 (
            .O(N__21981),
            .I(N__21975));
    Odrv4 I__2774 (
            .O(N__21978),
            .I(\u1.DMA_control.TxbufQ_8 ));
    Odrv4 I__2773 (
            .O(N__21975),
            .I(\u1.DMA_control.TxbufQ_8 ));
    InMux I__2772 (
            .O(N__21970),
            .I(N__21967));
    LocalMux I__2771 (
            .O(N__21967),
            .I(N__21964));
    Odrv4 I__2770 (
            .O(N__21964),
            .I(\u1.DMA_control.Td_0 ));
    InMux I__2769 (
            .O(N__21961),
            .I(N__21956));
    InMux I__2768 (
            .O(N__21960),
            .I(N__21952));
    InMux I__2767 (
            .O(N__21959),
            .I(N__21947));
    LocalMux I__2766 (
            .O(N__21956),
            .I(N__21944));
    InMux I__2765 (
            .O(N__21955),
            .I(N__21941));
    LocalMux I__2764 (
            .O(N__21952),
            .I(N__21937));
    CascadeMux I__2763 (
            .O(N__21951),
            .I(N__21934));
    CascadeMux I__2762 (
            .O(N__21950),
            .I(N__21931));
    LocalMux I__2761 (
            .O(N__21947),
            .I(N__21928));
    Span4Mux_v I__2760 (
            .O(N__21944),
            .I(N__21923));
    LocalMux I__2759 (
            .O(N__21941),
            .I(N__21923));
    InMux I__2758 (
            .O(N__21940),
            .I(N__21920));
    Span4Mux_v I__2757 (
            .O(N__21937),
            .I(N__21917));
    InMux I__2756 (
            .O(N__21934),
            .I(N__21914));
    InMux I__2755 (
            .O(N__21931),
            .I(N__21911));
    Span4Mux_v I__2754 (
            .O(N__21928),
            .I(N__21906));
    Span4Mux_v I__2753 (
            .O(N__21923),
            .I(N__21906));
    LocalMux I__2752 (
            .O(N__21920),
            .I(N__21903));
    Sp12to4 I__2751 (
            .O(N__21917),
            .I(N__21896));
    LocalMux I__2750 (
            .O(N__21914),
            .I(N__21896));
    LocalMux I__2749 (
            .O(N__21911),
            .I(N__21896));
    Span4Mux_h I__2748 (
            .O(N__21906),
            .I(N__21891));
    Span4Mux_v I__2747 (
            .O(N__21903),
            .I(N__21891));
    Odrv12 I__2746 (
            .O(N__21896),
            .I(wb_we_i_c));
    Odrv4 I__2745 (
            .O(N__21891),
            .I(wb_we_i_c));
    InMux I__2744 (
            .O(N__21886),
            .I(N__21880));
    InMux I__2743 (
            .O(N__21885),
            .I(N__21880));
    LocalMux I__2742 (
            .O(N__21880),
            .I(N__21877));
    Span4Mux_h I__2741 (
            .O(N__21877),
            .I(N__21874));
    Span4Mux_v I__2740 (
            .O(N__21874),
            .I(N__21870));
    InMux I__2739 (
            .O(N__21873),
            .I(N__21867));
    Sp12to4 I__2738 (
            .O(N__21870),
            .I(N__21862));
    LocalMux I__2737 (
            .O(N__21867),
            .I(N__21862));
    Span12Mux_v I__2736 (
            .O(N__21862),
            .I(N__21859));
    Odrv12 I__2735 (
            .O(N__21859),
            .I(wb_sel_i_c_3));
    CascadeMux I__2734 (
            .O(N__21856),
            .I(N__21853));
    InMux I__2733 (
            .O(N__21853),
            .I(N__21841));
    InMux I__2732 (
            .O(N__21852),
            .I(N__21841));
    InMux I__2731 (
            .O(N__21851),
            .I(N__21841));
    InMux I__2730 (
            .O(N__21850),
            .I(N__21841));
    LocalMux I__2729 (
            .O(N__21841),
            .I(N__21837));
    InMux I__2728 (
            .O(N__21840),
            .I(N__21834));
    Span4Mux_v I__2727 (
            .O(N__21837),
            .I(N__21831));
    LocalMux I__2726 (
            .O(N__21834),
            .I(N__21828));
    Span4Mux_h I__2725 (
            .O(N__21831),
            .I(N__21825));
    Span4Mux_v I__2724 (
            .O(N__21828),
            .I(N__21822));
    Span4Mux_v I__2723 (
            .O(N__21825),
            .I(N__21819));
    Span4Mux_v I__2722 (
            .O(N__21822),
            .I(N__21816));
    Span4Mux_v I__2721 (
            .O(N__21819),
            .I(N__21813));
    Span4Mux_v I__2720 (
            .O(N__21816),
            .I(N__21810));
    Odrv4 I__2719 (
            .O(N__21813),
            .I(N_1342));
    Odrv4 I__2718 (
            .O(N__21810),
            .I(N_1342));
    InMux I__2717 (
            .O(N__21805),
            .I(N__21800));
    InMux I__2716 (
            .O(N__21804),
            .I(N__21795));
    InMux I__2715 (
            .O(N__21803),
            .I(N__21795));
    LocalMux I__2714 (
            .O(N__21800),
            .I(N__21792));
    LocalMux I__2713 (
            .O(N__21795),
            .I(N__21789));
    Span4Mux_v I__2712 (
            .O(N__21792),
            .I(N__21786));
    Span12Mux_v I__2711 (
            .O(N__21789),
            .I(N__21783));
    Span4Mux_v I__2710 (
            .O(N__21786),
            .I(N__21780));
    Span12Mux_v I__2709 (
            .O(N__21783),
            .I(N__21777));
    Span4Mux_v I__2708 (
            .O(N__21780),
            .I(N__21774));
    Odrv12 I__2707 (
            .O(N__21777),
            .I(wb_sel_i_c_2));
    Odrv4 I__2706 (
            .O(N__21774),
            .I(wb_sel_i_c_2));
    InMux I__2705 (
            .O(N__21769),
            .I(N__21766));
    LocalMux I__2704 (
            .O(N__21766),
            .I(\u1.N_1435 ));
    IoInMux I__2703 (
            .O(N__21763),
            .I(N__21760));
    LocalMux I__2702 (
            .O(N__21760),
            .I(N__21757));
    Span4Mux_s3_v I__2701 (
            .O(N__21757),
            .I(N__21754));
    Span4Mux_h I__2700 (
            .O(N__21754),
            .I(N__21751));
    Sp12to4 I__2699 (
            .O(N__21751),
            .I(N__21748));
    Span12Mux_s11_v I__2698 (
            .O(N__21748),
            .I(N__21745));
    Span12Mux_h I__2697 (
            .O(N__21745),
            .I(N__21742));
    Odrv12 I__2696 (
            .O(N__21742),
            .I(dd_pad_o_c_10));
    CascadeMux I__2695 (
            .O(N__21739),
            .I(N__21736));
    InMux I__2694 (
            .O(N__21736),
            .I(N__21733));
    LocalMux I__2693 (
            .O(N__21733),
            .I(N__21730));
    Odrv4 I__2692 (
            .O(N__21730),
            .I(\u1.DMA_control.Td_3 ));
    InMux I__2691 (
            .O(N__21727),
            .I(N__21724));
    LocalMux I__2690 (
            .O(N__21724),
            .I(N__21721));
    Span4Mux_h I__2689 (
            .O(N__21721),
            .I(N__21718));
    Odrv4 I__2688 (
            .O(N__21718),
            .I(\u1.DMA_control.Td_4 ));
    InMux I__2687 (
            .O(N__21715),
            .I(N__21712));
    LocalMux I__2686 (
            .O(N__21712),
            .I(N__21709));
    Odrv4 I__2685 (
            .O(N__21709),
            .I(\u1.DMA_control.Td_7 ));
    CascadeMux I__2684 (
            .O(N__21706),
            .I(N__21702));
    InMux I__2683 (
            .O(N__21705),
            .I(N__21694));
    InMux I__2682 (
            .O(N__21702),
            .I(N__21694));
    InMux I__2681 (
            .O(N__21701),
            .I(N__21694));
    LocalMux I__2680 (
            .O(N__21694),
            .I(N__21690));
    InMux I__2679 (
            .O(N__21693),
            .I(N__21687));
    Odrv4 I__2678 (
            .O(N__21690),
            .I(N_1369));
    LocalMux I__2677 (
            .O(N__21687),
            .I(N_1369));
    InMux I__2676 (
            .O(N__21682),
            .I(N__21678));
    InMux I__2675 (
            .O(N__21681),
            .I(N__21675));
    LocalMux I__2674 (
            .O(N__21678),
            .I(N__21670));
    LocalMux I__2673 (
            .O(N__21675),
            .I(N__21670));
    Odrv4 I__2672 (
            .O(N__21670),
            .I(u1_PIO_control_gen_pingpong_iack));
    CascadeMux I__2671 (
            .O(N__21667),
            .I(\u0.N_1384_cascade_ ));
    CascadeMux I__2670 (
            .O(N__21664),
            .I(\u0.ack_o_i_i_1_cascade_ ));
    IoInMux I__2669 (
            .O(N__21661),
            .I(N__21658));
    LocalMux I__2668 (
            .O(N__21658),
            .I(N__21655));
    Span12Mux_s7_v I__2667 (
            .O(N__21655),
            .I(N__21652));
    Span12Mux_h I__2666 (
            .O(N__21652),
            .I(N__21649));
    Odrv12 I__2665 (
            .O(N__21649),
            .I(N_410_i));
    InMux I__2664 (
            .O(N__21646),
            .I(N__21638));
    InMux I__2663 (
            .O(N__21645),
            .I(N__21638));
    InMux I__2662 (
            .O(N__21644),
            .I(N__21635));
    InMux I__2661 (
            .O(N__21643),
            .I(N__21632));
    LocalMux I__2660 (
            .O(N__21638),
            .I(N_1360));
    LocalMux I__2659 (
            .O(N__21635),
            .I(N_1360));
    LocalMux I__2658 (
            .O(N__21632),
            .I(N_1360));
    IoInMux I__2657 (
            .O(N__21625),
            .I(N__21622));
    LocalMux I__2656 (
            .O(N__21622),
            .I(N__21619));
    Span12Mux_s6_v I__2655 (
            .O(N__21619),
            .I(N__21616));
    Span12Mux_h I__2654 (
            .O(N__21616),
            .I(N__21613));
    Odrv12 I__2653 (
            .O(N__21613),
            .I(N_288_i));
    InMux I__2652 (
            .O(N__21610),
            .I(N__21607));
    LocalMux I__2651 (
            .O(N__21607),
            .I(N__21604));
    Odrv4 I__2650 (
            .O(N__21604),
            .I(\u1.PIO_control.pong_d_10 ));
    CascadeMux I__2649 (
            .O(N__21601),
            .I(\u1.DMAtip_2_i_i_a2_0_1_cascade_ ));
    IoInMux I__2648 (
            .O(N__21598),
            .I(N__21595));
    LocalMux I__2647 (
            .O(N__21595),
            .I(N__21592));
    Span4Mux_s0_v I__2646 (
            .O(N__21592),
            .I(N__21589));
    Sp12to4 I__2645 (
            .O(N__21589),
            .I(N__21586));
    Span12Mux_h I__2644 (
            .O(N__21586),
            .I(N__21583));
    Span12Mux_v I__2643 (
            .O(N__21583),
            .I(N__21580));
    Odrv12 I__2642 (
            .O(N__21580),
            .I(dmackn_pad_o_c));
    InMux I__2641 (
            .O(N__21577),
            .I(N__21574));
    LocalMux I__2640 (
            .O(N__21574),
            .I(\u1.N_2150 ));
    InMux I__2639 (
            .O(N__21571),
            .I(N__21568));
    LocalMux I__2638 (
            .O(N__21568),
            .I(N__21565));
    Span4Mux_v I__2637 (
            .O(N__21565),
            .I(N__21562));
    Odrv4 I__2636 (
            .O(N__21562),
            .I(\u1.DMAtip_2_i_i_1 ));
    InMux I__2635 (
            .O(N__21559),
            .I(N__21556));
    LocalMux I__2634 (
            .O(N__21556),
            .I(N__21552));
    InMux I__2633 (
            .O(N__21555),
            .I(N__21549));
    Span4Mux_v I__2632 (
            .O(N__21552),
            .I(N__21543));
    LocalMux I__2631 (
            .O(N__21549),
            .I(N__21543));
    InMux I__2630 (
            .O(N__21548),
            .I(N__21540));
    Span4Mux_h I__2629 (
            .O(N__21543),
            .I(N__21537));
    LocalMux I__2628 (
            .O(N__21540),
            .I(\u1.Tdone_i ));
    Odrv4 I__2627 (
            .O(N__21537),
            .I(\u1.Tdone_i ));
    CascadeMux I__2626 (
            .O(N__21532),
            .I(\u1.N_2150_cascade_ ));
    InMux I__2625 (
            .O(N__21529),
            .I(N__21526));
    LocalMux I__2624 (
            .O(N__21526),
            .I(N__21523));
    Span4Mux_h I__2623 (
            .O(N__21523),
            .I(N__21519));
    InMux I__2622 (
            .O(N__21522),
            .I(N__21516));
    Odrv4 I__2621 (
            .O(N__21519),
            .I(\u1.N_1874 ));
    LocalMux I__2620 (
            .O(N__21516),
            .I(\u1.N_1874 ));
    InMux I__2619 (
            .O(N__21511),
            .I(N__21508));
    LocalMux I__2618 (
            .O(N__21508),
            .I(N__21505));
    Span4Mux_h I__2617 (
            .O(N__21505),
            .I(N__21502));
    Odrv4 I__2616 (
            .O(N__21502),
            .I(\u1.DMA_control.Tm_0 ));
    InMux I__2615 (
            .O(N__21499),
            .I(N__21494));
    CascadeMux I__2614 (
            .O(N__21498),
            .I(N__21491));
    InMux I__2613 (
            .O(N__21497),
            .I(N__21487));
    LocalMux I__2612 (
            .O(N__21494),
            .I(N__21484));
    InMux I__2611 (
            .O(N__21491),
            .I(N__21477));
    InMux I__2610 (
            .O(N__21490),
            .I(N__21477));
    LocalMux I__2609 (
            .O(N__21487),
            .I(N__21472));
    Span4Mux_h I__2608 (
            .O(N__21484),
            .I(N__21472));
    InMux I__2607 (
            .O(N__21483),
            .I(N__21469));
    InMux I__2606 (
            .O(N__21482),
            .I(N__21466));
    LocalMux I__2605 (
            .O(N__21477),
            .I(DMAtip));
    Odrv4 I__2604 (
            .O(N__21472),
            .I(DMAtip));
    LocalMux I__2603 (
            .O(N__21469),
            .I(DMAtip));
    LocalMux I__2602 (
            .O(N__21466),
            .I(DMAtip));
    InMux I__2601 (
            .O(N__21457),
            .I(N__21450));
    InMux I__2600 (
            .O(N__21456),
            .I(N__21450));
    InMux I__2599 (
            .O(N__21455),
            .I(N__21447));
    LocalMux I__2598 (
            .O(N__21450),
            .I(u0_gen_bc_dec_store_pp_full));
    LocalMux I__2597 (
            .O(N__21447),
            .I(u0_gen_bc_dec_store_pp_full));
    InMux I__2596 (
            .O(N__21442),
            .I(N__21439));
    LocalMux I__2595 (
            .O(N__21439),
            .I(N__21436));
    Span4Mux_h I__2594 (
            .O(N__21436),
            .I(N__21433));
    Odrv4 I__2593 (
            .O(N__21433),
            .I(\u1.DMA_control.Td_2 ));
    CascadeMux I__2592 (
            .O(N__21430),
            .I(N__21427));
    InMux I__2591 (
            .O(N__21427),
            .I(N__21420));
    InMux I__2590 (
            .O(N__21426),
            .I(N__21413));
    InMux I__2589 (
            .O(N__21425),
            .I(N__21413));
    InMux I__2588 (
            .O(N__21424),
            .I(N__21413));
    InMux I__2587 (
            .O(N__21423),
            .I(N__21410));
    LocalMux I__2586 (
            .O(N__21420),
            .I(N__21407));
    LocalMux I__2585 (
            .O(N__21413),
            .I(N__21404));
    LocalMux I__2584 (
            .O(N__21410),
            .I(N__21401));
    Span4Mux_v I__2583 (
            .O(N__21407),
            .I(N__21394));
    Span4Mux_v I__2582 (
            .O(N__21404),
            .I(N__21394));
    Span4Mux_h I__2581 (
            .O(N__21401),
            .I(N__21394));
    Span4Mux_h I__2580 (
            .O(N__21394),
            .I(N__21391));
    Odrv4 I__2579 (
            .O(N__21391),
            .I(DMA_dmarq));
    CascadeMux I__2578 (
            .O(N__21388),
            .I(\u1.c_state_RNIUC0A1Z0Z_1_cascade_ ));
    InMux I__2577 (
            .O(N__21385),
            .I(N__21382));
    LocalMux I__2576 (
            .O(N__21382),
            .I(N__21379));
    Odrv4 I__2575 (
            .O(N__21379),
            .I(\u1.DMAtip_2_i_i_a2_0_1 ));
    InMux I__2574 (
            .O(N__21376),
            .I(N__21370));
    InMux I__2573 (
            .O(N__21375),
            .I(N__21370));
    LocalMux I__2572 (
            .O(N__21370),
            .I(N__21367));
    Span4Mux_h I__2571 (
            .O(N__21367),
            .I(N__21362));
    InMux I__2570 (
            .O(N__21366),
            .I(N__21357));
    InMux I__2569 (
            .O(N__21365),
            .I(N__21357));
    Odrv4 I__2568 (
            .O(N__21362),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.val_c8_0_3 ));
    LocalMux I__2567 (
            .O(N__21357),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.val_c8_0_3 ));
    InMux I__2566 (
            .O(N__21352),
            .I(N__21349));
    LocalMux I__2565 (
            .O(N__21349),
            .I(N__21346));
    Span4Mux_v I__2564 (
            .O(N__21346),
            .I(N__21343));
    Odrv4 I__2563 (
            .O(N__21343),
            .I(\u1.PIO_control.pong_d_5 ));
    InMux I__2562 (
            .O(N__21340),
            .I(N__21337));
    LocalMux I__2561 (
            .O(N__21337),
            .I(N__21334));
    Odrv4 I__2560 (
            .O(N__21334),
            .I(\u1.PIO_control.ping_d_5 ));
    CascadeMux I__2559 (
            .O(N__21331),
            .I(\u1.N_1430_cascade_ ));
    IoInMux I__2558 (
            .O(N__21328),
            .I(N__21325));
    LocalMux I__2557 (
            .O(N__21325),
            .I(N__21322));
    Span4Mux_s0_v I__2556 (
            .O(N__21322),
            .I(N__21319));
    Odrv4 I__2555 (
            .O(N__21319),
            .I(dd_pad_o_c_5));
    InMux I__2554 (
            .O(N__21316),
            .I(N__21313));
    LocalMux I__2553 (
            .O(N__21313),
            .I(N__21310));
    Span4Mux_v I__2552 (
            .O(N__21310),
            .I(N__21307));
    Odrv4 I__2551 (
            .O(N__21307),
            .I(\u1.PIO_control.pong_d_6 ));
    InMux I__2550 (
            .O(N__21304),
            .I(N__21301));
    LocalMux I__2549 (
            .O(N__21301),
            .I(N__21298));
    Span12Mux_s7_v I__2548 (
            .O(N__21298),
            .I(N__21295));
    Odrv12 I__2547 (
            .O(N__21295),
            .I(\u1.PIO_control.ping_d_6 ));
    InMux I__2546 (
            .O(N__21292),
            .I(N__21289));
    LocalMux I__2545 (
            .O(N__21289),
            .I(N__21286));
    Span4Mux_v I__2544 (
            .O(N__21286),
            .I(N__21283));
    Odrv4 I__2543 (
            .O(N__21283),
            .I(\u1.PIO_control.pong_d_8 ));
    InMux I__2542 (
            .O(N__21280),
            .I(N__21277));
    LocalMux I__2541 (
            .O(N__21277),
            .I(N__21274));
    Span12Mux_s5_v I__2540 (
            .O(N__21274),
            .I(N__21271));
    Odrv12 I__2539 (
            .O(N__21271),
            .I(\u1.PIO_control.ping_d_8 ));
    InMux I__2538 (
            .O(N__21268),
            .I(N__21265));
    LocalMux I__2537 (
            .O(N__21265),
            .I(N__21262));
    Span4Mux_v I__2536 (
            .O(N__21262),
            .I(N__21259));
    Odrv4 I__2535 (
            .O(N__21259),
            .I(\u1.PIO_control.pong_d_7 ));
    InMux I__2534 (
            .O(N__21256),
            .I(N__21253));
    LocalMux I__2533 (
            .O(N__21253),
            .I(N__21250));
    Span12Mux_v I__2532 (
            .O(N__21250),
            .I(N__21247));
    Odrv12 I__2531 (
            .O(N__21247),
            .I(\u1.PIO_control.ping_d_7 ));
    IoInMux I__2530 (
            .O(N__21244),
            .I(N__21241));
    LocalMux I__2529 (
            .O(N__21241),
            .I(N__21238));
    Span4Mux_s2_v I__2528 (
            .O(N__21238),
            .I(N__21235));
    Odrv4 I__2527 (
            .O(N__21235),
            .I(dd_pad_o_c_13));
    InMux I__2526 (
            .O(N__21232),
            .I(N__21229));
    LocalMux I__2525 (
            .O(N__21229),
            .I(\u1.N_1431 ));
    IoInMux I__2524 (
            .O(N__21226),
            .I(N__21223));
    LocalMux I__2523 (
            .O(N__21223),
            .I(N__21220));
    Odrv4 I__2522 (
            .O(N__21220),
            .I(dd_pad_o_c_6));
    IoInMux I__2521 (
            .O(N__21217),
            .I(N__21214));
    LocalMux I__2520 (
            .O(N__21214),
            .I(N__21211));
    Span4Mux_s1_v I__2519 (
            .O(N__21211),
            .I(N__21208));
    Span4Mux_h I__2518 (
            .O(N__21208),
            .I(N__21205));
    Odrv4 I__2517 (
            .O(N__21205),
            .I(dd_pad_o_c_4));
    InMux I__2516 (
            .O(N__21202),
            .I(N__21199));
    LocalMux I__2515 (
            .O(N__21199),
            .I(N__21196));
    Span4Mux_v I__2514 (
            .O(N__21196),
            .I(N__21193));
    Odrv4 I__2513 (
            .O(N__21193),
            .I(\u1.PIO_control.dping_valid_3 ));
    InMux I__2512 (
            .O(N__21190),
            .I(N__21187));
    LocalMux I__2511 (
            .O(N__21187),
            .I(\u1.PIO_control.ping_d_15 ));
    InMux I__2510 (
            .O(N__21184),
            .I(N__21181));
    LocalMux I__2509 (
            .O(N__21181),
            .I(\u1.PIO_control.ping_d_2 ));
    InMux I__2508 (
            .O(N__21178),
            .I(N__21175));
    LocalMux I__2507 (
            .O(N__21175),
            .I(\u1.PIO_control.ping_d_3 ));
    InMux I__2506 (
            .O(N__21172),
            .I(N__21169));
    LocalMux I__2505 (
            .O(N__21169),
            .I(\u1.PIO_control.ping_d_4 ));
    CEMux I__2504 (
            .O(N__21166),
            .I(N__21154));
    CEMux I__2503 (
            .O(N__21165),
            .I(N__21154));
    CEMux I__2502 (
            .O(N__21164),
            .I(N__21154));
    CEMux I__2501 (
            .O(N__21163),
            .I(N__21154));
    GlobalMux I__2500 (
            .O(N__21154),
            .I(N__21151));
    gio2CtrlBuf I__2499 (
            .O(N__21151),
            .I(\u1.DMA_control.gen_DMAbuf_Txbuf.N_319_g ));
    InMux I__2498 (
            .O(N__21148),
            .I(N__21145));
    LocalMux I__2497 (
            .O(N__21145),
            .I(\u1.N_1359 ));
    CascadeMux I__2496 (
            .O(N__21142),
            .I(\u1.PIO_control.rpp_2_i_0_cascade_ ));
    CascadeMux I__2495 (
            .O(N__21139),
            .I(N__21131));
    InMux I__2494 (
            .O(N__21138),
            .I(N__21122));
    InMux I__2493 (
            .O(N__21137),
            .I(N__21122));
    InMux I__2492 (
            .O(N__21136),
            .I(N__21122));
    InMux I__2491 (
            .O(N__21135),
            .I(N__21117));
    InMux I__2490 (
            .O(N__21134),
            .I(N__21117));
    InMux I__2489 (
            .O(N__21131),
            .I(N__21114));
    InMux I__2488 (
            .O(N__21130),
            .I(N__21111));
    InMux I__2487 (
            .O(N__21129),
            .I(N__21108));
    LocalMux I__2486 (
            .O(N__21122),
            .I(N__21105));
    LocalMux I__2485 (
            .O(N__21117),
            .I(N__21100));
    LocalMux I__2484 (
            .O(N__21114),
            .I(N__21100));
    LocalMux I__2483 (
            .O(N__21111),
            .I(\u1.PIO_control.wpp ));
    LocalMux I__2482 (
            .O(N__21108),
            .I(\u1.PIO_control.wpp ));
    Odrv4 I__2481 (
            .O(N__21105),
            .I(\u1.PIO_control.wpp ));
    Odrv4 I__2480 (
            .O(N__21100),
            .I(\u1.PIO_control.wpp ));
    CascadeMux I__2479 (
            .O(N__21091),
            .I(N__21088));
    InMux I__2478 (
            .O(N__21088),
            .I(N__21085));
    LocalMux I__2477 (
            .O(N__21085),
            .I(N__21082));
    Odrv4 I__2476 (
            .O(N__21082),
            .I(\u1.PIO_control.pong_valid_3_0_a2_0 ));
    CascadeMux I__2475 (
            .O(N__21079),
            .I(N__21069));
    InMux I__2474 (
            .O(N__21078),
            .I(N__21061));
    InMux I__2473 (
            .O(N__21077),
            .I(N__21061));
    InMux I__2472 (
            .O(N__21076),
            .I(N__21061));
    InMux I__2471 (
            .O(N__21075),
            .I(N__21052));
    InMux I__2470 (
            .O(N__21074),
            .I(N__21052));
    InMux I__2469 (
            .O(N__21073),
            .I(N__21052));
    InMux I__2468 (
            .O(N__21072),
            .I(N__21052));
    InMux I__2467 (
            .O(N__21069),
            .I(N__21047));
    InMux I__2466 (
            .O(N__21068),
            .I(N__21047));
    LocalMux I__2465 (
            .O(N__21061),
            .I(N__21042));
    LocalMux I__2464 (
            .O(N__21052),
            .I(N__21042));
    LocalMux I__2463 (
            .O(N__21047),
            .I(u1_PIO_control_gen_pingpong_pong_valid));
    Odrv4 I__2462 (
            .O(N__21042),
            .I(u1_PIO_control_gen_pingpong_pong_valid));
    InMux I__2461 (
            .O(N__21037),
            .I(N__21033));
    InMux I__2460 (
            .O(N__21036),
            .I(N__21030));
    LocalMux I__2459 (
            .O(N__21033),
            .I(N__21027));
    LocalMux I__2458 (
            .O(N__21030),
            .I(\u1.PIO_control.dpong_valid ));
    Odrv4 I__2457 (
            .O(N__21027),
            .I(\u1.PIO_control.dpong_valid ));
    InMux I__2456 (
            .O(N__21022),
            .I(N__21016));
    InMux I__2455 (
            .O(N__21021),
            .I(N__21016));
    LocalMux I__2454 (
            .O(N__21016),
            .I(N__21011));
    CascadeMux I__2453 (
            .O(N__21015),
            .I(N__21008));
    CascadeMux I__2452 (
            .O(N__21014),
            .I(N__21004));
    Span4Mux_v I__2451 (
            .O(N__21011),
            .I(N__21001));
    InMux I__2450 (
            .O(N__21008),
            .I(N__20996));
    InMux I__2449 (
            .O(N__21007),
            .I(N__20996));
    InMux I__2448 (
            .O(N__21004),
            .I(N__20993));
    Odrv4 I__2447 (
            .O(N__21001),
            .I(\u1.DMAgoZ0 ));
    LocalMux I__2446 (
            .O(N__20996),
            .I(\u1.DMAgoZ0 ));
    LocalMux I__2445 (
            .O(N__20993),
            .I(\u1.DMAgoZ0 ));
    InMux I__2444 (
            .O(N__20986),
            .I(N__20983));
    LocalMux I__2443 (
            .O(N__20983),
            .I(\u1.DMA_control.hgo_2_i_0_0 ));
    InMux I__2442 (
            .O(N__20980),
            .I(N__20976));
    InMux I__2441 (
            .O(N__20979),
            .I(N__20973));
    LocalMux I__2440 (
            .O(N__20976),
            .I(\u1.DMA_control.hgo ));
    LocalMux I__2439 (
            .O(N__20973),
            .I(\u1.DMA_control.hgo ));
    InMux I__2438 (
            .O(N__20968),
            .I(N__20965));
    LocalMux I__2437 (
            .O(N__20965),
            .I(\u1.PIO_control.pong_valid_3_0_a2_0_1 ));
    InMux I__2436 (
            .O(N__20962),
            .I(N__20959));
    LocalMux I__2435 (
            .O(N__20959),
            .I(N__20956));
    Span4Mux_v I__2434 (
            .O(N__20956),
            .I(N__20953));
    Odrv4 I__2433 (
            .O(N__20953),
            .I(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.N_2138 ));
    CascadeMux I__2432 (
            .O(N__20950),
            .I(\u1.PIO_control.iack_7_u_0_0_1_cascade_ ));
    CascadeMux I__2431 (
            .O(N__20947),
            .I(\u1.PIO_control.iack_7_u_0_0_cascade_ ));
    InMux I__2430 (
            .O(N__20944),
            .I(N__20941));
    LocalMux I__2429 (
            .O(N__20941),
            .I(N__20937));
    InMux I__2428 (
            .O(N__20940),
            .I(N__20934));
    Span4Mux_v I__2427 (
            .O(N__20937),
            .I(N__20929));
    LocalMux I__2426 (
            .O(N__20934),
            .I(N__20929));
    Odrv4 I__2425 (
            .O(N__20929),
            .I(\u1.PIO_control.pong_we ));
    InMux I__2424 (
            .O(N__20926),
            .I(N__20923));
    LocalMux I__2423 (
            .O(N__20923),
            .I(N__20919));
    InMux I__2422 (
            .O(N__20922),
            .I(N__20916));
    Span4Mux_v I__2421 (
            .O(N__20919),
            .I(N__20911));
    LocalMux I__2420 (
            .O(N__20916),
            .I(N__20911));
    Odrv4 I__2419 (
            .O(N__20911),
            .I(\u1.PIO_control.ping_we ));
    InMux I__2418 (
            .O(N__20908),
            .I(N__20902));
    InMux I__2417 (
            .O(N__20907),
            .I(N__20902));
    LocalMux I__2416 (
            .O(N__20902),
            .I(\u1.PIO_control.N_1362 ));
    InMux I__2415 (
            .O(N__20899),
            .I(N__20896));
    LocalMux I__2414 (
            .O(N__20896),
            .I(N__20893));
    Odrv4 I__2413 (
            .O(N__20893),
            .I(\u1.PIO_control.iack_7_u_0_a2_1_1 ));
    InMux I__2412 (
            .O(N__20890),
            .I(N__20887));
    LocalMux I__2411 (
            .O(N__20887),
            .I(\u1.PIO_control.iack_7_u_0_a2_2_1 ));
    InMux I__2410 (
            .O(N__20884),
            .I(N__20880));
    InMux I__2409 (
            .O(N__20883),
            .I(N__20877));
    LocalMux I__2408 (
            .O(N__20880),
            .I(N__20874));
    LocalMux I__2407 (
            .O(N__20877),
            .I(N__20870));
    Span4Mux_v I__2406 (
            .O(N__20874),
            .I(N__20867));
    InMux I__2405 (
            .O(N__20873),
            .I(N__20864));
    Span4Mux_v I__2404 (
            .O(N__20870),
            .I(N__20861));
    Span4Mux_v I__2403 (
            .O(N__20867),
            .I(N__20856));
    LocalMux I__2402 (
            .O(N__20864),
            .I(N__20856));
    Odrv4 I__2401 (
            .O(N__20861),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.QiZ0Z_7 ));
    Odrv4 I__2400 (
            .O(N__20856),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.QiZ0Z_7 ));
    InMux I__2399 (
            .O(N__20851),
            .I(N__20847));
    InMux I__2398 (
            .O(N__20850),
            .I(N__20844));
    LocalMux I__2397 (
            .O(N__20847),
            .I(N__20841));
    LocalMux I__2396 (
            .O(N__20844),
            .I(N__20838));
    Odrv4 I__2395 (
            .O(N__20841),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.val_c7 ));
    Odrv12 I__2394 (
            .O(N__20838),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.val_c7 ));
    InMux I__2393 (
            .O(N__20833),
            .I(N__20830));
    LocalMux I__2392 (
            .O(N__20830),
            .I(N__20826));
    InMux I__2391 (
            .O(N__20829),
            .I(N__20823));
    Span4Mux_v I__2390 (
            .O(N__20826),
            .I(N__20820));
    LocalMux I__2389 (
            .O(N__20823),
            .I(N__20817));
    Odrv4 I__2388 (
            .O(N__20820),
            .I(\u1.N_1382 ));
    Odrv12 I__2387 (
            .O(N__20817),
            .I(\u1.N_1382 ));
    CascadeMux I__2386 (
            .O(N__20812),
            .I(\u1.PIOdone_i_cascade_ ));
    InMux I__2385 (
            .O(N__20809),
            .I(N__20806));
    LocalMux I__2384 (
            .O(N__20806),
            .I(N__20803));
    Span4Mux_h I__2383 (
            .O(N__20803),
            .I(N__20798));
    InMux I__2382 (
            .O(N__20802),
            .I(N__20793));
    InMux I__2381 (
            .O(N__20801),
            .I(N__20793));
    Odrv4 I__2380 (
            .O(N__20798),
            .I(\u1.N_1372 ));
    LocalMux I__2379 (
            .O(N__20793),
            .I(\u1.N_1372 ));
    InMux I__2378 (
            .O(N__20788),
            .I(N__20776));
    InMux I__2377 (
            .O(N__20787),
            .I(N__20776));
    InMux I__2376 (
            .O(N__20786),
            .I(N__20776));
    InMux I__2375 (
            .O(N__20785),
            .I(N__20776));
    LocalMux I__2374 (
            .O(N__20776),
            .I(N__20773));
    Odrv12 I__2373 (
            .O(N__20773),
            .I(\u1.PIOgoZ0 ));
    CascadeMux I__2372 (
            .O(N__20770),
            .I(N_468_cascade_));
    CascadeMux I__2371 (
            .O(N__20767),
            .I(\u1.PIO_control.N_2409_cascade_ ));
    CascadeMux I__2370 (
            .O(N__20764),
            .I(N__20761));
    InMux I__2369 (
            .O(N__20761),
            .I(N__20758));
    LocalMux I__2368 (
            .O(N__20758),
            .I(\u1.PIO_control.ping_valid_3_0_a2_0_1 ));
    CascadeMux I__2367 (
            .O(N__20755),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.val_c8_0_4_cascade_ ));
    CascadeMux I__2366 (
            .O(N__20752),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_1_sqmuxa_i_xZ0Z0_cascade_ ));
    InMux I__2365 (
            .O(N__20749),
            .I(N__20744));
    InMux I__2364 (
            .O(N__20748),
            .I(N__20739));
    InMux I__2363 (
            .O(N__20747),
            .I(N__20739));
    LocalMux I__2362 (
            .O(N__20744),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.val_c8_0_4 ));
    LocalMux I__2361 (
            .O(N__20739),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.val_c8_0_4 ));
    InMux I__2360 (
            .O(N__20734),
            .I(N__20731));
    LocalMux I__2359 (
            .O(N__20731),
            .I(N__20728));
    Odrv4 I__2358 (
            .O(N__20728),
            .I(\u1.sIORDYZ0 ));
    IoInMux I__2357 (
            .O(N__20725),
            .I(N__20722));
    LocalMux I__2356 (
            .O(N__20722),
            .I(N__20719));
    IoSpan4Mux I__2355 (
            .O(N__20719),
            .I(N__20716));
    Span4Mux_s3_v I__2354 (
            .O(N__20716),
            .I(N__20713));
    Span4Mux_v I__2353 (
            .O(N__20713),
            .I(N__20710));
    Span4Mux_h I__2352 (
            .O(N__20710),
            .I(N__20707));
    Span4Mux_v I__2351 (
            .O(N__20707),
            .I(N__20704));
    Span4Mux_h I__2350 (
            .O(N__20704),
            .I(N__20701));
    Odrv4 I__2349 (
            .O(N__20701),
            .I(da_pad_o_c_2));
    InMux I__2348 (
            .O(N__20698),
            .I(N__20693));
    InMux I__2347 (
            .O(N__20697),
            .I(N__20688));
    InMux I__2346 (
            .O(N__20696),
            .I(N__20688));
    LocalMux I__2345 (
            .O(N__20693),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.N_1358 ));
    LocalMux I__2344 (
            .O(N__20688),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.N_1358 ));
    CascadeMux I__2343 (
            .O(N__20683),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.N_1358_cascade_ ));
    CascadeMux I__2342 (
            .O(N__20680),
            .I(N__20677));
    InMux I__2341 (
            .O(N__20677),
            .I(N__20674));
    LocalMux I__2340 (
            .O(N__20674),
            .I(N__20669));
    InMux I__2339 (
            .O(N__20673),
            .I(N__20666));
    InMux I__2338 (
            .O(N__20672),
            .I(N__20663));
    Span4Mux_h I__2337 (
            .O(N__20669),
            .I(N__20660));
    LocalMux I__2336 (
            .O(N__20666),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.rciZ0 ));
    LocalMux I__2335 (
            .O(N__20663),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.rciZ0 ));
    Odrv4 I__2334 (
            .O(N__20660),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.rciZ0 ));
    CascadeMux I__2333 (
            .O(N__20653),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.N_1371_cascade_ ));
    CascadeMux I__2332 (
            .O(N__20650),
            .I(N__20647));
    InMux I__2331 (
            .O(N__20647),
            .I(N__20635));
    InMux I__2330 (
            .O(N__20646),
            .I(N__20635));
    InMux I__2329 (
            .O(N__20645),
            .I(N__20635));
    InMux I__2328 (
            .O(N__20644),
            .I(N__20635));
    LocalMux I__2327 (
            .O(N__20635),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.hold_goZ0 ));
    InMux I__2326 (
            .O(N__20632),
            .I(N__20620));
    InMux I__2325 (
            .O(N__20631),
            .I(N__20620));
    InMux I__2324 (
            .O(N__20630),
            .I(N__20620));
    InMux I__2323 (
            .O(N__20629),
            .I(N__20620));
    LocalMux I__2322 (
            .O(N__20620),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.busyZ0 ));
    InMux I__2321 (
            .O(N__20617),
            .I(N__20614));
    LocalMux I__2320 (
            .O(N__20614),
            .I(N__20611));
    Span4Mux_v I__2319 (
            .O(N__20611),
            .I(N__20608));
    Span4Mux_v I__2318 (
            .O(N__20608),
            .I(N__20605));
    Odrv4 I__2317 (
            .O(N__20605),
            .I(\u1.PIO_control.ping_d_9 ));
    InMux I__2316 (
            .O(N__20602),
            .I(N__20599));
    LocalMux I__2315 (
            .O(N__20599),
            .I(N__20596));
    Odrv4 I__2314 (
            .O(N__20596),
            .I(\u1.PIO_control.pong_d_15 ));
    InMux I__2313 (
            .O(N__20593),
            .I(N__20590));
    LocalMux I__2312 (
            .O(N__20590),
            .I(N__20587));
    Odrv4 I__2311 (
            .O(N__20587),
            .I(\u1.PIO_control.pong_d_4 ));
    InMux I__2310 (
            .O(N__20584),
            .I(N__20581));
    LocalMux I__2309 (
            .O(N__20581),
            .I(\u1.N_1436 ));
    IoInMux I__2308 (
            .O(N__20578),
            .I(N__20575));
    LocalMux I__2307 (
            .O(N__20575),
            .I(N__20572));
    Span4Mux_s1_v I__2306 (
            .O(N__20572),
            .I(N__20569));
    Span4Mux_h I__2305 (
            .O(N__20569),
            .I(N__20566));
    Odrv4 I__2304 (
            .O(N__20566),
            .I(dd_pad_o_c_15));
    InMux I__2303 (
            .O(N__20563),
            .I(N__20560));
    LocalMux I__2302 (
            .O(N__20560),
            .I(N__20555));
    CascadeMux I__2301 (
            .O(N__20559),
            .I(N__20552));
    InMux I__2300 (
            .O(N__20558),
            .I(N__20549));
    Span4Mux_h I__2299 (
            .O(N__20555),
            .I(N__20546));
    InMux I__2298 (
            .O(N__20552),
            .I(N__20543));
    LocalMux I__2297 (
            .O(N__20549),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.Qi_6 ));
    Odrv4 I__2296 (
            .O(N__20546),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.Qi_6 ));
    LocalMux I__2295 (
            .O(N__20543),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.Qi_6 ));
    InMux I__2294 (
            .O(N__20536),
            .I(N__20533));
    LocalMux I__2293 (
            .O(N__20533),
            .I(N__20530));
    Span4Mux_h I__2292 (
            .O(N__20530),
            .I(N__20525));
    InMux I__2291 (
            .O(N__20529),
            .I(N__20522));
    InMux I__2290 (
            .O(N__20528),
            .I(N__20519));
    Odrv4 I__2289 (
            .O(N__20525),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.Qi_5 ));
    LocalMux I__2288 (
            .O(N__20522),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.Qi_5 ));
    LocalMux I__2287 (
            .O(N__20519),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.Qi_5 ));
    CascadeMux I__2286 (
            .O(N__20512),
            .I(N__20509));
    InMux I__2285 (
            .O(N__20509),
            .I(N__20506));
    LocalMux I__2284 (
            .O(N__20506),
            .I(N__20502));
    InMux I__2283 (
            .O(N__20505),
            .I(N__20498));
    Span4Mux_h I__2282 (
            .O(N__20502),
            .I(N__20495));
    InMux I__2281 (
            .O(N__20501),
            .I(N__20492));
    LocalMux I__2280 (
            .O(N__20498),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.Qi_7 ));
    Odrv4 I__2279 (
            .O(N__20495),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.Qi_7 ));
    LocalMux I__2278 (
            .O(N__20492),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.Qi_7 ));
    InMux I__2277 (
            .O(N__20485),
            .I(N__20482));
    LocalMux I__2276 (
            .O(N__20482),
            .I(N__20479));
    Span4Mux_h I__2275 (
            .O(N__20479),
            .I(N__20474));
    InMux I__2274 (
            .O(N__20478),
            .I(N__20471));
    InMux I__2273 (
            .O(N__20477),
            .I(N__20468));
    Odrv4 I__2272 (
            .O(N__20474),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.Qi_2 ));
    LocalMux I__2271 (
            .O(N__20471),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.Qi_2 ));
    LocalMux I__2270 (
            .O(N__20468),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.Qi_2 ));
    InMux I__2269 (
            .O(N__20461),
            .I(N__20458));
    LocalMux I__2268 (
            .O(N__20458),
            .I(N__20455));
    Span4Mux_h I__2267 (
            .O(N__20455),
            .I(N__20450));
    InMux I__2266 (
            .O(N__20454),
            .I(N__20447));
    InMux I__2265 (
            .O(N__20453),
            .I(N__20444));
    Odrv4 I__2264 (
            .O(N__20450),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.Qi_4 ));
    LocalMux I__2263 (
            .O(N__20447),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.Qi_4 ));
    LocalMux I__2262 (
            .O(N__20444),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.Qi_4 ));
    InMux I__2261 (
            .O(N__20437),
            .I(N__20434));
    LocalMux I__2260 (
            .O(N__20434),
            .I(N__20431));
    Span4Mux_h I__2259 (
            .O(N__20431),
            .I(N__20426));
    InMux I__2258 (
            .O(N__20430),
            .I(N__20423));
    InMux I__2257 (
            .O(N__20429),
            .I(N__20420));
    Odrv4 I__2256 (
            .O(N__20426),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.Qi_3 ));
    LocalMux I__2255 (
            .O(N__20423),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.Qi_3 ));
    LocalMux I__2254 (
            .O(N__20420),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.Qi_3 ));
    CascadeMux I__2253 (
            .O(N__20413),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.val_c8_0_4_cascade_ ));
    InMux I__2252 (
            .O(N__20410),
            .I(N__20407));
    LocalMux I__2251 (
            .O(N__20407),
            .I(N__20404));
    Span4Mux_v I__2250 (
            .O(N__20404),
            .I(N__20399));
    InMux I__2249 (
            .O(N__20403),
            .I(N__20396));
    InMux I__2248 (
            .O(N__20402),
            .I(N__20393));
    Odrv4 I__2247 (
            .O(N__20399),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.Qi_1 ));
    LocalMux I__2246 (
            .O(N__20396),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.Qi_1 ));
    LocalMux I__2245 (
            .O(N__20393),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.Qi_1 ));
    InMux I__2244 (
            .O(N__20386),
            .I(N__20383));
    LocalMux I__2243 (
            .O(N__20383),
            .I(N__20377));
    InMux I__2242 (
            .O(N__20382),
            .I(N__20370));
    InMux I__2241 (
            .O(N__20381),
            .I(N__20370));
    InMux I__2240 (
            .O(N__20380),
            .I(N__20370));
    Odrv4 I__2239 (
            .O(N__20377),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.rci ));
    LocalMux I__2238 (
            .O(N__20370),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.rci ));
    CascadeMux I__2237 (
            .O(N__20365),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.val_c8_0_5_cascade_ ));
    InMux I__2236 (
            .O(N__20362),
            .I(N__20358));
    InMux I__2235 (
            .O(N__20361),
            .I(N__20355));
    LocalMux I__2234 (
            .O(N__20358),
            .I(N__20352));
    LocalMux I__2233 (
            .O(N__20355),
            .I(N__20349));
    Span4Mux_v I__2232 (
            .O(N__20352),
            .I(N__20342));
    Span4Mux_v I__2231 (
            .O(N__20349),
            .I(N__20342));
    InMux I__2230 (
            .O(N__20348),
            .I(N__20339));
    InMux I__2229 (
            .O(N__20347),
            .I(N__20336));
    Odrv4 I__2228 (
            .O(N__20342),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.Qi_0 ));
    LocalMux I__2227 (
            .O(N__20339),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.Qi_0 ));
    LocalMux I__2226 (
            .O(N__20336),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.Qi_0 ));
    InMux I__2225 (
            .O(N__20329),
            .I(N__20326));
    LocalMux I__2224 (
            .O(N__20326),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.busy_3_i_0 ));
    InMux I__2223 (
            .O(N__20323),
            .I(N__20320));
    LocalMux I__2222 (
            .O(N__20320),
            .I(N__20317));
    Odrv4 I__2221 (
            .O(N__20317),
            .I(\u1.PIO_control.pong_d_2 ));
    CascadeMux I__2220 (
            .O(N__20314),
            .I(\u1.N_1428_cascade_ ));
    IoInMux I__2219 (
            .O(N__20311),
            .I(N__20308));
    LocalMux I__2218 (
            .O(N__20308),
            .I(N__20305));
    Span4Mux_s2_v I__2217 (
            .O(N__20305),
            .I(N__20302));
    Span4Mux_h I__2216 (
            .O(N__20302),
            .I(N__20299));
    Odrv4 I__2215 (
            .O(N__20299),
            .I(dd_pad_o_c_2));
    InMux I__2214 (
            .O(N__20296),
            .I(N__20293));
    LocalMux I__2213 (
            .O(N__20293),
            .I(N__20290));
    Odrv12 I__2212 (
            .O(N__20290),
            .I(\u1.PIO_control.pong_d_3 ));
    CascadeMux I__2211 (
            .O(N__20287),
            .I(\u1.N_1449_cascade_ ));
    IoInMux I__2210 (
            .O(N__20284),
            .I(N__20281));
    LocalMux I__2209 (
            .O(N__20281),
            .I(N__20278));
    Span4Mux_s1_v I__2208 (
            .O(N__20278),
            .I(N__20275));
    Span4Mux_h I__2207 (
            .O(N__20275),
            .I(N__20272));
    Span4Mux_v I__2206 (
            .O(N__20272),
            .I(N__20269));
    Odrv4 I__2205 (
            .O(N__20269),
            .I(dd_pad_o_c_3));
    InMux I__2204 (
            .O(N__20266),
            .I(N__20260));
    InMux I__2203 (
            .O(N__20265),
            .I(N__20257));
    InMux I__2202 (
            .O(N__20264),
            .I(N__20252));
    InMux I__2201 (
            .O(N__20263),
            .I(N__20252));
    LocalMux I__2200 (
            .O(N__20260),
            .I(N__20246));
    LocalMux I__2199 (
            .O(N__20257),
            .I(N__20241));
    LocalMux I__2198 (
            .O(N__20252),
            .I(N__20241));
    InMux I__2197 (
            .O(N__20251),
            .I(N__20234));
    InMux I__2196 (
            .O(N__20250),
            .I(N__20234));
    InMux I__2195 (
            .O(N__20249),
            .I(N__20234));
    Span4Mux_v I__2194 (
            .O(N__20246),
            .I(N__20229));
    Span4Mux_v I__2193 (
            .O(N__20241),
            .I(N__20229));
    LocalMux I__2192 (
            .O(N__20234),
            .I(\u1.Tfw ));
    Odrv4 I__2191 (
            .O(N__20229),
            .I(\u1.Tfw ));
    CascadeMux I__2190 (
            .O(N__20224),
            .I(N__20221));
    InMux I__2189 (
            .O(N__20221),
            .I(N__20218));
    LocalMux I__2188 (
            .O(N__20218),
            .I(\u1.DMA_control.iDMA_req_2_0_0_a2_1 ));
    InMux I__2187 (
            .O(N__20215),
            .I(N__20212));
    LocalMux I__2186 (
            .O(N__20212),
            .I(\u1.DMA_control.N_1769 ));
    IoInMux I__2185 (
            .O(N__20209),
            .I(N__20206));
    LocalMux I__2184 (
            .O(N__20206),
            .I(N__20203));
    Span4Mux_s3_h I__2183 (
            .O(N__20203),
            .I(N__20200));
    Sp12to4 I__2182 (
            .O(N__20200),
            .I(N__20197));
    Span12Mux_v I__2181 (
            .O(N__20197),
            .I(N__20193));
    InMux I__2180 (
            .O(N__20196),
            .I(N__20190));
    Odrv12 I__2179 (
            .O(N__20193),
            .I(DMA_req_c));
    LocalMux I__2178 (
            .O(N__20190),
            .I(DMA_req_c));
    CascadeMux I__2177 (
            .O(N__20185),
            .I(\u1.DMA_control.iDMA_req_2_0_0_a2_0_2_cascade_ ));
    InMux I__2176 (
            .O(N__20182),
            .I(N__20176));
    InMux I__2175 (
            .O(N__20181),
            .I(N__20176));
    LocalMux I__2174 (
            .O(N__20176),
            .I(N__20173));
    Span4Mux_v I__2173 (
            .O(N__20173),
            .I(N__20170));
    Sp12to4 I__2172 (
            .O(N__20170),
            .I(N__20167));
    Span12Mux_s6_h I__2171 (
            .O(N__20167),
            .I(N__20164));
    Span12Mux_v I__2170 (
            .O(N__20164),
            .I(N__20161));
    Span12Mux_h I__2169 (
            .O(N__20161),
            .I(N__20158));
    Span12Mux_h I__2168 (
            .O(N__20158),
            .I(N__20155));
    Odrv12 I__2167 (
            .O(N__20155),
            .I(DMA_Ack_c));
    InMux I__2166 (
            .O(N__20152),
            .I(N__20146));
    InMux I__2165 (
            .O(N__20151),
            .I(N__20146));
    LocalMux I__2164 (
            .O(N__20146),
            .I(N__20143));
    Span4Mux_v I__2163 (
            .O(N__20143),
            .I(N__20140));
    Span4Mux_v I__2162 (
            .O(N__20140),
            .I(N__20137));
    Odrv4 I__2161 (
            .O(N__20137),
            .I(irq));
    InMux I__2160 (
            .O(N__20134),
            .I(N__20131));
    LocalMux I__2159 (
            .O(N__20131),
            .I(N__20128));
    Odrv4 I__2158 (
            .O(N__20128),
            .I(\u0.dirq ));
    InMux I__2157 (
            .O(N__20125),
            .I(N__20122));
    LocalMux I__2156 (
            .O(N__20122),
            .I(N__20119));
    Odrv4 I__2155 (
            .O(N__20119),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.DIOR_RNO_1_0 ));
    InMux I__2154 (
            .O(N__20116),
            .I(N__20113));
    LocalMux I__2153 (
            .O(N__20113),
            .I(N__20110));
    Odrv4 I__2152 (
            .O(N__20110),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.DIOR_RNOZ0Z_0 ));
    InMux I__2151 (
            .O(N__20107),
            .I(N__20102));
    InMux I__2150 (
            .O(N__20106),
            .I(N__20097));
    InMux I__2149 (
            .O(N__20105),
            .I(N__20097));
    LocalMux I__2148 (
            .O(N__20102),
            .I(N__20094));
    LocalMux I__2147 (
            .O(N__20097),
            .I(N__20091));
    Odrv12 I__2146 (
            .O(N__20094),
            .I(\u1.DMAdior ));
    Odrv4 I__2145 (
            .O(N__20091),
            .I(\u1.DMAdior ));
    InMux I__2144 (
            .O(N__20086),
            .I(N__20082));
    InMux I__2143 (
            .O(N__20085),
            .I(N__20079));
    LocalMux I__2142 (
            .O(N__20082),
            .I(N__20073));
    LocalMux I__2141 (
            .O(N__20079),
            .I(N__20073));
    InMux I__2140 (
            .O(N__20078),
            .I(N__20070));
    Span4Mux_h I__2139 (
            .O(N__20073),
            .I(N__20065));
    LocalMux I__2138 (
            .O(N__20070),
            .I(N__20065));
    Odrv4 I__2137 (
            .O(N__20065),
            .I(\u1.DMA_control.igo ));
    InMux I__2136 (
            .O(N__20062),
            .I(N__20054));
    InMux I__2135 (
            .O(N__20061),
            .I(N__20054));
    InMux I__2134 (
            .O(N__20060),
            .I(N__20049));
    InMux I__2133 (
            .O(N__20059),
            .I(N__20049));
    LocalMux I__2132 (
            .O(N__20054),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.rci ));
    LocalMux I__2131 (
            .O(N__20049),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.rci ));
    InMux I__2130 (
            .O(N__20044),
            .I(N__20034));
    InMux I__2129 (
            .O(N__20043),
            .I(N__20034));
    InMux I__2128 (
            .O(N__20042),
            .I(N__20034));
    InMux I__2127 (
            .O(N__20041),
            .I(N__20031));
    LocalMux I__2126 (
            .O(N__20034),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.Tmdone_i_i ));
    LocalMux I__2125 (
            .O(N__20031),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.Tmdone_i_i ));
    InMux I__2124 (
            .O(N__20026),
            .I(N__20023));
    LocalMux I__2123 (
            .O(N__20023),
            .I(N__20015));
    InMux I__2122 (
            .O(N__20022),
            .I(N__20010));
    InMux I__2121 (
            .O(N__20021),
            .I(N__20010));
    InMux I__2120 (
            .O(N__20020),
            .I(N__20003));
    InMux I__2119 (
            .O(N__20019),
            .I(N__20003));
    InMux I__2118 (
            .O(N__20018),
            .I(N__20003));
    Odrv4 I__2117 (
            .O(N__20015),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.Tddone_i ));
    LocalMux I__2116 (
            .O(N__20010),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.Tddone_i ));
    LocalMux I__2115 (
            .O(N__20003),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.Tddone_i ));
    CascadeMux I__2114 (
            .O(N__19996),
            .I(N__19992));
    CascadeMux I__2113 (
            .O(N__19995),
            .I(N__19989));
    InMux I__2112 (
            .O(N__19992),
            .I(N__19984));
    InMux I__2111 (
            .O(N__19989),
            .I(N__19984));
    LocalMux I__2110 (
            .O(N__19984),
            .I(N__19978));
    InMux I__2109 (
            .O(N__19983),
            .I(N__19975));
    InMux I__2108 (
            .O(N__19982),
            .I(N__19972));
    InMux I__2107 (
            .O(N__19981),
            .I(N__19969));
    Span4Mux_h I__2106 (
            .O(N__19978),
            .I(N__19966));
    LocalMux I__2105 (
            .O(N__19975),
            .I(N__19963));
    LocalMux I__2104 (
            .O(N__19972),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.rci_0 ));
    LocalMux I__2103 (
            .O(N__19969),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.rci_0 ));
    Odrv4 I__2102 (
            .O(N__19966),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.rci_0 ));
    Odrv4 I__2101 (
            .O(N__19963),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.rci_0 ));
    InMux I__2100 (
            .O(N__19954),
            .I(N__19951));
    LocalMux I__2099 (
            .O(N__19951),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_s_7 ));
    CascadeMux I__2098 (
            .O(N__19948),
            .I(N__19944));
    InMux I__2097 (
            .O(N__19947),
            .I(N__19941));
    InMux I__2096 (
            .O(N__19944),
            .I(N__19938));
    LocalMux I__2095 (
            .O(N__19941),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.QiZ0Z_7 ));
    LocalMux I__2094 (
            .O(N__19938),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.QiZ0Z_7 ));
    InMux I__2093 (
            .O(N__19933),
            .I(N__19930));
    LocalMux I__2092 (
            .O(N__19930),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_s_1 ));
    InMux I__2091 (
            .O(N__19927),
            .I(N__19923));
    InMux I__2090 (
            .O(N__19926),
            .I(N__19920));
    LocalMux I__2089 (
            .O(N__19923),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.QiZ0Z_1 ));
    LocalMux I__2088 (
            .O(N__19920),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.QiZ0Z_1 ));
    InMux I__2087 (
            .O(N__19915),
            .I(N__19908));
    InMux I__2086 (
            .O(N__19914),
            .I(N__19908));
    InMux I__2085 (
            .O(N__19913),
            .I(N__19905));
    LocalMux I__2084 (
            .O(N__19908),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.val_c8_0_3 ));
    LocalMux I__2083 (
            .O(N__19905),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.val_c8_0_3 ));
    InMux I__2082 (
            .O(N__19900),
            .I(N__19897));
    LocalMux I__2081 (
            .O(N__19897),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_s_3 ));
    InMux I__2080 (
            .O(N__19894),
            .I(N__19890));
    InMux I__2079 (
            .O(N__19893),
            .I(N__19887));
    LocalMux I__2078 (
            .O(N__19890),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.QiZ0Z_3 ));
    LocalMux I__2077 (
            .O(N__19887),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.QiZ0Z_3 ));
    CascadeMux I__2076 (
            .O(N__19882),
            .I(N__19879));
    InMux I__2075 (
            .O(N__19879),
            .I(N__19876));
    LocalMux I__2074 (
            .O(N__19876),
            .I(N__19873));
    Span4Mux_h I__2073 (
            .O(N__19873),
            .I(N__19870));
    Span4Mux_s0_h I__2072 (
            .O(N__19870),
            .I(N__19867));
    Odrv4 I__2071 (
            .O(N__19867),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_s_0 ));
    InMux I__2070 (
            .O(N__19864),
            .I(N__19861));
    LocalMux I__2069 (
            .O(N__19861),
            .I(N__19856));
    InMux I__2068 (
            .O(N__19860),
            .I(N__19851));
    InMux I__2067 (
            .O(N__19859),
            .I(N__19848));
    Span4Mux_h I__2066 (
            .O(N__19856),
            .I(N__19845));
    InMux I__2065 (
            .O(N__19855),
            .I(N__19840));
    InMux I__2064 (
            .O(N__19854),
            .I(N__19840));
    LocalMux I__2063 (
            .O(N__19851),
            .I(N__19835));
    LocalMux I__2062 (
            .O(N__19848),
            .I(N__19835));
    Odrv4 I__2061 (
            .O(N__19845),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.Qi_0_0 ));
    LocalMux I__2060 (
            .O(N__19840),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.Qi_0_0 ));
    Odrv4 I__2059 (
            .O(N__19835),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.Qi_0_0 ));
    InMux I__2058 (
            .O(N__19828),
            .I(N__19808));
    InMux I__2057 (
            .O(N__19827),
            .I(N__19808));
    InMux I__2056 (
            .O(N__19826),
            .I(N__19808));
    InMux I__2055 (
            .O(N__19825),
            .I(N__19808));
    InMux I__2054 (
            .O(N__19824),
            .I(N__19808));
    InMux I__2053 (
            .O(N__19823),
            .I(N__19808));
    InMux I__2052 (
            .O(N__19822),
            .I(N__19803));
    InMux I__2051 (
            .O(N__19821),
            .I(N__19803));
    LocalMux I__2050 (
            .O(N__19808),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.N_2415_i ));
    LocalMux I__2049 (
            .O(N__19803),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.N_2415_i ));
    InMux I__2048 (
            .O(N__19798),
            .I(N__19795));
    LocalMux I__2047 (
            .O(N__19795),
            .I(N__19792));
    Odrv4 I__2046 (
            .O(N__19792),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_s_4 ));
    CascadeMux I__2045 (
            .O(N__19789),
            .I(N__19786));
    InMux I__2044 (
            .O(N__19786),
            .I(N__19783));
    LocalMux I__2043 (
            .O(N__19783),
            .I(N__19779));
    InMux I__2042 (
            .O(N__19782),
            .I(N__19776));
    Odrv4 I__2041 (
            .O(N__19779),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.QiZ0Z_4 ));
    LocalMux I__2040 (
            .O(N__19776),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.QiZ0Z_4 ));
    CEMux I__2039 (
            .O(N__19771),
            .I(N__19767));
    CEMux I__2038 (
            .O(N__19770),
            .I(N__19764));
    LocalMux I__2037 (
            .O(N__19767),
            .I(N__19761));
    LocalMux I__2036 (
            .O(N__19764),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qie_0_iZ0 ));
    Odrv4 I__2035 (
            .O(N__19761),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qie_0_iZ0 ));
    InMux I__2034 (
            .O(N__19756),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_cry_2 ));
    InMux I__2033 (
            .O(N__19753),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_cry_3 ));
    InMux I__2032 (
            .O(N__19750),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_cry_4 ));
    InMux I__2031 (
            .O(N__19747),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_cry_5 ));
    InMux I__2030 (
            .O(N__19744),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_cry_6 ));
    InMux I__2029 (
            .O(N__19741),
            .I(N__19738));
    LocalMux I__2028 (
            .O(N__19738),
            .I(N__19735));
    Span4Mux_s3_h I__2027 (
            .O(N__19735),
            .I(N__19730));
    InMux I__2026 (
            .O(N__19734),
            .I(N__19725));
    InMux I__2025 (
            .O(N__19733),
            .I(N__19725));
    Odrv4 I__2024 (
            .O(N__19730),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.val_c8_0_4 ));
    LocalMux I__2023 (
            .O(N__19725),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.val_c8_0_4 ));
    InMux I__2022 (
            .O(N__19720),
            .I(N__19717));
    LocalMux I__2021 (
            .O(N__19717),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_s_2 ));
    CascadeMux I__2020 (
            .O(N__19714),
            .I(N__19711));
    InMux I__2019 (
            .O(N__19711),
            .I(N__19707));
    InMux I__2018 (
            .O(N__19710),
            .I(N__19704));
    LocalMux I__2017 (
            .O(N__19707),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.QiZ0Z_2 ));
    LocalMux I__2016 (
            .O(N__19704),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.QiZ0Z_2 ));
    InMux I__2015 (
            .O(N__19699),
            .I(N__19696));
    LocalMux I__2014 (
            .O(N__19696),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_s_5 ));
    InMux I__2013 (
            .O(N__19693),
            .I(N__19689));
    InMux I__2012 (
            .O(N__19692),
            .I(N__19686));
    LocalMux I__2011 (
            .O(N__19689),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.QiZ0Z_5 ));
    LocalMux I__2010 (
            .O(N__19686),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.QiZ0Z_5 ));
    InMux I__2009 (
            .O(N__19681),
            .I(N__19678));
    LocalMux I__2008 (
            .O(N__19678),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_s_6 ));
    CascadeMux I__2007 (
            .O(N__19675),
            .I(N__19672));
    InMux I__2006 (
            .O(N__19672),
            .I(N__19668));
    InMux I__2005 (
            .O(N__19671),
            .I(N__19665));
    LocalMux I__2004 (
            .O(N__19668),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.QiZ0Z_6 ));
    LocalMux I__2003 (
            .O(N__19665),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.QiZ0Z_6 ));
    CascadeMux I__2002 (
            .O(N__19660),
            .I(N__19657));
    InMux I__2001 (
            .O(N__19657),
            .I(N__19653));
    InMux I__2000 (
            .O(N__19656),
            .I(N__19650));
    LocalMux I__1999 (
            .O(N__19653),
            .I(\u1.PIOdior ));
    LocalMux I__1998 (
            .O(N__19650),
            .I(\u1.PIOdior ));
    IoInMux I__1997 (
            .O(N__19645),
            .I(N__19642));
    LocalMux I__1996 (
            .O(N__19642),
            .I(N__19639));
    Span4Mux_s3_v I__1995 (
            .O(N__19639),
            .I(N__19636));
    Span4Mux_h I__1994 (
            .O(N__19636),
            .I(N__19633));
    Sp12to4 I__1993 (
            .O(N__19633),
            .I(N__19630));
    Span12Mux_v I__1992 (
            .O(N__19630),
            .I(N__19627));
    Span12Mux_h I__1991 (
            .O(N__19627),
            .I(N__19624));
    Odrv12 I__1990 (
            .O(N__19624),
            .I(diorn_pad_o_c));
    InMux I__1989 (
            .O(N__19621),
            .I(N__19618));
    LocalMux I__1988 (
            .O(N__19618),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.DIOR_RNOZ0Z_1 ));
    CascadeMux I__1987 (
            .O(N__19615),
            .I(\u1.PIO_control.N_1450_cascade_ ));
    CascadeMux I__1986 (
            .O(N__19612),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.DIOW_RNOZ0Z_1_cascade_ ));
    CascadeMux I__1985 (
            .O(N__19609),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.N_1378_cascade_ ));
    InMux I__1984 (
            .O(N__19606),
            .I(N__19603));
    LocalMux I__1983 (
            .O(N__19603),
            .I(N__19600));
    Span4Mux_v I__1982 (
            .O(N__19600),
            .I(N__19596));
    InMux I__1981 (
            .O(N__19599),
            .I(N__19593));
    Odrv4 I__1980 (
            .O(N__19596),
            .I(\u1.PIOdiow ));
    LocalMux I__1979 (
            .O(N__19593),
            .I(\u1.PIOdiow ));
    InMux I__1978 (
            .O(N__19588),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_cry_0 ));
    InMux I__1977 (
            .O(N__19585),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_cry_1 ));
    InMux I__1976 (
            .O(N__19582),
            .I(N__19579));
    LocalMux I__1975 (
            .O(N__19579),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qilde_i_sxZ0 ));
    CascadeMux I__1974 (
            .O(N__19576),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.rci_3_i_a0_4_cascade_ ));
    CascadeMux I__1973 (
            .O(N__19573),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qilde_i_sxZ0_cascade_ ));
    CEMux I__1972 (
            .O(N__19570),
            .I(N__19567));
    LocalMux I__1971 (
            .O(N__19567),
            .I(N__19564));
    Span4Mux_s3_h I__1970 (
            .O(N__19564),
            .I(N__19561));
    Odrv4 I__1969 (
            .O(N__19561),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.N_1083 ));
    InMux I__1968 (
            .O(N__19558),
            .I(N__19555));
    LocalMux I__1967 (
            .O(N__19555),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.rci_3_i_a0_5 ));
    CascadeMux I__1966 (
            .O(N__19552),
            .I(N__19549));
    InMux I__1965 (
            .O(N__19549),
            .I(N__19546));
    LocalMux I__1964 (
            .O(N__19546),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.rci_3_i_a0_6 ));
    CascadeMux I__1963 (
            .O(N__19543),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.N_1377_cascade_ ));
    InMux I__1962 (
            .O(N__19540),
            .I(N__19537));
    LocalMux I__1961 (
            .O(N__19537),
            .I(N__19534));
    Span4Mux_v I__1960 (
            .O(N__19534),
            .I(N__19531));
    Odrv4 I__1959 (
            .O(N__19531),
            .I(iordy_pad_i_c));
    InMux I__1958 (
            .O(N__19528),
            .I(N__19525));
    LocalMux I__1957 (
            .O(N__19525),
            .I(N__19522));
    Odrv12 I__1956 (
            .O(N__19522),
            .I(\u1.cIORDY ));
    InMux I__1955 (
            .O(N__19519),
            .I(N__19516));
    LocalMux I__1954 (
            .O(N__19516),
            .I(N__19513));
    Span4Mux_v I__1953 (
            .O(N__19513),
            .I(N__19510));
    Span4Mux_h I__1952 (
            .O(N__19510),
            .I(N__19507));
    Odrv4 I__1951 (
            .O(N__19507),
            .I(\u1.PIO_control.pong_d_9 ));
    CascadeMux I__1950 (
            .O(N__19504),
            .I(\u1.N_1434_cascade_ ));
    IoInMux I__1949 (
            .O(N__19501),
            .I(N__19498));
    LocalMux I__1948 (
            .O(N__19498),
            .I(N__19495));
    Span12Mux_s9_v I__1947 (
            .O(N__19495),
            .I(N__19492));
    Odrv12 I__1946 (
            .O(N__19492),
            .I(dd_pad_o_c_9));
    InMux I__1945 (
            .O(N__19489),
            .I(N__19483));
    InMux I__1944 (
            .O(N__19488),
            .I(N__19483));
    LocalMux I__1943 (
            .O(N__19483),
            .I(\u1.N_1387 ));
    CascadeMux I__1942 (
            .O(N__19480),
            .I(N__19477));
    InMux I__1941 (
            .O(N__19477),
            .I(N__19473));
    InMux I__1940 (
            .O(N__19476),
            .I(N__19470));
    LocalMux I__1939 (
            .O(N__19473),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.QiZ0Z_6 ));
    LocalMux I__1938 (
            .O(N__19470),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.QiZ0Z_6 ));
    InMux I__1937 (
            .O(N__19465),
            .I(N__19461));
    InMux I__1936 (
            .O(N__19464),
            .I(N__19458));
    LocalMux I__1935 (
            .O(N__19461),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.QiZ0Z_5 ));
    LocalMux I__1934 (
            .O(N__19458),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.QiZ0Z_5 ));
    InMux I__1933 (
            .O(N__19453),
            .I(N__19450));
    LocalMux I__1932 (
            .O(N__19450),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.val_c8_a0_3 ));
    CascadeMux I__1931 (
            .O(N__19447),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.val_c8_a0_3_cascade_ ));
    InMux I__1930 (
            .O(N__19444),
            .I(N__19441));
    LocalMux I__1929 (
            .O(N__19441),
            .I(N__19435));
    InMux I__1928 (
            .O(N__19440),
            .I(N__19430));
    InMux I__1927 (
            .O(N__19439),
            .I(N__19430));
    InMux I__1926 (
            .O(N__19438),
            .I(N__19427));
    Odrv4 I__1925 (
            .O(N__19435),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.Qi_0 ));
    LocalMux I__1924 (
            .O(N__19430),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.Qi_0 ));
    LocalMux I__1923 (
            .O(N__19427),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.Qi_0 ));
    CascadeMux I__1922 (
            .O(N__19420),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.N_2415_i_xZ0Z1_cascade_ ));
    InMux I__1921 (
            .O(N__19417),
            .I(N__19414));
    LocalMux I__1920 (
            .O(N__19414),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.val_c8_a0_4 ));
    InMux I__1919 (
            .O(N__19411),
            .I(N__19408));
    LocalMux I__1918 (
            .O(N__19408),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.DIOW_RNO_1_0 ));
    InMux I__1917 (
            .O(N__19405),
            .I(N__19402));
    LocalMux I__1916 (
            .O(N__19402),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.DIOW_RNOZ0Z_0 ));
    InMux I__1915 (
            .O(N__19399),
            .I(N__19394));
    InMux I__1914 (
            .O(N__19398),
            .I(N__19391));
    InMux I__1913 (
            .O(N__19397),
            .I(N__19388));
    LocalMux I__1912 (
            .O(N__19394),
            .I(\u1.DMAdiow ));
    LocalMux I__1911 (
            .O(N__19391),
            .I(\u1.DMAdiow ));
    LocalMux I__1910 (
            .O(N__19388),
            .I(\u1.DMAdiow ));
    CascadeMux I__1909 (
            .O(N__19381),
            .I(\u1.N_1395_cascade_ ));
    IoInMux I__1908 (
            .O(N__19378),
            .I(N__19375));
    LocalMux I__1907 (
            .O(N__19375),
            .I(N__19372));
    IoSpan4Mux I__1906 (
            .O(N__19372),
            .I(N__19369));
    IoSpan4Mux I__1905 (
            .O(N__19369),
            .I(N__19366));
    Span4Mux_s1_v I__1904 (
            .O(N__19366),
            .I(N__19363));
    Span4Mux_v I__1903 (
            .O(N__19363),
            .I(N__19360));
    Span4Mux_v I__1902 (
            .O(N__19360),
            .I(N__19357));
    Odrv4 I__1901 (
            .O(N__19357),
            .I(dd_padoe_o_c));
    CascadeMux I__1900 (
            .O(N__19354),
            .I(\u1.N_1387_cascade_ ));
    InMux I__1899 (
            .O(N__19351),
            .I(N__19347));
    InMux I__1898 (
            .O(N__19350),
            .I(N__19344));
    LocalMux I__1897 (
            .O(N__19347),
            .I(\u1.PIOoe ));
    LocalMux I__1896 (
            .O(N__19344),
            .I(\u1.PIOoe ));
    CascadeMux I__1895 (
            .O(N__19339),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.Tddone_i_cascade_ ));
    IoInMux I__1894 (
            .O(N__19336),
            .I(N__19333));
    LocalMux I__1893 (
            .O(N__19333),
            .I(N__19330));
    Span4Mux_s2_h I__1892 (
            .O(N__19330),
            .I(N__19327));
    Sp12to4 I__1891 (
            .O(N__19327),
            .I(N__19324));
    Span12Mux_s9_v I__1890 (
            .O(N__19324),
            .I(N__19321));
    Odrv12 I__1889 (
            .O(N__19321),
            .I(diown_pad_o_c));
    InMux I__1888 (
            .O(N__19318),
            .I(N__19314));
    InMux I__1887 (
            .O(N__19317),
            .I(N__19311));
    LocalMux I__1886 (
            .O(N__19314),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.QiZ0Z_3 ));
    LocalMux I__1885 (
            .O(N__19311),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.QiZ0Z_3 ));
    CascadeMux I__1884 (
            .O(N__19306),
            .I(N__19302));
    InMux I__1883 (
            .O(N__19305),
            .I(N__19299));
    InMux I__1882 (
            .O(N__19302),
            .I(N__19296));
    LocalMux I__1881 (
            .O(N__19299),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.QiZ0Z_2 ));
    LocalMux I__1880 (
            .O(N__19296),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.QiZ0Z_2 ));
    CascadeMux I__1879 (
            .O(N__19291),
            .I(N__19287));
    CascadeMux I__1878 (
            .O(N__19290),
            .I(N__19284));
    InMux I__1877 (
            .O(N__19287),
            .I(N__19281));
    InMux I__1876 (
            .O(N__19284),
            .I(N__19278));
    LocalMux I__1875 (
            .O(N__19281),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.QiZ0Z_4 ));
    LocalMux I__1874 (
            .O(N__19278),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.QiZ0Z_4 ));
    InMux I__1873 (
            .O(N__19273),
            .I(N__19269));
    InMux I__1872 (
            .O(N__19272),
            .I(N__19266));
    LocalMux I__1871 (
            .O(N__19269),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.QiZ0Z_1 ));
    LocalMux I__1870 (
            .O(N__19266),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.QiZ0Z_1 ));
    CascadeMux I__1869 (
            .O(N__19261),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.val_c8_a0_4_cascade_ ));
    CascadeMux I__1868 (
            .O(N__19258),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.Tmdone_i_i_cascade_ ));
    InMux I__1867 (
            .O(N__19255),
            .I(N__19252));
    LocalMux I__1866 (
            .O(N__19252),
            .I(N__19249));
    Span4Mux_h I__1865 (
            .O(N__19249),
            .I(N__19246));
    Odrv4 I__1864 (
            .O(N__19246),
            .I(\u1.DMA_control.Teoc_1 ));
    InMux I__1863 (
            .O(N__19243),
            .I(N__19240));
    LocalMux I__1862 (
            .O(N__19240),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_s_1 ));
    InMux I__1861 (
            .O(N__19237),
            .I(N__19233));
    InMux I__1860 (
            .O(N__19236),
            .I(N__19230));
    LocalMux I__1859 (
            .O(N__19233),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.QiZ0Z_1 ));
    LocalMux I__1858 (
            .O(N__19230),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.QiZ0Z_1 ));
    InMux I__1857 (
            .O(N__19225),
            .I(N__19222));
    LocalMux I__1856 (
            .O(N__19222),
            .I(N__19219));
    Odrv4 I__1855 (
            .O(N__19219),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_s_3 ));
    InMux I__1854 (
            .O(N__19216),
            .I(N__19213));
    LocalMux I__1853 (
            .O(N__19213),
            .I(N__19209));
    InMux I__1852 (
            .O(N__19212),
            .I(N__19206));
    Odrv4 I__1851 (
            .O(N__19209),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.QiZ0Z_3 ));
    LocalMux I__1850 (
            .O(N__19206),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.QiZ0Z_3 ));
    InMux I__1849 (
            .O(N__19201),
            .I(N__19198));
    LocalMux I__1848 (
            .O(N__19198),
            .I(N__19195));
    Span4Mux_h I__1847 (
            .O(N__19195),
            .I(N__19192));
    Odrv4 I__1846 (
            .O(N__19192),
            .I(\u1.DMA_control.Teoc_4 ));
    InMux I__1845 (
            .O(N__19189),
            .I(N__19186));
    LocalMux I__1844 (
            .O(N__19186),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_s_4 ));
    CascadeMux I__1843 (
            .O(N__19183),
            .I(N__19180));
    InMux I__1842 (
            .O(N__19180),
            .I(N__19176));
    InMux I__1841 (
            .O(N__19179),
            .I(N__19173));
    LocalMux I__1840 (
            .O(N__19176),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.QiZ0Z_4 ));
    LocalMux I__1839 (
            .O(N__19173),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.QiZ0Z_4 ));
    InMux I__1838 (
            .O(N__19168),
            .I(N__19165));
    LocalMux I__1837 (
            .O(N__19165),
            .I(N__19162));
    Span4Mux_h I__1836 (
            .O(N__19162),
            .I(N__19159));
    Odrv4 I__1835 (
            .O(N__19159),
            .I(\u1.DMA_control.Teoc_5 ));
    InMux I__1834 (
            .O(N__19156),
            .I(N__19153));
    LocalMux I__1833 (
            .O(N__19153),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_s_5 ));
    InMux I__1832 (
            .O(N__19150),
            .I(N__19146));
    InMux I__1831 (
            .O(N__19149),
            .I(N__19143));
    LocalMux I__1830 (
            .O(N__19146),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.QiZ0Z_5 ));
    LocalMux I__1829 (
            .O(N__19143),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.QiZ0Z_5 ));
    InMux I__1828 (
            .O(N__19138),
            .I(N__19120));
    InMux I__1827 (
            .O(N__19137),
            .I(N__19120));
    InMux I__1826 (
            .O(N__19136),
            .I(N__19120));
    InMux I__1825 (
            .O(N__19135),
            .I(N__19120));
    InMux I__1824 (
            .O(N__19134),
            .I(N__19120));
    InMux I__1823 (
            .O(N__19133),
            .I(N__19115));
    InMux I__1822 (
            .O(N__19132),
            .I(N__19115));
    InMux I__1821 (
            .O(N__19131),
            .I(N__19112));
    LocalMux I__1820 (
            .O(N__19120),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_1_sqmuxa_i ));
    LocalMux I__1819 (
            .O(N__19115),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_1_sqmuxa_i ));
    LocalMux I__1818 (
            .O(N__19112),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_1_sqmuxa_i ));
    InMux I__1817 (
            .O(N__19105),
            .I(N__19102));
    LocalMux I__1816 (
            .O(N__19102),
            .I(N__19099));
    Span4Mux_h I__1815 (
            .O(N__19099),
            .I(N__19096));
    Odrv4 I__1814 (
            .O(N__19096),
            .I(\u1.DMA_control.Teoc_6 ));
    InMux I__1813 (
            .O(N__19093),
            .I(N__19090));
    LocalMux I__1812 (
            .O(N__19090),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_s_6 ));
    CascadeMux I__1811 (
            .O(N__19087),
            .I(N__19083));
    InMux I__1810 (
            .O(N__19086),
            .I(N__19080));
    InMux I__1809 (
            .O(N__19083),
            .I(N__19077));
    LocalMux I__1808 (
            .O(N__19080),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.QiZ0Z_6 ));
    LocalMux I__1807 (
            .O(N__19077),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.QiZ0Z_6 ));
    CEMux I__1806 (
            .O(N__19072),
            .I(N__19067));
    CEMux I__1805 (
            .O(N__19071),
            .I(N__19064));
    CEMux I__1804 (
            .O(N__19070),
            .I(N__19061));
    LocalMux I__1803 (
            .O(N__19067),
            .I(N__19058));
    LocalMux I__1802 (
            .O(N__19064),
            .I(N__19055));
    LocalMux I__1801 (
            .O(N__19061),
            .I(N__19052));
    Odrv4 I__1800 (
            .O(N__19058),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qie_0_iZ0 ));
    Odrv4 I__1799 (
            .O(N__19055),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qie_0_iZ0 ));
    Odrv4 I__1798 (
            .O(N__19052),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qie_0_iZ0 ));
    IoInMux I__1797 (
            .O(N__19045),
            .I(N__19042));
    LocalMux I__1796 (
            .O(N__19042),
            .I(N__19039));
    Span4Mux_s2_v I__1795 (
            .O(N__19039),
            .I(N__19036));
    Sp12to4 I__1794 (
            .O(N__19036),
            .I(N__19033));
    Span12Mux_h I__1793 (
            .O(N__19033),
            .I(N__19030));
    Odrv12 I__1792 (
            .O(N__19030),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.rd_dstrb ));
    CascadeMux I__1791 (
            .O(N__19027),
            .I(N__19024));
    InMux I__1790 (
            .O(N__19024),
            .I(N__19021));
    LocalMux I__1789 (
            .O(N__19021),
            .I(N__19017));
    InMux I__1788 (
            .O(N__19020),
            .I(N__19014));
    Odrv4 I__1787 (
            .O(N__19017),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.QiZ0Z_3 ));
    LocalMux I__1786 (
            .O(N__19014),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.QiZ0Z_3 ));
    InMux I__1785 (
            .O(N__19009),
            .I(N__19006));
    LocalMux I__1784 (
            .O(N__19006),
            .I(N__19002));
    InMux I__1783 (
            .O(N__19005),
            .I(N__18999));
    Odrv4 I__1782 (
            .O(N__19002),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.QiZ0Z_1 ));
    LocalMux I__1781 (
            .O(N__18999),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.QiZ0Z_1 ));
    CascadeMux I__1780 (
            .O(N__18994),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNIPRNIZ0Z_0_cascade_ ));
    InMux I__1779 (
            .O(N__18991),
            .I(N__18987));
    CascadeMux I__1778 (
            .O(N__18990),
            .I(N__18984));
    LocalMux I__1777 (
            .O(N__18987),
            .I(N__18981));
    InMux I__1776 (
            .O(N__18984),
            .I(N__18978));
    Odrv4 I__1775 (
            .O(N__18981),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.QiZ0Z_6 ));
    LocalMux I__1774 (
            .O(N__18978),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.QiZ0Z_6 ));
    InMux I__1773 (
            .O(N__18973),
            .I(N__18970));
    LocalMux I__1772 (
            .O(N__18970),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.val_c7_0_3 ));
    InMux I__1771 (
            .O(N__18967),
            .I(N__18964));
    LocalMux I__1770 (
            .O(N__18964),
            .I(N__18961));
    Span4Mux_h I__1769 (
            .O(N__18961),
            .I(N__18958));
    Odrv4 I__1768 (
            .O(N__18958),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_s_2 ));
    InMux I__1767 (
            .O(N__18955),
            .I(N__18952));
    LocalMux I__1766 (
            .O(N__18952),
            .I(N__18949));
    Span4Mux_s2_h I__1765 (
            .O(N__18949),
            .I(N__18945));
    InMux I__1764 (
            .O(N__18948),
            .I(N__18942));
    Odrv4 I__1763 (
            .O(N__18945),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.QiZ0Z_2 ));
    LocalMux I__1762 (
            .O(N__18942),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.QiZ0Z_2 ));
    CascadeMux I__1761 (
            .O(N__18937),
            .I(N__18934));
    InMux I__1760 (
            .O(N__18934),
            .I(N__18931));
    LocalMux I__1759 (
            .O(N__18931),
            .I(N__18928));
    Span4Mux_v I__1758 (
            .O(N__18928),
            .I(N__18925));
    Odrv4 I__1757 (
            .O(N__18925),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_s_4 ));
    InMux I__1756 (
            .O(N__18922),
            .I(N__18919));
    LocalMux I__1755 (
            .O(N__18919),
            .I(N__18916));
    Span4Mux_s2_h I__1754 (
            .O(N__18916),
            .I(N__18912));
    InMux I__1753 (
            .O(N__18915),
            .I(N__18909));
    Odrv4 I__1752 (
            .O(N__18912),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.QiZ0Z_4 ));
    LocalMux I__1751 (
            .O(N__18909),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.QiZ0Z_4 ));
    InMux I__1750 (
            .O(N__18904),
            .I(N__18901));
    LocalMux I__1749 (
            .O(N__18901),
            .I(N__18898));
    Span4Mux_h I__1748 (
            .O(N__18898),
            .I(N__18895));
    Odrv4 I__1747 (
            .O(N__18895),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_s_0 ));
    InMux I__1746 (
            .O(N__18892),
            .I(N__18889));
    LocalMux I__1745 (
            .O(N__18889),
            .I(N__18885));
    InMux I__1744 (
            .O(N__18888),
            .I(N__18882));
    Span4Mux_v I__1743 (
            .O(N__18885),
            .I(N__18879));
    LocalMux I__1742 (
            .O(N__18882),
            .I(N__18876));
    IoSpan4Mux I__1741 (
            .O(N__18879),
            .I(N__18872));
    Span4Mux_s2_h I__1740 (
            .O(N__18876),
            .I(N__18869));
    InMux I__1739 (
            .O(N__18875),
            .I(N__18866));
    Odrv4 I__1738 (
            .O(N__18872),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.QiZ0Z_0 ));
    Odrv4 I__1737 (
            .O(N__18869),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.QiZ0Z_0 ));
    LocalMux I__1736 (
            .O(N__18866),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.QiZ0Z_0 ));
    InMux I__1735 (
            .O(N__18859),
            .I(N__18828));
    InMux I__1734 (
            .O(N__18858),
            .I(N__18828));
    InMux I__1733 (
            .O(N__18857),
            .I(N__18828));
    InMux I__1732 (
            .O(N__18856),
            .I(N__18828));
    InMux I__1731 (
            .O(N__18855),
            .I(N__18828));
    InMux I__1730 (
            .O(N__18854),
            .I(N__18828));
    InMux I__1729 (
            .O(N__18853),
            .I(N__18828));
    InMux I__1728 (
            .O(N__18852),
            .I(N__18828));
    InMux I__1727 (
            .O(N__18851),
            .I(N__18819));
    InMux I__1726 (
            .O(N__18850),
            .I(N__18819));
    InMux I__1725 (
            .O(N__18849),
            .I(N__18819));
    InMux I__1724 (
            .O(N__18848),
            .I(N__18819));
    InMux I__1723 (
            .O(N__18847),
            .I(N__18812));
    InMux I__1722 (
            .O(N__18846),
            .I(N__18812));
    InMux I__1721 (
            .O(N__18845),
            .I(N__18812));
    LocalMux I__1720 (
            .O(N__18828),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.N_1545 ));
    LocalMux I__1719 (
            .O(N__18819),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.N_1545 ));
    LocalMux I__1718 (
            .O(N__18812),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.N_1545 ));
    InMux I__1717 (
            .O(N__18805),
            .I(N__18802));
    LocalMux I__1716 (
            .O(N__18802),
            .I(N__18799));
    Span4Mux_v I__1715 (
            .O(N__18799),
            .I(N__18796));
    Odrv4 I__1714 (
            .O(N__18796),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_s_5 ));
    InMux I__1713 (
            .O(N__18793),
            .I(N__18790));
    LocalMux I__1712 (
            .O(N__18790),
            .I(N__18787));
    Span4Mux_s2_h I__1711 (
            .O(N__18787),
            .I(N__18783));
    InMux I__1710 (
            .O(N__18786),
            .I(N__18780));
    Odrv4 I__1709 (
            .O(N__18783),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.QiZ0Z_5 ));
    LocalMux I__1708 (
            .O(N__18780),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.QiZ0Z_5 ));
    CEMux I__1707 (
            .O(N__18775),
            .I(N__18772));
    LocalMux I__1706 (
            .O(N__18772),
            .I(N__18768));
    CEMux I__1705 (
            .O(N__18771),
            .I(N__18765));
    Span4Mux_h I__1704 (
            .O(N__18768),
            .I(N__18762));
    LocalMux I__1703 (
            .O(N__18765),
            .I(N__18759));
    Span4Mux_s0_h I__1702 (
            .O(N__18762),
            .I(N__18756));
    Odrv4 I__1701 (
            .O(N__18759),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.N_290 ));
    Odrv4 I__1700 (
            .O(N__18756),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.N_290 ));
    InMux I__1699 (
            .O(N__18751),
            .I(N__18748));
    LocalMux I__1698 (
            .O(N__18748),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_1_sqmuxa_i_x0_0 ));
    InMux I__1697 (
            .O(N__18745),
            .I(N__18742));
    LocalMux I__1696 (
            .O(N__18742),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_s_6 ));
    InMux I__1695 (
            .O(N__18739),
            .I(N__18736));
    LocalMux I__1694 (
            .O(N__18736),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_s_7 ));
    CascadeMux I__1693 (
            .O(N__18733),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.val_c8_cascade_ ));
    CascadeMux I__1692 (
            .O(N__18730),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.N_1545_cascade_ ));
    InMux I__1691 (
            .O(N__18727),
            .I(N__18724));
    LocalMux I__1690 (
            .O(N__18724),
            .I(N__18721));
    Odrv4 I__1689 (
            .O(N__18721),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_s_1 ));
    InMux I__1688 (
            .O(N__18718),
            .I(N__18715));
    LocalMux I__1687 (
            .O(N__18715),
            .I(N__18712));
    Span4Mux_h I__1686 (
            .O(N__18712),
            .I(N__18709));
    Odrv4 I__1685 (
            .O(N__18709),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_s_6 ));
    InMux I__1684 (
            .O(N__18706),
            .I(N__18703));
    LocalMux I__1683 (
            .O(N__18703),
            .I(N__18700));
    Odrv12 I__1682 (
            .O(N__18700),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_s_7 ));
    InMux I__1681 (
            .O(N__18697),
            .I(N__18694));
    LocalMux I__1680 (
            .O(N__18694),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.val_c8_0_3 ));
    InMux I__1679 (
            .O(N__18691),
            .I(N__18688));
    LocalMux I__1678 (
            .O(N__18688),
            .I(N__18685));
    Odrv4 I__1677 (
            .O(N__18685),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_s_3 ));
    InMux I__1676 (
            .O(N__18682),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_cry_6 ));
    InMux I__1675 (
            .O(N__18679),
            .I(N__18676));
    LocalMux I__1674 (
            .O(N__18676),
            .I(N__18672));
    InMux I__1673 (
            .O(N__18675),
            .I(N__18669));
    Span4Mux_h I__1672 (
            .O(N__18672),
            .I(N__18664));
    LocalMux I__1671 (
            .O(N__18669),
            .I(N__18664));
    Span4Mux_v I__1670 (
            .O(N__18664),
            .I(N__18661));
    Odrv4 I__1669 (
            .O(N__18661),
            .I(wb_cyc_i_c));
    CascadeMux I__1668 (
            .O(N__18658),
            .I(N__18654));
    InMux I__1667 (
            .O(N__18657),
            .I(N__18651));
    InMux I__1666 (
            .O(N__18654),
            .I(N__18648));
    LocalMux I__1665 (
            .O(N__18651),
            .I(N__18645));
    LocalMux I__1664 (
            .O(N__18648),
            .I(N__18642));
    Span4Mux_v I__1663 (
            .O(N__18645),
            .I(N__18639));
    Span4Mux_v I__1662 (
            .O(N__18642),
            .I(N__18636));
    Odrv4 I__1661 (
            .O(N__18639),
            .I(wb_stb_i_c));
    Odrv4 I__1660 (
            .O(N__18636),
            .I(wb_stb_i_c));
    InMux I__1659 (
            .O(N__18631),
            .I(N__18628));
    LocalMux I__1658 (
            .O(N__18628),
            .I(N__18625));
    Odrv4 I__1657 (
            .O(N__18625),
            .I(\u1.cINTRQ ));
    InMux I__1656 (
            .O(N__18622),
            .I(N__18619));
    LocalMux I__1655 (
            .O(N__18619),
            .I(N__18616));
    Span4Mux_h I__1654 (
            .O(N__18616),
            .I(N__18613));
    Odrv4 I__1653 (
            .O(N__18613),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_s_0 ));
    InMux I__1652 (
            .O(N__18610),
            .I(N__18607));
    LocalMux I__1651 (
            .O(N__18607),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_s_1 ));
    InMux I__1650 (
            .O(N__18604),
            .I(N__18601));
    LocalMux I__1649 (
            .O(N__18601),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_s_2 ));
    InMux I__1648 (
            .O(N__18598),
            .I(N__18595));
    LocalMux I__1647 (
            .O(N__18595),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_s_3 ));
    InMux I__1646 (
            .O(N__18592),
            .I(N__18589));
    LocalMux I__1645 (
            .O(N__18589),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_s_4 ));
    InMux I__1644 (
            .O(N__18586),
            .I(N__18583));
    LocalMux I__1643 (
            .O(N__18583),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_s_5 ));
    InMux I__1642 (
            .O(N__18580),
            .I(N__18577));
    LocalMux I__1641 (
            .O(N__18577),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_s_1 ));
    InMux I__1640 (
            .O(N__18574),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_cry_0 ));
    InMux I__1639 (
            .O(N__18571),
            .I(N__18568));
    LocalMux I__1638 (
            .O(N__18568),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_s_2 ));
    InMux I__1637 (
            .O(N__18565),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_cry_1 ));
    InMux I__1636 (
            .O(N__18562),
            .I(N__18559));
    LocalMux I__1635 (
            .O(N__18559),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_s_3 ));
    InMux I__1634 (
            .O(N__18556),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_cry_2 ));
    InMux I__1633 (
            .O(N__18553),
            .I(N__18550));
    LocalMux I__1632 (
            .O(N__18550),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_s_4 ));
    InMux I__1631 (
            .O(N__18547),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_cry_3 ));
    InMux I__1630 (
            .O(N__18544),
            .I(N__18541));
    LocalMux I__1629 (
            .O(N__18541),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_s_5 ));
    InMux I__1628 (
            .O(N__18538),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_cry_4 ));
    InMux I__1627 (
            .O(N__18535),
            .I(N__18532));
    LocalMux I__1626 (
            .O(N__18532),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_s_6 ));
    InMux I__1625 (
            .O(N__18529),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_cry_5 ));
    CascadeMux I__1624 (
            .O(N__18526),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.N_2413_iZ0_cascade_ ));
    InMux I__1623 (
            .O(N__18523),
            .I(N__18520));
    LocalMux I__1622 (
            .O(N__18520),
            .I(N__18517));
    Span4Mux_v I__1621 (
            .O(N__18517),
            .I(N__18514));
    Odrv4 I__1620 (
            .O(N__18514),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_s_0 ));
    InMux I__1619 (
            .O(N__18511),
            .I(N__18508));
    LocalMux I__1618 (
            .O(N__18508),
            .I(\u1.DMA_control.Tm_2 ));
    InMux I__1617 (
            .O(N__18505),
            .I(N__18501));
    InMux I__1616 (
            .O(N__18504),
            .I(N__18498));
    LocalMux I__1615 (
            .O(N__18501),
            .I(N__18493));
    LocalMux I__1614 (
            .O(N__18498),
            .I(N__18493));
    Odrv4 I__1613 (
            .O(N__18493),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.QiZ0Z_2 ));
    InMux I__1612 (
            .O(N__18490),
            .I(N__18487));
    LocalMux I__1611 (
            .O(N__18487),
            .I(N__18484));
    Odrv4 I__1610 (
            .O(N__18484),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_s_2 ));
    InMux I__1609 (
            .O(N__18481),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_cry_1 ));
    InMux I__1608 (
            .O(N__18478),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_cry_2 ));
    InMux I__1607 (
            .O(N__18475),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_cry_3 ));
    InMux I__1606 (
            .O(N__18472),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_cry_4 ));
    InMux I__1605 (
            .O(N__18469),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_cry_5 ));
    InMux I__1604 (
            .O(N__18466),
            .I(N__18462));
    InMux I__1603 (
            .O(N__18465),
            .I(N__18459));
    LocalMux I__1602 (
            .O(N__18462),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.QiZ0Z_7 ));
    LocalMux I__1601 (
            .O(N__18459),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.QiZ0Z_7 ));
    InMux I__1600 (
            .O(N__18454),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_cry_6 ));
    InMux I__1599 (
            .O(N__18451),
            .I(N__18448));
    LocalMux I__1598 (
            .O(N__18448),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_s_7 ));
    InMux I__1597 (
            .O(N__18445),
            .I(N__18442));
    LocalMux I__1596 (
            .O(N__18442),
            .I(N__18439));
    Odrv4 I__1595 (
            .O(N__18439),
            .I(\u1.DMA_control.Teoc_0 ));
    InMux I__1594 (
            .O(N__18436),
            .I(N__18433));
    LocalMux I__1593 (
            .O(N__18433),
            .I(N__18430));
    Odrv12 I__1592 (
            .O(N__18430),
            .I(\u1.DMA_control.Teoc_2 ));
    CascadeMux I__1591 (
            .O(N__18427),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.val_c7_0_3_cascade_ ));
    CascadeMux I__1590 (
            .O(N__18424),
            .I(\u1.Tdone_i_cascade_ ));
    InMux I__1589 (
            .O(N__18421),
            .I(N__18418));
    LocalMux I__1588 (
            .O(N__18418),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNIDE5P1Z0Z_0 ));
    CascadeMux I__1587 (
            .O(N__18415),
            .I(N__18410));
    InMux I__1586 (
            .O(N__18414),
            .I(N__18407));
    InMux I__1585 (
            .O(N__18413),
            .I(N__18402));
    InMux I__1584 (
            .O(N__18410),
            .I(N__18402));
    LocalMux I__1583 (
            .O(N__18407),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.rciZ0 ));
    LocalMux I__1582 (
            .O(N__18402),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.rciZ0 ));
    InMux I__1581 (
            .O(N__18397),
            .I(N__18394));
    LocalMux I__1580 (
            .O(N__18394),
            .I(\u1.DMA_control.dTfw ));
    InMux I__1579 (
            .O(N__18391),
            .I(N__18386));
    InMux I__1578 (
            .O(N__18390),
            .I(N__18383));
    InMux I__1577 (
            .O(N__18389),
            .I(N__18380));
    LocalMux I__1576 (
            .O(N__18386),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.QiZ0Z_0 ));
    LocalMux I__1575 (
            .O(N__18383),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.QiZ0Z_0 ));
    LocalMux I__1574 (
            .O(N__18380),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.QiZ0Z_0 ));
    InMux I__1573 (
            .O(N__18373),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_cry_0 ));
    InMux I__1572 (
            .O(N__18370),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_cry_3 ));
    InMux I__1571 (
            .O(N__18367),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_cry_4 ));
    InMux I__1570 (
            .O(N__18364),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_cry_5 ));
    InMux I__1569 (
            .O(N__18361),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_cry_6 ));
    InMux I__1568 (
            .O(N__18358),
            .I(N__18355));
    LocalMux I__1567 (
            .O(N__18355),
            .I(\u1.DMA_control.Teoc_7 ));
    InMux I__1566 (
            .O(N__18352),
            .I(N__18349));
    LocalMux I__1565 (
            .O(N__18349),
            .I(N__18346));
    Span4Mux_v I__1564 (
            .O(N__18346),
            .I(N__18343));
    Odrv4 I__1563 (
            .O(N__18343),
            .I(intrq_pad_i_c));
    InMux I__1562 (
            .O(N__18340),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_cry_0 ));
    InMux I__1561 (
            .O(N__18337),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_cry_1 ));
    InMux I__1560 (
            .O(N__18334),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_cry_2 ));
    InMux I__1559 (
            .O(N__18331),
            .I(N__18328));
    LocalMux I__1558 (
            .O(N__18328),
            .I(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_s_0 ));
    InMux I__1557 (
            .O(N__18325),
            .I(N__18322));
    LocalMux I__1556 (
            .O(N__18322),
            .I(N__18319));
    Span12Mux_v I__1555 (
            .O(N__18319),
            .I(N__18316));
    Odrv12 I__1554 (
            .O(N__18316),
            .I(\u1.cDMARQ ));
    InMux I__1553 (
            .O(N__18313),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_cry_4 ));
    InMux I__1552 (
            .O(N__18310),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_cry_5 ));
    InMux I__1551 (
            .O(N__18307),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_cry_6 ));
    CascadeMux I__1550 (
            .O(N__18304),
            .I(CONSTANT_ONE_NET_cascade_));
    InMux I__1549 (
            .O(N__18301),
            .I(N__18298));
    LocalMux I__1548 (
            .O(N__18298),
            .I(N__18295));
    Span4Mux_v I__1547 (
            .O(N__18295),
            .I(N__18292));
    Odrv4 I__1546 (
            .O(N__18292),
            .I(arst_i_c));
    IoInMux I__1545 (
            .O(N__18289),
            .I(N__18286));
    LocalMux I__1544 (
            .O(N__18286),
            .I(N__18283));
    IoSpan4Mux I__1543 (
            .O(N__18283),
            .I(N__18280));
    IoSpan4Mux I__1542 (
            .O(N__18280),
            .I(N__18277));
    IoSpan4Mux I__1541 (
            .O(N__18277),
            .I(N__18274));
    Odrv4 I__1540 (
            .O(N__18274),
            .I(arst_i_c_i));
    InMux I__1539 (
            .O(N__18271),
            .I(N__18268));
    LocalMux I__1538 (
            .O(N__18268),
            .I(N__18265));
    Span4Mux_v I__1537 (
            .O(N__18265),
            .I(N__18262));
    Span4Mux_v I__1536 (
            .O(N__18262),
            .I(N__18259));
    Odrv4 I__1535 (
            .O(N__18259),
            .I(dmarq_pad_i_c));
    InMux I__1534 (
            .O(N__18256),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_cry_0 ));
    InMux I__1533 (
            .O(N__18253),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_cry_1 ));
    InMux I__1532 (
            .O(N__18250),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_cry_2 ));
    InMux I__1531 (
            .O(N__18247),
            .I(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_cry_3 ));
    defparam IN_MUX_bfv_12_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_18_0_));
    defparam IN_MUX_bfv_7_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_17_0_));
    defparam IN_MUX_bfv_2_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_17_0_));
    defparam IN_MUX_bfv_1_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_18_0_));
    defparam IN_MUX_bfv_2_24_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_24_0_));
    defparam IN_MUX_bfv_4_20_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_20_0_));
    defparam IN_MUX_bfv_2_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_21_0_));
    ICE_GB \u1.DMA_control.gen_DMAbuf_Txbuf.valid_RNI2KL74_0  (
            .USERSIGNALTOGLOBALBUFFER(N__24073),
            .GLOBALBUFFEROUTPUT(\u1.DMA_control.gen_DMAbuf_Txbuf.N_319_g ));
    ICE_GB \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.dstrb_RNIBHHI_0  (
            .USERSIGNALTOGLOBALBUFFER(N__19045),
            .GLOBALBUFFEROUTPUT(\u1.DMA_control.rd_dstrb_g ));
    ICE_GB arst_i_ibuf_RNI7B6A_0 (
            .USERSIGNALTOGLOBALBUFFER(N__18289),
            .GLOBALBUFFEROUTPUT(arst_i_c_i_g));
    VCC VCC (
            .Y(VCCG0));
    ICE_GB N_77_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__50593),
            .GLOBALBUFFEROUTPUT(N_77_g));
    ICE_GB N_448_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__43798),
            .GLOBALBUFFEROUTPUT(N_448_g));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam arst_i_ibuf_RNI7B6A_LC_1_7_5.C_ON=1'b0;
    defparam arst_i_ibuf_RNI7B6A_LC_1_7_5.SEQ_MODE=4'b0000;
    defparam arst_i_ibuf_RNI7B6A_LC_1_7_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 arst_i_ibuf_RNI7B6A_LC_1_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18301),
            .lcout(arst_i_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.synch_incoming_cDMARQ_LC_1_13_4 .C_ON=1'b0;
    defparam \u1.synch_incoming_cDMARQ_LC_1_13_4 .SEQ_MODE=4'b1000;
    defparam \u1.synch_incoming_cDMARQ_LC_1_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.synch_incoming_cDMARQ_LC_1_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18271),
            .lcout(\u1.cDMARQ ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54118),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_cry_c_0_LC_1_18_0 .C_ON=1'b1;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_cry_c_0_LC_1_18_0 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_cry_c_0_LC_1_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_cry_c_0_LC_1_18_0  (
            .in0(_gnd_net_),
            .in1(N__18888),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_18_0_),
            .carryout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNO_0_1_LC_1_18_1 .C_ON=1'b1;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNO_0_1_LC_1_18_1 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNO_0_1_LC_1_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNO_0_1_LC_1_18_1  (
            .in0(_gnd_net_),
            .in1(N__19009),
            .in2(N__28575),
            .in3(N__18256),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_s_1 ),
            .ltout(),
            .carryin(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_cry_0 ),
            .carryout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNO_0_2_LC_1_18_2 .C_ON=1'b1;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNO_0_2_LC_1_18_2 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNO_0_2_LC_1_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNO_0_2_LC_1_18_2  (
            .in0(_gnd_net_),
            .in1(N__18955),
            .in2(N__28577),
            .in3(N__18253),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_s_2 ),
            .ltout(),
            .carryin(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_cry_1 ),
            .carryout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNO_0_3_LC_1_18_3 .C_ON=1'b1;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNO_0_3_LC_1_18_3 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNO_0_3_LC_1_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNO_0_3_LC_1_18_3  (
            .in0(_gnd_net_),
            .in1(N__28500),
            .in2(N__19027),
            .in3(N__18250),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_s_3 ),
            .ltout(),
            .carryin(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_cry_2 ),
            .carryout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNO_0_4_LC_1_18_4 .C_ON=1'b1;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNO_0_4_LC_1_18_4 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNO_0_4_LC_1_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNO_0_4_LC_1_18_4  (
            .in0(_gnd_net_),
            .in1(N__18922),
            .in2(N__28578),
            .in3(N__18247),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_s_4 ),
            .ltout(),
            .carryin(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_cry_3 ),
            .carryout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNO_0_5_LC_1_18_5 .C_ON=1'b1;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNO_0_5_LC_1_18_5 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNO_0_5_LC_1_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNO_0_5_LC_1_18_5  (
            .in0(_gnd_net_),
            .in1(N__18793),
            .in2(N__28576),
            .in3(N__18313),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_s_5 ),
            .ltout(),
            .carryin(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_cry_4 ),
            .carryout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNO_0_6_LC_1_18_6 .C_ON=1'b1;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNO_0_6_LC_1_18_6 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNO_0_6_LC_1_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNO_0_6_LC_1_18_6  (
            .in0(_gnd_net_),
            .in1(N__18991),
            .in2(N__28579),
            .in3(N__18310),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_s_6 ),
            .ltout(),
            .carryin(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_cry_5 ),
            .carryout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNO_0_7_LC_1_18_7 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNO_0_7_LC_1_18_7 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNO_0_7_LC_1_18_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNO_0_7_LC_1_18_7  (
            .in0(_gnd_net_),
            .in1(N__20873),
            .in2(_gnd_net_),
            .in3(N__18307),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_s_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_pong_d_9_LC_1_19_0 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_pong_d_9_LC_1_19_0 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_pong_d_9_LC_1_19_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.PIO_control.gen_pingpong_pong_d_9_LC_1_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36019),
            .lcout(\u1.PIO_control.pong_d_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54111),
            .ce(N__24884),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_pong_we_LC_1_19_1 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_pong_we_LC_1_19_1 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_pong_we_LC_1_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.PIO_control.gen_pingpong_pong_we_LC_1_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21940),
            .lcout(\u1.PIO_control.pong_we ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54111),
            .ce(N__24884),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNO_0_0_LC_1_20_1 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNO_0_0_LC_1_20_1 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNO_0_0_LC_1_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNO_0_0_LC_1_20_1  (
            .in0(_gnd_net_),
            .in1(N__28423),
            .in2(_gnd_net_),
            .in3(N__19444),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_s_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_7_LC_1_20_2 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_7_LC_1_20_2 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_7_LC_1_20_2 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_7_LC_1_20_2  (
            .in0(N__19133),
            .in1(N__18358),
            .in2(N__52242),
            .in3(N__18451),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.QiZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54114),
            .ce(N__19070),
            .sr(N__53308));
    defparam CONSTANT_ONE_LUT4_LC_1_20_3.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_1_20_3.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_1_20_3.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_1_20_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(CONSTANT_ONE_NET_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNO_0_0_LC_1_20_4 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNO_0_0_LC_1_20_4 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNO_0_0_LC_1_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNO_0_0_LC_1_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18304),
            .in3(N__19864),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_s_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_0_LC_1_20_5 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_0_LC_1_20_5 .SEQ_MODE=4'b1011;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_0_LC_1_20_5 .LUT_INIT=16'b1111101011001100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_0_LC_1_20_5  (
            .in0(N__18445),
            .in1(N__18331),
            .in2(N__52241),
            .in3(N__19132),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.QiZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54114),
            .ce(N__19070),
            .sr(N__53308));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNO_0_0_LC_1_20_6 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNO_0_0_LC_1_20_6 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNO_0_0_LC_1_20_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNO_0_0_LC_1_20_6  (
            .in0(N__28424),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18892),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_s_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_RNO_0_0_LC_1_20_7 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_RNO_0_0_LC_1_20_7 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_RNO_0_0_LC_1_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_RNO_0_0_LC_1_20_7  (
            .in0(_gnd_net_),
            .in1(N__28425),
            .in2(_gnd_net_),
            .in3(N__20361),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_s_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNO_0_0_LC_1_21_4 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNO_0_0_LC_1_21_4 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNO_0_0_LC_1_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNO_0_0_LC_1_21_4  (
            .in0(_gnd_net_),
            .in1(N__28426),
            .in2(_gnd_net_),
            .in3(N__18391),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_s_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.sDMARQ_LC_1_21_5 .C_ON=1'b0;
    defparam \u1.sDMARQ_LC_1_21_5 .SEQ_MODE=4'b1000;
    defparam \u1.sDMARQ_LC_1_21_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.sDMARQ_LC_1_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18325),
            .lcout(DMA_dmarq),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54119),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev0_Tm_0_LC_1_22_0 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Tm_0_LC_1_22_0 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev0_Tm_0_LC_1_22_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.DMA_dev0_Tm_0_LC_1_22_0  (
            .in0(N__49549),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51849),
            .lcout(DMA_dev0_Tm_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54125),
            .ce(N__39723),
            .sr(N__53316));
    defparam \u0.DMA_dev0_Td_7_LC_1_22_2 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Td_7_LC_1_22_2 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev0_Td_7_LC_1_22_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.DMA_dev0_Td_7_LC_1_22_2  (
            .in0(N__34568),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51841),
            .lcout(DMA_dev0_Td_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54125),
            .ce(N__39723),
            .sr(N__53316));
    defparam \u0.DMA_dev0_Teoc_7_LC_1_22_3 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Teoc_7_LC_1_22_3 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev0_Teoc_7_LC_1_22_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.DMA_dev0_Teoc_7_LC_1_22_3  (
            .in0(N__51848),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40487),
            .lcout(DMA_dev0_Teoc_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54125),
            .ce(N__39723),
            .sr(N__53316));
    defparam \u0.DMA_dev0_Teoc_0_LC_1_22_4 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Teoc_0_LC_1_22_4 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev0_Teoc_0_LC_1_22_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \u0.DMA_dev0_Teoc_0_LC_1_22_4  (
            .in0(_gnd_net_),
            .in1(N__39878),
            .in2(_gnd_net_),
            .in3(N__51842),
            .lcout(DMA_dev0_Teoc_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54125),
            .ce(N__39723),
            .sr(N__53316));
    defparam \u0.DMA_dev0_Teoc_1_LC_1_22_5 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Teoc_1_LC_1_22_5 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev0_Teoc_1_LC_1_22_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.DMA_dev0_Teoc_1_LC_1_22_5  (
            .in0(N__51843),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40812),
            .lcout(DMA_dev0_Teoc_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54125),
            .ce(N__39723),
            .sr(N__53316));
    defparam \u0.DMA_dev0_Teoc_2_LC_1_22_6 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Teoc_2_LC_1_22_6 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev0_Teoc_2_LC_1_22_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.DMA_dev0_Teoc_2_LC_1_22_6  (
            .in0(N__44205),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51844),
            .lcout(DMA_dev0_Teoc_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54125),
            .ce(N__39723),
            .sr(N__53316));
    defparam \u0.DMA_dev0_Teoc_6_LC_1_22_7 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Teoc_6_LC_1_22_7 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev0_Teoc_6_LC_1_22_7 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \u0.DMA_dev0_Teoc_6_LC_1_22_7  (
            .in0(N__47794),
            .in1(_gnd_net_),
            .in2(N__52051),
            .in3(_gnd_net_),
            .lcout(DMA_dev0_Teoc_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54125),
            .ce(N__39723),
            .sr(N__53316));
    defparam \u1.PIO_control.PIO_access_control.q_12_LC_1_23_1 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.q_12_LC_1_23_1 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.q_12_LC_1_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.PIO_control.PIO_access_control.q_12_LC_1_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25221),
            .lcout(PIOq_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54130),
            .ce(N__45926),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.q_14_LC_1_23_2 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.q_14_LC_1_23_2 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.q_14_LC_1_23_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.PIO_control.PIO_access_control.q_14_LC_1_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32850),
            .lcout(PIOq_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54130),
            .ce(N__45926),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_pong_d_2_LC_1_27_4 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_pong_d_2_LC_1_27_4 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_pong_d_2_LC_1_27_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.PIO_control.gen_pingpong_pong_d_2_LC_1_27_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34264),
            .lcout(\u1.PIO_control.pong_d_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54162),
            .ce(N__24894),
            .sr(_gnd_net_));
    defparam \u0.ack_o_i_i_o2_LC_2_7_4 .C_ON=1'b0;
    defparam \u0.ack_o_i_i_o2_LC_2_7_4 .SEQ_MODE=4'b0000;
    defparam \u0.ack_o_i_i_o2_LC_2_7_4 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \u0.ack_o_i_i_o2_LC_2_7_4  (
            .in0(N__22818),
            .in1(N__18675),
            .in2(N__18658),
            .in3(N__22770),
            .lcout(N_1342),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.synch_incoming_cINTRQ_LC_2_11_6 .C_ON=1'b0;
    defparam \u1.synch_incoming_cINTRQ_LC_2_11_6 .SEQ_MODE=4'b1000;
    defparam \u1.synch_incoming_cINTRQ_LC_2_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.synch_incoming_cINTRQ_LC_2_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18352),
            .lcout(\u1.cINTRQ ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54137),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_cry_c_0_LC_2_17_0 .C_ON=1'b1;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_cry_c_0_LC_2_17_0 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_cry_c_0_LC_2_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_cry_c_0_LC_2_17_0  (
            .in0(_gnd_net_),
            .in1(N__20347),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_17_0_),
            .carryout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_RNO_0_1_LC_2_17_1 .C_ON=1'b1;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_RNO_0_1_LC_2_17_1 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_RNO_0_1_LC_2_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_RNO_0_1_LC_2_17_1  (
            .in0(_gnd_net_),
            .in1(N__20402),
            .in2(N__28647),
            .in3(N__18340),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_s_1 ),
            .ltout(),
            .carryin(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_cry_0 ),
            .carryout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_RNO_0_2_LC_2_17_2 .C_ON=1'b1;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_RNO_0_2_LC_2_17_2 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_RNO_0_2_LC_2_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_RNO_0_2_LC_2_17_2  (
            .in0(_gnd_net_),
            .in1(N__20477),
            .in2(N__28650),
            .in3(N__18337),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_s_2 ),
            .ltout(),
            .carryin(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_cry_1 ),
            .carryout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_RNO_0_3_LC_2_17_3 .C_ON=1'b1;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_RNO_0_3_LC_2_17_3 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_RNO_0_3_LC_2_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_RNO_0_3_LC_2_17_3  (
            .in0(_gnd_net_),
            .in1(N__20429),
            .in2(N__28648),
            .in3(N__18334),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_s_3 ),
            .ltout(),
            .carryin(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_cry_2 ),
            .carryout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_RNO_0_4_LC_2_17_4 .C_ON=1'b1;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_RNO_0_4_LC_2_17_4 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_RNO_0_4_LC_2_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_RNO_0_4_LC_2_17_4  (
            .in0(_gnd_net_),
            .in1(N__20453),
            .in2(N__28651),
            .in3(N__18370),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_s_4 ),
            .ltout(),
            .carryin(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_cry_3 ),
            .carryout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_RNO_0_5_LC_2_17_5 .C_ON=1'b1;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_RNO_0_5_LC_2_17_5 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_RNO_0_5_LC_2_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_RNO_0_5_LC_2_17_5  (
            .in0(_gnd_net_),
            .in1(N__20529),
            .in2(N__28649),
            .in3(N__18367),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_s_5 ),
            .ltout(),
            .carryin(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_cry_4 ),
            .carryout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_RNO_0_6_LC_2_17_6 .C_ON=1'b1;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_RNO_0_6_LC_2_17_6 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_RNO_0_6_LC_2_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_RNO_0_6_LC_2_17_6  (
            .in0(_gnd_net_),
            .in1(N__20558),
            .in2(N__28652),
            .in3(N__18364),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_s_6 ),
            .ltout(),
            .carryin(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_cry_5 ),
            .carryout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_RNO_0_7_LC_2_17_7 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_RNO_0_7_LC_2_17_7 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_RNO_0_7_LC_2_17_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_RNO_0_7_LC_2_17_7  (
            .in0(_gnd_net_),
            .in1(N__20505),
            .in2(_gnd_net_),
            .in3(N__18361),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_s_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_2_LC_2_18_4 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_2_LC_2_18_4 .SEQ_MODE=4'b1011;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_2_LC_2_18_4 .LUT_INIT=16'b1111101011001100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_2_LC_2_18_4  (
            .in0(N__18436),
            .in1(N__18490),
            .in2(N__52769),
            .in3(N__19131),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.QiZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54112),
            .ce(N__19072),
            .sr(N__53305));
    defparam \u1.c_state_RNIV4MT_0_LC_2_19_2 .C_ON=1'b0;
    defparam \u1.c_state_RNIV4MT_0_LC_2_19_2 .SEQ_MODE=4'b0000;
    defparam \u1.c_state_RNIV4MT_0_LC_2_19_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \u1.c_state_RNIV4MT_0_LC_2_19_2  (
            .in0(_gnd_net_),
            .in1(N__24447),
            .in2(_gnd_net_),
            .in3(N__24406),
            .lcout(\u1.N_1382 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_1_sqmuxa_i_ns_LC_2_19_3 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_1_sqmuxa_i_ns_LC_2_19_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_1_sqmuxa_i_ns_LC_2_19_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_1_sqmuxa_i_ns_LC_2_19_3  (
            .in0(N__52601),
            .in1(N__19741),
            .in2(_gnd_net_),
            .in3(N__18751),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_1_sqmuxa_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_Teoc_7_LC_2_19_4 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_Teoc_7_LC_2_19_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.DMA_timing_ctrl_Teoc_7_LC_2_19_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_Teoc_7_LC_2_19_4  (
            .in0(N__40408),
            .in1(N__40434),
            .in2(_gnd_net_),
            .in3(N__36290),
            .lcout(\u1.DMA_control.Teoc_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54115),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNIHI1O1_2_LC_2_20_0 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNIHI1O1_2_LC_2_20_0 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNIHI1O1_2_LC_2_20_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNIHI1O1_2_LC_2_20_0  (
            .in0(N__19149),
            .in1(N__19179),
            .in2(N__19087),
            .in3(N__18505),
            .lcout(),
            .ltout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.val_c7_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNIDG7V3_7_LC_2_20_1 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNIDG7V3_7_LC_2_20_1 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNIDG7V3_7_LC_2_20_1 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNIDG7V3_7_LC_2_20_1  (
            .in0(_gnd_net_),
            .in1(N__18466),
            .in2(N__18427),
            .in3(N__18421),
            .lcout(\u1.Tdone_i ),
            .ltout(\u1.Tdone_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.Tfw_LC_2_20_2 .C_ON=1'b0;
    defparam \u1.DMA_control.Tfw_LC_2_20_2 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.Tfw_LC_2_20_2 .LUT_INIT=16'b0011001100100000;
    LogicCell40 \u1.DMA_control.Tfw_LC_2_20_2  (
            .in0(N__20251),
            .in1(N__51565),
            .in2(N__18424),
            .in3(N__21022),
            .lcout(\u1.Tfw ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54120),
            .ce(),
            .sr(N__53312));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.rci_LC_2_20_3 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.rci_LC_2_20_3 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.rci_LC_2_20_3 .LUT_INIT=16'b0000100000001111;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.rci_LC_2_20_3  (
            .in0(N__18414),
            .in1(N__21548),
            .in2(N__51839),
            .in3(N__20022),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.rciZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54120),
            .ce(),
            .sr(N__53312));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNIDE5P1_0_LC_2_20_4 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNIDE5P1_0_LC_2_20_4 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNIDE5P1_0_LC_2_20_4 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNIDE5P1_0_LC_2_20_4  (
            .in0(N__19216),
            .in1(N__19237),
            .in2(N__18415),
            .in3(N__18390),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNIDE5P1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qie_0_i_LC_2_20_5 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qie_0_i_LC_2_20_5 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qie_0_i_LC_2_20_5 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qie_0_i_LC_2_20_5  (
            .in0(N__51560),
            .in1(N__18413),
            .in2(_gnd_net_),
            .in3(N__20021),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qie_0_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_igo_LC_2_20_6 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_igo_LC_2_20_6 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.DMA_timing_ctrl_igo_LC_2_20_6 .LUT_INIT=16'b0000111100000100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_igo_LC_2_20_6  (
            .in0(N__20250),
            .in1(N__18397),
            .in2(N__51840),
            .in3(N__21021),
            .lcout(\u1.DMA_control.igo ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54120),
            .ce(),
            .sr(N__53312));
    defparam \u1.DMA_control.DMA_timing_ctrl_dTfw_LC_2_20_7 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_dTfw_LC_2_20_7 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.DMA_timing_ctrl_dTfw_LC_2_20_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_dTfw_LC_2_20_7  (
            .in0(N__51564),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20249),
            .lcout(\u1.DMA_control.dTfw ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54120),
            .ce(),
            .sr(N__53312));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_cry_c_0_LC_2_21_0 .C_ON=1'b1;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_cry_c_0_LC_2_21_0 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_cry_c_0_LC_2_21_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_cry_c_0_LC_2_21_0  (
            .in0(_gnd_net_),
            .in1(N__18389),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_21_0_),
            .carryout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNO_0_1_LC_2_21_1 .C_ON=1'b1;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNO_0_1_LC_2_21_1 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNO_0_1_LC_2_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNO_0_1_LC_2_21_1  (
            .in0(_gnd_net_),
            .in1(N__19236),
            .in2(N__28507),
            .in3(N__18373),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_s_1 ),
            .ltout(),
            .carryin(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_cry_0 ),
            .carryout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNO_0_2_LC_2_21_2 .C_ON=1'b1;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNO_0_2_LC_2_21_2 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNO_0_2_LC_2_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNO_0_2_LC_2_21_2  (
            .in0(_gnd_net_),
            .in1(N__18504),
            .in2(N__28510),
            .in3(N__18481),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_s_2 ),
            .ltout(),
            .carryin(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_cry_1 ),
            .carryout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNO_0_3_LC_2_21_3 .C_ON=1'b1;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNO_0_3_LC_2_21_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNO_0_3_LC_2_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNO_0_3_LC_2_21_3  (
            .in0(_gnd_net_),
            .in1(N__19212),
            .in2(N__28508),
            .in3(N__18478),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_s_3 ),
            .ltout(),
            .carryin(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_cry_2 ),
            .carryout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNO_0_4_LC_2_21_4 .C_ON=1'b1;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNO_0_4_LC_2_21_4 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNO_0_4_LC_2_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNO_0_4_LC_2_21_4  (
            .in0(_gnd_net_),
            .in1(N__28447),
            .in2(N__19183),
            .in3(N__18475),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_s_4 ),
            .ltout(),
            .carryin(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_cry_3 ),
            .carryout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNO_0_5_LC_2_21_5 .C_ON=1'b1;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNO_0_5_LC_2_21_5 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNO_0_5_LC_2_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNO_0_5_LC_2_21_5  (
            .in0(_gnd_net_),
            .in1(N__19150),
            .in2(N__28509),
            .in3(N__18472),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_s_5 ),
            .ltout(),
            .carryin(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_cry_4 ),
            .carryout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNO_0_6_LC_2_21_6 .C_ON=1'b1;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNO_0_6_LC_2_21_6 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNO_0_6_LC_2_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNO_0_6_LC_2_21_6  (
            .in0(_gnd_net_),
            .in1(N__19086),
            .in2(N__28511),
            .in3(N__18469),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_s_6 ),
            .ltout(),
            .carryin(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_cry_5 ),
            .carryout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNO_0_7_LC_2_21_7 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNO_0_7_LC_2_21_7 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNO_0_7_LC_2_21_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_RNO_0_7_LC_2_21_7  (
            .in0(_gnd_net_),
            .in1(N__18465),
            .in2(_gnd_net_),
            .in3(N__18454),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_s_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_Teoc_0_LC_2_22_0 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_Teoc_0_LC_2_22_0 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.DMA_timing_ctrl_Teoc_0_LC_2_22_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_Teoc_0_LC_2_22_0  (
            .in0(N__54522),
            .in1(N__46638),
            .in2(_gnd_net_),
            .in3(N__36283),
            .lcout(\u1.DMA_control.Teoc_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54131),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_Teoc_1_LC_2_22_1 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_Teoc_1_LC_2_22_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.DMA_timing_ctrl_Teoc_1_LC_2_22_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_Teoc_1_LC_2_22_1  (
            .in0(N__36284),
            .in1(N__49158),
            .in2(_gnd_net_),
            .in3(N__40761),
            .lcout(\u1.DMA_control.Teoc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54131),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_Teoc_2_LC_2_22_2 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_Teoc_2_LC_2_22_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.DMA_timing_ctrl_Teoc_2_LC_2_22_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_Teoc_2_LC_2_22_2  (
            .in0(N__44337),
            .in1(N__44139),
            .in2(_gnd_net_),
            .in3(N__36285),
            .lcout(\u1.DMA_control.Teoc_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54131),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_Tm_2_LC_2_22_3 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_Tm_2_LC_2_22_3 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.DMA_timing_ctrl_Tm_2_LC_2_22_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_Tm_2_LC_2_22_3  (
            .in0(N__36289),
            .in1(N__31684),
            .in2(_gnd_net_),
            .in3(N__31210),
            .lcout(\u1.DMA_control.Tm_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54131),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_Teoc_4_LC_2_22_4 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_Teoc_4_LC_2_22_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.DMA_timing_ctrl_Teoc_4_LC_2_22_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_Teoc_4_LC_2_22_4  (
            .in0(N__36852),
            .in1(N__46702),
            .in2(_gnd_net_),
            .in3(N__36286),
            .lcout(\u1.DMA_control.Teoc_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54131),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_Teoc_5_LC_2_22_5 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_Teoc_5_LC_2_22_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.DMA_timing_ctrl_Teoc_5_LC_2_22_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_Teoc_5_LC_2_22_5  (
            .in0(N__36287),
            .in1(N__43888),
            .in2(_gnd_net_),
            .in3(N__43854),
            .lcout(\u1.DMA_control.Teoc_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54131),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_Teoc_6_LC_2_22_6 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_Teoc_6_LC_2_22_6 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.DMA_timing_ctrl_Teoc_6_LC_2_22_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_Teoc_6_LC_2_22_6  (
            .in0(N__47884),
            .in1(N__47919),
            .in2(_gnd_net_),
            .in3(N__36288),
            .lcout(\u1.DMA_control.Teoc_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54131),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_1_LC_2_23_0 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_1_LC_2_23_0 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_1_LC_2_23_0 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_1_LC_2_23_0  (
            .in0(N__24637),
            .in1(N__18580),
            .in2(N__51853),
            .in3(N__22216),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.QiZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54138),
            .ce(N__22158),
            .sr(N__53322));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.N_2413_i_LC_2_23_1 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.N_2413_i_LC_2_23_1 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.N_2413_i_LC_2_23_1 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.N_2413_i_LC_2_23_1  (
            .in0(N__51584),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20078),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.N_2413_iZ0 ),
            .ltout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.N_2413_iZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_0_LC_2_23_2 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_0_LC_2_23_2 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_0_LC_2_23_2 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_0_LC_2_23_2  (
            .in0(N__51594),
            .in1(N__21511),
            .in2(N__18526),
            .in3(N__18523),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.Qi_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54138),
            .ce(N__22158),
            .sr(N__53322));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_2_LC_2_23_3 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_2_LC_2_23_3 .SEQ_MODE=4'b1011;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_2_LC_2_23_3 .LUT_INIT=16'b1111110110101000;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_2_LC_2_23_3  (
            .in0(N__22217),
            .in1(N__18511),
            .in2(N__51850),
            .in3(N__18571),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.QiZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54138),
            .ce(N__22158),
            .sr(N__53322));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_3_LC_2_23_4 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_3_LC_2_23_4 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_3_LC_2_23_4 .LUT_INIT=16'b0011101100001000;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_3_LC_2_23_4  (
            .in0(N__31834),
            .in1(N__22218),
            .in2(N__51854),
            .in3(N__18562),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.QiZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54138),
            .ce(N__22158),
            .sr(N__53322));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_4_LC_2_23_5 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_4_LC_2_23_5 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_4_LC_2_23_5 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_4_LC_2_23_5  (
            .in0(N__22219),
            .in1(N__31822),
            .in2(N__51851),
            .in3(N__18553),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.QiZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54138),
            .ce(N__22158),
            .sr(N__53322));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_5_LC_2_23_6 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_5_LC_2_23_6 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_5_LC_2_23_6 .LUT_INIT=16'b0011101100001000;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_5_LC_2_23_6  (
            .in0(N__31810),
            .in1(N__22220),
            .in2(N__51855),
            .in3(N__18544),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.QiZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54138),
            .ce(N__22158),
            .sr(N__53322));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_6_LC_2_23_7 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_6_LC_2_23_7 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_6_LC_2_23_7 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_6_LC_2_23_7  (
            .in0(N__22221),
            .in1(N__31795),
            .in2(N__51852),
            .in3(N__18535),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.QiZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54138),
            .ce(N__22158),
            .sr(N__53322));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_cry_c_0_LC_2_24_0 .C_ON=1'b1;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_cry_c_0_LC_2_24_0 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_cry_c_0_LC_2_24_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_cry_c_0_LC_2_24_0  (
            .in0(_gnd_net_),
            .in1(N__19438),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_24_0_),
            .carryout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNO_0_1_LC_2_24_1 .C_ON=1'b1;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNO_0_1_LC_2_24_1 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNO_0_1_LC_2_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNO_0_1_LC_2_24_1  (
            .in0(_gnd_net_),
            .in1(N__19273),
            .in2(N__28682),
            .in3(N__18574),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_s_1 ),
            .ltout(),
            .carryin(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_cry_0 ),
            .carryout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNO_0_2_LC_2_24_2 .C_ON=1'b1;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNO_0_2_LC_2_24_2 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNO_0_2_LC_2_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNO_0_2_LC_2_24_2  (
            .in0(_gnd_net_),
            .in1(N__28633),
            .in2(N__19306),
            .in3(N__18565),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_s_2 ),
            .ltout(),
            .carryin(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_cry_1 ),
            .carryout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNO_0_3_LC_2_24_3 .C_ON=1'b1;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNO_0_3_LC_2_24_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNO_0_3_LC_2_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNO_0_3_LC_2_24_3  (
            .in0(_gnd_net_),
            .in1(N__19318),
            .in2(N__28683),
            .in3(N__18556),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_s_3 ),
            .ltout(),
            .carryin(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_cry_2 ),
            .carryout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNO_0_4_LC_2_24_4 .C_ON=1'b1;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNO_0_4_LC_2_24_4 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNO_0_4_LC_2_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNO_0_4_LC_2_24_4  (
            .in0(_gnd_net_),
            .in1(N__28637),
            .in2(N__19290),
            .in3(N__18547),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_s_4 ),
            .ltout(),
            .carryin(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_cry_3 ),
            .carryout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNO_0_5_LC_2_24_5 .C_ON=1'b1;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNO_0_5_LC_2_24_5 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNO_0_5_LC_2_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNO_0_5_LC_2_24_5  (
            .in0(_gnd_net_),
            .in1(N__19465),
            .in2(N__28684),
            .in3(N__18538),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_s_5 ),
            .ltout(),
            .carryin(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_cry_4 ),
            .carryout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNO_0_6_LC_2_24_6 .C_ON=1'b1;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNO_0_6_LC_2_24_6 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNO_0_6_LC_2_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNO_0_6_LC_2_24_6  (
            .in0(_gnd_net_),
            .in1(N__28641),
            .in2(N__19480),
            .in3(N__18529),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_s_6 ),
            .ltout(),
            .carryin(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_cry_5 ),
            .carryout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNO_0_7_LC_2_24_7 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNO_0_7_LC_2_24_7 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNO_0_7_LC_2_24_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNO_0_7_LC_2_24_7  (
            .in0(_gnd_net_),
            .in1(N__22183),
            .in2(_gnd_net_),
            .in3(N__18682),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_s_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.gen_bc_dec_un1_piosel_LC_3_7_7 .C_ON=1'b0;
    defparam \u0.gen_bc_dec_un1_piosel_LC_3_7_7 .SEQ_MODE=4'b0000;
    defparam \u0.gen_bc_dec_un1_piosel_LC_3_7_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \u0.gen_bc_dec_un1_piosel_LC_3_7_7  (
            .in0(_gnd_net_),
            .in1(N__18679),
            .in2(_gnd_net_),
            .in3(N__18657),
            .lcout(\u0.un1_piosel ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.irq_LC_3_14_6 .C_ON=1'b0;
    defparam \u1.irq_LC_3_14_6 .SEQ_MODE=4'b1000;
    defparam \u1.irq_LC_3_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.irq_LC_3_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18631),
            .lcout(irq),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54126),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_0_LC_3_17_0 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_0_LC_3_17_0 .SEQ_MODE=4'b1011;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_0_LC_3_17_0 .LUT_INIT=16'b1111101111001000;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_0_LC_3_17_0  (
            .in0(N__29662),
            .in1(N__18852),
            .in2(N__52577),
            .in3(N__18622),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.Qi_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54110),
            .ce(N__19570),
            .sr(N__53306));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_1_LC_3_17_1 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_1_LC_3_17_1 .SEQ_MODE=4'b1011;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_1_LC_3_17_1 .LUT_INIT=16'b1111110110101000;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_1_LC_3_17_1  (
            .in0(N__18853),
            .in1(N__29527),
            .in2(N__52573),
            .in3(N__18610),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.Qi_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54110),
            .ce(N__19570),
            .sr(N__53306));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_2_LC_3_17_2 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_2_LC_3_17_2 .SEQ_MODE=4'b1011;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_2_LC_3_17_2 .LUT_INIT=16'b1111101111001000;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_2_LC_3_17_2  (
            .in0(N__27481),
            .in1(N__18854),
            .in2(N__52578),
            .in3(N__18604),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.Qi_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54110),
            .ce(N__19570),
            .sr(N__53306));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_3_LC_3_17_3 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_3_LC_3_17_3 .SEQ_MODE=4'b1010;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_3_LC_3_17_3 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_3_LC_3_17_3  (
            .in0(N__18855),
            .in1(N__29482),
            .in2(N__52574),
            .in3(N__18598),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.Qi_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54110),
            .ce(N__19570),
            .sr(N__53306));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_4_LC_3_17_4 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_4_LC_3_17_4 .SEQ_MODE=4'b1011;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_4_LC_3_17_4 .LUT_INIT=16'b1111101111001000;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_4_LC_3_17_4  (
            .in0(N__29134),
            .in1(N__18856),
            .in2(N__52579),
            .in3(N__18592),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.Qi_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54110),
            .ce(N__19570),
            .sr(N__53306));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_5_LC_3_17_5 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_5_LC_3_17_5 .SEQ_MODE=4'b1010;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_5_LC_3_17_5 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_5_LC_3_17_5  (
            .in0(N__18857),
            .in1(N__27565),
            .in2(N__52575),
            .in3(N__18586),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.Qi_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54110),
            .ce(N__19570),
            .sr(N__53306));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_6_LC_3_17_6 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_6_LC_3_17_6 .SEQ_MODE=4'b1010;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_6_LC_3_17_6 .LUT_INIT=16'b0011101100001000;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_6_LC_3_17_6  (
            .in0(N__26203),
            .in1(N__18858),
            .in2(N__52580),
            .in3(N__18745),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.Qi_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54110),
            .ce(N__19570),
            .sr(N__53306));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_7_LC_3_17_7 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_7_LC_3_17_7 .SEQ_MODE=4'b1010;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_7_LC_3_17_7 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_7_LC_3_17_7  (
            .in0(N__18859),
            .in1(N__26176),
            .in2(N__52576),
            .in3(N__18739),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.Qi_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54110),
            .ce(N__19570),
            .sr(N__53306));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNIJBHR_0_LC_3_18_0 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNIJBHR_0_LC_3_18_0 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNIJBHR_0_LC_3_18_0 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNIJBHR_0_LC_3_18_0  (
            .in0(N__24724),
            .in1(N__24669),
            .in2(N__28954),
            .in3(N__18697),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.val_c8 ),
            .ltout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.val_c8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.hT2done_RNIFNDQ1_LC_3_18_1 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.hT2done_RNIFNDQ1_LC_3_18_1 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.hT2done_RNIFNDQ1_LC_3_18_1 .LUT_INIT=16'b1111111100100011;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.hT2done_RNIFNDQ1_LC_3_18_1  (
            .in0(N__24599),
            .in1(N__24515),
            .in2(N__18733),
            .in3(N__52588),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.N_1545 ),
            .ltout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.N_1545_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_1_LC_3_18_2 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_1_LC_3_18_2 .SEQ_MODE=4'b1011;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_1_LC_3_18_2 .LUT_INIT=16'b1110111111100000;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_1_LC_3_18_2  (
            .in0(N__52581),
            .in1(N__29506),
            .in2(N__18730),
            .in3(N__18727),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.QiZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54116),
            .ce(N__18775),
            .sr(N__53309));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_6_LC_3_18_3 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_6_LC_3_18_3 .SEQ_MODE=4'b1010;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_6_LC_3_18_3 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_6_LC_3_18_3  (
            .in0(N__18846),
            .in1(N__29116),
            .in2(N__52768),
            .in3(N__18718),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.QiZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54116),
            .ce(N__18775),
            .sr(N__53309));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_7_LC_3_18_4 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_7_LC_3_18_4 .SEQ_MODE=4'b1010;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_7_LC_3_18_4 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_7_LC_3_18_4  (
            .in0(N__27583),
            .in1(N__18706),
            .in2(N__52693),
            .in3(N__18847),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.QiZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54116),
            .ce(N__18775),
            .sr(N__53309));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNI2MD5_1_LC_3_18_5 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNI2MD5_1_LC_3_18_5 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNI2MD5_1_LC_3_18_5 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNI2MD5_1_LC_3_18_5  (
            .in0(N__28821),
            .in1(N__28857),
            .in2(_gnd_net_),
            .in3(N__28920),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.val_c8_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_3_LC_3_18_6 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_3_LC_3_18_6 .SEQ_MODE=4'b1010;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_3_LC_3_18_6 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_3_LC_3_18_6  (
            .in0(N__26623),
            .in1(N__18691),
            .in2(N__52692),
            .in3(N__18845),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.QiZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54116),
            .ce(N__18775),
            .sr(N__53309));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qilde_i_LC_3_18_7 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qilde_i_LC_3_18_7 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qilde_i_LC_3_18_7 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qilde_i_LC_3_18_7  (
            .in0(N__24546),
            .in1(N__24516),
            .in2(_gnd_net_),
            .in3(N__19582),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.N_290 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNIPRNI_0_LC_3_19_0 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNIPRNI_0_LC_3_19_0 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNIPRNI_0_LC_3_19_0 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNIPRNI_0_LC_3_19_0  (
            .in0(N__19020),
            .in1(N__19005),
            .in2(N__20680),
            .in3(N__18875),
            .lcout(),
            .ltout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNIPRNIZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNIMTBN_0_LC_3_19_1 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNIMTBN_0_LC_3_19_1 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNIMTBN_0_LC_3_19_1 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNIMTBN_0_LC_3_19_1  (
            .in0(N__28583),
            .in1(_gnd_net_),
            .in2(N__18994),
            .in3(N__18973),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.val_c7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNIT1K4_2_LC_3_19_2 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNIT1K4_2_LC_3_19_2 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNIT1K4_2_LC_3_19_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNIT1K4_2_LC_3_19_2  (
            .in0(N__18786),
            .in1(N__18915),
            .in2(N__18990),
            .in3(N__18948),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.val_c7_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_2_LC_3_19_3 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_2_LC_3_19_3 .SEQ_MODE=4'b1010;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_2_LC_3_19_3 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_2_LC_3_19_3  (
            .in0(N__26641),
            .in1(N__18967),
            .in2(N__52771),
            .in3(N__18849),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.QiZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54121),
            .ce(N__18771),
            .sr(N__53313));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_4_LC_3_19_4 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_4_LC_3_19_4 .SEQ_MODE=4'b1010;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_4_LC_3_19_4 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_4_LC_3_19_4  (
            .in0(N__18850),
            .in1(N__52732),
            .in2(N__18937),
            .in3(N__26608),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.QiZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54121),
            .ce(N__18771),
            .sr(N__53313));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_0_LC_3_19_5 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_0_LC_3_19_5 .SEQ_MODE=4'b1010;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_0_LC_3_19_5 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_0_LC_3_19_5  (
            .in0(N__27493),
            .in1(N__18904),
            .in2(N__52770),
            .in3(N__18848),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.QiZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54121),
            .ce(N__18771),
            .sr(N__53313));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_5_LC_3_19_6 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_5_LC_3_19_6 .SEQ_MODE=4'b1010;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_5_LC_3_19_6 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_5_LC_3_19_6  (
            .in0(N__18851),
            .in1(N__26590),
            .in2(N__52772),
            .in3(N__18805),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.QiZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54121),
            .ce(N__18771),
            .sr(N__53313));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_1_sqmuxa_i_x0_LC_3_20_0 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_1_sqmuxa_i_x0_LC_3_20_0 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_1_sqmuxa_i_x0_LC_3_20_0 .LUT_INIT=16'b1111000011110010;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_1_sqmuxa_i_x0_LC_3_20_0  (
            .in0(N__19983),
            .in1(N__19860),
            .in2(N__52695),
            .in3(N__19913),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_1_sqmuxa_i_x0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_1_LC_3_20_2 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_1_LC_3_20_2 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_1_LC_3_20_2 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_1_LC_3_20_2  (
            .in0(N__19255),
            .in1(N__19243),
            .in2(N__52694),
            .in3(N__19134),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.QiZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54127),
            .ce(N__19071),
            .sr(N__53317));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_3_LC_3_20_4 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_3_LC_3_20_4 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_3_LC_3_20_4 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_3_LC_3_20_4  (
            .in0(N__27544),
            .in1(N__19225),
            .in2(N__52696),
            .in3(N__19135),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.QiZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54127),
            .ce(N__19071),
            .sr(N__53317));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_4_LC_3_20_5 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_4_LC_3_20_5 .SEQ_MODE=4'b1011;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_4_LC_3_20_5 .LUT_INIT=16'b1111110110101000;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_4_LC_3_20_5  (
            .in0(N__19136),
            .in1(N__19201),
            .in2(N__52773),
            .in3(N__19189),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.QiZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54127),
            .ce(N__19071),
            .sr(N__53317));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_5_LC_3_20_6 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_5_LC_3_20_6 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_5_LC_3_20_6 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_5_LC_3_20_6  (
            .in0(N__19168),
            .in1(N__19156),
            .in2(N__52697),
            .in3(N__19137),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.QiZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54127),
            .ce(N__19071),
            .sr(N__53317));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_6_LC_3_20_7 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_6_LC_3_20_7 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_6_LC_3_20_7 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.Qi_6_LC_3_20_7  (
            .in0(N__19138),
            .in1(N__19105),
            .in2(N__52774),
            .in3(N__19093),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.eoc_cnt.cnt.QiZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54127),
            .ce(N__19071),
            .sr(N__53317));
    defparam \u0.PIO_cmdport_T2_RNINM6Q3_5_LC_3_21_0 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_T2_RNINM6Q3_5_LC_3_21_0 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_cmdport_T2_RNINM6Q3_5_LC_3_21_0 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \u0.PIO_cmdport_T2_RNINM6Q3_5_LC_3_21_0  (
            .in0(N__23653),
            .in1(N__48144),
            .in2(N__48332),
            .in3(N__29644),
            .lcout(\u0.dat_o_0_0_2_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.dstrb_RNIBHHI_LC_3_21_1 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.dstrb_RNIBHHI_LC_3_21_1 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.dstrb_RNIBHHI_LC_3_21_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.dstrb_RNIBHHI_LC_3_21_1  (
            .in0(_gnd_net_),
            .in1(N__22493),
            .in2(_gnd_net_),
            .in3(N__23651),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.rd_dstrb ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.dstrb_LC_3_21_2 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.dstrb_LC_3_21_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.dstrb_LC_3_21_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.dstrb_LC_3_21_2  (
            .in0(N__19855),
            .in1(N__19734),
            .in2(N__19996),
            .in3(N__19915),
            .lcout(\u1.DMA_control.dstrb ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54132),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.DIOW_RNO_1_LC_3_21_3 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.DIOW_RNO_1_LC_3_21_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.DIOW_RNO_1_LC_3_21_3 .LUT_INIT=16'b0000111000001100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.DIOW_RNO_1_LC_3_21_3  (
            .in0(N__19398),
            .in1(N__23652),
            .in2(N__52609),
            .in3(N__20020),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.DIOW_RNO_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNIM65O1_0_LC_3_21_4 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNIM65O1_0_LC_3_21_4 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNIM65O1_0_LC_3_21_4 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNIM65O1_0_LC_3_21_4  (
            .in0(N__19854),
            .in1(N__19733),
            .in2(N__19995),
            .in3(N__19914),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.Tddone_i ),
            .ltout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.Tddone_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.DIOR_RNO_0_LC_3_21_5 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.DIOR_RNO_0_LC_3_21_5 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.DIOR_RNO_0_LC_3_21_5 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.DIOR_RNO_0_LC_3_21_5  (
            .in0(N__20105),
            .in1(_gnd_net_),
            .in2(N__19339),
            .in3(N__52602),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.DIOR_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.DIOR_RNO_1_LC_3_21_6 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.DIOR_RNO_1_LC_3_21_6 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.DIOR_RNO_1_LC_3_21_6 .LUT_INIT=16'b0000100000001111;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.DIOR_RNO_1_LC_3_21_6  (
            .in0(N__20019),
            .in1(N__20106),
            .in2(N__52698),
            .in3(N__23654),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.DIOR_RNO_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.DIOW_RNO_0_LC_3_21_7 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.DIOW_RNO_0_LC_3_21_7 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.DIOW_RNO_0_LC_3_21_7 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.DIOW_RNO_0_LC_3_21_7  (
            .in0(N__52436),
            .in1(N__19397),
            .in2(_gnd_net_),
            .in3(N__20018),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.DIOW_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DIOWn_LC_3_22_0 .C_ON=1'b0;
    defparam \u1.DIOWn_LC_3_22_0 .SEQ_MODE=4'b1011;
    defparam \u1.DIOWn_LC_3_22_0 .LUT_INIT=16'b1111010011110111;
    LogicCell40 \u1.DIOWn_LC_3_22_0  (
            .in0(N__19606),
            .in1(N__36668),
            .in2(N__52788),
            .in3(N__19399),
            .lcout(diown_pad_o_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54139),
            .ce(),
            .sr(N__53323));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNIIK4B1_1_LC_3_22_1 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNIIK4B1_1_LC_3_22_1 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNIIK4B1_1_LC_3_22_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNIIK4B1_1_LC_3_22_1  (
            .in0(N__19317),
            .in1(N__19305),
            .in2(N__19291),
            .in3(N__19272),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.val_c8_a0_4 ),
            .ltout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.val_c8_a0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNI71R53_0_LC_3_22_2 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNI71R53_0_LC_3_22_2 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNI71R53_0_LC_3_22_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNI71R53_0_LC_3_22_2  (
            .in0(N__19440),
            .in1(N__20060),
            .in2(N__19261),
            .in3(N__19453),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.Tmdone_i_i ),
            .ltout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.Tmdone_i_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qie_0_i_LC_3_22_3 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qie_0_i_LC_3_22_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qie_0_i_LC_3_22_3 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qie_0_i_LC_3_22_3  (
            .in0(_gnd_net_),
            .in1(N__52780),
            .in2(N__19258),
            .in3(N__19981),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qie_0_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNI8QB01_7_LC_3_22_4 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNI8QB01_7_LC_3_22_4 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNI8QB01_7_LC_3_22_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_RNI8QB01_7_LC_3_22_4  (
            .in0(N__22179),
            .in1(N__19476),
            .in2(_gnd_net_),
            .in3(N__19464),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.val_c8_a0_3 ),
            .ltout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.val_c8_a0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.N_2415_i_x1_LC_3_22_5 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.N_2415_i_x1_LC_3_22_5 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.N_2415_i_x1_LC_3_22_5 .LUT_INIT=16'b1100110011101100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.N_2415_i_x1_LC_3_22_5  (
            .in0(N__20059),
            .in1(N__52779),
            .in2(N__19447),
            .in3(N__19439),
            .lcout(),
            .ltout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.N_2415_i_xZ0Z1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.N_2415_i_ns_LC_3_22_6 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.N_2415_i_ns_LC_3_22_6 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.N_2415_i_ns_LC_3_22_6 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.N_2415_i_ns_LC_3_22_6  (
            .in0(N__52778),
            .in1(_gnd_net_),
            .in2(N__19420),
            .in3(N__19417),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.N_2415_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.DIOW_LC_3_22_7 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.DIOW_LC_3_22_7 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.DIOW_LC_3_22_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.DIOW_LC_3_22_7  (
            .in0(N__20041),
            .in1(N__19411),
            .in2(_gnd_net_),
            .in3(N__19405),
            .lcout(\u1.DMAdiow ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54139),
            .ce(),
            .sr(N__53323));
    defparam \u1.PIOtip_LC_3_23_0 .C_ON=1'b0;
    defparam \u1.PIOtip_LC_3_23_0 .SEQ_MODE=4'b1010;
    defparam \u1.PIOtip_LC_3_23_0 .LUT_INIT=16'b0101000001010001;
    LogicCell40 \u1.PIOtip_LC_3_23_0  (
            .in0(N__19489),
            .in1(N__20833),
            .in2(N__36694),
            .in3(N__20801),
            .lcout(PIOtip),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54146),
            .ce(),
            .sr(N__53327));
    defparam \u1.DDoe_RNO_0_LC_3_23_1 .C_ON=1'b0;
    defparam \u1.DDoe_RNO_0_LC_3_23_1 .SEQ_MODE=4'b0000;
    defparam \u1.DDoe_RNO_0_LC_3_23_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \u1.DDoe_RNO_0_LC_3_23_1  (
            .in0(N__19350),
            .in1(N__36662),
            .in2(_gnd_net_),
            .in3(N__21499),
            .lcout(),
            .ltout(\u1.N_1395_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DDoe_LC_3_23_2 .C_ON=1'b0;
    defparam \u1.DDoe_LC_3_23_2 .SEQ_MODE=4'b1010;
    defparam \u1.DDoe_LC_3_23_2 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \u1.DDoe_LC_3_23_2  (
            .in0(N__36664),
            .in1(N__52782),
            .in2(N__19381),
            .in3(N__23650),
            .lcout(dd_padoe_o_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54146),
            .ce(),
            .sr(N__53327));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNIU87U_7_LC_3_23_3 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNIU87U_7_LC_3_23_3 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNIU87U_7_LC_3_23_3 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNIU87U_7_LC_3_23_3  (
            .in0(N__52783),
            .in1(N__20883),
            .in2(_gnd_net_),
            .in3(N__20850),
            .lcout(\u1.N_1387 ),
            .ltout(\u1.N_1387_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.oe_LC_3_23_4 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.oe_LC_3_23_4 .SEQ_MODE=4'b1010;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.oe_LC_3_23_4 .LUT_INIT=16'b0000101100001010;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.oe_LC_3_23_4  (
            .in0(N__19351),
            .in1(N__23284),
            .in2(N__19354),
            .in3(N__26364),
            .lcout(\u1.PIOoe ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54146),
            .ce(),
            .sr(N__53327));
    defparam \u1.PIO_control.gen_pingpong_pong_d_RNIL3IN_9_LC_3_23_5 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_pong_d_RNIL3IN_9_LC_3_23_5 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.gen_pingpong_pong_d_RNIL3IN_9_LC_3_23_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.PIO_control.gen_pingpong_pong_d_RNIL3IN_9_LC_3_23_5  (
            .in0(N__19519),
            .in1(N__20617),
            .in2(_gnd_net_),
            .in3(N__26929),
            .lcout(),
            .ltout(\u1.N_1434_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DDo_9_LC_3_23_6 .C_ON=1'b0;
    defparam \u1.DDo_9_LC_3_23_6 .SEQ_MODE=4'b1010;
    defparam \u1.DDo_9_LC_3_23_6 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \u1.DDo_9_LC_3_23_6  (
            .in0(N__36663),
            .in1(N__52781),
            .in2(N__19504),
            .in3(N__23896),
            .lcout(dd_pad_o_c_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54146),
            .ce(),
            .sr(N__53327));
    defparam \u1.c_state_0_LC_3_23_7 .C_ON=1'b0;
    defparam \u1.c_state_0_LC_3_23_7 .SEQ_MODE=4'b1010;
    defparam \u1.c_state_0_LC_3_23_7 .LUT_INIT=16'b0000000000110001;
    LogicCell40 \u1.c_state_0_LC_3_23_7  (
            .in0(N__20802),
            .in1(N__24405),
            .in2(N__24445),
            .in3(N__19488),
            .lcout(\u1.c_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54146),
            .ce(),
            .sr(N__53327));
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_30_LC_3_24_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_30_LC_3_24_0 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_30_LC_3_24_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Txbuf.Q_30_LC_3_24_0  (
            .in0(N__47795),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23862),
            .lcout(\u1.DMA_control.TxbufQ_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54152),
            .ce(N__21163),
            .sr(N__53331));
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_21_LC_3_24_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_21_LC_3_24_1 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_21_LC_3_24_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Txbuf.Q_21_LC_3_24_1  (
            .in0(N__23859),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38047),
            .lcout(\u1.DMA_control.TxbufQ_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54152),
            .ce(N__21163),
            .sr(N__53331));
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_31_LC_3_24_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_31_LC_3_24_2 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_31_LC_3_24_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Txbuf.Q_31_LC_3_24_2  (
            .in0(N__40488),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23863),
            .lcout(\u1.DMA_control.TxbufQ_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54152),
            .ce(N__21163),
            .sr(N__53331));
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_5_LC_3_24_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_5_LC_3_24_3 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_5_LC_3_24_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Txbuf.Q_5_LC_3_24_3  (
            .in0(N__23864),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46288),
            .lcout(\u1.DMA_control.TxbufQ_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54152),
            .ce(N__21163),
            .sr(N__53331));
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_6_LC_3_24_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_6_LC_3_24_4 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_6_LC_3_24_4 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Txbuf.Q_6_LC_3_24_4  (
            .in0(N__39480),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23865),
            .lcout(\u1.DMA_control.TxbufQ_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54152),
            .ce(N__21163),
            .sr(N__53331));
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_2_LC_3_24_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_2_LC_3_24_5 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_2_LC_3_24_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Txbuf.Q_2_LC_3_24_5  (
            .in0(N__23861),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34276),
            .lcout(\u1.DMA_control.TxbufQ_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54152),
            .ce(N__21163),
            .sr(N__53331));
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_1_LC_3_24_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_1_LC_3_24_6 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_1_LC_3_24_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Txbuf.Q_1_LC_3_24_6  (
            .in0(N__39358),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23858),
            .lcout(\u1.DMA_control.TxbufQ_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54152),
            .ce(N__21163),
            .sr(N__53331));
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_25_LC_3_24_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_25_LC_3_24_7 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_25_LC_3_24_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Txbuf.Q_25_LC_3_24_7  (
            .in0(N__23860),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40839),
            .lcout(\u1.DMA_control.TxbufQ_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54152),
            .ce(N__21163),
            .sr(N__53331));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__18_LC_3_25_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__18_LC_3_25_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__18_LC_3_25_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__18_LC_3_25_1  (
            .in0(N__30432),
            .in1(N__30286),
            .in2(_gnd_net_),
            .in3(N__42962),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54163),
            .ce(N__41833),
            .sr(_gnd_net_));
    defparam \u0.CtrlReg_20_LC_3_26_1 .C_ON=1'b0;
    defparam \u0.CtrlReg_20_LC_3_26_1 .SEQ_MODE=4'b1010;
    defparam \u0.CtrlReg_20_LC_3_26_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.CtrlReg_20_LC_3_26_1  (
            .in0(N__34780),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52789),
            .lcout(\u0.CtrlRegZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54174),
            .ce(N__53641),
            .sr(N__53346));
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_2_LC_3_27_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_2_LC_3_27_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_2_LC_3_27_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_readDlw_2_LC_3_27_1  (
            .in0(N__32298),
            .in1(N__32336),
            .in2(_gnd_net_),
            .in3(N__42961),
            .lcout(\u1.DMA_control.readDlw_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54186),
            .ce(N__36327),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_2_LC_3_30_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_2_LC_3_30_0 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_2_LC_3_30_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_readDfw_2_LC_3_30_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30460),
            .lcout(\u1.DMA_control.readDfw_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54225),
            .ce(N__36325),
            .sr(_gnd_net_));
    defparam \u1.synch_incoming_cIORDY_LC_4_10_6 .C_ON=1'b0;
    defparam \u1.synch_incoming_cIORDY_LC_4_10_6 .SEQ_MODE=4'b1000;
    defparam \u1.synch_incoming_cIORDY_LC_4_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.synch_incoming_cIORDY_LC_4_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19540),
            .lcout(\u1.cIORDY ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54164),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.sIORDY_LC_4_16_0 .C_ON=1'b0;
    defparam \u1.sIORDY_LC_4_16_0 .SEQ_MODE=4'b1000;
    defparam \u1.sIORDY_LC_4_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.sIORDY_LC_4_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19528),
            .lcout(\u1.sIORDYZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54122),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.gen_regs_un1_ena_i_0_a2_0_LC_4_16_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.gen_regs_un1_ena_i_0_a2_0_LC_4_16_1 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.gen_regs_un1_ena_i_0_a2_0_LC_4_16_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.gen_regs_un1_ena_i_0_a2_0_LC_4_16_1  (
            .in0(N__21805),
            .in1(N__21840),
            .in2(_gnd_net_),
            .in3(N__21873),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.N_2138 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.c_state_1_LC_4_17_4 .C_ON=1'b0;
    defparam \u1.c_state_1_LC_4_17_4 .SEQ_MODE=4'b1010;
    defparam \u1.c_state_1_LC_4_17_4 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \u1.c_state_1_LC_4_17_4  (
            .in0(N__20266),
            .in1(N__21555),
            .in2(N__24364),
            .in3(N__21529),
            .lcout(\u1.c_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54113),
            .ce(),
            .sr(N__53310));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qilde_i_sx_LC_4_18_0 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qilde_i_sx_LC_4_18_0 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qilde_i_sx_LC_4_18_0 .LUT_INIT=16'b1111111111110010;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qilde_i_sx_LC_4_18_0  (
            .in0(N__24587),
            .in1(N__24502),
            .in2(N__52459),
            .in3(N__20672),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qilde_i_sxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.hT2done_LC_4_18_1 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.hT2done_LC_4_18_1 .SEQ_MODE=4'b1010;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.hT2done_LC_4_18_1 .LUT_INIT=16'b0010001000000010;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.hT2done_LC_4_18_1  (
            .in0(N__24505),
            .in1(N__52253),
            .in2(N__24561),
            .in3(N__24589),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.hT2doneZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54123),
            .ce(),
            .sr(N__53314));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.rci_RNO_1_LC_4_18_2 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.rci_RNO_1_LC_4_18_2 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.rci_RNO_1_LC_4_18_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.rci_RNO_1_LC_4_18_2  (
            .in0(N__20430),
            .in1(N__20501),
            .in2(N__20559),
            .in3(N__20478),
            .lcout(),
            .ltout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.rci_3_i_a0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.rci_RNO_0_LC_4_18_3 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.rci_RNO_0_LC_4_18_3 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.rci_RNO_0_LC_4_18_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.rci_RNO_0_LC_4_18_3  (
            .in0(N__20381),
            .in1(N__19558),
            .in2(N__19576),
            .in3(N__20348),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.rci_3_i_a0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qilde_i_sx_LC_4_18_4 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qilde_i_sx_LC_4_18_4 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qilde_i_sx_LC_4_18_4 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qilde_i_sx_LC_4_18_4  (
            .in0(N__24588),
            .in1(N__20380),
            .in2(N__52460),
            .in3(N__24503),
            .lcout(),
            .ltout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qilde_i_sxZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qilde_i_LC_4_18_5 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qilde_i_LC_4_18_5 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qilde_i_LC_4_18_5 .LUT_INIT=16'b1111000111110001;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qilde_i_LC_4_18_5  (
            .in0(N__24504),
            .in1(N__24547),
            .in2(N__19573),
            .in3(_gnd_net_),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.N_1083 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.rci_RNO_2_LC_4_18_6 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.rci_RNO_2_LC_4_18_6 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.rci_RNO_2_LC_4_18_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.rci_RNO_2_LC_4_18_6  (
            .in0(N__20528),
            .in1(N__20454),
            .in2(_gnd_net_),
            .in3(N__20403),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.rci_3_i_a0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.rci_LC_4_18_7 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.rci_LC_4_18_7 .SEQ_MODE=4'b1010;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.rci_LC_4_18_7 .LUT_INIT=16'b0000001000110011;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.rci_LC_4_18_7  (
            .in0(N__20382),
            .in1(N__52252),
            .in2(N__19552),
            .in3(N__20698),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.rci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54123),
            .ce(),
            .sr(N__53314));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.DIOR_RNO_0_LC_4_19_0 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.DIOR_RNO_0_LC_4_19_0 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.DIOR_RNO_0_LC_4_19_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.DIOR_RNO_0_LC_4_19_0  (
            .in0(N__28584),
            .in1(N__19621),
            .in2(_gnd_net_),
            .in3(N__21375),
            .lcout(),
            .ltout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.N_1377_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.DIOR_LC_4_19_1 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.DIOR_LC_4_19_1 .SEQ_MODE=4'b1010;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.DIOR_LC_4_19_1 .LUT_INIT=16'b0010001100000011;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.DIOR_LC_4_19_1  (
            .in0(N__19656),
            .in1(N__52245),
            .in2(N__19543),
            .in3(N__20696),
            .lcout(\u1.PIOdior ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54128),
            .ce(),
            .sr(N__53318));
    defparam \u1.DIORn_LC_4_19_2 .C_ON=1'b0;
    defparam \u1.DIORn_LC_4_19_2 .SEQ_MODE=4'b1011;
    defparam \u1.DIORn_LC_4_19_2 .LUT_INIT=16'b1100111111011101;
    LogicCell40 \u1.DIORn_LC_4_19_2  (
            .in0(N__20107),
            .in1(N__52262),
            .in2(N__19660),
            .in3(N__36730),
            .lcout(diorn_pad_o_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54128),
            .ce(),
            .sr(N__53318));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.DIOR_RNO_1_LC_4_19_3 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.DIOR_RNO_1_LC_4_19_3 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.DIOR_RNO_1_LC_4_19_3 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.DIOR_RNO_1_LC_4_19_3  (
            .in0(N__26078),
            .in1(N__20747),
            .in2(N__23257),
            .in3(N__26344),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.DIOR_RNOZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_pong_we_RNI38NC_LC_4_19_4 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_pong_we_RNI38NC_LC_4_19_4 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.gen_pingpong_pong_we_RNI38NC_LC_4_19_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.PIO_control.gen_pingpong_pong_we_RNI38NC_LC_4_19_4  (
            .in0(N__20940),
            .in1(N__20922),
            .in2(_gnd_net_),
            .in3(N__26896),
            .lcout(\u1.PIO_control.N_1450 ),
            .ltout(\u1.PIO_control.N_1450_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.DIOW_RNO_1_LC_4_19_5 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.DIOW_RNO_1_LC_4_19_5 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.DIOW_RNO_1_LC_4_19_5 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.DIOW_RNO_1_LC_4_19_5  (
            .in0(N__26079),
            .in1(N__20748),
            .in2(N__19615),
            .in3(N__23256),
            .lcout(),
            .ltout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.DIOW_RNOZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.DIOW_RNO_0_LC_4_19_6 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.DIOW_RNO_0_LC_4_19_6 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.DIOW_RNO_0_LC_4_19_6 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.DIOW_RNO_0_LC_4_19_6  (
            .in0(N__28585),
            .in1(_gnd_net_),
            .in2(N__19612),
            .in3(N__21376),
            .lcout(),
            .ltout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.N_1378_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.DIOW_LC_4_19_7 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.DIOW_LC_4_19_7 .SEQ_MODE=4'b1010;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.DIOW_LC_4_19_7 .LUT_INIT=16'b0100010100000101;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.DIOW_LC_4_19_7  (
            .in0(N__52263),
            .in1(N__19599),
            .in2(N__19609),
            .in3(N__20697),
            .lcout(\u1.PIOdiow ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54128),
            .ce(),
            .sr(N__53318));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_cry_c_0_LC_4_20_0 .C_ON=1'b1;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_cry_c_0_LC_4_20_0 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_cry_c_0_LC_4_20_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_cry_c_0_LC_4_20_0  (
            .in0(_gnd_net_),
            .in1(N__19859),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_20_0_),
            .carryout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNO_0_1_LC_4_20_1 .C_ON=1'b1;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNO_0_1_LC_4_20_1 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNO_0_1_LC_4_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNO_0_1_LC_4_20_1  (
            .in0(_gnd_net_),
            .in1(N__19927),
            .in2(N__28580),
            .in3(N__19588),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_s_1 ),
            .ltout(),
            .carryin(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_cry_0 ),
            .carryout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNO_0_2_LC_4_20_2 .C_ON=1'b1;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNO_0_2_LC_4_20_2 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNO_0_2_LC_4_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNO_0_2_LC_4_20_2  (
            .in0(_gnd_net_),
            .in1(N__28515),
            .in2(N__19714),
            .in3(N__19585),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_s_2 ),
            .ltout(),
            .carryin(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_cry_1 ),
            .carryout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNO_0_3_LC_4_20_3 .C_ON=1'b1;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNO_0_3_LC_4_20_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNO_0_3_LC_4_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNO_0_3_LC_4_20_3  (
            .in0(_gnd_net_),
            .in1(N__19894),
            .in2(N__28581),
            .in3(N__19756),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_s_3 ),
            .ltout(),
            .carryin(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_cry_2 ),
            .carryout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNO_0_4_LC_4_20_4 .C_ON=1'b1;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNO_0_4_LC_4_20_4 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNO_0_4_LC_4_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNO_0_4_LC_4_20_4  (
            .in0(_gnd_net_),
            .in1(N__28519),
            .in2(N__19789),
            .in3(N__19753),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_s_4 ),
            .ltout(),
            .carryin(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_cry_3 ),
            .carryout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNO_0_5_LC_4_20_5 .C_ON=1'b1;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNO_0_5_LC_4_20_5 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNO_0_5_LC_4_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNO_0_5_LC_4_20_5  (
            .in0(_gnd_net_),
            .in1(N__19693),
            .in2(N__28582),
            .in3(N__19750),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_s_5 ),
            .ltout(),
            .carryin(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_cry_4 ),
            .carryout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNO_0_6_LC_4_20_6 .C_ON=1'b1;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNO_0_6_LC_4_20_6 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNO_0_6_LC_4_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNO_0_6_LC_4_20_6  (
            .in0(_gnd_net_),
            .in1(N__28523),
            .in2(N__19675),
            .in3(N__19747),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_s_6 ),
            .ltout(),
            .carryin(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_cry_5 ),
            .carryout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNO_0_7_LC_4_20_7 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNO_0_7_LC_4_20_7 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNO_0_7_LC_4_20_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNO_0_7_LC_4_20_7  (
            .in0(_gnd_net_),
            .in1(N__19947),
            .in2(_gnd_net_),
            .in3(N__19744),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_s_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNIO59K_7_LC_4_21_0 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNIO59K_7_LC_4_21_0 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNIO59K_7_LC_4_21_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNIO59K_7_LC_4_21_0  (
            .in0(N__19671),
            .in1(N__19692),
            .in2(N__19948),
            .in3(N__19710),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.val_c8_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_2_LC_4_21_1 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_2_LC_4_21_1 .SEQ_MODE=4'b1011;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_2_LC_4_21_1 .LUT_INIT=16'b1111101011001100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_2_LC_4_21_1  (
            .in0(N__21442),
            .in1(N__19720),
            .in2(N__52607),
            .in3(N__19824),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.QiZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54140),
            .ce(N__19770),
            .sr(N__53324));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_5_LC_4_21_2 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_5_LC_4_21_2 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_5_LC_4_21_2 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_5_LC_4_21_2  (
            .in0(N__19826),
            .in1(N__23971),
            .in2(N__52461),
            .in3(N__19699),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.QiZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54140),
            .ce(N__19770),
            .sr(N__53324));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_6_LC_4_21_3 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_6_LC_4_21_3 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_6_LC_4_21_3 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_6_LC_4_21_3  (
            .in0(N__31630),
            .in1(N__19681),
            .in2(N__52608),
            .in3(N__19827),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.QiZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54140),
            .ce(N__19770),
            .sr(N__53324));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_7_LC_4_21_4 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_7_LC_4_21_4 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_7_LC_4_21_4 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_7_LC_4_21_4  (
            .in0(N__19828),
            .in1(N__21715),
            .in2(N__52462),
            .in3(N__19954),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.QiZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54140),
            .ce(N__19770),
            .sr(N__53324));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_1_LC_4_21_5 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_1_LC_4_21_5 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_1_LC_4_21_5 .LUT_INIT=16'b0000110010101010;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_1_LC_4_21_5  (
            .in0(N__19933),
            .in1(N__26512),
            .in2(N__52606),
            .in3(N__19823),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.QiZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54140),
            .ce(N__19770),
            .sr(N__53324));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNI3L6F_1_LC_4_21_6 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNI3L6F_1_LC_4_21_6 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNI3L6F_1_LC_4_21_6 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_RNI3L6F_1_LC_4_21_6  (
            .in0(N__19782),
            .in1(N__19893),
            .in2(_gnd_net_),
            .in3(N__19926),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.val_c8_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_3_LC_4_21_7 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_3_LC_4_21_7 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_3_LC_4_21_7 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_3_LC_4_21_7  (
            .in0(N__19900),
            .in1(N__52255),
            .in2(N__21739),
            .in3(N__19825),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.QiZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54140),
            .ce(N__19770),
            .sr(N__53324));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_0_LC_4_22_0 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_0_LC_4_22_0 .SEQ_MODE=4'b1011;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_0_LC_4_22_0 .LUT_INIT=16'b1110111011110000;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_0_LC_4_22_0  (
            .in0(N__21970),
            .in1(N__52463),
            .in2(N__19882),
            .in3(N__19821),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.Qi_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54147),
            .ce(N__19771),
            .sr(N__53328));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_4_LC_4_22_1 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_4_LC_4_22_1 .SEQ_MODE=4'b1011;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_4_LC_4_22_1 .LUT_INIT=16'b1111110110101000;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.Qi_4_LC_4_22_1  (
            .in0(N__19822),
            .in1(N__21727),
            .in2(N__52623),
            .in3(N__19798),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.cnt.QiZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54147),
            .ce(N__19771),
            .sr(N__53328));
    defparam \u1.DMA_control.gen_DMA_req_hgo_RNO_0_LC_4_22_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_req_hgo_RNO_0_LC_4_22_2 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMA_req_hgo_RNO_0_LC_4_22_2 .LUT_INIT=16'b1100110111001100;
    LogicCell40 \u1.DMA_control.gen_DMA_req_hgo_RNO_0_LC_4_22_2  (
            .in0(N__20263),
            .in1(N__52467),
            .in2(N__21014),
            .in3(N__22494),
            .lcout(\u1.DMA_control.hgo_2_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMAtip_RNO_0_LC_4_22_3 .C_ON=1'b0;
    defparam \u1.DMAtip_RNO_0_LC_4_22_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMAtip_RNO_0_LC_4_22_3 .LUT_INIT=16'b0011001100010001;
    LogicCell40 \u1.DMAtip_RNO_0_LC_4_22_3  (
            .in0(N__21424),
            .in1(N__20264),
            .in2(_gnd_net_),
            .in3(N__23659),
            .lcout(\u1.DMAtip_2_i_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_req_iDMA_req_RNO_2_LC_4_22_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_req_iDMA_req_RNO_2_LC_4_22_4 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMA_req_iDMA_req_RNO_2_LC_4_22_4 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \u1.DMA_control.gen_DMA_req_iDMA_req_RNO_2_LC_4_22_4  (
            .in0(N__23658),
            .in1(N__52469),
            .in2(N__24972),
            .in3(N__21426),
            .lcout(),
            .ltout(\u1.DMA_control.iDMA_req_2_0_0_a2_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_req_iDMA_req_RNO_0_LC_4_22_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_req_iDMA_req_RNO_0_LC_4_22_5 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMA_req_iDMA_req_RNO_0_LC_4_22_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \u1.DMA_control.gen_DMA_req_iDMA_req_RNO_0_LC_4_22_5  (
            .in0(N__20979),
            .in1(N__20181),
            .in2(N__20185),
            .in3(N__31443),
            .lcout(\u1.DMA_control.N_1769 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_req_iDMA_req_RNO_1_LC_4_22_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_req_iDMA_req_RNO_1_LC_4_22_6 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMA_req_iDMA_req_RNO_1_LC_4_22_6 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \u1.DMA_control.gen_DMA_req_iDMA_req_RNO_1_LC_4_22_6  (
            .in0(N__20182),
            .in1(_gnd_net_),
            .in2(N__24973),
            .in3(N__52468),
            .lcout(\u1.DMA_control.iDMA_req_2_0_0_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.sDMARQ_RNIBPTG1_LC_4_22_7 .C_ON=1'b0;
    defparam \u1.sDMARQ_RNIBPTG1_LC_4_22_7 .SEQ_MODE=4'b0000;
    defparam \u1.sDMARQ_RNIBPTG1_LC_4_22_7 .LUT_INIT=16'b1000100011111111;
    LogicCell40 \u1.sDMARQ_RNIBPTG1_LC_4_22_7  (
            .in0(N__21425),
            .in1(N__24964),
            .in2(_gnd_net_),
            .in3(N__21148),
            .lcout(\u1.N_1372 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.register_block_gen_stat_reg_int_LC_4_23_0 .C_ON=1'b0;
    defparam \u0.register_block_gen_stat_reg_int_LC_4_23_0 .SEQ_MODE=4'b1010;
    defparam \u0.register_block_gen_stat_reg_int_LC_4_23_0 .LUT_INIT=16'b0000110000001110;
    LogicCell40 \u0.register_block_gen_stat_reg_int_LC_4_23_0  (
            .in0(N__20152),
            .in1(N__37079),
            .in2(N__26026),
            .in3(N__20134),
            .lcout(wb_inta_o_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54153),
            .ce(),
            .sr(N__53332));
    defparam \u0.register_block_gen_stat_reg_dirq_LC_4_23_1 .C_ON=1'b0;
    defparam \u0.register_block_gen_stat_reg_dirq_LC_4_23_1 .SEQ_MODE=4'b1010;
    defparam \u0.register_block_gen_stat_reg_dirq_LC_4_23_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \u0.register_block_gen_stat_reg_dirq_LC_4_23_1  (
            .in0(_gnd_net_),
            .in1(N__52470),
            .in2(_gnd_net_),
            .in3(N__20151),
            .lcout(\u0.dirq ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54153),
            .ce(),
            .sr(N__53332));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.DIOR_LC_4_23_2 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.DIOR_LC_4_23_2 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.DIOR_LC_4_23_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.DIOR_LC_4_23_2  (
            .in0(N__20042),
            .in1(N__20125),
            .in2(_gnd_net_),
            .in3(N__20116),
            .lcout(\u1.DMAdior ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54153),
            .ce(),
            .sr(N__53332));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.rci_LC_4_23_3 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.rci_LC_4_23_3 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.rci_LC_4_23_3 .LUT_INIT=16'b0000110000001110;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.rci_LC_4_23_3  (
            .in0(N__20062),
            .in1(N__20086),
            .in2(N__52629),
            .in3(N__20043),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.rci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54153),
            .ce(),
            .sr(N__53332));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qie_0_i_LC_4_23_4 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qie_0_i_LC_4_23_4 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qie_0_i_LC_4_23_4 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qie_0_i_LC_4_23_4  (
            .in0(N__52471),
            .in1(N__20085),
            .in2(_gnd_net_),
            .in3(N__20061),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qie_0_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.rci_LC_4_23_5 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.rci_LC_4_23_5 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.rci_LC_4_23_5 .LUT_INIT=16'b0000111000001100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.td_cnt.rci_LC_4_23_5  (
            .in0(N__19982),
            .in1(N__20044),
            .in2(N__52628),
            .in3(N__20026),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.rci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54153),
            .ce(),
            .sr(N__53332));
    defparam \u1.DMA_control.RxWr_LC_4_23_6 .C_ON=1'b0;
    defparam \u1.DMA_control.RxWr_LC_4_23_6 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.RxWr_LC_4_23_6 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \u1.DMA_control.RxWr_LC_4_23_6  (
            .in0(N__52472),
            .in1(N__20265),
            .in2(_gnd_net_),
            .in3(N__36331),
            .lcout(\u1.DMA_control.RxWrZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54153),
            .ce(),
            .sr(N__53332));
    defparam \u1.DMA_control.gen_DMA_req_iDMA_req_LC_4_23_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_req_iDMA_req_LC_4_23_7 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMA_req_iDMA_req_LC_4_23_7 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \u1.DMA_control.gen_DMA_req_iDMA_req_LC_4_23_7  (
            .in0(N__23404),
            .in1(N__20196),
            .in2(N__20224),
            .in3(N__20215),
            .lcout(DMA_req_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54153),
            .ce(),
            .sr(N__53332));
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_26_LC_4_24_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_26_LC_4_24_0 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_26_LC_4_24_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Txbuf.Q_26_LC_4_24_0  (
            .in0(N__23836),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44206),
            .lcout(\u1.DMA_control.TxbufQ_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54165),
            .ce(N__21164),
            .sr(N__53340));
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_3_LC_4_24_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_3_LC_4_24_1 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_3_LC_4_24_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Txbuf.Q_3_LC_4_24_1  (
            .in0(_gnd_net_),
            .in1(N__37369),
            .in2(_gnd_net_),
            .in3(N__23837),
            .lcout(\u1.DMA_control.TxbufQ_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54165),
            .ce(N__21164),
            .sr(N__53340));
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_18_LC_4_24_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_18_LC_4_24_2 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_18_LC_4_24_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Txbuf.Q_18_LC_4_24_2  (
            .in0(N__23834),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35020),
            .lcout(\u1.DMA_control.TxbufQ_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54165),
            .ce(N__21164),
            .sr(N__53340));
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_0_LC_4_24_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_0_LC_4_24_3 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_0_LC_4_24_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Txbuf.Q_0_LC_4_24_3  (
            .in0(N__49545),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23833),
            .lcout(\u1.DMA_control.TxbufQ_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54165),
            .ce(N__21164),
            .sr(N__53340));
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_7_LC_4_24_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_7_LC_4_24_4 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_7_LC_4_24_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Txbuf.Q_7_LC_4_24_4  (
            .in0(N__23839),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39657),
            .lcout(\u1.DMA_control.TxbufQ_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54165),
            .ce(N__21164),
            .sr(N__53340));
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_20_LC_4_24_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_20_LC_4_24_5 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_20_LC_4_24_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Txbuf.Q_20_LC_4_24_5  (
            .in0(N__34788),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23835),
            .lcout(\u1.DMA_control.TxbufQ_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54165),
            .ce(N__21164),
            .sr(N__53340));
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_4_LC_4_24_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_4_LC_4_24_6 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_4_LC_4_24_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Txbuf.Q_4_LC_4_24_6  (
            .in0(N__23838),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37226),
            .lcout(\u1.DMA_control.TxbufQ_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54165),
            .ce(N__21164),
            .sr(N__53340));
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_8_LC_4_24_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_8_LC_4_24_7 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_8_LC_4_24_7 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Txbuf.Q_8_LC_4_24_7  (
            .in0(N__54466),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23840),
            .lcout(\u1.DMA_control.TxbufQ_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54165),
            .ce(N__21164),
            .sr(N__53340));
    defparam \u1.PIO_control.gen_pingpong_pong_d_15_LC_4_25_0 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_pong_d_15_LC_4_25_0 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_pong_d_15_LC_4_25_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \u1.PIO_control.gen_pingpong_pong_d_15_LC_4_25_0  (
            .in0(N__34570),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\u1.PIO_control.pong_d_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54175),
            .ce(N__24882),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_pong_d_3_LC_4_25_2 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_pong_d_3_LC_4_25_2 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_pong_d_3_LC_4_25_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.PIO_control.gen_pingpong_pong_d_3_LC_4_25_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37370),
            .lcout(\u1.PIO_control.pong_d_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54175),
            .ce(N__24882),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_pong_d_4_LC_4_25_3 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_pong_d_4_LC_4_25_3 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_pong_d_4_LC_4_25_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \u1.PIO_control.gen_pingpong_pong_d_4_LC_4_25_3  (
            .in0(N__37245),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\u1.PIO_control.pong_d_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54175),
            .ce(N__24882),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_pong_d_5_LC_4_25_4 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_pong_d_5_LC_4_25_4 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_pong_d_5_LC_4_25_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \u1.PIO_control.gen_pingpong_pong_d_5_LC_4_25_4  (
            .in0(N__46303),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\u1.PIO_control.pong_d_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54175),
            .ce(N__24882),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_pong_d_6_LC_4_25_5 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_pong_d_6_LC_4_25_5 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_pong_d_6_LC_4_25_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \u1.PIO_control.gen_pingpong_pong_d_6_LC_4_25_5  (
            .in0(N__39487),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\u1.PIO_control.pong_d_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54175),
            .ce(N__24882),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_pong_d_7_LC_4_25_6 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_pong_d_7_LC_4_25_6 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_pong_d_7_LC_4_25_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.PIO_control.gen_pingpong_pong_d_7_LC_4_25_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39661),
            .lcout(\u1.PIO_control.pong_d_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54175),
            .ce(N__24882),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_pong_d_8_LC_4_25_7 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_pong_d_8_LC_4_25_7 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_pong_d_8_LC_4_25_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.PIO_control.gen_pingpong_pong_d_8_LC_4_25_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54467),
            .lcout(\u1.PIO_control.pong_d_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54175),
            .ce(N__24882),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_22_LC_4_26_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_22_LC_4_26_0 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_22_LC_4_26_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Txbuf.Q_22_LC_4_26_0  (
            .in0(_gnd_net_),
            .in1(N__38149),
            .in2(_gnd_net_),
            .in3(N__23878),
            .lcout(\u1.DMA_control.TxbufQ_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54187),
            .ce(N__21166),
            .sr(N__53353));
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_11_LC_4_26_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_11_LC_4_26_1 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_11_LC_4_26_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Txbuf.Q_11_LC_4_26_1  (
            .in0(N__23872),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43639),
            .lcout(\u1.DMA_control.TxbufQ_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54187),
            .ce(N__21166),
            .sr(N__53353));
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_10_LC_4_26_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_10_LC_4_26_2 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_10_LC_4_26_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Txbuf.Q_10_LC_4_26_2  (
            .in0(_gnd_net_),
            .in1(N__40122),
            .in2(_gnd_net_),
            .in3(N__23871),
            .lcout(\u1.DMA_control.TxbufQ_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54187),
            .ce(N__21166),
            .sr(N__53353));
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_19_LC_4_26_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_19_LC_4_26_3 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_19_LC_4_26_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Txbuf.Q_19_LC_4_26_3  (
            .in0(N__23877),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34333),
            .lcout(\u1.DMA_control.TxbufQ_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54187),
            .ce(N__21166),
            .sr(N__53353));
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_12_LC_4_26_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_12_LC_4_26_4 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_12_LC_4_26_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Txbuf.Q_12_LC_4_26_4  (
            .in0(_gnd_net_),
            .in1(N__36938),
            .in2(_gnd_net_),
            .in3(N__23873),
            .lcout(\u1.DMA_control.TxbufQ_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54187),
            .ce(N__21166),
            .sr(N__53353));
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_13_LC_4_26_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_13_LC_4_26_5 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_13_LC_4_26_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Txbuf.Q_13_LC_4_26_5  (
            .in0(N__23874),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34708),
            .lcout(\u1.DMA_control.TxbufQ_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54187),
            .ce(N__21166),
            .sr(N__53353));
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_14_LC_4_26_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_14_LC_4_26_6 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_14_LC_4_26_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Txbuf.Q_14_LC_4_26_6  (
            .in0(N__44006),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23875),
            .lcout(\u1.DMA_control.TxbufQ_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54187),
            .ce(N__21166),
            .sr(N__53353));
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_15_LC_4_26_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_15_LC_4_26_7 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_15_LC_4_26_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Txbuf.Q_15_LC_4_26_7  (
            .in0(N__23876),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34523),
            .lcout(\u1.DMA_control.TxbufQ_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54187),
            .ce(N__21166),
            .sr(N__53353));
    defparam \u1.PIO_control.gen_pingpong_pong_d_RNI7LHN_2_LC_4_27_1 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_pong_d_RNI7LHN_2_LC_4_27_1 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.gen_pingpong_pong_d_RNI7LHN_2_LC_4_27_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.PIO_control.gen_pingpong_pong_d_RNI7LHN_2_LC_4_27_1  (
            .in0(N__20323),
            .in1(N__21184),
            .in2(_gnd_net_),
            .in3(N__26919),
            .lcout(),
            .ltout(\u1.N_1428_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DDo_2_LC_4_27_2 .C_ON=1'b0;
    defparam \u1.DDo_2_LC_4_27_2 .SEQ_MODE=4'b1010;
    defparam \u1.DDo_2_LC_4_27_2 .LUT_INIT=16'b0101000001000100;
    LogicCell40 \u1.DDo_2_LC_4_27_2  (
            .in0(N__52630),
            .in1(N__25819),
            .in2(N__20314),
            .in3(N__36740),
            .lcout(dd_pad_o_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54198),
            .ce(),
            .sr(N__53359));
    defparam \u1.PIO_control.gen_pingpong_pong_d_RNI9NHN_3_LC_4_27_3 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_pong_d_RNI9NHN_3_LC_4_27_3 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.gen_pingpong_pong_d_RNI9NHN_3_LC_4_27_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.PIO_control.gen_pingpong_pong_d_RNI9NHN_3_LC_4_27_3  (
            .in0(N__20296),
            .in1(N__21178),
            .in2(_gnd_net_),
            .in3(N__26920),
            .lcout(),
            .ltout(\u1.N_1449_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DDo_3_LC_4_27_4 .C_ON=1'b0;
    defparam \u1.DDo_3_LC_4_27_4 .SEQ_MODE=4'b1010;
    defparam \u1.DDo_3_LC_4_27_4 .LUT_INIT=16'b0101000001000100;
    LogicCell40 \u1.DDo_3_LC_4_27_4  (
            .in0(N__52631),
            .in1(N__25747),
            .in2(N__20287),
            .in3(N__36741),
            .lcout(dd_pad_o_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54198),
            .ce(),
            .sr(N__53359));
    defparam \u1.PIO_control.gen_pingpong_pong_d_RNIF6CJ_15_LC_4_27_5 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_pong_d_RNIF6CJ_15_LC_4_27_5 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.gen_pingpong_pong_d_RNIF6CJ_15_LC_4_27_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.PIO_control.gen_pingpong_pong_d_RNIF6CJ_15_LC_4_27_5  (
            .in0(N__20602),
            .in1(N__21190),
            .in2(_gnd_net_),
            .in3(N__26918),
            .lcout(\u1.N_1436 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_pong_d_RNIBPHN_4_LC_4_27_7 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_pong_d_RNIBPHN_4_LC_4_27_7 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.gen_pingpong_pong_d_RNIBPHN_4_LC_4_27_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.PIO_control.gen_pingpong_pong_d_RNIBPHN_4_LC_4_27_7  (
            .in0(N__20593),
            .in1(N__21172),
            .in2(_gnd_net_),
            .in3(N__26917),
            .lcout(\u1.N_1429 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DDo_15_LC_4_28_4 .C_ON=1'b0;
    defparam \u1.DDo_15_LC_4_28_4 .SEQ_MODE=4'b1010;
    defparam \u1.DDo_15_LC_4_28_4 .LUT_INIT=16'b0000111000000010;
    LogicCell40 \u1.DDo_15_LC_4_28_4  (
            .in0(N__25411),
            .in1(N__36742),
            .in2(N__52707),
            .in3(N__20584),
            .lcout(dd_pad_o_c_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54211),
            .ce(),
            .sr(N__53368));
    defparam \u1.PIO_control.PIO_access_control.q_11_LC_5_15_6 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.q_11_LC_5_15_6 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.q_11_LC_5_15_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \u1.PIO_control.PIO_access_control.q_11_LC_5_15_6  (
            .in0(N__33111),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(PIOq_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54133),
            .ce(N__45908),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_RNIGUSK_7_LC_5_16_0 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_RNIGUSK_7_LC_5_16_0 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_RNIGUSK_7_LC_5_16_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_RNIGUSK_7_LC_5_16_0  (
            .in0(N__20563),
            .in1(N__20536),
            .in2(N__20512),
            .in3(N__20485),
            .lcout(),
            .ltout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.val_c8_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_RNI5EI41_1_LC_5_16_1 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_RNI5EI41_1_LC_5_16_1 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_RNI5EI41_1_LC_5_16_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.eoc_cnt.cnt.Qi_RNI5EI41_1_LC_5_16_1  (
            .in0(N__20461),
            .in1(N__20437),
            .in2(N__20413),
            .in3(N__20410),
            .lcout(),
            .ltout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.val_c8_0_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.busy_LC_5_16_2 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.busy_LC_5_16_2 .SEQ_MODE=4'b1010;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.busy_LC_5_16_2 .LUT_INIT=16'b0011001100110001;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.busy_LC_5_16_2  (
            .in0(N__20386),
            .in1(N__20329),
            .in2(N__20365),
            .in3(N__20362),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.busyZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54129),
            .ce(),
            .sr(N__53307));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.busy_RNO_0_LC_5_16_3 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.busy_RNO_0_LC_5_16_3 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.busy_RNO_0_LC_5_16_3 .LUT_INIT=16'b1111000011110001;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.busy_RNO_0_LC_5_16_3  (
            .in0(N__20786),
            .in1(N__20645),
            .in2(N__52194),
            .in3(N__20630),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.busy_3_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.hold_go_LC_5_16_4 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.hold_go_LC_5_16_4 .SEQ_MODE=4'b1010;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.hold_go_LC_5_16_4 .LUT_INIT=16'b0010001000100000;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.hold_go_LC_5_16_4  (
            .in0(N__20632),
            .in1(N__52007),
            .in2(N__20650),
            .in3(N__20788),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.hold_goZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54129),
            .ce(),
            .sr(N__53307));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qilde_i_o3_LC_5_16_5 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qilde_i_o3_LC_5_16_5 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qilde_i_o3_LC_5_16_5 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qilde_i_o3_LC_5_16_5  (
            .in0(N__20785),
            .in1(N__20644),
            .in2(_gnd_net_),
            .in3(N__20629),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.N_1371 ),
            .ltout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.N_1371_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qilde_i_LC_5_16_6 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qilde_i_LC_5_16_6 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qilde_i_LC_5_16_6 .LUT_INIT=16'b1111111111001111;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qilde_i_LC_5_16_6  (
            .in0(_gnd_net_),
            .in1(N__52011),
            .in2(N__20653),
            .in3(N__23252),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.N_1071 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_1_sqmuxa_i_1_LC_5_16_7 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_1_sqmuxa_i_1_LC_5_16_7 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_1_sqmuxa_i_1_LC_5_16_7 .LUT_INIT=16'b1111000011111110;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_1_sqmuxa_i_1_LC_5_16_7  (
            .in0(N__20787),
            .in1(N__20646),
            .in2(N__52195),
            .in3(N__20631),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.N_1073 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_ping_d_6_LC_5_17_0 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_ping_d_6_LC_5_17_0 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_ping_d_6_LC_5_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.PIO_control.gen_pingpong_ping_d_6_LC_5_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39476),
            .lcout(\u1.PIO_control.ping_d_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54117),
            .ce(N__25086),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_ping_d_7_LC_5_17_1 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_ping_d_7_LC_5_17_1 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_ping_d_7_LC_5_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.PIO_control.gen_pingpong_ping_d_7_LC_5_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39649),
            .lcout(\u1.PIO_control.ping_d_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54117),
            .ce(N__25086),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_ping_d_8_LC_5_17_2 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_ping_d_8_LC_5_17_2 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_ping_d_8_LC_5_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.PIO_control.gen_pingpong_ping_d_8_LC_5_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54475),
            .lcout(\u1.PIO_control.ping_d_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54117),
            .ce(N__25086),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_ping_d_9_LC_5_17_3 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_ping_d_9_LC_5_17_3 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_ping_d_9_LC_5_17_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \u1.PIO_control.gen_pingpong_ping_d_9_LC_5_17_3  (
            .in0(N__35994),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\u1.PIO_control.ping_d_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54117),
            .ce(N__25086),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_ping_we_LC_5_17_4 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_ping_we_LC_5_17_4 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_ping_we_LC_5_17_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \u1.PIO_control.gen_pingpong_ping_we_LC_5_17_4  (
            .in0(N__21961),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\u1.PIO_control.ping_we ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54117),
            .ce(N__25086),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNI84QB_7_LC_5_18_0 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNI84QB_7_LC_5_18_0 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNI84QB_7_LC_5_18_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNI84QB_7_LC_5_18_0  (
            .in0(N__23025),
            .in1(N__23046),
            .in2(N__24784),
            .in3(N__23109),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.val_c8_0_4 ),
            .ltout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.val_c8_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNIAJPR_0_LC_5_18_1 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNIAJPR_0_LC_5_18_1 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNIAJPR_0_LC_5_18_1 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNIAJPR_0_LC_5_18_1  (
            .in0(N__21366),
            .in1(N__23238),
            .in2(N__20755),
            .in3(N__26069),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.T1done_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_1_sqmuxa_i_x0_LC_5_18_2 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_1_sqmuxa_i_x0_LC_5_18_2 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_1_sqmuxa_i_x0_LC_5_18_2 .LUT_INIT=16'b1100110011011100;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_1_sqmuxa_i_x0_LC_5_18_2  (
            .in0(N__26068),
            .in1(N__52200),
            .in2(N__23251),
            .in3(N__21365),
            .lcout(),
            .ltout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_1_sqmuxa_i_xZ0Z0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_1_sqmuxa_i_ns_LC_5_18_3 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_1_sqmuxa_i_ns_LC_5_18_3 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_1_sqmuxa_i_ns_LC_5_18_3 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_1_sqmuxa_i_ns_LC_5_18_3  (
            .in0(N__52199),
            .in1(_gnd_net_),
            .in2(N__20752),
            .in3(N__20749),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_1_sqmuxa_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev1_Td_RNIORB59_0_LC_5_18_5 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Td_RNIORB59_0_LC_5_18_5 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev1_Td_RNIORB59_0_LC_5_18_5 .LUT_INIT=16'b1111111011101110;
    LogicCell40 \u0.DMA_dev1_Td_RNIORB59_0_LC_5_18_5  (
            .in0(N__31153),
            .in1(N__31462),
            .in2(N__21430),
            .in3(N__46602),
            .lcout(\u0.dat_o_0_0_6_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.iordy_done_LC_5_18_6 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.iordy_done_LC_5_18_6 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.iordy_done_LC_5_18_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.iordy_done_LC_5_18_6  (
            .in0(_gnd_net_),
            .in1(N__20734),
            .in2(_gnd_net_),
            .in3(N__26545),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.iordy_done_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DA_2_LC_5_19_0 .C_ON=1'b0;
    defparam \u1.DA_2_LC_5_19_0 .SEQ_MODE=4'b1010;
    defparam \u1.DA_2_LC_5_19_0 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \u1.DA_2_LC_5_19_0  (
            .in0(N__26233),
            .in1(N__26855),
            .in2(N__52426),
            .in3(N__26253),
            .lcout(da_pad_o_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54134),
            .ce(),
            .sr(N__53320));
    defparam \u1.PIO_control.SelDev_RNO_1_LC_5_19_1 .C_ON=1'b0;
    defparam \u1.PIO_control.SelDev_RNO_1_LC_5_19_1 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.SelDev_RNO_1_LC_5_19_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.PIO_control.SelDev_RNO_1_LC_5_19_1  (
            .in0(N__26853),
            .in1(N__26252),
            .in2(_gnd_net_),
            .in3(N__26232),
            .lcout(\u1.PIO_control.un3_idone_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.hT2done_RNIHFNK1_LC_5_19_2 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.hT2done_RNIHFNK1_LC_5_19_2 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.hT2done_RNIHFNK1_LC_5_19_2 .LUT_INIT=16'b1010111110101110;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.hT2done_RNIHFNK1_LC_5_19_2  (
            .in0(N__24511),
            .in1(N__24676),
            .in2(N__24603),
            .in3(N__24688),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.N_1358 ),
            .ltout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.N_1358_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.rci_LC_5_19_3 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.rci_LC_5_19_3 .SEQ_MODE=4'b1010;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.rci_LC_5_19_3 .LUT_INIT=16'b0100010100000101;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.rci_LC_5_19_3  (
            .in0(N__52205),
            .in1(N__20673),
            .in2(N__20683),
            .in3(N__26295),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.rciZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54134),
            .ce(),
            .sr(N__53320));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNI01HO_7_LC_5_19_4 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNI01HO_7_LC_5_19_4 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNI01HO_7_LC_5_19_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.dhold_cnt.cnt.Qi_RNI01HO_7_LC_5_19_4  (
            .in0(N__20884),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20851),
            .lcout(\u1.PIOdone_i ),
            .ltout(\u1.PIOdone_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIOgo_LC_5_19_5 .C_ON=1'b0;
    defparam \u1.PIOgo_LC_5_19_5 .SEQ_MODE=4'b1010;
    defparam \u1.PIOgo_LC_5_19_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \u1.PIOgo_LC_5_19_5  (
            .in0(N__20829),
            .in1(N__52204),
            .in2(N__20812),
            .in3(N__20809),
            .lcout(\u1.PIOgoZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54134),
            .ce(),
            .sr(N__53320));
    defparam \u1.PIO_control.gen_pingpong_pong_valid_LC_5_19_6 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_pong_valid_LC_5_19_6 .SEQ_MODE=4'b1010;
    defparam \u1.PIO_control.gen_pingpong_pong_valid_LC_5_19_6 .LUT_INIT=16'b1110111011100000;
    LogicCell40 \u1.PIO_control.gen_pingpong_pong_valid_LC_5_19_6  (
            .in0(N__26297),
            .in1(N__26856),
            .in2(N__21091),
            .in3(N__20968),
            .lcout(u1_PIO_control_gen_pingpong_pong_valid),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54134),
            .ce(),
            .sr(N__53320));
    defparam \u1.PIO_control.gen_pingpong_ping_valid_LC_5_19_7 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_ping_valid_LC_5_19_7 .SEQ_MODE=4'b1010;
    defparam \u1.PIO_control.gen_pingpong_ping_valid_LC_5_19_7 .LUT_INIT=16'b1111110001010100;
    LogicCell40 \u1.PIO_control.gen_pingpong_ping_valid_LC_5_19_7  (
            .in0(N__26854),
            .in1(N__21202),
            .in2(N__20764),
            .in3(N__26296),
            .lcout(u1_PIO_control_gen_pingpong_ping_valid),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54134),
            .ce(),
            .sr(N__53320));
    defparam \u0.CtrlReg_RNI0DNL2_4_LC_5_20_0 .C_ON=1'b0;
    defparam \u0.CtrlReg_RNI0DNL2_4_LC_5_20_0 .SEQ_MODE=4'b0000;
    defparam \u0.CtrlReg_RNI0DNL2_4_LC_5_20_0 .LUT_INIT=16'b1000000011000000;
    LogicCell40 \u0.CtrlReg_RNI0DNL2_4_LC_5_20_0  (
            .in0(N__23511),
            .in1(N__46594),
            .in2(N__21079),
            .in3(N__27744),
            .lcout(\u0.N_1969 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_ping_valid_RNIOA821_LC_5_20_1 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_ping_valid_RNIOA821_LC_5_20_1 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.gen_pingpong_ping_valid_RNIOA821_LC_5_20_1 .LUT_INIT=16'b0011001110111011;
    LogicCell40 \u1.PIO_control.gen_pingpong_ping_valid_RNIOA821_LC_5_20_1  (
            .in0(N__27743),
            .in1(N__21068),
            .in2(_gnd_net_),
            .in3(N__23510),
            .lcout(),
            .ltout(N_468_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.gen_bc_dec_store_pp_full_LC_5_20_2 .C_ON=1'b0;
    defparam \u0.gen_bc_dec_store_pp_full_LC_5_20_2 .SEQ_MODE=4'b1000;
    defparam \u0.gen_bc_dec_store_pp_full_LC_5_20_2 .LUT_INIT=16'b0000111100001110;
    LogicCell40 \u0.gen_bc_dec_store_pp_full_LC_5_20_2  (
            .in0(N__21457),
            .in1(N__21497),
            .in2(N__20770),
            .in3(N__21701),
            .lcout(u0_gen_bc_dec_store_pp_full),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54141),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_gen_sel_strb_dsel_3_0_a2_1_LC_5_20_3 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_gen_sel_strb_dsel_3_0_a2_1_LC_5_20_3 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.gen_pingpong_gen_sel_strb_dsel_3_0_a2_1_LC_5_20_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \u1.PIO_control.gen_pingpong_gen_sel_strb_dsel_3_0_a2_1_LC_5_20_3  (
            .in0(N__52254),
            .in1(N__21456),
            .in2(N__21706),
            .in3(N__21483),
            .lcout(\u1.PIO_control.N_2409 ),
            .ltout(\u1.PIO_control.N_2409_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_ping_valid_RNO_0_LC_5_20_4 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_ping_valid_RNO_0_LC_5_20_4 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.gen_pingpong_ping_valid_RNO_0_LC_5_20_4 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \u1.PIO_control.gen_pingpong_ping_valid_RNO_0_LC_5_20_4  (
            .in0(N__21137),
            .in1(N__23151),
            .in2(N__20767),
            .in3(N__38340),
            .lcout(\u1.PIO_control.ping_valid_3_0_a2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_pong_valid_RNO_1_LC_5_20_5 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_pong_valid_RNO_1_LC_5_20_5 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.gen_pingpong_pong_valid_RNO_1_LC_5_20_5 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \u1.PIO_control.gen_pingpong_pong_valid_RNO_1_LC_5_20_5  (
            .in0(N__38339),
            .in1(N__21138),
            .in2(N__23155),
            .in3(N__23166),
            .lcout(\u1.PIO_control.pong_valid_3_0_a2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.gen_regs_un1_ena_i_0_a2_sx_LC_5_20_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.gen_regs_un1_ena_i_0_a2_sx_LC_5_20_6 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.gen_regs_un1_ena_i_0_a2_sx_LC_5_20_6 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.gen_regs_un1_ena_i_0_a2_sx_LC_5_20_6  (
            .in0(N__47262),
            .in1(N__21955),
            .in2(_gnd_net_),
            .in3(N__20962),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.un1_ena_i_0_a2_sx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_wpp_RNIKPCQ2_LC_5_20_7 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_wpp_RNIKPCQ2_LC_5_20_7 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.gen_pingpong_wpp_RNIKPCQ2_LC_5_20_7 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \u1.PIO_control.gen_pingpong_wpp_RNIKPCQ2_LC_5_20_7  (
            .in0(N__21705),
            .in1(N__21643),
            .in2(N__23526),
            .in3(N__21136),
            .lcout(\u1.PIO_control.ping_we_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_iack_RNO_3_LC_5_21_0 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_iack_RNO_3_LC_5_21_0 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.gen_pingpong_iack_RNO_3_LC_5_21_0 .LUT_INIT=16'b0001101100010001;
    LogicCell40 \u1.PIO_control.gen_pingpong_iack_RNO_3_LC_5_21_0  (
            .in0(N__26890),
            .in1(N__21037),
            .in2(N__23525),
            .in3(N__23469),
            .lcout(),
            .ltout(\u1.PIO_control.iack_7_u_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_iack_RNO_0_LC_5_21_1 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_iack_RNO_0_LC_5_21_1 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.gen_pingpong_iack_RNO_0_LC_5_21_1 .LUT_INIT=16'b1100000000000100;
    LogicCell40 \u1.PIO_control.gen_pingpong_iack_RNO_0_LC_5_21_1  (
            .in0(N__21075),
            .in1(N__20907),
            .in2(N__20950),
            .in3(N__26891),
            .lcout(),
            .ltout(\u1.PIO_control.iack_7_u_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_iack_LC_5_21_2 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_iack_LC_5_21_2 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_iack_LC_5_21_2 .LUT_INIT=16'b1111010111110100;
    LogicCell40 \u1.PIO_control.gen_pingpong_iack_LC_5_21_2  (
            .in0(N__20908),
            .in1(N__20890),
            .in2(N__20947),
            .in3(N__20899),
            .lcout(u1_PIO_control_gen_pingpong_iack),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54148),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_pong_we_RNILH6S_LC_5_21_3 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_pong_we_RNILH6S_LC_5_21_3 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.gen_pingpong_pong_we_RNILH6S_LC_5_21_3 .LUT_INIT=16'b0011111101011111;
    LogicCell40 \u1.PIO_control.gen_pingpong_pong_we_RNILH6S_LC_5_21_3  (
            .in0(N__20944),
            .in1(N__20926),
            .in2(N__27745),
            .in3(N__26889),
            .lcout(\u1.PIO_control.N_1362 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_iack_RNO_1_LC_5_21_4 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_iack_RNO_1_LC_5_21_4 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.gen_pingpong_iack_RNO_1_LC_5_21_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \u1.PIO_control.gen_pingpong_iack_RNO_1_LC_5_21_4  (
            .in0(N__23514),
            .in1(N__21135),
            .in2(N__21950),
            .in3(N__23470),
            .lcout(\u1.PIO_control.iack_7_u_0_a2_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_iack_RNO_2_LC_5_21_5 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_iack_RNO_2_LC_5_21_5 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.gen_pingpong_iack_RNO_2_LC_5_21_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \u1.PIO_control.gen_pingpong_iack_RNO_2_LC_5_21_5  (
            .in0(N__21074),
            .in1(N__21129),
            .in2(N__21951),
            .in3(N__21036),
            .lcout(\u1.PIO_control.iack_7_u_0_a2_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_dsel_RNO_0_LC_5_21_6 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_dsel_RNO_0_LC_5_21_6 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.gen_pingpong_dsel_RNO_0_LC_5_21_6 .LUT_INIT=16'b0100010001110111;
    LogicCell40 \u1.PIO_control.gen_pingpong_dsel_RNO_0_LC_5_21_6  (
            .in0(N__23513),
            .in1(N__21134),
            .in2(_gnd_net_),
            .in3(N__21073),
            .lcout(\u1.PIO_control.dsel_3_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_ping_valid_RNIBNER_LC_5_21_7 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_ping_valid_RNIBNER_LC_5_21_7 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.gen_pingpong_ping_valid_RNIBNER_LC_5_21_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.PIO_control.gen_pingpong_ping_valid_RNIBNER_LC_5_21_7  (
            .in0(N__21072),
            .in1(N__23512),
            .in2(_gnd_net_),
            .in3(N__26888),
            .lcout(\u1.N_1359 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_gen_pp_rpp_2_i_0_LC_5_22_0 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_gen_pp_rpp_2_i_0_LC_5_22_0 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.gen_pingpong_gen_pp_rpp_2_i_0_LC_5_22_0 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \u1.PIO_control.gen_pingpong_gen_pp_rpp_2_i_0_LC_5_22_0  (
            .in0(N__52444),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27742),
            .lcout(\u1.PIO_control.rpp_2_i_0 ),
            .ltout(\u1.PIO_control.rpp_2_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_wpp_LC_5_22_1 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_wpp_LC_5_22_1 .SEQ_MODE=4'b1010;
    defparam \u1.PIO_control.gen_pingpong_wpp_LC_5_22_1 .LUT_INIT=16'b0000011000001010;
    LogicCell40 \u1.PIO_control.gen_pingpong_wpp_LC_5_22_1  (
            .in0(N__21130),
            .in1(N__21959),
            .in2(N__21142),
            .in3(N__21681),
            .lcout(\u1.PIO_control.wpp ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54154),
            .ce(),
            .sr(N__53333));
    defparam \u1.PIO_control.gen_pingpong_wpp_RNIQ9MF2_LC_5_22_2 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_wpp_RNIQ9MF2_LC_5_22_2 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.gen_pingpong_wpp_RNIQ9MF2_LC_5_22_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \u1.PIO_control.gen_pingpong_wpp_RNIQ9MF2_LC_5_22_2  (
            .in0(N__21076),
            .in1(N__21693),
            .in2(N__21139),
            .in3(N__21644),
            .lcout(\u1.PIO_control.pong_we_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_pong_valid_RNO_0_LC_5_22_3 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_pong_valid_RNO_0_LC_5_22_3 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.gen_pingpong_pong_valid_RNO_0_LC_5_22_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \u1.PIO_control.gen_pingpong_pong_valid_RNO_0_LC_5_22_3  (
            .in0(_gnd_net_),
            .in1(N__52445),
            .in2(_gnd_net_),
            .in3(N__21077),
            .lcout(\u1.PIO_control.pong_valid_3_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_dpong_valid_LC_5_22_4 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_dpong_valid_LC_5_22_4 .SEQ_MODE=4'b1010;
    defparam \u1.PIO_control.gen_pingpong_dpong_valid_LC_5_22_4 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \u1.PIO_control.gen_pingpong_dpong_valid_LC_5_22_4  (
            .in0(N__21078),
            .in1(_gnd_net_),
            .in2(N__52610),
            .in3(_gnd_net_),
            .lcout(\u1.PIO_control.dpong_valid ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54154),
            .ce(),
            .sr(N__53333));
    defparam \u1.DMAgo_LC_5_22_5 .C_ON=1'b0;
    defparam \u1.DMAgo_LC_5_22_5 .SEQ_MODE=4'b1010;
    defparam \u1.DMAgo_LC_5_22_5 .LUT_INIT=16'b1111010000000000;
    LogicCell40 \u1.DMAgo_LC_5_22_5  (
            .in0(N__23662),
            .in1(N__23335),
            .in2(N__23317),
            .in3(N__21385),
            .lcout(\u1.DMAgoZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54154),
            .ce(),
            .sr(N__53333));
    defparam \u1.DMA_control.TxRd_LC_5_22_6 .C_ON=1'b0;
    defparam \u1.DMA_control.TxRd_LC_5_22_6 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.TxRd_LC_5_22_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \u1.DMA_control.TxRd_LC_5_22_6  (
            .in0(N__52440),
            .in1(N__21007),
            .in2(_gnd_net_),
            .in3(N__23660),
            .lcout(\u1.DMA_control.TxRdZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54154),
            .ce(),
            .sr(N__53333));
    defparam \u1.DMA_control.gen_DMA_req_hgo_LC_5_22_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_req_hgo_LC_5_22_7 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMA_req_hgo_LC_5_22_7 .LUT_INIT=16'b0000000011111000;
    LogicCell40 \u1.DMA_control.gen_DMA_req_hgo_LC_5_22_7  (
            .in0(N__23661),
            .in1(N__20980),
            .in2(N__21015),
            .in3(N__20986),
            .lcout(\u1.DMA_control.hgo ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54154),
            .ce(),
            .sr(N__53333));
    defparam \u0.PIO_dport1_Teoc_3_LC_5_23_5 .C_ON=1'b0;
    defparam \u0.PIO_dport1_Teoc_3_LC_5_23_5 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport1_Teoc_3_LC_5_23_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.PIO_dport1_Teoc_3_LC_5_23_5  (
            .in0(N__37687),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52450),
            .lcout(PIO_dport1_Teoc_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54166),
            .ce(N__39208),
            .sr(N__53341));
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_23_LC_5_24_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_23_LC_5_24_0 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_23_LC_5_24_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Txbuf.Q_23_LC_5_24_0  (
            .in0(N__44819),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23827),
            .lcout(\u1.DMA_control.TxbufQ_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54176),
            .ce(N__21165),
            .sr(N__53347));
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_24_LC_5_24_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_24_LC_5_24_1 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_24_LC_5_24_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Txbuf.Q_24_LC_5_24_1  (
            .in0(N__23828),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39879),
            .lcout(\u1.DMA_control.TxbufQ_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54176),
            .ce(N__21165),
            .sr(N__53347));
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_17_LC_5_24_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_17_LC_5_24_2 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_17_LC_5_24_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Txbuf.Q_17_LC_5_24_2  (
            .in0(N__45117),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23826),
            .lcout(\u1.DMA_control.TxbufQ_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54176),
            .ce(N__21165),
            .sr(N__53347));
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_27_LC_5_24_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_27_LC_5_24_3 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_27_LC_5_24_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Txbuf.Q_27_LC_5_24_3  (
            .in0(N__23829),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37674),
            .lcout(\u1.DMA_control.TxbufQ_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54176),
            .ce(N__21165),
            .sr(N__53347));
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_16_LC_5_24_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_16_LC_5_24_4 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_16_LC_5_24_4 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Txbuf.Q_16_LC_5_24_4  (
            .in0(N__40994),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23825),
            .lcout(\u1.DMA_control.TxbufQ_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54176),
            .ce(N__21165),
            .sr(N__53347));
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_28_LC_5_24_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_28_LC_5_24_5 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_28_LC_5_24_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Txbuf.Q_28_LC_5_24_5  (
            .in0(N__23830),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46150),
            .lcout(\u1.DMA_control.TxbufQ_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54176),
            .ce(N__21165),
            .sr(N__53347));
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_9_LC_5_24_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_9_LC_5_24_6 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_9_LC_5_24_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Txbuf.Q_9_LC_5_24_6  (
            .in0(N__36017),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23832),
            .lcout(\u1.DMA_control.TxbufQ_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54176),
            .ce(N__21165),
            .sr(N__53347));
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_29_LC_5_24_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_29_LC_5_24_7 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.Q_29_LC_5_24_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Txbuf.Q_29_LC_5_24_7  (
            .in0(N__23831),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49348),
            .lcout(\u1.DMA_control.TxbufQ_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54176),
            .ce(N__21165),
            .sr(N__53347));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__29_LC_5_25_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__29_LC_5_25_0 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__29_LC_5_25_0 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__29_LC_5_25_0  (
            .in0(N__42974),
            .in1(N__33594),
            .in2(N__33461),
            .in3(_gnd_net_),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54188),
            .ce(N__41853),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__6_LC_5_25_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__6_LC_5_25_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__6_LC_5_25_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__6_LC_5_25_1  (
            .in0(N__32830),
            .in1(N__32706),
            .in2(_gnd_net_),
            .in3(N__42975),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54188),
            .ce(N__41853),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_ping_valid_RNIE0EK_LC_5_25_2 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_ping_valid_RNIE0EK_LC_5_25_2 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.gen_pingpong_ping_valid_RNIE0EK_LC_5_25_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u1.PIO_control.gen_pingpong_ping_valid_RNIE0EK_LC_5_25_2  (
            .in0(N__52449),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23524),
            .lcout(\u1.PIO_control.dping_valid_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_ping_d_12_LC_5_26_0 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_ping_d_12_LC_5_26_0 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_ping_d_12_LC_5_26_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \u1.PIO_control.gen_pingpong_ping_d_12_LC_5_26_0  (
            .in0(N__36961),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\u1.PIO_control.ping_d_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54199),
            .ce(N__25085),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_ping_d_13_LC_5_26_1 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_ping_d_13_LC_5_26_1 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_ping_d_13_LC_5_26_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \u1.PIO_control.gen_pingpong_ping_d_13_LC_5_26_1  (
            .in0(N__34699),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\u1.PIO_control.ping_d_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54199),
            .ce(N__25085),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_ping_d_14_LC_5_26_2 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_ping_d_14_LC_5_26_2 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_ping_d_14_LC_5_26_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.PIO_control.gen_pingpong_ping_d_14_LC_5_26_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44028),
            .lcout(\u1.PIO_control.ping_d_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54199),
            .ce(N__25085),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_ping_d_15_LC_5_26_3 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_ping_d_15_LC_5_26_3 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_ping_d_15_LC_5_26_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.PIO_control.gen_pingpong_ping_d_15_LC_5_26_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34569),
            .lcout(\u1.PIO_control.ping_d_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54199),
            .ce(N__25085),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_ping_d_2_LC_5_26_4 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_ping_d_2_LC_5_26_4 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_ping_d_2_LC_5_26_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.PIO_control.gen_pingpong_ping_d_2_LC_5_26_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34271),
            .lcout(\u1.PIO_control.ping_d_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54199),
            .ce(N__25085),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_ping_d_3_LC_5_26_5 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_ping_d_3_LC_5_26_5 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_ping_d_3_LC_5_26_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.PIO_control.gen_pingpong_ping_d_3_LC_5_26_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37377),
            .lcout(\u1.PIO_control.ping_d_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54199),
            .ce(N__25085),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_ping_d_4_LC_5_26_6 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_ping_d_4_LC_5_26_6 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_ping_d_4_LC_5_26_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.PIO_control.gen_pingpong_ping_d_4_LC_5_26_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37246),
            .lcout(\u1.PIO_control.ping_d_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54199),
            .ce(N__25085),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_ping_d_5_LC_5_26_7 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_ping_d_5_LC_5_26_7 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_ping_d_5_LC_5_26_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.PIO_control.gen_pingpong_ping_d_5_LC_5_26_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46302),
            .lcout(\u1.PIO_control.ping_d_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54199),
            .ce(N__25085),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_0_LC_5_27_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_0_LC_5_27_0 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_0_LC_5_27_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDlw_0_LC_5_27_0  (
            .in0(N__22629),
            .in1(N__22608),
            .in2(_gnd_net_),
            .in3(N__42952),
            .lcout(\u1.DMA_control.writeDlw_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54212),
            .ce(N__25549),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_1_LC_5_27_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_1_LC_5_27_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_1_LC_5_27_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDlw_1_LC_5_27_1  (
            .in0(N__42951),
            .in1(N__23922),
            .in2(_gnd_net_),
            .in3(N__23956),
            .lcout(\u1.DMA_control.writeDlw_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54212),
            .ce(N__25549),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_3_LC_5_27_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_3_LC_5_27_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_3_LC_5_27_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDlw_3_LC_5_27_2  (
            .in0(N__22410),
            .in1(N__22090),
            .in2(_gnd_net_),
            .in3(N__42955),
            .lcout(\u1.DMA_control.writeDlw_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54212),
            .ce(N__25549),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_11_LC_5_27_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_11_LC_5_27_3 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_11_LC_5_27_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDlw_11_LC_5_27_3  (
            .in0(N__42948),
            .in1(N__25761),
            .in2(_gnd_net_),
            .in3(N__25803),
            .lcout(\u1.DMA_control.writeDlw_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54212),
            .ce(N__25549),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_12_LC_5_27_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_12_LC_5_27_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_12_LC_5_27_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDlw_12_LC_5_27_4  (
            .in0(N__25317),
            .in1(N__25728),
            .in2(_gnd_net_),
            .in3(N__42953),
            .lcout(\u1.DMA_control.writeDlw_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54212),
            .ce(N__25549),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_13_LC_5_27_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_13_LC_5_27_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_13_LC_5_27_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDlw_13_LC_5_27_5  (
            .in0(N__42949),
            .in1(_gnd_net_),
            .in2(N__22291),
            .in3(N__22575),
            .lcout(\u1.DMA_control.writeDlw_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54212),
            .ce(N__25549),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_14_LC_5_27_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_14_LC_5_27_6 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_14_LC_5_27_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDlw_14_LC_5_27_6  (
            .in0(N__22719),
            .in1(N__22242),
            .in2(_gnd_net_),
            .in3(N__42954),
            .lcout(\u1.DMA_control.writeDlw_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54212),
            .ce(N__25549),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_15_LC_5_27_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_15_LC_5_27_7 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_15_LC_5_27_7 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDlw_15_LC_5_27_7  (
            .in0(N__42950),
            .in1(_gnd_net_),
            .in2(N__22687),
            .in3(N__22653),
            .lcout(\u1.DMA_control.writeDlw_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54212),
            .ce(N__25549),
            .sr(_gnd_net_));
    defparam \u1.DDo_4_LC_5_28_5 .C_ON=1'b0;
    defparam \u1.DDo_4_LC_5_28_5 .SEQ_MODE=4'b1010;
    defparam \u1.DDo_4_LC_5_28_5 .LUT_INIT=16'b0000111000000010;
    LogicCell40 \u1.DDo_4_LC_5_28_5  (
            .in0(N__25306),
            .in1(N__36777),
            .in2(N__52708),
            .in3(N__24987),
            .lcout(dd_pad_o_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54226),
            .ce(),
            .sr(N__53378));
    defparam \u1.PIO_control.gen_pingpong_pong_d_RNIDRHN_5_LC_5_29_1 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_pong_d_RNIDRHN_5_LC_5_29_1 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.gen_pingpong_pong_d_RNIDRHN_5_LC_5_29_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.PIO_control.gen_pingpong_pong_d_RNIDRHN_5_LC_5_29_1  (
            .in0(N__21352),
            .in1(N__21340),
            .in2(_gnd_net_),
            .in3(N__26895),
            .lcout(),
            .ltout(\u1.N_1430_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DDo_5_LC_5_29_2 .C_ON=1'b0;
    defparam \u1.DDo_5_LC_5_29_2 .SEQ_MODE=4'b1010;
    defparam \u1.DDo_5_LC_5_29_2 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \u1.DDo_5_LC_5_29_2  (
            .in0(N__36775),
            .in1(N__52627),
            .in2(N__21331),
            .in3(N__22552),
            .lcout(dd_pad_o_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54237),
            .ce(),
            .sr(N__53383));
    defparam \u1.PIO_control.gen_pingpong_pong_d_RNIFTHN_6_LC_5_29_3 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_pong_d_RNIFTHN_6_LC_5_29_3 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.gen_pingpong_pong_d_RNIFTHN_6_LC_5_29_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.PIO_control.gen_pingpong_pong_d_RNIFTHN_6_LC_5_29_3  (
            .in0(N__21316),
            .in1(N__21304),
            .in2(_gnd_net_),
            .in3(N__26892),
            .lcout(\u1.N_1431 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_pong_d_RNIJ1IN_8_LC_5_29_5 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_pong_d_RNIJ1IN_8_LC_5_29_5 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.gen_pingpong_pong_d_RNIJ1IN_8_LC_5_29_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.PIO_control.gen_pingpong_pong_d_RNIJ1IN_8_LC_5_29_5  (
            .in0(N__21292),
            .in1(N__21280),
            .in2(_gnd_net_),
            .in3(N__26894),
            .lcout(\u1.N_1433 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_pong_d_RNIHVHN_7_LC_5_29_7 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_pong_d_RNIHVHN_7_LC_5_29_7 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.gen_pingpong_pong_d_RNIHVHN_7_LC_5_29_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.PIO_control.gen_pingpong_pong_d_RNIHVHN_7_LC_5_29_7  (
            .in0(N__21268),
            .in1(N__21256),
            .in2(_gnd_net_),
            .in3(N__26893),
            .lcout(\u1.N_1432 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DDo_13_LC_5_30_0 .C_ON=1'b0;
    defparam \u1.DDo_13_LC_5_30_0 .SEQ_MODE=4'b1010;
    defparam \u1.DDo_13_LC_5_30_0 .LUT_INIT=16'b0000111000000010;
    LogicCell40 \u1.DDo_13_LC_5_30_0  (
            .in0(N__22336),
            .in1(N__36779),
            .in2(N__52761),
            .in3(N__22951),
            .lcout(dd_pad_o_c_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54252),
            .ce(),
            .sr(N__53389));
    defparam \u1.DDo_6_LC_5_30_6 .C_ON=1'b0;
    defparam \u1.DDo_6_LC_5_30_6 .SEQ_MODE=4'b1010;
    defparam \u1.DDo_6_LC_5_30_6 .LUT_INIT=16'b0000111000000010;
    LogicCell40 \u1.DDo_6_LC_5_30_6  (
            .in0(N__22705),
            .in1(N__36780),
            .in2(N__52762),
            .in3(N__21232),
            .lcout(dd_pad_o_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54252),
            .ce(),
            .sr(N__53389));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_0_LC_6_16_2 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_0_LC_6_16_2 .SEQ_MODE=4'b1010;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_0_LC_6_16_2 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_0_LC_6_16_2  (
            .in0(N__24616),
            .in1(N__26038),
            .in2(N__52305),
            .in3(N__24822),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.Qi_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54135),
            .ce(N__24752),
            .sr(N__53311));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_1_LC_6_17_2 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_1_LC_6_17_2 .SEQ_MODE=4'b1011;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_1_LC_6_17_2 .LUT_INIT=16'b1111101111001000;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_1_LC_6_17_2  (
            .in0(N__26527),
            .in1(N__24823),
            .in2(N__52196),
            .in3(N__23119),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.QiZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54124),
            .ce(N__24759),
            .sr(N__53319));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_2_LC_6_17_3 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_2_LC_6_17_3 .SEQ_MODE=4'b1011;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_2_LC_6_17_3 .LUT_INIT=16'b1111110110101000;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_2_LC_6_17_3  (
            .in0(N__24824),
            .in1(N__24475),
            .in2(N__52306),
            .in3(N__23098),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.QiZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54124),
            .ce(N__24759),
            .sr(N__53319));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_3_LC_6_17_4 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_3_LC_6_17_4 .SEQ_MODE=4'b1010;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_3_LC_6_17_4 .LUT_INIT=16'b0011101100001000;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_3_LC_6_17_4  (
            .in0(N__26161),
            .in1(N__24825),
            .in2(N__52197),
            .in3(N__23077),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.QiZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54124),
            .ce(N__24759),
            .sr(N__53319));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_4_LC_6_17_5 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_4_LC_6_17_5 .SEQ_MODE=4'b1010;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_4_LC_6_17_5 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_4_LC_6_17_5  (
            .in0(N__24826),
            .in1(N__24466),
            .in2(N__52307),
            .in3(N__23056),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.QiZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54124),
            .ce(N__24759),
            .sr(N__53319));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_5_LC_6_17_6 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_5_LC_6_17_6 .SEQ_MODE=4'b1010;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_5_LC_6_17_6 .LUT_INIT=16'b0011101100001000;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_5_LC_6_17_6  (
            .in0(N__26188),
            .in1(N__24827),
            .in2(N__52198),
            .in3(N__23035),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.QiZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54124),
            .ce(N__24759),
            .sr(N__53319));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_6_LC_6_17_7 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_6_LC_6_17_7 .SEQ_MODE=4'b1010;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_6_LC_6_17_7 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_6_LC_6_17_7  (
            .in0(N__24828),
            .in1(N__27373),
            .in2(N__52308),
            .in3(N__23296),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.QiZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54124),
            .ce(N__24759),
            .sr(N__53319));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qie_0_i_LC_6_18_2 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qie_0_i_LC_6_18_2 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qie_0_i_LC_6_18_2 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qie_0_i_LC_6_18_2  (
            .in0(N__52502),
            .in1(N__23199),
            .in2(_gnd_net_),
            .in3(N__24715),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qie_0_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNIVBR8_1_LC_6_18_3 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNIVBR8_1_LC_6_18_3 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNIVBR8_1_LC_6_18_3 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNIVBR8_1_LC_6_18_3  (
            .in0(N__23067),
            .in1(N__23088),
            .in2(_gnd_net_),
            .in3(N__23130),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.val_c8_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_2_LC_6_18_6 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_2_LC_6_18_6 .SEQ_MODE=4'b1011;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_2_LC_6_18_6 .LUT_INIT=16'b1111101011001100;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_2_LC_6_18_6  (
            .in0(N__27439),
            .in1(N__28870),
            .in2(N__52636),
            .in3(N__26450),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.QiZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54136),
            .ce(N__26427),
            .sr(N__53321));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_5_LC_6_18_7 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_5_LC_6_18_7 .SEQ_MODE=4'b1010;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_5_LC_6_18_7 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_5_LC_6_18_7  (
            .in0(N__26451),
            .in1(N__52501),
            .in2(N__28765),
            .in3(N__27526),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.QiZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54136),
            .ce(N__26427),
            .sr(N__53321));
    defparam \u1.PIO_control.gen_pingpong_pong_a_2_LC_6_19_0 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_pong_a_2_LC_6_19_0 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_pong_a_2_LC_6_19_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.PIO_control.gen_pingpong_pong_a_2_LC_6_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53068),
            .lcout(\u1.pong_a_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54142),
            .ce(N__24883),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_pong_d_0_LC_6_19_1 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_pong_d_0_LC_6_19_1 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_pong_d_0_LC_6_19_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \u1.PIO_control.gen_pingpong_pong_d_0_LC_6_19_1  (
            .in0(N__49533),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\u1.PIO_control.pong_d_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54142),
            .ce(N__24883),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_pong_d_1_LC_6_19_2 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_pong_d_1_LC_6_19_2 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_pong_d_1_LC_6_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.PIO_control.gen_pingpong_pong_d_1_LC_6_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39345),
            .lcout(\u1.PIO_control.pong_d_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54142),
            .ce(N__24883),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_pong_d_10_LC_6_19_3 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_pong_d_10_LC_6_19_3 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_pong_d_10_LC_6_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.PIO_control.gen_pingpong_pong_d_10_LC_6_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40172),
            .lcout(\u1.PIO_control.pong_d_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54142),
            .ce(N__24883),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_pong_d_11_LC_6_19_4 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_pong_d_11_LC_6_19_4 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_pong_d_11_LC_6_19_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \u1.PIO_control.gen_pingpong_pong_d_11_LC_6_19_4  (
            .in0(N__43676),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\u1.PIO_control.pong_d_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54142),
            .ce(N__24883),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_pong_d_12_LC_6_19_5 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_pong_d_12_LC_6_19_5 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_pong_d_12_LC_6_19_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \u1.PIO_control.gen_pingpong_pong_d_12_LC_6_19_5  (
            .in0(N__36951),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\u1.PIO_control.pong_d_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54142),
            .ce(N__24883),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_pong_d_13_LC_6_19_6 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_pong_d_13_LC_6_19_6 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_pong_d_13_LC_6_19_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \u1.PIO_control.gen_pingpong_pong_d_13_LC_6_19_6  (
            .in0(N__34698),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\u1.PIO_control.pong_d_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54142),
            .ce(N__24883),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_pong_d_14_LC_6_19_7 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_pong_d_14_LC_6_19_7 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_pong_d_14_LC_6_19_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \u1.PIO_control.gen_pingpong_pong_d_14_LC_6_19_7  (
            .in0(N__44015),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\u1.PIO_control.pong_d_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54142),
            .ce(N__24883),
            .sr(_gnd_net_));
    defparam \u1.c_state_RNIUC0A1_1_LC_6_20_0 .C_ON=1'b0;
    defparam \u1.c_state_RNIUC0A1_1_LC_6_20_0 .SEQ_MODE=4'b0000;
    defparam \u1.c_state_RNIUC0A1_1_LC_6_20_0 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \u1.c_state_RNIUC0A1_1_LC_6_20_0  (
            .in0(N__24953),
            .in1(N__24404),
            .in2(N__52494),
            .in3(N__21423),
            .lcout(),
            .ltout(\u1.c_state_RNIUC0A1Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.c_state_RNITERO1_0_LC_6_20_1 .C_ON=1'b0;
    defparam \u1.c_state_RNITERO1_0_LC_6_20_1 .SEQ_MODE=4'b0000;
    defparam \u1.c_state_RNITERO1_0_LC_6_20_1 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \u1.c_state_RNITERO1_0_LC_6_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21388),
            .in3(N__24446),
            .lcout(\u1.DMAtip_2_i_i_a2_0_1 ),
            .ltout(\u1.DMAtip_2_i_i_a2_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.valid_RNIGA8B4_LC_6_20_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.valid_RNIGA8B4_LC_6_20_2 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.valid_RNIGA8B4_LC_6_20_2 .LUT_INIT=16'b1111000001000000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Txbuf.valid_RNIGA8B4_LC_6_20_2  (
            .in0(N__23656),
            .in1(N__23328),
            .in2(N__21601),
            .in3(N__23307),
            .lcout(\u1.N_1874 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_cmdport_T2_RNIAION3_7_LC_6_20_3 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_T2_RNIAION3_7_LC_6_20_3 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_cmdport_T2_RNIAION3_7_LC_6_20_3 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \u0.PIO_cmdport_T2_RNIAION3_7_LC_6_20_3  (
            .in0(N__46593),
            .in1(N__48145),
            .in2(N__21498),
            .in3(N__29619),
            .lcout(\u0.dat_o_0_0_3_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMACKn_LC_6_20_4 .C_ON=1'b0;
    defparam \u1.DMACKn_LC_6_20_4 .SEQ_MODE=4'b1011;
    defparam \u1.DMACKn_LC_6_20_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \u1.DMACKn_LC_6_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21577),
            .lcout(dmackn_pad_o_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54149),
            .ce(),
            .sr(N__53329));
    defparam \u1.DMAtip_RNIHESH_LC_6_20_6 .C_ON=1'b0;
    defparam \u1.DMAtip_RNIHESH_LC_6_20_6 .SEQ_MODE=4'b0000;
    defparam \u1.DMAtip_RNIHESH_LC_6_20_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u1.DMAtip_RNIHESH_LC_6_20_6  (
            .in0(N__52301),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21490),
            .lcout(\u1.N_2150 ),
            .ltout(\u1.N_2150_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMAtip_LC_6_20_7 .C_ON=1'b0;
    defparam \u1.DMAtip_LC_6_20_7 .SEQ_MODE=4'b1010;
    defparam \u1.DMAtip_LC_6_20_7 .LUT_INIT=16'b1111111111010000;
    LogicCell40 \u1.DMAtip_LC_6_20_7  (
            .in0(N__21571),
            .in1(N__21559),
            .in2(N__21532),
            .in3(N__21522),
            .lcout(DMAtip),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54149),
            .ce(),
            .sr(N__53329));
    defparam \u0.PIO_dport1_T1_RNIC3004_0_LC_6_21_0 .C_ON=1'b0;
    defparam \u0.PIO_dport1_T1_RNIC3004_0_LC_6_21_0 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport1_T1_RNIC3004_0_LC_6_21_0 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \u0.PIO_dport1_T1_RNIC3004_0_LC_6_21_0  (
            .in0(N__46984),
            .in1(N__54673),
            .in2(N__23578),
            .in3(N__26005),
            .lcout(\u0.dat_o_0_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_Tm_0_LC_6_21_1 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_Tm_0_LC_6_21_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.DMA_timing_ctrl_Tm_0_LC_6_21_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_Tm_0_LC_6_21_1  (
            .in0(N__36231),
            .in1(N__23574),
            .in2(_gnd_net_),
            .in3(N__41160),
            .lcout(\u1.DMA_control.Tm_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54155),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.gen_bc_dec_store_pp_full_RNIRR9R_LC_6_21_2 .C_ON=1'b0;
    defparam \u0.gen_bc_dec_store_pp_full_RNIRR9R_LC_6_21_2 .SEQ_MODE=4'b0000;
    defparam \u0.gen_bc_dec_store_pp_full_RNIRR9R_LC_6_21_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \u0.gen_bc_dec_store_pp_full_RNIRR9R_LC_6_21_2  (
            .in0(N__21482),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21455),
            .lcout(N_1360),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_Td_2_LC_6_21_4 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_Td_2_LC_6_21_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.DMA_timing_ctrl_Td_2_LC_6_21_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_Td_2_LC_6_21_4  (
            .in0(N__43560),
            .in1(N__40056),
            .in2(_gnd_net_),
            .in3(N__36227),
            .lcout(\u1.DMA_control.Td_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54155),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_Td_3_LC_6_21_5 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_Td_3_LC_6_21_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.DMA_timing_ctrl_Td_3_LC_6_21_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_Td_3_LC_6_21_5  (
            .in0(N__36228),
            .in1(N__31288),
            .in2(_gnd_net_),
            .in3(N__43752),
            .lcout(\u1.DMA_control.Td_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54155),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_Td_4_LC_6_21_6 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_Td_4_LC_6_21_6 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.DMA_timing_ctrl_Td_4_LC_6_21_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_Td_4_LC_6_21_6  (
            .in0(N__31561),
            .in1(N__29682),
            .in2(_gnd_net_),
            .in3(N__36229),
            .lcout(\u1.DMA_control.Td_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54155),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_Td_7_LC_6_21_7 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_Td_7_LC_6_21_7 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.DMA_timing_ctrl_Td_7_LC_6_21_7 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_Td_7_LC_6_21_7  (
            .in0(N__36230),
            .in1(_gnd_net_),
            .in2(N__31365),
            .in3(N__24924),
            .lcout(\u1.DMA_control.Td_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54155),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.rty_o_i_o2_LC_6_22_0 .C_ON=1'b0;
    defparam \u0.rty_o_i_o2_LC_6_22_0 .SEQ_MODE=4'b0000;
    defparam \u0.rty_o_i_o2_LC_6_22_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \u0.rty_o_i_o2_LC_6_22_0  (
            .in0(_gnd_net_),
            .in1(N__47517),
            .in2(_gnd_net_),
            .in3(N__21852),
            .lcout(N_1369),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.err_o_i_o3_LC_6_22_1 .C_ON=1'b0;
    defparam \u0.err_o_i_o3_LC_6_22_1 .SEQ_MODE=4'b0000;
    defparam \u0.err_o_i_o3_LC_6_22_1 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \u0.err_o_i_o3_LC_6_22_1  (
            .in0(N__47516),
            .in1(N__21885),
            .in2(_gnd_net_),
            .in3(N__21803),
            .lcout(\u0.N_1384 ),
            .ltout(\u0.N_1384_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.CtrlReg_RNIR8PJ1_7_LC_6_22_2 .C_ON=1'b0;
    defparam \u0.CtrlReg_RNIR8PJ1_7_LC_6_22_2 .SEQ_MODE=4'b0000;
    defparam \u0.CtrlReg_RNIR8PJ1_7_LC_6_22_2 .LUT_INIT=16'b0010111100001111;
    LogicCell40 \u0.CtrlReg_RNIR8PJ1_7_LC_6_22_2  (
            .in0(N__47512),
            .in1(N__21682),
            .in2(N__21667),
            .in3(N__38326),
            .lcout(),
            .ltout(\u0.ack_o_i_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.CtrlReg_RNIL9JM3_7_LC_6_22_3 .C_ON=1'b0;
    defparam \u0.CtrlReg_RNIL9JM3_7_LC_6_22_3 .SEQ_MODE=4'b0000;
    defparam \u0.CtrlReg_RNIL9JM3_7_LC_6_22_3 .LUT_INIT=16'b0000000100000101;
    LogicCell40 \u0.CtrlReg_RNIL9JM3_7_LC_6_22_3  (
            .in0(N__21850),
            .in1(N__47511),
            .in2(N__21664),
            .in3(N__21645),
            .lcout(N_410_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.gen_bc_dec_store_pp_full_RNIQ0Q22_LC_6_22_4 .C_ON=1'b0;
    defparam \u0.gen_bc_dec_store_pp_full_RNIQ0Q22_LC_6_22_4 .SEQ_MODE=4'b0000;
    defparam \u0.gen_bc_dec_store_pp_full_RNIQ0Q22_LC_6_22_4 .LUT_INIT=16'b0010000000100000;
    LogicCell40 \u0.gen_bc_dec_store_pp_full_RNIQ0Q22_LC_6_22_4  (
            .in0(N__21646),
            .in1(N__21851),
            .in2(N__47518),
            .in3(_gnd_net_),
            .lcout(N_288_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_ping_d_RNI5SB31_10_LC_6_22_5 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_ping_d_RNI5SB31_10_LC_6_22_5 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.gen_pingpong_ping_d_RNI5SB31_10_LC_6_22_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.PIO_control.gen_pingpong_ping_d_RNI5SB31_10_LC_6_22_5  (
            .in0(N__21610),
            .in1(N__25114),
            .in2(_gnd_net_),
            .in3(N__26921),
            .lcout(\u1.N_1435 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_Td_0_LC_6_22_6 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_Td_0_LC_6_22_6 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.DMA_timing_ctrl_Td_0_LC_6_22_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_Td_0_LC_6_22_6  (
            .in0(N__23424),
            .in1(N__31333),
            .in2(_gnd_net_),
            .in3(N__36257),
            .lcout(\u1.DMA_control.Td_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54167),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.valid_3_0_0_a2_2_LC_6_22_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.valid_3_0_0_a2_2_LC_6_22_7 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.valid_3_0_0_a2_2_LC_6_22_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Txbuf.valid_3_0_0_a2_2_LC_6_22_7  (
            .in0(N__21960),
            .in1(N__21886),
            .in2(N__21856),
            .in3(N__21804),
            .lcout(N_2140),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DDo_10_LC_6_23_2 .C_ON=1'b0;
    defparam \u1.DDo_10_LC_6_23_2 .SEQ_MODE=4'b1010;
    defparam \u1.DDo_10_LC_6_23_2 .LUT_INIT=16'b0000111000000010;
    LogicCell40 \u1.DDo_10_LC_6_23_2  (
            .in0(N__22429),
            .in1(N__36698),
            .in2(N__52709),
            .in3(N__21769),
            .lcout(dd_pad_o_c_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54177),
            .ce(),
            .sr(N__53348));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_2_LC_6_24_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_2_LC_6_24_0 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_2_LC_6_24_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDlw_2_LC_6_24_0  (
            .in0(N__22446),
            .in1(N__24006),
            .in2(_gnd_net_),
            .in3(N__42980),
            .lcout(\u1.DMA_control.writeDlw_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54189),
            .ce(N__25607),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_10_LC_6_24_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_10_LC_6_24_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_10_LC_6_24_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDlw_10_LC_6_24_1  (
            .in0(N__42976),
            .in1(N__25845),
            .in2(_gnd_net_),
            .in3(N__25881),
            .lcout(\u1.DMA_control.writeDlw_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54189),
            .ce(N__25607),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_4_LC_6_24_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_4_LC_6_24_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_4_LC_6_24_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDlw_4_LC_6_24_2  (
            .in0(N__22380),
            .in1(N__22062),
            .in2(_gnd_net_),
            .in3(N__42981),
            .lcout(\u1.DMA_control.writeDlw_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54189),
            .ce(N__25607),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_5_LC_6_24_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_5_LC_6_24_3 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_5_LC_6_24_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDlw_5_LC_6_24_3  (
            .in0(N__42977),
            .in1(N__22350),
            .in2(_gnd_net_),
            .in3(N__24039),
            .lcout(\u1.DMA_control.writeDlw_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54189),
            .ce(N__25607),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_6_LC_6_24_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_6_LC_6_24_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_6_LC_6_24_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDlw_6_LC_6_24_4  (
            .in0(N__22320),
            .in1(N__22035),
            .in2(_gnd_net_),
            .in3(N__42982),
            .lcout(\u1.DMA_control.writeDlw_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54189),
            .ce(N__25607),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_7_LC_6_24_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_7_LC_6_24_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_7_LC_6_24_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDlw_7_LC_6_24_5  (
            .in0(N__42978),
            .in1(N__25647),
            .in2(_gnd_net_),
            .in3(N__25674),
            .lcout(\u1.DMA_control.writeDlw_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54189),
            .ce(N__25607),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_8_LC_6_24_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_8_LC_6_24_6 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_8_LC_6_24_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDlw_8_LC_6_24_6  (
            .in0(N__21987),
            .in1(N__22135),
            .in2(_gnd_net_),
            .in3(N__42983),
            .lcout(\u1.DMA_control.writeDlw_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54189),
            .ce(N__25607),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_9_LC_6_24_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_9_LC_6_24_7 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDlw_9_LC_6_24_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDlw_9_LC_6_24_7  (
            .in0(N__42979),
            .in1(_gnd_net_),
            .in2(N__22470),
            .in3(N__22114),
            .lcout(\u1.DMA_control.writeDlw_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54189),
            .ce(N__25607),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_7_LC_6_25_0 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_7_LC_6_25_0 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_7_LC_6_25_0 .LUT_INIT=16'b0011101100001000;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.Qi_7_LC_6_25_0  (
            .in0(N__36103),
            .in1(N__22228),
            .in2(N__52611),
            .in3(N__22195),
            .lcout(\u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.tm_cnt.cnt.QiZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54200),
            .ce(N__22162),
            .sr(N__53360));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_0_LC_6_25_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_0_LC_6_25_1 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_0_LC_6_25_1 .LUT_INIT=16'b0000001101010011;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_0_LC_6_25_1  (
            .in0(N__22134),
            .in1(N__22123),
            .in2(N__25585),
            .in3(N__42740),
            .lcout(\u1.DMA_control.writeDfw_6_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_1_LC_6_25_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_1_LC_6_25_2 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_1_LC_6_25_2 .LUT_INIT=16'b0001000100001111;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_1_LC_6_25_2  (
            .in0(N__42739),
            .in1(N__22113),
            .in2(N__22102),
            .in3(N__25528),
            .lcout(\u1.DMA_control.writeDfw_6_i_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_11_LC_6_25_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_11_LC_6_25_4 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_11_LC_6_25_4 .LUT_INIT=16'b0001000100001111;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_11_LC_6_25_4  (
            .in0(N__42738),
            .in1(N__22086),
            .in2(N__22075),
            .in3(N__25527),
            .lcout(\u1.DMA_control.writeDfw_6_i_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_12_LC_6_25_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_12_LC_6_25_5 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_12_LC_6_25_5 .LUT_INIT=16'b0000001101000111;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_12_LC_6_25_5  (
            .in0(N__22063),
            .in1(N__25529),
            .in2(N__22048),
            .in3(N__42741),
            .lcout(\u1.DMA_control.writeDfw_6_i_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_14_LC_6_25_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_14_LC_6_25_7 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_14_LC_6_25_7 .LUT_INIT=16'b0000001101000111;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_14_LC_6_25_7  (
            .in0(N__22036),
            .in1(N__25530),
            .in2(N__22015),
            .in3(N__42742),
            .lcout(\u1.DMA_control.writeDfw_6_i_m3_i_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_0_LC_6_26_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_0_LC_6_26_0 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_0_LC_6_26_0 .LUT_INIT=16'b0011000100110011;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDfw_0_LC_6_26_0  (
            .in0(N__25567),
            .in1(N__22000),
            .in2(N__21994),
            .in3(N__42811),
            .lcout(\u1.DMAd_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54213),
            .ce(N__25381),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.dstrb_RNI1KRS_LC_6_26_1 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.dstrb_RNI1KRS_LC_6_26_1 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.dstrb_RNI1KRS_LC_6_26_1 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_DMA_timing_ctrl.dstrb_RNI1KRS_LC_6_26_1  (
            .in0(N__25550),
            .in1(N__22504),
            .in2(_gnd_net_),
            .in3(N__23657),
            .lcout(\u1.DMA_control.N_53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_1_LC_6_26_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_1_LC_6_26_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_1_LC_6_26_2 .LUT_INIT=16'b0011001100010011;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDfw_1_LC_6_26_2  (
            .in0(N__25570),
            .in1(N__22477),
            .in2(N__42984),
            .in3(N__22471),
            .lcout(\u1.DMAd_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54213),
            .ce(N__25381),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_10_LC_6_26_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_10_LC_6_26_3 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_10_LC_6_26_3 .LUT_INIT=16'b0000000011110111;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDfw_10_LC_6_26_3  (
            .in0(N__42807),
            .in1(N__25571),
            .in2(N__22453),
            .in3(N__23977),
            .lcout(\u1.DMAd_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54213),
            .ce(N__25381),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_11_LC_6_26_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_11_LC_6_26_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_11_LC_6_26_4 .LUT_INIT=16'b0011000100110011;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDfw_11_LC_6_26_4  (
            .in0(N__25568),
            .in1(N__22420),
            .in2(N__22414),
            .in3(N__42812),
            .lcout(\u1.DMAd_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54213),
            .ce(N__25381),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_12_LC_6_26_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_12_LC_6_26_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_12_LC_6_26_5 .LUT_INIT=16'b0000000011110111;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDfw_12_LC_6_26_5  (
            .in0(N__42808),
            .in1(N__25572),
            .in2(N__22387),
            .in3(N__22363),
            .lcout(\u1.DMAd_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54213),
            .ce(N__25381),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_13_LC_6_26_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_13_LC_6_26_6 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_13_LC_6_26_6 .LUT_INIT=16'b0000000011110111;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDfw_13_LC_6_26_6  (
            .in0(N__25569),
            .in1(N__42810),
            .in2(N__22357),
            .in3(N__24025),
            .lcout(\u1.DMAd_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54213),
            .ce(N__25381),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_14_LC_6_26_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_14_LC_6_26_7 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_14_LC_6_26_7 .LUT_INIT=16'b0000000011110111;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDfw_14_LC_6_26_7  (
            .in0(N__42809),
            .in1(N__25573),
            .in2(N__22324),
            .in3(N__22297),
            .lcout(\u1.DMAd_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54213),
            .ce(N__25381),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_5_LC_6_27_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_5_LC_6_27_0 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_5_LC_6_27_0 .LUT_INIT=16'b0000001101000111;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_5_LC_6_27_0  (
            .in0(N__22287),
            .in1(N__25551),
            .in2(N__22270),
            .in3(N__42502),
            .lcout(\u1.DMA_control.writeDfw_6_i_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_6_LC_6_27_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_6_LC_6_27_1 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_6_LC_6_27_1 .LUT_INIT=16'b0000001101010011;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_6_LC_6_27_1  (
            .in0(N__42503),
            .in1(N__22258),
            .in2(N__25608),
            .in3(N__22246),
            .lcout(),
            .ltout(\u1.DMA_control.writeDfw_6_i_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_6_LC_6_27_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_6_LC_6_27_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_6_LC_6_27_2 .LUT_INIT=16'b0000101100001111;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDfw_6_LC_6_27_2  (
            .in0(N__22726),
            .in1(N__25561),
            .in2(N__22708),
            .in3(N__42507),
            .lcout(\u1.DMAd_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54227),
            .ce(N__25391),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_7_LC_6_27_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_7_LC_6_27_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_7_LC_6_27_3 .LUT_INIT=16'b0000001101010011;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_7_LC_6_27_3  (
            .in0(N__42504),
            .in1(N__22696),
            .in2(N__25609),
            .in3(N__22686),
            .lcout(),
            .ltout(\u1.DMA_control.writeDfw_6_i_0_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_7_LC_6_27_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_7_LC_6_27_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_7_LC_6_27_4 .LUT_INIT=16'b0000101100001111;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDfw_7_LC_6_27_4  (
            .in0(N__22663),
            .in1(N__25562),
            .in2(N__22642),
            .in3(N__42508),
            .lcout(\u1.DMAd_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54227),
            .ce(N__25391),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_8_LC_6_27_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_8_LC_6_27_5 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_8_LC_6_27_5 .LUT_INIT=16'b0000001101010011;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_8_LC_6_27_5  (
            .in0(N__42505),
            .in1(N__22639),
            .in2(N__25610),
            .in3(N__22630),
            .lcout(),
            .ltout(\u1.DMA_control.writeDfw_6_i_0_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_8_LC_6_27_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_8_LC_6_27_6 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_8_LC_6_27_6 .LUT_INIT=16'b0000101100001111;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDfw_8_LC_6_27_6  (
            .in0(N__22609),
            .in1(N__25563),
            .in2(N__22585),
            .in3(N__42509),
            .lcout(\u1.DMAd_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54227),
            .ce(N__25391),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_5_LC_6_27_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_5_LC_6_27_7 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_5_LC_6_27_7 .LUT_INIT=16'b0000000011011111;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDfw_5_LC_6_27_7  (
            .in0(N__42506),
            .in1(N__22582),
            .in2(N__25611),
            .in3(N__22558),
            .lcout(\u1.DMAd_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54227),
            .ce(N__25391),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_ping_d_RNI7UB31_11_LC_6_28_1 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_ping_d_RNI7UB31_11_LC_6_28_1 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.gen_pingpong_ping_d_RNI7UB31_11_LC_6_28_1 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \u1.PIO_control.gen_pingpong_ping_d_RNI7UB31_11_LC_6_28_1  (
            .in0(N__22543),
            .in1(N__25102),
            .in2(N__26928),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\u1.N_1448_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DDo_11_LC_6_28_2 .C_ON=1'b0;
    defparam \u1.DDo_11_LC_6_28_2 .SEQ_MODE=4'b1010;
    defparam \u1.DDo_11_LC_6_28_2 .LUT_INIT=16'b0101000001000100;
    LogicCell40 \u1.DDo_11_LC_6_28_2  (
            .in0(N__52710),
            .in1(N__22531),
            .in2(N__22522),
            .in3(N__36778),
            .lcout(dd_pad_o_c_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54238),
            .ce(),
            .sr(N__53384));
    defparam \u1.PIO_control.gen_pingpong_ping_d_RNI90C31_12_LC_6_28_3 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_ping_d_RNI90C31_12_LC_6_28_3 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.gen_pingpong_ping_d_RNI90C31_12_LC_6_28_3 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \u1.PIO_control.gen_pingpong_ping_d_RNI90C31_12_LC_6_28_3  (
            .in0(N__23014),
            .in1(N__23002),
            .in2(N__26927),
            .in3(_gnd_net_),
            .lcout(\u1.N_1447 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_ping_d_RNID4C31_14_LC_6_28_5 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_ping_d_RNID4C31_14_LC_6_28_5 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.gen_pingpong_ping_d_RNID4C31_14_LC_6_28_5 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \u1.PIO_control.gen_pingpong_ping_d_RNID4C31_14_LC_6_28_5  (
            .in0(N__22993),
            .in1(N__22981),
            .in2(N__26926),
            .in3(_gnd_net_),
            .lcout(\u1.N_1445 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_ping_d_RNIB2C31_13_LC_6_28_7 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_ping_d_RNIB2C31_13_LC_6_28_7 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.gen_pingpong_ping_d_RNIB2C31_13_LC_6_28_7 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \u1.PIO_control.gen_pingpong_ping_d_RNIB2C31_13_LC_6_28_7  (
            .in0(N__22972),
            .in1(N__22960),
            .in2(N__26925),
            .in3(_gnd_net_),
            .lcout(\u1.N_1446 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DDo_12_LC_6_29_2 .C_ON=1'b0;
    defparam \u1.DDo_12_LC_6_29_2 .SEQ_MODE=4'b1010;
    defparam \u1.DDo_12_LC_6_29_2 .LUT_INIT=16'b0000111000000010;
    LogicCell40 \u1.DDo_12_LC_6_29_2  (
            .in0(N__22942),
            .in1(N__36776),
            .in2(N__52767),
            .in3(N__22933),
            .lcout(dd_pad_o_c_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54253),
            .ce(),
            .sr(N__53390));
    defparam \u1.DDo_14_LC_6_29_5 .C_ON=1'b0;
    defparam \u1.DDo_14_LC_6_29_5 .SEQ_MODE=4'b1010;
    defparam \u1.DDo_14_LC_6_29_5 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \u1.DDo_14_LC_6_29_5  (
            .in0(N__22915),
            .in1(N__22909),
            .in2(N__52699),
            .in3(N__36781),
            .lcout(dd_pad_o_c_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54253),
            .ce(),
            .sr(N__53390));
    defparam \u1.DDo_8_LC_6_29_7 .C_ON=1'b0;
    defparam \u1.DDo_8_LC_6_29_7 .SEQ_MODE=4'b1010;
    defparam \u1.DDo_8_LC_6_29_7 .LUT_INIT=16'b0000111000000010;
    LogicCell40 \u1.DDo_8_LC_6_29_7  (
            .in0(N__22888),
            .in1(N__36782),
            .in2(N__52700),
            .in3(N__22879),
            .lcout(dd_pad_o_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54253),
            .ce(),
            .sr(N__53390));
    defparam \u1.DDo_7_LC_6_30_0 .C_ON=1'b0;
    defparam \u1.DDo_7_LC_6_30_0 .SEQ_MODE=4'b1010;
    defparam \u1.DDo_7_LC_6_30_0 .LUT_INIT=16'b0000111000000010;
    LogicCell40 \u1.DDo_7_LC_6_30_0  (
            .in0(N__22861),
            .in1(N__36783),
            .in2(N__52787),
            .in3(N__22852),
            .lcout(dd_pad_o_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54265),
            .ce(),
            .sr(N__53393));
    defparam \u0.N_284_i_LC_7_14_2 .C_ON=1'b0;
    defparam \u0.N_284_i_LC_7_14_2 .SEQ_MODE=4'b0000;
    defparam \u0.N_284_i_LC_7_14_2 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \u0.N_284_i_LC_7_14_2  (
            .in0(N__22837),
            .in1(N__22822),
            .in2(N__22795),
            .in3(N__22780),
            .lcout(N_284_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev0_Td_RNIQ5H22_0_LC_7_14_6 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Td_RNIQ5H22_0_LC_7_14_6 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev0_Td_RNIQ5H22_0_LC_7_14_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \u0.DMA_dev0_Td_RNIQ5H22_0_LC_7_14_6  (
            .in0(_gnd_net_),
            .in1(N__48604),
            .in2(_gnd_net_),
            .in3(N__23425),
            .lcout(\u0.N_1736 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport0_T1_2_LC_7_16_3 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T1_2_LC_7_16_3 .SEQ_MODE=4'b1011;
    defparam \u0.PIO_dport0_T1_2_LC_7_16_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \u0.PIO_dport0_T1_2_LC_7_16_3  (
            .in0(_gnd_net_),
            .in1(N__34243),
            .in2(_gnd_net_),
            .in3(N__52115),
            .lcout(PIO_dport0_T1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54143),
            .ce(N__49383),
            .sr(N__53315));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_cry_c_0_LC_7_17_0 .C_ON=1'b1;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_cry_c_0_LC_7_17_0 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_cry_c_0_LC_7_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_cry_c_0_LC_7_17_0  (
            .in0(_gnd_net_),
            .in1(N__26056),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_17_0_),
            .carryout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNO_0_1_LC_7_17_1 .C_ON=1'b1;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNO_0_1_LC_7_17_1 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNO_0_1_LC_7_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNO_0_1_LC_7_17_1  (
            .in0(_gnd_net_),
            .in1(N__23131),
            .in2(N__28699),
            .in3(N__23113),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_s_1 ),
            .ltout(),
            .carryin(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_cry_0 ),
            .carryout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNO_0_2_LC_7_17_2 .C_ON=1'b1;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNO_0_2_LC_7_17_2 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNO_0_2_LC_7_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNO_0_2_LC_7_17_2  (
            .in0(_gnd_net_),
            .in1(N__23110),
            .in2(N__28703),
            .in3(N__23092),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_s_2 ),
            .ltout(),
            .carryin(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_cry_1 ),
            .carryout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNO_0_3_LC_7_17_3 .C_ON=1'b1;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNO_0_3_LC_7_17_3 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNO_0_3_LC_7_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNO_0_3_LC_7_17_3  (
            .in0(_gnd_net_),
            .in1(N__23089),
            .in2(N__28700),
            .in3(N__23071),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_s_3 ),
            .ltout(),
            .carryin(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_cry_2 ),
            .carryout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNO_0_4_LC_7_17_4 .C_ON=1'b1;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNO_0_4_LC_7_17_4 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNO_0_4_LC_7_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNO_0_4_LC_7_17_4  (
            .in0(_gnd_net_),
            .in1(N__23068),
            .in2(N__28704),
            .in3(N__23050),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_s_4 ),
            .ltout(),
            .carryin(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_cry_3 ),
            .carryout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNO_0_5_LC_7_17_5 .C_ON=1'b1;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNO_0_5_LC_7_17_5 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNO_0_5_LC_7_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNO_0_5_LC_7_17_5  (
            .in0(_gnd_net_),
            .in1(N__23047),
            .in2(N__28701),
            .in3(N__23029),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_s_5 ),
            .ltout(),
            .carryin(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_cry_4 ),
            .carryout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNO_0_6_LC_7_17_6 .C_ON=1'b1;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNO_0_6_LC_7_17_6 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNO_0_6_LC_7_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNO_0_6_LC_7_17_6  (
            .in0(_gnd_net_),
            .in1(N__23026),
            .in2(N__28705),
            .in3(N__23290),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_s_6 ),
            .ltout(),
            .carryin(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_cry_5 ),
            .carryout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNO_0_7_LC_7_17_7 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNO_0_7_LC_7_17_7 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNO_0_7_LC_7_17_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNO_0_7_LC_7_17_7  (
            .in0(_gnd_net_),
            .in1(N__24783),
            .in2(_gnd_net_),
            .in3(N__23287),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_s_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_1_LC_7_18_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_1_LC_7_18_0 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_1_LC_7_18_0 .LUT_INIT=16'b0001000101010000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_1_LC_7_18_0  (
            .in0(N__23866),
            .in1(N__27970),
            .in2(N__45253),
            .in3(N__23366),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54144),
            .ce(),
            .sr(N__53325));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_2_LC_7_18_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_2_LC_7_18_1 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_2_LC_7_18_1 .LUT_INIT=16'b0000000011001010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_2_LC_7_18_1  (
            .in0(N__49802),
            .in1(N__45210),
            .in2(N__23367),
            .in3(N__23867),
            .lcout(\u1.DMA_control.rd_ptr_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54144),
            .ce(),
            .sr(N__53325));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_3_LC_7_18_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_3_LC_7_18_2 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_3_LC_7_18_2 .LUT_INIT=16'b0101000001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_3_LC_7_18_2  (
            .in0(N__23868),
            .in1(N__48709),
            .in2(N__49835),
            .in3(N__23362),
            .lcout(u1_DMA_control_gen_DMAbuf_Rxbuf_rd_ptr_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54144),
            .ce(),
            .sr(N__53325));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.msb_LC_7_18_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.msb_LC_7_18_3 .SEQ_MODE=4'b1011;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.msb_LC_7_18_3 .LUT_INIT=16'b1110111111101100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.msb_LC_7_18_3  (
            .in0(N__48708),
            .in1(N__23869),
            .in2(N__23368),
            .in3(N__23347),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.drd_ptr_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54144),
            .ce(),
            .sr(N__53325));
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.valid_LC_7_18_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.valid_LC_7_18_4 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.valid_LC_7_18_4 .LUT_INIT=16'b0100010101000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Txbuf.valid_LC_7_18_4  (
            .in0(N__23870),
            .in1(N__23674),
            .in2(N__25630),
            .in3(N__31429),
            .lcout(DMATxFull),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54144),
            .ce(),
            .sr(N__53325));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.rci_LC_7_18_5 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.rci_LC_7_18_5 .SEQ_MODE=4'b1010;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.rci_LC_7_18_5 .LUT_INIT=16'b0000101100000011;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.rci_LC_7_18_5  (
            .in0(N__23206),
            .in1(N__23280),
            .in2(N__52493),
            .in3(N__23237),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.rci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54144),
            .ce(),
            .sr(N__53325));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.rci_LC_7_18_6 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.rci_LC_7_18_6 .SEQ_MODE=4'b1010;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.rci_LC_7_18_6 .LUT_INIT=16'b0000101100000011;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.rci_LC_7_18_6  (
            .in0(N__24560),
            .in1(N__23205),
            .in2(N__52635),
            .in3(N__24716),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.rciZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54144),
            .ce(),
            .sr(N__53325));
    defparam \u1.PIO_control.gen_pingpong_dsel_LC_7_18_7 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_dsel_LC_7_18_7 .SEQ_MODE=4'b1010;
    defparam \u1.PIO_control.gen_pingpong_dsel_LC_7_18_7 .LUT_INIT=16'b1110101000000000;
    LogicCell40 \u1.PIO_control.gen_pingpong_dsel_LC_7_18_7  (
            .in0(N__23145),
            .in1(N__38335),
            .in2(N__23188),
            .in3(N__23173),
            .lcout(\u1.PIO_control.dsel ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54144),
            .ce(),
            .sr(N__53325));
    defparam \u1.PIO_control.PIO_access_control.q_10_LC_7_19_0 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.q_10_LC_7_19_0 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.q_10_LC_7_19_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \u1.PIO_control.PIO_access_control.q_10_LC_7_19_0  (
            .in0(N__32297),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(PIOq_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54150),
            .ce(N__45873),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIAKTN_0_3_LC_7_19_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIAKTN_0_3_LC_7_19_1 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIAKTN_0_3_LC_7_19_1 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIAKTN_0_3_LC_7_19_1  (
            .in0(N__48706),
            .in1(N__23450),
            .in2(N__49834),
            .in3(N__23715),
            .lcout(),
            .ltout(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.un1_ena_i_0_o3_sx_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIV9B91_1_LC_7_19_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIV9B91_1_LC_7_19_2 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIV9B91_1_LC_7_19_2 .LUT_INIT=16'b1111001111111100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIV9B91_1_LC_7_19_2  (
            .in0(_gnd_net_),
            .in1(N__45181),
            .in2(N__23407),
            .in3(N__24320),
            .lcout(N_1364),
            .ltout(N_1364_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.dat_o_i_i_2_10_LC_7_19_3 .C_ON=1'b0;
    defparam \u0.dat_o_i_i_2_10_LC_7_19_3 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_i_i_2_10_LC_7_19_3 .LUT_INIT=16'b1000111110001000;
    LogicCell40 \u0.dat_o_i_i_2_10_LC_7_19_3  (
            .in0(N__47493),
            .in1(N__23392),
            .in2(N__23386),
            .in3(N__46603),
            .lcout(\u0.dat_o_i_i_2Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIAKTN_3_LC_7_19_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIAKTN_3_LC_7_19_4 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIAKTN_3_LC_7_19_4 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIAKTN_3_LC_7_19_4  (
            .in0(N__23716),
            .in1(N__49801),
            .in2(N__23455),
            .in3(N__48707),
            .lcout(),
            .ltout(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.un1_ena_i_0_o3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI497L4_1_LC_7_19_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI497L4_1_LC_7_19_5 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI497L4_1_LC_7_19_5 .LUT_INIT=16'b0000000011110110;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI497L4_1_LC_7_19_5  (
            .in0(N__24321),
            .in1(N__45182),
            .in2(N__23383),
            .in3(N__23380),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.N_2092 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.msb_RNI832T_LC_7_19_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.msb_RNI832T_LC_7_19_6 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.msb_RNI832T_LC_7_19_6 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.msb_RNI832T_LC_7_19_6  (
            .in0(N__23714),
            .in1(N__48705),
            .in2(N__23454),
            .in3(N__23346),
            .lcout(\u1.DMA_control.N_1346 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.valid_RNI9BM61_LC_7_19_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.valid_RNI9BM61_LC_7_19_7 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.valid_RNI9BM61_LC_7_19_7 .LUT_INIT=16'b1101111000010010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Txbuf.valid_RNI9BM61_LC_7_19_7  (
            .in0(N__49797),
            .in1(N__23655),
            .in2(N__24322),
            .in3(N__31425),
            .lcout(\u1.DMA_control.gen_DMAbuf_Txbuf.N_1341 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.register_block_gen_DMA_dev0_reg_un6_sel_dma_dev0_i_0_LC_7_20_0 .C_ON=1'b0;
    defparam \u0.register_block_gen_DMA_dev0_reg_un6_sel_dma_dev0_i_0_LC_7_20_0 .SEQ_MODE=4'b0000;
    defparam \u0.register_block_gen_DMA_dev0_reg_un6_sel_dma_dev0_i_0_LC_7_20_0 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \u0.register_block_gen_DMA_dev0_reg_un6_sel_dma_dev0_i_0_LC_7_20_0  (
            .in0(N__48599),
            .in1(N__52510),
            .in2(_gnd_net_),
            .in3(N__50822),
            .lcout(\u0.N_444 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev0_Td_0_LC_7_20_1 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Td_0_LC_7_20_1 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev0_Td_0_LC_7_20_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.DMA_dev0_Td_0_LC_7_20_1  (
            .in0(N__54468),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52503),
            .lcout(DMA_dev0_Td_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54156),
            .ce(N__39693),
            .sr(N__53334));
    defparam \u0.DMA_dev0_Td_1_LC_7_20_2 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Td_1_LC_7_20_2 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev0_Td_1_LC_7_20_2 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \u0.DMA_dev0_Td_1_LC_7_20_2  (
            .in0(N__36010),
            .in1(N__52504),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(DMA_dev0_Td_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54156),
            .ce(N__39693),
            .sr(N__53334));
    defparam \u0.DMA_dev0_Td_2_LC_7_20_3 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Td_2_LC_7_20_3 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev0_Td_2_LC_7_20_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.DMA_dev0_Td_2_LC_7_20_3  (
            .in0(N__52505),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40167),
            .lcout(DMA_dev0_Td_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54156),
            .ce(N__39693),
            .sr(N__53334));
    defparam \u0.DMA_dev0_Td_3_LC_7_20_4 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Td_3_LC_7_20_4 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev0_Td_3_LC_7_20_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \u0.DMA_dev0_Td_3_LC_7_20_4  (
            .in0(_gnd_net_),
            .in1(N__52506),
            .in2(_gnd_net_),
            .in3(N__43671),
            .lcout(DMA_dev0_Td_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54156),
            .ce(N__39693),
            .sr(N__53334));
    defparam \u0.DMA_dev0_Td_4_LC_7_20_5 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Td_4_LC_7_20_5 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev0_Td_4_LC_7_20_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.DMA_dev0_Td_4_LC_7_20_5  (
            .in0(N__52507),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36981),
            .lcout(DMA_dev0_Td_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54156),
            .ce(N__39693),
            .sr(N__53334));
    defparam \u0.DMA_dev0_Td_5_LC_7_20_6 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Td_5_LC_7_20_6 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev0_Td_5_LC_7_20_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \u0.DMA_dev0_Td_5_LC_7_20_6  (
            .in0(_gnd_net_),
            .in1(N__52508),
            .in2(_gnd_net_),
            .in3(N__34703),
            .lcout(DMA_dev0_Td_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54156),
            .ce(N__39693),
            .sr(N__53334));
    defparam \u0.DMA_dev0_Td_6_LC_7_20_7 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Td_6_LC_7_20_7 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev0_Td_6_LC_7_20_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.DMA_dev0_Td_6_LC_7_20_7  (
            .in0(N__52509),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44035),
            .lcout(DMA_dev0_Td_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54156),
            .ce(N__39693),
            .sr(N__53334));
    defparam \u0.DMA_dev1_Tm_1_LC_7_21_0 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Tm_1_LC_7_21_0 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev1_Tm_1_LC_7_21_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.DMA_dev1_Tm_1_LC_7_21_0  (
            .in0(N__52517),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39354),
            .lcout(DMA_dev1_Tm_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54168),
            .ce(N__39544),
            .sr(N__53342));
    defparam \u0.DMA_dev1_Tm_2_LC_7_21_1 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Tm_2_LC_7_21_1 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev1_Tm_2_LC_7_21_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.DMA_dev1_Tm_2_LC_7_21_1  (
            .in0(N__34272),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52518),
            .lcout(DMA_dev1_Tm_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54168),
            .ce(N__39544),
            .sr(N__53342));
    defparam \u0.DMA_dev1_Teoc_0_LC_7_21_2 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Teoc_0_LC_7_21_2 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev1_Teoc_0_LC_7_21_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.DMA_dev1_Teoc_0_LC_7_21_2  (
            .in0(N__52512),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39883),
            .lcout(DMA_dev1_Teoc_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54168),
            .ce(N__39544),
            .sr(N__53342));
    defparam \u0.DMA_dev1_Teoc_1_LC_7_21_3 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Teoc_1_LC_7_21_3 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev1_Teoc_1_LC_7_21_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \u0.DMA_dev1_Teoc_1_LC_7_21_3  (
            .in0(_gnd_net_),
            .in1(N__40854),
            .in2(_gnd_net_),
            .in3(N__52513),
            .lcout(DMA_dev1_Teoc_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54168),
            .ce(N__39544),
            .sr(N__53342));
    defparam \u0.DMA_dev1_Teoc_2_LC_7_21_4 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Teoc_2_LC_7_21_4 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev1_Teoc_2_LC_7_21_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.DMA_dev1_Teoc_2_LC_7_21_4  (
            .in0(N__52514),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44218),
            .lcout(DMA_dev1_Teoc_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54168),
            .ce(N__39544),
            .sr(N__53342));
    defparam \u0.DMA_dev1_Teoc_4_LC_7_21_5 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Teoc_4_LC_7_21_5 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev1_Teoc_4_LC_7_21_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \u0.DMA_dev1_Teoc_4_LC_7_21_5  (
            .in0(_gnd_net_),
            .in1(N__46149),
            .in2(_gnd_net_),
            .in3(N__52515),
            .lcout(DMA_dev1_Teoc_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54168),
            .ce(N__39544),
            .sr(N__53342));
    defparam \u0.DMA_dev1_Tm_0_LC_7_21_6 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Tm_0_LC_7_21_6 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev1_Tm_0_LC_7_21_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.DMA_dev1_Tm_0_LC_7_21_6  (
            .in0(N__52516),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49534),
            .lcout(DMA_dev1_Tm_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54168),
            .ce(N__39544),
            .sr(N__53342));
    defparam \u0.DMA_dev1_Td_7_LC_7_21_7 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Td_7_LC_7_21_7 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev1_Td_7_LC_7_21_7 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.DMA_dev1_Td_7_LC_7_21_7  (
            .in0(N__34549),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52511),
            .lcout(DMA_dev1_Td_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54168),
            .ce(N__39544),
            .sr(N__53342));
    defparam \u1.DA_1_LC_7_22_0 .C_ON=1'b0;
    defparam \u1.DA_1_LC_7_22_0 .SEQ_MODE=4'b1010;
    defparam \u1.DA_1_LC_7_22_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u1.DA_1_LC_7_22_0  (
            .in0(N__52637),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25030),
            .lcout(da_pad_o_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54178),
            .ce(),
            .sr(N__53349));
    defparam \u1.RESETn_LC_7_22_1 .C_ON=1'b0;
    defparam \u1.RESETn_LC_7_22_1 .SEQ_MODE=4'b1010;
    defparam \u1.RESETn_LC_7_22_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \u1.RESETn_LC_7_22_1  (
            .in0(_gnd_net_),
            .in1(N__43286),
            .in2(_gnd_net_),
            .in3(N__52639),
            .lcout(resetn_pad_o_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54178),
            .ce(),
            .sr(N__53349));
    defparam \u1.PIO_control.gen_pingpong_dping_valid_LC_7_22_2 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_dping_valid_LC_7_22_2 .SEQ_MODE=4'b1010;
    defparam \u1.PIO_control.gen_pingpong_dping_valid_LC_7_22_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u1.PIO_control.gen_pingpong_dping_valid_LC_7_22_2  (
            .in0(N__52638),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23527),
            .lcout(\u1.PIO_control.dping_valid ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54178),
            .ce(),
            .sr(N__53349));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_fast_3_LC_7_22_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_fast_3_LC_7_22_6 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_fast_3_LC_7_22_6 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_fast_3_LC_7_22_6  (
            .in0(N__24181),
            .in1(N__23824),
            .in2(N__24257),
            .in3(N__23439),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.iQ_fast_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54178),
            .ce(),
            .sr(N__53349));
    defparam \u0.CtrlReg_0_LC_7_23_0 .C_ON=1'b0;
    defparam \u0.CtrlReg_0_LC_7_23_0 .SEQ_MODE=4'b1011;
    defparam \u0.CtrlReg_0_LC_7_23_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \u0.CtrlReg_0_LC_7_23_0  (
            .in0(_gnd_net_),
            .in1(N__52640),
            .in2(_gnd_net_),
            .in3(N__49544),
            .lcout(IDEctrl_rst),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54190),
            .ce(N__53514),
            .sr(N__53354));
    defparam \u0.CtrlReg_13_LC_7_23_1 .C_ON=1'b0;
    defparam \u0.CtrlReg_13_LC_7_23_1 .SEQ_MODE=4'b1010;
    defparam \u0.CtrlReg_13_LC_7_23_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.CtrlReg_13_LC_7_23_1  (
            .in0(N__34704),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52645),
            .lcout(DMActrl_dir),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54190),
            .ce(N__53514),
            .sr(N__53354));
    defparam \u0.CtrlReg_15_LC_7_23_2 .C_ON=1'b0;
    defparam \u0.CtrlReg_15_LC_7_23_2 .SEQ_MODE=4'b1010;
    defparam \u0.CtrlReg_15_LC_7_23_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \u0.CtrlReg_15_LC_7_23_2  (
            .in0(_gnd_net_),
            .in1(N__52641),
            .in2(_gnd_net_),
            .in3(N__34550),
            .lcout(DMActrl_DMAen),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54190),
            .ce(N__53514),
            .sr(N__53354));
    defparam \u0.CtrlReg_4_LC_7_23_3 .C_ON=1'b0;
    defparam \u0.CtrlReg_4_LC_7_23_3 .SEQ_MODE=4'b1010;
    defparam \u0.CtrlReg_4_LC_7_23_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.CtrlReg_4_LC_7_23_3  (
            .in0(N__37233),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52646),
            .lcout(IDEctrl_ppen),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54190),
            .ce(N__53514),
            .sr(N__53354));
    defparam \u0.CtrlReg_5_LC_7_23_4 .C_ON=1'b0;
    defparam \u0.CtrlReg_5_LC_7_23_4 .SEQ_MODE=4'b1010;
    defparam \u0.CtrlReg_5_LC_7_23_4 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.CtrlReg_5_LC_7_23_4  (
            .in0(N__46264),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52642),
            .lcout(IDEctrl_FATR0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54190),
            .ce(N__53514),
            .sr(N__53354));
    defparam \u0.CtrlReg_6_LC_7_23_5 .C_ON=1'b0;
    defparam \u0.CtrlReg_6_LC_7_23_5 .SEQ_MODE=4'b1010;
    defparam \u0.CtrlReg_6_LC_7_23_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.CtrlReg_6_LC_7_23_5  (
            .in0(N__39471),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52647),
            .lcout(IDEctrl_FATR1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54190),
            .ce(N__53514),
            .sr(N__53354));
    defparam \u0.CtrlReg_7_LC_7_23_6 .C_ON=1'b0;
    defparam \u0.CtrlReg_7_LC_7_23_6 .SEQ_MODE=4'b1010;
    defparam \u0.CtrlReg_7_LC_7_23_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \u0.CtrlReg_7_LC_7_23_6  (
            .in0(_gnd_net_),
            .in1(N__52643),
            .in2(_gnd_net_),
            .in3(N__39650),
            .lcout(IDEctrl_IDEen),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54190),
            .ce(N__53514),
            .sr(N__53354));
    defparam \u0.CtrlReg_9_LC_7_23_7 .C_ON=1'b0;
    defparam \u0.CtrlReg_9_LC_7_23_7 .SEQ_MODE=4'b1010;
    defparam \u0.CtrlReg_9_LC_7_23_7 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \u0.CtrlReg_9_LC_7_23_7  (
            .in0(N__52644),
            .in1(_gnd_net_),
            .in2(N__36018),
            .in3(_gnd_net_),
            .lcout(DMActrl_BeLeC1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54190),
            .ce(N__53514),
            .sr(N__53354));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_RNIM9N61_5_3_LC_7_24_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_RNIM9N61_5_3_LC_7_24_0 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_RNIM9N61_5_3_LC_7_24_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_RNIM9N61_5_3_LC_7_24_0  (
            .in0(N__24108),
            .in1(N__24147),
            .in2(N__24261),
            .in3(N__24300),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_awe0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_2_LC_7_24_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_2_LC_7_24_1 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_2_LC_7_24_1 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_2_LC_7_24_1  (
            .in0(N__24301),
            .in1(N__24251),
            .in2(N__24168),
            .in3(N__23753),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.wr_ptr_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54201),
            .ce(),
            .sr(N__53361));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_RNO_0_1_LC_7_24_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_RNO_0_1_LC_7_24_2 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_RNO_0_1_LC_7_24_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_RNO_0_1_LC_7_24_2  (
            .in0(_gnd_net_),
            .in1(N__24106),
            .in2(_gnd_net_),
            .in3(N__24146),
            .lcout(),
            .ltout(\u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.N_1385_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_1_LC_7_24_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_1_LC_7_24_3 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_1_LC_7_24_3 .LUT_INIT=16'b0000000000101110;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_1_LC_7_24_3  (
            .in0(N__24303),
            .in1(N__24252),
            .in2(N__23881),
            .in3(N__23752),
            .lcout(\u1.DMA_control.wr_ptr_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54201),
            .ce(),
            .sr(N__53361));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_3_LC_7_24_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_3_LC_7_24_4 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_3_LC_7_24_4 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_3_LC_7_24_4  (
            .in0(N__23754),
            .in1(N__24107),
            .in2(N__24262),
            .in3(N__24148),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.wr_ptr_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54201),
            .ce(),
            .sr(N__53361));
    defparam \u1.DMA_control.N_101_i_i_o2_LC_7_24_5 .C_ON=1'b0;
    defparam \u1.DMA_control.N_101_i_i_o2_LC_7_24_5 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.N_101_i_i_o2_LC_7_24_5 .LUT_INIT=16'b1110111011101110;
    LogicCell40 \u1.DMA_control.N_101_i_i_o2_LC_7_24_5  (
            .in0(N__52651),
            .in1(N__43285),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\u1.DMA_control.N_1326 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_fast_2_LC_7_24_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_fast_2_LC_7_24_7 .SEQ_MODE=4'b1010;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_fast_2_LC_7_24_7 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_fast_2_LC_7_24_7  (
            .in0(N__24302),
            .in1(N__23755),
            .in2(N__23713),
            .in3(N__24256),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.iQ_fast_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54201),
            .ce(),
            .sr(N__53361));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIG7GT_18_LC_7_25_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIG7GT_18_LC_7_25_0 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIG7GT_18_LC_7_25_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIG7GT_18_LC_7_25_0  (
            .in0(N__45337),
            .in1(N__23689),
            .in2(_gnd_net_),
            .in3(N__24646),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIG7GTZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__2_LC_7_25_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__2_LC_7_25_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__2_LC_7_25_2 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__2_LC_7_25_2  (
            .in0(N__30479),
            .in1(N__30337),
            .in2(N__42964),
            .in3(_gnd_net_),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54214),
            .ce(N__41798),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNII9GT_19_LC_7_25_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNII9GT_19_LC_7_25_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNII9GT_19_LC_7_25_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNII9GT_19_LC_7_25_3  (
            .in0(N__27280),
            .in1(N__23680),
            .in2(_gnd_net_),
            .in3(N__45338),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNII9GTZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__19_LC_7_25_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__19_LC_7_25_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__19_LC_7_25_4 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__19_LC_7_25_4  (
            .in0(N__36552),
            .in1(_gnd_net_),
            .in2(N__42963),
            .in3(N__36436),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54214),
            .ce(N__41798),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.valid_RNIM6GI3_LC_7_25_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.valid_RNIM6GI3_LC_7_25_5 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.valid_RNIM6GI3_LC_7_25_5 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Txbuf.valid_RNIM6GI3_LC_7_25_5  (
            .in0(N__50831),
            .in1(N__47245),
            .in2(_gnd_net_),
            .in3(N__31442),
            .lcout(\u1.DMA_control.gen_DMAbuf_Txbuf.N_1602 ),
            .ltout(\u1.DMA_control.gen_DMAbuf_Txbuf.N_1602_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.valid_RNI2KL74_LC_7_25_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.valid_RNI2KL74_LC_7_25_6 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.valid_RNI2KL74_LC_7_25_6 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Txbuf.valid_RNI2KL74_LC_7_25_6  (
            .in0(N__52652),
            .in1(_gnd_net_),
            .in2(N__24076),
            .in3(N__43290),
            .lcout(\u1.DMA_control.gen_DMAbuf_Txbuf.N_319 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__3_LC_7_25_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__3_LC_7_25_7 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__3_LC_7_25_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__3_LC_7_25_7  (
            .in0(N__36437),
            .in1(N__42746),
            .in2(_gnd_net_),
            .in3(N__36553),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54214),
            .ce(N__41798),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_13_LC_7_26_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_13_LC_7_26_0 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_13_LC_7_26_0 .LUT_INIT=16'b0000001101010011;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_13_LC_7_26_0  (
            .in0(N__42767),
            .in1(N__24055),
            .in2(N__25622),
            .in3(N__24043),
            .lcout(\u1.DMA_control.writeDfw_6_i_m2_i_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNIA9TN_6_LC_7_26_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNIA9TN_6_LC_7_26_1 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNIA9TN_6_LC_7_26_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNIA9TN_6_LC_7_26_1  (
            .in0(N__45339),
            .in1(N__24019),
            .in2(_gnd_net_),
            .in3(N__25924),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNIA9TNZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_10_LC_7_26_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_10_LC_7_26_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_10_LC_7_26_3 .LUT_INIT=16'b0000001101010011;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_10_LC_7_26_3  (
            .in0(N__24007),
            .in1(N__23986),
            .in2(N__25619),
            .in3(N__42784),
            .lcout(\u1.DMA_control.writeDfw_6_i_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_Td_5_LC_7_26_5 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_Td_5_LC_7_26_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.DMA_timing_ctrl_Td_5_LC_7_26_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_Td_5_LC_7_26_5  (
            .in0(N__31533),
            .in1(N__25047),
            .in2(_gnd_net_),
            .in3(N__36291),
            .lcout(\u1.DMA_control.Td_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54228),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_9_LC_7_27_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_9_LC_7_27_0 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_9_LC_7_27_0 .LUT_INIT=16'b0001000100001111;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_9_LC_7_27_0  (
            .in0(N__42711),
            .in1(N__23955),
            .in2(N__23938),
            .in3(N__25620),
            .lcout(),
            .ltout(\u1.DMA_control.writeDfw_6_i_0_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_9_LC_7_27_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_9_LC_7_27_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_9_LC_7_27_1 .LUT_INIT=16'b0000110100001111;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDfw_9_LC_7_27_1  (
            .in0(N__25621),
            .in1(N__23926),
            .in2(N__23899),
            .in3(N__42712),
            .lcout(\u1.DMAd_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54239),
            .ce(N__25395),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_RNIM9N61_0_3_LC_7_27_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_RNIM9N61_0_3_LC_7_27_2 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_RNIM9N61_0_3_LC_7_27_2 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_RNIM9N61_0_3_LC_7_27_2  (
            .in0(N__24122),
            .in1(N__24169),
            .in2(N__24259),
            .in3(N__24306),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_awe5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_RNIM9N61_1_3_LC_7_27_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_RNIM9N61_1_3_LC_7_27_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_RNIM9N61_1_3_LC_7_27_3 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_RNIM9N61_1_3_LC_7_27_3  (
            .in0(N__24304),
            .in1(N__24239),
            .in2(N__24182),
            .in3(N__24123),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_awe4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_RNIM9N61_2_3_LC_7_27_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_RNIM9N61_2_3_LC_7_27_4 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_RNIM9N61_2_3_LC_7_27_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_RNIM9N61_2_3_LC_7_27_4  (
            .in0(N__24124),
            .in1(N__24173),
            .in2(N__24260),
            .in3(N__24308),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_awe3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_RNIM9N61_3_LC_7_27_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_RNIM9N61_3_LC_7_27_5 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_RNIM9N61_3_LC_7_27_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_RNIM9N61_3_LC_7_27_5  (
            .in0(N__24307),
            .in1(N__24243),
            .in2(N__24183),
            .in3(N__24126),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_awe6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_RNIM9N61_3_3_LC_7_27_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_RNIM9N61_3_3_LC_7_27_6 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_RNIM9N61_3_3_LC_7_27_6 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_RNIM9N61_3_3_LC_7_27_6  (
            .in0(N__24125),
            .in1(N__24174),
            .in2(N__24258),
            .in3(N__24305),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_awe2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_RNIM9N61_4_3_LC_7_27_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_RNIM9N61_4_3_LC_7_27_7 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_RNIM9N61_4_3_LC_7_27_7 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.wr_ptr_lfsr.iQ_RNIM9N61_4_3_LC_7_27_7  (
            .in0(N__24309),
            .in1(N__24247),
            .in2(N__24184),
            .in3(N__24127),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_awe1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI099K_21_LC_7_28_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI099K_21_LC_7_28_0 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI099K_21_LC_7_28_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI099K_21_LC_7_28_0  (
            .in0(N__27256),
            .in1(N__24088),
            .in2(_gnd_net_),
            .in3(N__45492),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI099KZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__21_LC_7_28_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__21_LC_7_28_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__21_LC_7_28_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__21_LC_7_28_1  (
            .in0(N__42852),
            .in1(N__35669),
            .in2(_gnd_net_),
            .in3(N__35558),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54254),
            .ce(N__30766),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__5_LC_7_28_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__5_LC_7_28_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__5_LC_7_28_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__5_LC_7_28_2  (
            .in0(N__35559),
            .in1(N__35670),
            .in2(_gnd_net_),
            .in3(N__42855),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54254),
            .ce(N__30766),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI4N4N_5_LC_7_28_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI4N4N_5_LC_7_28_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI4N4N_5_LC_7_28_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI4N4N_5_LC_7_28_3  (
            .in0(N__45494),
            .in1(N__25933),
            .in2(_gnd_net_),
            .in3(N__24082),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI4N4NZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI0J4N_3_LC_7_28_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI0J4N_3_LC_7_28_4 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI0J4N_3_LC_7_28_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI0J4N_3_LC_7_28_4  (
            .in0(N__24352),
            .in1(N__25891),
            .in2(_gnd_net_),
            .in3(N__45493),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI0J4NZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__3_LC_7_28_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__3_LC_7_28_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__3_LC_7_28_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__3_LC_7_28_5  (
            .in0(N__42853),
            .in1(_gnd_net_),
            .in2(N__36439),
            .in3(N__36551),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54254),
            .ce(N__30766),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__19_LC_7_28_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__19_LC_7_28_6 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__19_LC_7_28_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__19_LC_7_28_6  (
            .in0(N__36550),
            .in1(N__36431),
            .in2(_gnd_net_),
            .in3(N__42854),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54254),
            .ce(N__30766),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIEL7K_19_LC_7_28_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIEL7K_19_LC_7_28_7 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIEL7K_19_LC_7_28_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIEL7K_19_LC_7_28_7  (
            .in0(N__45495),
            .in1(N__27244),
            .in2(_gnd_net_),
            .in3(N__24346),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIEL7KZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIQPOD1_6_LC_7_29_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIQPOD1_6_LC_7_29_2 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIQPOD1_6_LC_7_29_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIQPOD1_6_LC_7_29_2  (
            .in0(N__24328),
            .in1(N__24340),
            .in2(_gnd_net_),
            .in3(N__50052),
            .lcout(),
            .ltout(mem_mem_ram6__RNIQPOD1_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.dat_o_0_0_a2_1_6_LC_7_29_3 .C_ON=1'b0;
    defparam \u0.dat_o_0_0_a2_1_6_LC_7_29_3 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_0_0_a2_1_6_LC_7_29_3 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \u0.dat_o_0_0_a2_1_6_LC_7_29_3  (
            .in0(N__47255),
            .in1(N__31237),
            .in2(N__24331),
            .in3(N__48813),
            .lcout(\u0.N_1971 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__6_LC_7_29_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__6_LC_7_29_6 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__6_LC_7_29_6 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__6_LC_7_29_6  (
            .in0(_gnd_net_),
            .in1(N__42763),
            .in2(N__32716),
            .in3(N__32820),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54266),
            .ce(N__41246),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__22_LC_7_29_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__22_LC_7_29_7 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__22_LC_7_29_7 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__22_LC_7_29_7  (
            .in0(N__32819),
            .in1(N__32707),
            .in2(N__42966),
            .in3(_gnd_net_),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54266),
            .ce(N__41246),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport0_T2_3_LC_7_30_1 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T2_3_LC_7_30_1 .SEQ_MODE=4'b1011;
    defparam \u0.PIO_dport0_T2_3_LC_7_30_1 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \u0.PIO_dport0_T2_3_LC_7_30_1  (
            .in0(N__43627),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52763),
            .lcout(PIO_dport0_T2_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54276),
            .ce(N__49384),
            .sr(N__53399));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__18_LC_7_31_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__18_LC_7_31_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__18_LC_7_31_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__18_LC_7_31_4  (
            .in0(N__30480),
            .in1(N__30309),
            .in2(_gnd_net_),
            .in3(N__42960),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54286),
            .ce(N__28291),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_Tm_1_LC_9_13_7 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_Tm_1_LC_9_13_7 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.DMA_timing_ctrl_Tm_1_LC_9_13_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_Tm_1_LC_9_13_7  (
            .in0(N__31762),
            .in1(N__44691),
            .in2(_gnd_net_),
            .in3(N__36282),
            .lcout(\u1.DMA_control.Tm_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54191),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_cmdport_T1_2_LC_9_14_5 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_T1_2_LC_9_14_5 .SEQ_MODE=4'b1011;
    defparam \u0.PIO_cmdport_T1_2_LC_9_14_5 .LUT_INIT=16'b1110111011101110;
    LogicCell40 \u0.PIO_cmdport_T1_2_LC_9_14_5  (
            .in0(N__51907),
            .in1(N__34241),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(PIO_cmdport_T1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54179),
            .ce(N__49699),
            .sr(N__53335));
    defparam \u1.PIO_control.PIO_access_control.T1_0_LC_9_16_1 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T1_0_LC_9_16_1 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.T1_0_LC_9_16_1 .LUT_INIT=16'b0000000010111011;
    LogicCell40 \u1.PIO_control.PIO_access_control.T1_0_LC_9_16_1  (
            .in0(N__49417),
            .in1(N__29090),
            .in2(_gnd_net_),
            .in3(N__25981),
            .lcout(\u1.PIO_control.PIO_access_control.T1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54157),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dstrb_LC_9_16_5 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dstrb_LC_9_16_5 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.dstrb_LC_9_16_5 .LUT_INIT=16'b0000000010111011;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.dstrb_LC_9_16_5  (
            .in0(N__24607),
            .in1(N__24565),
            .in2(_gnd_net_),
            .in3(N__24520),
            .lcout(\u1.PIO_control.PIO_access_control.dstrb ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54157),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T1_2_LC_9_17_0 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T1_2_LC_9_17_0 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.T1_2_LC_9_17_0 .LUT_INIT=16'b0000000010111011;
    LogicCell40 \u1.PIO_control.PIO_access_control.T1_2_LC_9_17_0  (
            .in0(N__31701),
            .in1(N__29061),
            .in2(_gnd_net_),
            .in3(N__26149),
            .lcout(\u1.PIO_control.PIO_access_control.T1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54145),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T1_4_LC_9_17_1 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T1_4_LC_9_17_1 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.T1_4_LC_9_17_1 .LUT_INIT=16'b0000000011011101;
    LogicCell40 \u1.PIO_control.PIO_access_control.T1_4_LC_9_17_1  (
            .in0(N__29062),
            .in1(N__36064),
            .in2(_gnd_net_),
            .in3(N__24652),
            .lcout(\u1.PIO_control.PIO_access_control.T1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54145),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.c_state_RNO_0_1_LC_9_17_3 .C_ON=1'b0;
    defparam \u1.c_state_RNO_0_1_LC_9_17_3 .SEQ_MODE=4'b0000;
    defparam \u1.c_state_RNO_0_1_LC_9_17_3 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \u1.c_state_RNO_0_1_LC_9_17_3  (
            .in0(N__52106),
            .in1(N__24454),
            .in2(_gnd_net_),
            .in3(N__24403),
            .lcout(\u1.c_state_ns_i_i_i_a2_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.dat_o_0_a2_i_a2_4_16_LC_9_17_5 .C_ON=1'b0;
    defparam \u0.dat_o_0_a2_i_a2_4_16_LC_9_17_5 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_0_a2_i_a2_4_16_LC_9_17_5 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \u0.dat_o_0_a2_i_a2_4_16_LC_9_17_5  (
            .in0(N__47735),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53066),
            .lcout(\u0.N_2101 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_7_LC_9_18_0 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_7_LC_9_18_0 .SEQ_MODE=4'b1010;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_7_LC_9_18_0 .LUT_INIT=16'b0011101100001000;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_7_LC_9_18_0  (
            .in0(N__27343),
            .in1(N__24835),
            .in2(N__52243),
            .in3(N__24796),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.QiZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54158),
            .ce(N__24760),
            .sr(N__53336));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNI9LFI_1_LC_9_18_1 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNI9LFI_1_LC_9_18_1 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNI9LFI_1_LC_9_18_1 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNI9LFI_1_LC_9_18_1  (
            .in0(N__28850),
            .in1(N__28814),
            .in2(N__24723),
            .in3(N__28913),
            .lcout(),
            .ltout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNI9LFIZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNI7F9K_0_LC_9_18_2 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNI7F9K_0_LC_9_18_2 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNI7F9K_0_LC_9_18_2 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNI7F9K_0_LC_9_18_2  (
            .in0(N__28706),
            .in1(_gnd_net_),
            .in2(N__24691),
            .in3(N__28943),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.Qi_RNI7F9K_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNO_0_0_LC_9_18_3 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNO_0_0_LC_9_18_3 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNO_0_0_LC_9_18_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNO_0_0_LC_9_18_3  (
            .in0(N__28944),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28707),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_s_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNICS77_7_LC_9_18_4 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNICS77_7_LC_9_18_4 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNICS77_7_LC_9_18_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNICS77_7_LC_9_18_4  (
            .in0(N__28743),
            .in1(N__28782),
            .in2(N__29562),
            .in3(N__28884),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.val_c8_0_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T1_RNO_0_4_LC_9_18_6 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T1_RNO_0_4_LC_9_18_6 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.T1_RNO_0_4_LC_9_18_6 .LUT_INIT=16'b0011101100001010;
    LogicCell40 \u1.PIO_control.PIO_access_control.T1_RNO_0_4_LC_9_18_6  (
            .in0(N__29257),
            .in1(N__27772),
            .in2(N__29872),
            .in3(N__29388),
            .lcout(\u1.PIO_control.PIO_access_control.it1_1_iv_0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_pong_a_1_LC_9_19_1 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_pong_a_1_LC_9_19_1 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_pong_a_1_LC_9_19_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \u1.PIO_control.gen_pingpong_pong_a_1_LC_9_19_1  (
            .in0(N__47700),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\u1.PIO_control.pong_a_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54169),
            .ce(N__24895),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_pong_a_RNIV0V01_1_LC_9_19_2 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_pong_a_RNIV0V01_1_LC_9_19_2 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.gen_pingpong_pong_a_RNIV0V01_1_LC_9_19_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.PIO_control.gen_pingpong_pong_a_RNIV0V01_1_LC_9_19_2  (
            .in0(N__26575),
            .in1(N__26273),
            .in2(_gnd_net_),
            .in3(N__26794),
            .lcout(\u1.N_1423 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_pong_a_RNI914A1_0_LC_9_19_3 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_pong_a_RNI914A1_0_LC_9_19_3 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.gen_pingpong_pong_a_RNI914A1_0_LC_9_19_3 .LUT_INIT=16'b1110111011100100;
    LogicCell40 \u1.PIO_control.gen_pingpong_pong_a_RNI914A1_0_LC_9_19_3  (
            .in0(N__26793),
            .in1(N__26415),
            .in2(N__26404),
            .in3(N__26991),
            .lcout(),
            .ltout(\u1.PIO_control.pong_a_RNI914A1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_pong_a_RNIL58K2_3_LC_9_19_4 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_pong_a_RNIL58K2_3_LC_9_19_4 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.gen_pingpong_pong_a_RNIL58K2_3_LC_9_19_4 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \u1.PIO_control.gen_pingpong_pong_a_RNIL58K2_3_LC_9_19_4  (
            .in0(_gnd_net_),
            .in1(N__27006),
            .in2(N__24904),
            .in3(N__24901),
            .lcout(\u1.PIO_control.N_1315 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_pong_a_3_LC_9_19_5 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_pong_a_3_LC_9_19_5 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_pong_a_3_LC_9_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.PIO_control.gen_pingpong_pong_a_3_LC_9_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50458),
            .lcout(\u1.PIO_control.pong_a_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54169),
            .ce(N__24895),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_ping_a_RNIQNVQ_0_LC_9_19_6 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_ping_a_RNIQNVQ_0_LC_9_19_6 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.gen_pingpong_ping_a_RNIQNVQ_0_LC_9_19_6 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \u1.PIO_control.gen_pingpong_ping_a_RNIQNVQ_0_LC_9_19_6  (
            .in0(N__26990),
            .in1(N__26399),
            .in2(_gnd_net_),
            .in3(N__26792),
            .lcout(\u1.PIO_control.ping_a_RNIQNVQ_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_pong_a_0_LC_9_19_7 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_pong_a_0_LC_9_19_7 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_pong_a_0_LC_9_19_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \u1.PIO_control.gen_pingpong_pong_a_0_LC_9_19_7  (
            .in0(N__50573),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\u1.pong_a_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54169),
            .ce(N__24895),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_ping_a_0_LC_9_20_0 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_ping_a_0_LC_9_20_0 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_ping_a_0_LC_9_20_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \u1.PIO_control.gen_pingpong_ping_a_0_LC_9_20_0  (
            .in0(N__50574),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\u1.ping_a_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54180),
            .ce(N__25087),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_ping_a_1_LC_9_20_1 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_ping_a_1_LC_9_20_1 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_ping_a_1_LC_9_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.PIO_control.gen_pingpong_ping_a_1_LC_9_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47737),
            .lcout(\u1.PIO_control.ping_a_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54180),
            .ce(N__25087),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_ping_a_2_LC_9_20_2 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_ping_a_2_LC_9_20_2 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_ping_a_2_LC_9_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.PIO_control.gen_pingpong_ping_a_2_LC_9_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53067),
            .lcout(\u1.ping_a_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54180),
            .ce(N__25087),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_ping_a_3_LC_9_20_3 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_ping_a_3_LC_9_20_3 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_ping_a_3_LC_9_20_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \u1.PIO_control.gen_pingpong_ping_a_3_LC_9_20_3  (
            .in0(N__50459),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\u1.PIO_control.ping_a_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54180),
            .ce(N__25087),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_ping_d_0_LC_9_20_4 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_ping_d_0_LC_9_20_4 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_ping_d_0_LC_9_20_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.PIO_control.gen_pingpong_ping_d_0_LC_9_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49526),
            .lcout(\u1.PIO_control.ping_d_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54180),
            .ce(N__25087),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_ping_d_1_LC_9_20_5 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_ping_d_1_LC_9_20_5 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_ping_d_1_LC_9_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.PIO_control.gen_pingpong_ping_d_1_LC_9_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39353),
            .lcout(\u1.PIO_control.ping_d_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54180),
            .ce(N__25087),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_ping_d_10_LC_9_20_6 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_ping_d_10_LC_9_20_6 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_ping_d_10_LC_9_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.PIO_control.gen_pingpong_ping_d_10_LC_9_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40168),
            .lcout(\u1.PIO_control.ping_d_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54180),
            .ce(N__25087),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_ping_d_11_LC_9_20_7 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_ping_d_11_LC_9_20_7 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.gen_pingpong_ping_d_11_LC_9_20_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \u1.PIO_control.gen_pingpong_ping_d_11_LC_9_20_7  (
            .in0(N__43672),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\u1.PIO_control.ping_d_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54180),
            .ce(N__25087),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev1_Td_RNI9BOI3_3_LC_9_21_0 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Td_RNI9BOI3_3_LC_9_21_0 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev1_Td_RNI9BOI3_3_LC_9_21_0 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \u0.DMA_dev1_Td_RNI9BOI3_3_LC_9_21_0  (
            .in0(N__54714),
            .in1(N__31287),
            .in2(N__50767),
            .in3(N__27427),
            .lcout(\u0.dat_o_0_0_3_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev1_Td_RNIDFOI3_5_LC_9_21_1 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Td_RNIDFOI3_5_LC_9_21_1 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev1_Td_RNIDFOI3_5_LC_9_21_1 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \u0.DMA_dev1_Td_RNIDFOI3_5_LC_9_21_1  (
            .in0(N__31537),
            .in1(N__54715),
            .in2(N__34597),
            .in3(N__50765),
            .lcout(\u0.dat_o_0_0_3_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport1_T2_RNIDFO24_5_LC_9_21_3 .C_ON=1'b0;
    defparam \u0.PIO_dport1_T2_RNIDFO24_5_LC_9_21_3 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport1_T2_RNIDFO24_5_LC_9_21_3 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \u0.PIO_dport1_T2_RNIDFO24_5_LC_9_21_3  (
            .in0(N__46979),
            .in1(N__31507),
            .in2(N__25054),
            .in3(N__48598),
            .lcout(\u0.dat_o_0_0_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.SelDev_RNO_0_LC_9_21_4 .C_ON=1'b0;
    defparam \u1.PIO_control.SelDev_RNO_0_LC_9_21_4 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.SelDev_RNO_0_LC_9_21_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \u1.PIO_control.SelDev_RNO_0_LC_9_21_4  (
            .in0(N__25026),
            .in1(N__26365),
            .in2(N__25012),
            .in3(N__26683),
            .lcout(),
            .ltout(\u1.PIO_control.SelDev_e_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.SelDev_LC_9_21_5 .C_ON=1'b0;
    defparam \u1.PIO_control.SelDev_LC_9_21_5 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.SelDev_LC_9_21_5 .LUT_INIT=16'b1100110010101100;
    LogicCell40 \u1.PIO_control.SelDev_LC_9_21_5  (
            .in0(N__24997),
            .in1(N__36208),
            .in2(N__24976),
            .in3(N__26308),
            .lcout(\u1.SelDev ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54192),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.CtrlReg_RNIMPDE2_15_LC_9_22_0 .C_ON=1'b0;
    defparam \u0.CtrlReg_RNIMPDE2_15_LC_9_22_0 .SEQ_MODE=4'b0000;
    defparam \u0.CtrlReg_RNIMPDE2_15_LC_9_22_0 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \u0.CtrlReg_RNIMPDE2_15_LC_9_22_0  (
            .in0(N__25144),
            .in1(N__48333),
            .in2(N__47510),
            .in3(N__24971),
            .lcout(),
            .ltout(\u0.dat_o_0_0_2_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev0_Td_RNIM4E99_7_LC_9_22_1 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Td_RNIM4E99_7_LC_9_22_1 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev0_Td_RNIM4E99_7_LC_9_22_1 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \u0.DMA_dev0_Td_RNIM4E99_7_LC_9_22_1  (
            .in0(N__25156),
            .in1(N__48566),
            .in2(N__24931),
            .in3(N__24928),
            .lcout(),
            .ltout(\u0.dat_o_0_0_5_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev1_Td_RNI1H6KI_7_LC_9_22_2 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Td_RNI1H6KI_7_LC_9_22_2 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev1_Td_RNI1H6KI_7_LC_9_22_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \u0.DMA_dev1_Td_RNI1H6KI_7_LC_9_22_2  (
            .in0(N__25198),
            .in1(N__31348),
            .in2(N__25186),
            .in3(N__34384),
            .lcout(wb_dat_o_c_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIAVA71_15_LC_9_22_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIAVA71_15_LC_9_22_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIAVA71_15_LC_9_22_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIAVA71_15_LC_9_22_3  (
            .in0(N__27097),
            .in1(N__27109),
            .in2(_gnd_net_),
            .in3(N__49915),
            .lcout(),
            .ltout(mem_mem_ram6__RNIAVA71_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.dat_o_0_0_a2_0_15_LC_9_22_4 .C_ON=1'b0;
    defparam \u0.dat_o_0_0_a2_0_15_LC_9_22_4 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_0_0_a2_0_15_LC_9_22_4 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \u0.dat_o_0_0_a2_0_15_LC_9_22_4  (
            .in0(N__25150),
            .in1(N__47220),
            .in2(N__25159),
            .in3(N__48829),
            .lcout(\u0.N_2029 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIQGDM1_2_LC_9_22_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIQGDM1_2_LC_9_22_5 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIQGDM1_2_LC_9_22_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIQGDM1_2_LC_9_22_5  (
            .in0(N__28039),
            .in1(N__25957),
            .in2(_gnd_net_),
            .in3(N__49916),
            .lcout(iQ_RNIQGDM1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.q_15_LC_9_22_6 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.q_15_LC_9_22_6 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.q_15_LC_9_22_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \u1.PIO_control.PIO_access_control.q_15_LC_9_22_6  (
            .in0(N__32382),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(PIOq_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54202),
            .ce(N__45880),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIA1EM1_2_LC_9_23_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIA1EM1_2_LC_9_23_0 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIA1EM1_2_LC_9_23_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIA1EM1_2_LC_9_23_0  (
            .in0(N__50037),
            .in1(N__25138),
            .in2(_gnd_net_),
            .in3(N__25120),
            .lcout(),
            .ltout(iQ_RNIA1EM1_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.dat_o_i_0_a2_19_LC_9_23_1 .C_ON=1'b0;
    defparam \u0.dat_o_i_0_a2_19_LC_9_23_1 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_i_0_a2_19_LC_9_23_1 .LUT_INIT=16'b0010001000001010;
    LogicCell40 \u0.dat_o_i_0_a2_19_LC_9_23_1  (
            .in0(N__50467),
            .in1(N__25276),
            .in2(N__25123),
            .in3(N__48858),
            .lcout(\u0.N_1724 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.CtrlReg_19_LC_9_23_2 .C_ON=1'b0;
    defparam \u0.CtrlReg_19_LC_9_23_2 .SEQ_MODE=4'b1010;
    defparam \u0.CtrlReg_19_LC_9_23_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.CtrlReg_19_LC_9_23_2  (
            .in0(N__34358),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52244),
            .lcout(\u0.CtrlRegZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54215),
            .ce(N__53513),
            .sr(N__53369));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIA1VQ_19_LC_9_23_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIA1VQ_19_LC_9_23_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIA1VQ_19_LC_9_23_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIA1VQ_19_LC_9_23_3  (
            .in0(N__45340),
            .in1(N__27211),
            .in2(_gnd_net_),
            .in3(N__27151),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIA1VQZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIMBB71_19_LC_9_23_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIMBB71_19_LC_9_23_4 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIMBB71_19_LC_9_23_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIMBB71_19_LC_9_23_4  (
            .in0(N__50036),
            .in1(N__28093),
            .in2(_gnd_net_),
            .in3(N__25294),
            .lcout(mem_mem_ram6__RNIMBB71_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.CtrlReg_RNI9DKU1_19_LC_9_23_5 .C_ON=1'b0;
    defparam \u0.CtrlReg_RNI9DKU1_19_LC_9_23_5 .SEQ_MODE=4'b0000;
    defparam \u0.CtrlReg_RNI9DKU1_19_LC_9_23_5 .LUT_INIT=16'b0100010011110100;
    LogicCell40 \u0.CtrlReg_RNI9DKU1_19_LC_9_23_5  (
            .in0(N__25270),
            .in1(N__44995),
            .in2(N__44935),
            .in3(N__29599),
            .lcout(),
            .ltout(\u0.dat_o_i_0_2_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport0_T4_RNI59JO9_3_LC_9_23_6 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T4_RNI59JO9_3_LC_9_23_6 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport0_T4_RNI59JO9_3_LC_9_23_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \u0.PIO_dport0_T4_RNI59JO9_3_LC_9_23_6  (
            .in0(N__49645),
            .in1(N__34426),
            .in2(N__25264),
            .in3(N__25261),
            .lcout(N_327_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_12_LC_9_24_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_12_LC_9_24_0 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_12_LC_9_24_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_readDlw_12_LC_9_24_0  (
            .in0(N__25230),
            .in1(N__29810),
            .in2(_gnd_net_),
            .in3(N__42956),
            .lcout(\u1.DMA_control.readDlw_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54229),
            .ce(N__36326),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_12_LC_9_24_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_12_LC_9_24_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_12_LC_9_24_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_readDfw_12_LC_9_24_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32162),
            .lcout(\u1.DMA_control.readDfw_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54229),
            .ce(N__36326),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_4_LC_9_24_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_4_LC_9_24_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_4_LC_9_24_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_readDlw_4_LC_9_24_2  (
            .in0(N__25231),
            .in1(N__29811),
            .in2(_gnd_net_),
            .in3(N__42958),
            .lcout(\u1.DMA_control.readDlw_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54229),
            .ce(N__36326),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_4_LC_9_24_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_4_LC_9_24_3 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_4_LC_9_24_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_readDfw_4_LC_9_24_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30979),
            .lcout(\u1.DMA_control.readDfw_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54229),
            .ce(N__36326),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_13_LC_9_24_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_13_LC_9_24_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_13_LC_9_24_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_readDlw_13_LC_9_24_4  (
            .in0(N__31862),
            .in1(N__34025),
            .in2(_gnd_net_),
            .in3(N__42957),
            .lcout(\u1.DMA_control.readDlw_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54229),
            .ce(N__36326),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_13_LC_9_24_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_13_LC_9_24_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_13_LC_9_24_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_readDfw_13_LC_9_24_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33524),
            .lcout(\u1.DMA_control.readDfw_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54229),
            .ce(N__36326),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_5_LC_9_24_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_5_LC_9_24_6 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_5_LC_9_24_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_readDlw_5_LC_9_24_6  (
            .in0(N__31863),
            .in1(N__34026),
            .in2(_gnd_net_),
            .in3(N__42959),
            .lcout(\u1.DMA_control.readDlw_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54229),
            .ce(N__36326),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI2RHT_20_LC_9_25_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI2RHT_20_LC_9_25_0 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI2RHT_20_LC_9_25_0 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI2RHT_20_LC_9_25_0  (
            .in0(N__25345),
            .in1(N__25354),
            .in2(N__45549),
            .in3(_gnd_net_),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI2RHTZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__20_LC_9_25_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__20_LC_9_25_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__20_LC_9_25_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__20_LC_9_25_1  (
            .in0(N__30954),
            .in1(N__30861),
            .in2(_gnd_net_),
            .in3(N__42735),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54240),
            .ce(N__41854),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__4_LC_9_25_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__4_LC_9_25_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__4_LC_9_25_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__4_LC_9_25_2  (
            .in0(N__42734),
            .in1(N__30955),
            .in2(_gnd_net_),
            .in3(N__30862),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54240),
            .ce(N__41854),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI4THT_21_LC_9_25_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI4THT_21_LC_9_25_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI4THT_21_LC_9_25_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI4THT_21_LC_9_25_3  (
            .in0(N__25900),
            .in1(N__45430),
            .in2(_gnd_net_),
            .in3(N__25339),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI4THTZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__21_LC_9_25_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__21_LC_9_25_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__21_LC_9_25_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__21_LC_9_25_4  (
            .in0(N__42733),
            .in1(N__35603),
            .in2(_gnd_net_),
            .in3(N__35548),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54240),
            .ce(N__41854),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__5_LC_9_25_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__5_LC_9_25_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__5_LC_9_25_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__5_LC_9_25_5  (
            .in0(N__35549),
            .in1(N__35604),
            .in2(_gnd_net_),
            .in3(N__42737),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54240),
            .ce(N__41854),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI6VHT_22_LC_9_25_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI6VHT_22_LC_9_25_6 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI6VHT_22_LC_9_25_6 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI6VHT_22_LC_9_25_6  (
            .in0(N__25333),
            .in1(N__25912),
            .in2(N__45550),
            .in3(_gnd_net_),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI6VHTZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__22_LC_9_25_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__22_LC_9_25_7 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__22_LC_9_25_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__22_LC_9_25_7  (
            .in0(N__32789),
            .in1(N__32683),
            .in2(_gnd_net_),
            .in3(N__42736),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54240),
            .ce(N__41854),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_4_LC_9_26_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_4_LC_9_26_0 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_4_LC_9_26_0 .LUT_INIT=16'b0000000011110111;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDfw_4_LC_9_26_0  (
            .in0(N__42244),
            .in1(N__25623),
            .in2(N__25327),
            .in3(N__25693),
            .lcout(\u1.DMAd_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54255),
            .ce(N__25396),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_2_LC_9_26_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_2_LC_9_26_1 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_2_LC_9_26_1 .LUT_INIT=16'b0000001101000111;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_2_LC_9_26_1  (
            .in0(N__25882),
            .in1(N__25613),
            .in2(N__25861),
            .in3(N__42240),
            .lcout(),
            .ltout(\u1.DMA_control.writeDfw_6_i_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_2_LC_9_26_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_2_LC_9_26_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_2_LC_9_26_2 .LUT_INIT=16'b0000110100001111;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDfw_2_LC_9_26_2  (
            .in0(N__42242),
            .in1(N__25846),
            .in2(N__25822),
            .in3(N__25624),
            .lcout(\u1.DMAd_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54255),
            .ce(N__25396),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_3_LC_9_26_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_3_LC_9_26_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_3_LC_9_26_3 .LUT_INIT=16'b0000001101000111;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_3_LC_9_26_3  (
            .in0(N__25804),
            .in1(N__25614),
            .in2(N__25783),
            .in3(N__42241),
            .lcout(),
            .ltout(\u1.DMA_control.writeDfw_6_i_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_3_LC_9_26_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_3_LC_9_26_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_3_LC_9_26_4 .LUT_INIT=16'b0000110100001111;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDfw_3_LC_9_26_4  (
            .in0(N__42243),
            .in1(N__25768),
            .in2(N__25750),
            .in3(N__25625),
            .lcout(\u1.DMAd_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54255),
            .ce(N__25396),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_4_LC_9_26_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_4_LC_9_26_5 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_4_LC_9_26_5 .LUT_INIT=16'b0000001101000111;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_4_LC_9_26_5  (
            .in0(N__25732),
            .in1(N__25612),
            .in2(N__25708),
            .in3(N__42238),
            .lcout(\u1.DMA_control.writeDfw_6_i_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_15_LC_9_26_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_15_LC_9_26_6 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_15_LC_9_26_6 .LUT_INIT=16'b0000001101010011;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDfw_RNO_0_15_LC_9_26_6  (
            .in0(N__42239),
            .in1(N__25687),
            .in2(N__25629),
            .in3(N__25675),
            .lcout(),
            .ltout(\u1.DMA_control.writeDfw_6_i_m3_i_0_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_15_LC_9_26_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_15_LC_9_26_7 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_writeDfw_15_LC_9_26_7 .LUT_INIT=16'b0000101100001111;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_writeDfw_15_LC_9_26_7  (
            .in0(N__25654),
            .in1(N__25618),
            .in2(N__25414),
            .in3(N__42245),
            .lcout(\u1.DMAd_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54255),
            .ce(N__25396),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__20_LC_9_27_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__20_LC_9_27_0 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__20_LC_9_27_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__20_LC_9_27_0  (
            .in0(N__31001),
            .in1(N__30891),
            .in2(_gnd_net_),
            .in3(N__42374),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54267),
            .ce(N__28260),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__2_LC_9_27_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__2_LC_9_27_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__2_LC_9_27_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__2_LC_9_27_1  (
            .in0(N__42371),
            .in1(N__30433),
            .in2(_gnd_net_),
            .in3(N__30339),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54267),
            .ce(N__28260),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__4_LC_9_27_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__4_LC_9_27_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__4_LC_9_27_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__4_LC_9_27_2  (
            .in0(N__31002),
            .in1(N__30892),
            .in2(_gnd_net_),
            .in3(N__42375),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54267),
            .ce(N__28260),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__23_LC_9_27_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__23_LC_9_27_3 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__23_LC_9_27_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__23_LC_9_27_3  (
            .in0(N__42370),
            .in1(N__38849),
            .in2(_gnd_net_),
            .in3(N__38743),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54267),
            .ce(N__28260),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__14_LC_9_27_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__14_LC_9_27_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__14_LC_9_27_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__14_LC_9_27_4  (
            .in0(N__33061),
            .in1(N__32973),
            .in2(_gnd_net_),
            .in3(N__42373),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54267),
            .ce(N__28260),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__30_LC_9_27_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__30_LC_9_27_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__30_LC_9_27_5 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__30_LC_9_27_5  (
            .in0(N__42372),
            .in1(N__33062),
            .in2(N__32980),
            .in3(_gnd_net_),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54267),
            .ce(N__28260),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__5_LC_9_27_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__5_LC_9_27_6 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__5_LC_9_27_6 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__5_LC_9_27_6  (
            .in0(N__35551),
            .in1(_gnd_net_),
            .in2(N__35664),
            .in3(N__42376),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54267),
            .ce(N__28260),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__21_LC_9_27_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__21_LC_9_27_7 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__21_LC_9_27_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__21_LC_9_27_7  (
            .in0(N__42369),
            .in1(N__35638),
            .in2(_gnd_net_),
            .in3(N__35550),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54267),
            .ce(N__28260),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__3_LC_9_28_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__3_LC_9_28_0 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__3_LC_9_28_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__3_LC_9_28_0  (
            .in0(N__36426),
            .in1(N__36538),
            .in2(_gnd_net_),
            .in3(N__42381),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54277),
            .ce(N__28137),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__29_LC_9_28_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__29_LC_9_28_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__29_LC_9_28_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__29_LC_9_28_1  (
            .in0(N__42378),
            .in1(N__33530),
            .in2(_gnd_net_),
            .in3(N__33424),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54277),
            .ce(N__28137),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__4_LC_9_28_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__4_LC_9_28_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__4_LC_9_28_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__4_LC_9_28_2  (
            .in0(N__30900),
            .in1(N__31004),
            .in2(_gnd_net_),
            .in3(N__42382),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54277),
            .ce(N__28137),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__20_LC_9_28_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__20_LC_9_28_3 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__20_LC_9_28_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__20_LC_9_28_3  (
            .in0(N__42377),
            .in1(N__31003),
            .in2(_gnd_net_),
            .in3(N__30899),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54277),
            .ce(N__28137),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__14_LC_9_28_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__14_LC_9_28_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__14_LC_9_28_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__14_LC_9_28_4  (
            .in0(N__33074),
            .in1(N__32969),
            .in2(_gnd_net_),
            .in3(N__42380),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54277),
            .ce(N__28137),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__30_LC_9_28_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__30_LC_9_28_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__30_LC_9_28_5 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__30_LC_9_28_5  (
            .in0(N__42379),
            .in1(N__33075),
            .in2(N__32979),
            .in3(_gnd_net_),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54277),
            .ce(N__28137),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__5_LC_9_28_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__5_LC_9_28_6 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__5_LC_9_28_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__5_LC_9_28_6  (
            .in0(N__35665),
            .in1(N__35552),
            .in2(_gnd_net_),
            .in3(N__42383),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54277),
            .ce(N__28137),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__15_LC_9_29_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__15_LC_9_29_0 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__15_LC_9_29_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__15_LC_9_29_0  (
            .in0(N__32610),
            .in1(N__32492),
            .in2(_gnd_net_),
            .in3(N__42494),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54287),
            .ce(N__28292),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__31_LC_9_29_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__31_LC_9_29_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__31_LC_9_29_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__31_LC_9_29_1  (
            .in0(N__42493),
            .in1(_gnd_net_),
            .in2(N__32497),
            .in3(N__32611),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54287),
            .ce(N__28292),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__6_LC_9_29_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__6_LC_9_29_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__6_LC_9_29_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__6_LC_9_29_2  (
            .in0(N__32712),
            .in1(N__32826),
            .in2(_gnd_net_),
            .in3(N__42495),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54287),
            .ce(N__28292),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__22_LC_9_29_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__22_LC_9_29_3 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__22_LC_9_29_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__22_LC_9_29_3  (
            .in0(N__42492),
            .in1(N__32825),
            .in2(_gnd_net_),
            .in3(N__32711),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54287),
            .ce(N__28292),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__7_LC_9_29_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__7_LC_9_29_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__7_LC_9_29_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__7_LC_9_29_4  (
            .in0(N__38850),
            .in1(N__38749),
            .in2(_gnd_net_),
            .in3(N__42496),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54287),
            .ce(N__28292),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__13_LC_9_29_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__13_LC_9_29_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__13_LC_9_29_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__13_LC_9_29_5  (
            .in0(N__42491),
            .in1(N__33562),
            .in2(_gnd_net_),
            .in3(N__33425),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54287),
            .ce(N__28292),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__8_LC_9_29_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__8_LC_9_29_6 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__8_LC_9_29_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__8_LC_9_29_6  (
            .in0(N__38530),
            .in1(N__38625),
            .in2(_gnd_net_),
            .in3(N__42497),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54287),
            .ce(N__28292),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI2B9K_22_LC_9_30_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI2B9K_22_LC_9_30_0 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI2B9K_22_LC_9_30_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI2B9K_22_LC_9_30_0  (
            .in0(N__45683),
            .in1(N__25975),
            .in2(_gnd_net_),
            .in3(N__27265),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI2B9KZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__22_LC_9_30_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__22_LC_9_30_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__22_LC_9_30_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__22_LC_9_30_1  (
            .in0(N__42499),
            .in1(N__32822),
            .in2(_gnd_net_),
            .in3(N__32714),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54298),
            .ce(N__30787),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__6_LC_9_30_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__6_LC_9_30_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__6_LC_9_30_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__6_LC_9_30_2  (
            .in0(N__32715),
            .in1(N__32823),
            .in2(_gnd_net_),
            .in3(N__42501),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54298),
            .ce(N__30787),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI2DBK_31_LC_9_30_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI2DBK_31_LC_9_30_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI2DBK_31_LC_9_30_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI2DBK_31_LC_9_30_3  (
            .in0(N__25969),
            .in1(N__28162),
            .in2(_gnd_net_),
            .in3(N__45684),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI2DBKZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__31_LC_9_30_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__31_LC_9_30_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__31_LC_9_30_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__31_LC_9_30_4  (
            .in0(N__32490),
            .in1(N__32609),
            .in2(_gnd_net_),
            .in3(N__42500),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54298),
            .ce(N__30787),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__15_LC_9_30_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__15_LC_9_30_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__15_LC_9_30_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__15_LC_9_30_5  (
            .in0(N__42498),
            .in1(N__32608),
            .in2(_gnd_net_),
            .in3(N__32489),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54298),
            .ce(N__30787),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI6D7K_15_LC_9_30_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI6D7K_15_LC_9_30_6 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI6D7K_15_LC_9_30_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI6D7K_15_LC_9_30_6  (
            .in0(N__45686),
            .in1(N__28174),
            .in2(_gnd_net_),
            .in3(N__25963),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI6D7KZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI2L4N_4_LC_9_30_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI2L4N_4_LC_9_30_7 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI2L4N_4_LC_9_30_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI2L4N_4_LC_9_30_7  (
            .in0(N__28222),
            .in1(N__25942),
            .in2(_gnd_net_),
            .in3(N__45685),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI2L4NZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__28_LC_9_31_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__28_LC_9_31_6 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__28_LC_9_31_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__28_LC_9_31_6  (
            .in0(N__32184),
            .in1(N__32074),
            .in2(_gnd_net_),
            .in3(N__43028),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54306),
            .ce(N__28294),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev1_Td_RNIABGKG_5_LC_9_32_6 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Td_RNIABGKG_5_LC_9_32_6 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev1_Td_RNIABGKG_5_LC_9_32_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \u0.DMA_dev1_Td_RNIABGKG_5_LC_9_32_6  (
            .in0(N__34069),
            .in1(N__26137),
            .in2(N__26125),
            .in3(N__26113),
            .lcout(wb_dat_o_c_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_cmdport_T1_1_LC_10_14_0 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_T1_1_LC_10_14_0 .SEQ_MODE=4'b1011;
    defparam \u0.PIO_cmdport_T1_1_LC_10_14_0 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \u0.PIO_cmdport_T1_1_LC_10_14_0  (
            .in0(N__51946),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39337),
            .lcout(PIO_cmdport_T1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54182),
            .ce(N__49696),
            .sr(N__53338));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNO_0_0_LC_10_15_5 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNO_0_0_LC_10_15_5 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNO_0_0_LC_10_15_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_RNO_0_0_LC_10_15_5  (
            .in0(N__28702),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26080),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t1_cnt.cnt.Qi_s_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport0_T2_RNIP0VR3_4_LC_10_16_0 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T2_RNIP0VR3_4_LC_10_16_0 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport0_T2_RNIP0VR3_4_LC_10_16_0 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \u0.PIO_dport0_T2_RNIP0VR3_4_LC_10_16_0  (
            .in0(N__46983),
            .in1(N__50766),
            .in2(N__28354),
            .in3(N__27364),
            .lcout(\u0.dat_o_0_0_3_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport1_T2_4_LC_10_16_3 .C_ON=1'b0;
    defparam \u0.PIO_dport1_T2_4_LC_10_16_3 .SEQ_MODE=4'b1011;
    defparam \u0.PIO_dport1_T2_4_LC_10_16_3 .LUT_INIT=16'b1110111011101110;
    LogicCell40 \u0.PIO_dport1_T2_4_LC_10_16_3  (
            .in0(N__51783),
            .in1(N__36985),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(PIO_dport1_T2_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54160),
            .ce(N__39154),
            .sr(N__53326));
    defparam \u0.register_block_gen_stat_reg_int_RNO_0_LC_10_16_5 .C_ON=1'b0;
    defparam \u0.register_block_gen_stat_reg_int_RNO_0_LC_10_16_5 .SEQ_MODE=4'b0000;
    defparam \u0.register_block_gen_stat_reg_int_RNO_0_LC_10_16_5 .LUT_INIT=16'b1111111101000000;
    LogicCell40 \u0.register_block_gen_stat_reg_int_RNO_0_LC_10_16_5  (
            .in0(N__49501),
            .in1(N__46601),
            .in2(N__50863),
            .in3(N__52105),
            .lcout(\u0.int_3_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport1_T1_0_LC_10_16_6 .C_ON=1'b0;
    defparam \u0.PIO_dport1_T1_0_LC_10_16_6 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport1_T1_0_LC_10_16_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \u0.PIO_dport1_T1_0_LC_10_16_6  (
            .in0(_gnd_net_),
            .in1(N__51782),
            .in2(_gnd_net_),
            .in3(N__49500),
            .lcout(PIO_dport1_T1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54160),
            .ce(N__39154),
            .sr(N__53326));
    defparam \u1.PIO_control.PIO_access_control.T1_RNO_0_0_LC_10_16_7 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T1_RNO_0_0_LC_10_16_7 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.T1_RNO_0_0_LC_10_16_7 .LUT_INIT=16'b0101110100001100;
    LogicCell40 \u1.PIO_control.PIO_access_control.T1_RNO_0_0_LC_10_16_7  (
            .in0(N__36570),
            .in1(N__29256),
            .in2(N__25998),
            .in3(N__29451),
            .lcout(\u1.PIO_control.PIO_access_control.it1_1_iv_i_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.Teoc_RNO_0_6_LC_10_17_0 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.Teoc_RNO_0_6_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.Teoc_RNO_0_6_LC_10_17_0 .LUT_INIT=16'b0111001101010000;
    LogicCell40 \u1.PIO_control.PIO_access_control.Teoc_RNO_0_6_LC_10_17_0  (
            .in0(N__47955),
            .in1(N__46767),
            .in2(N__29463),
            .in3(N__29031),
            .lcout(),
            .ltout(\u1.PIO_control.PIO_access_control.iteoc_1_iv_0_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.Teoc_6_LC_10_17_1 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.Teoc_6_LC_10_17_1 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.Teoc_6_LC_10_17_1 .LUT_INIT=16'b0000110000001111;
    LogicCell40 \u1.PIO_control.PIO_access_control.Teoc_6_LC_10_17_1  (
            .in0(_gnd_net_),
            .in1(N__46798),
            .in2(N__26206),
            .in3(N__29255),
            .lcout(\u1.PIO_control.PIO_access_control.TeocZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54151),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T1_5_LC_10_17_2 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T1_5_LC_10_17_2 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.T1_5_LC_10_17_2 .LUT_INIT=16'b0000000011011101;
    LogicCell40 \u1.PIO_control.PIO_access_control.T1_5_LC_10_17_2  (
            .in0(N__29254),
            .in1(N__31899),
            .in2(_gnd_net_),
            .in3(N__26479),
            .lcout(\u1.PIO_control.PIO_access_control.T1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54151),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.Teoc_7_LC_10_17_3 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.Teoc_7_LC_10_17_3 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.Teoc_7_LC_10_17_3 .LUT_INIT=16'b0000000011011101;
    LogicCell40 \u1.PIO_control.PIO_access_control.Teoc_7_LC_10_17_3  (
            .in0(N__29033),
            .in1(N__40305),
            .in2(_gnd_net_),
            .in3(N__26653),
            .lcout(\u1.PIO_control.PIO_access_control.TeocZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54151),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T1_RNO_0_3_LC_10_17_5 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T1_RNO_0_3_LC_10_17_5 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.T1_RNO_0_3_LC_10_17_5 .LUT_INIT=16'b0101110100001100;
    LogicCell40 \u1.PIO_control.PIO_access_control.T1_RNO_0_3_LC_10_17_5  (
            .in0(N__27807),
            .in1(N__29253),
            .in2(N__34975),
            .in3(N__29441),
            .lcout(),
            .ltout(\u1.PIO_control.PIO_access_control.it1_1_iv_i_i_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T1_3_LC_10_17_6 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T1_3_LC_10_17_6 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.T1_3_LC_10_17_6 .LUT_INIT=16'b0000101000001111;
    LogicCell40 \u1.PIO_control.PIO_access_control.T1_3_LC_10_17_6  (
            .in0(N__31647),
            .in1(_gnd_net_),
            .in2(N__26164),
            .in3(N__29032),
            .lcout(\u1.PIO_control.PIO_access_control.T1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54151),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T1_RNO_0_2_LC_10_17_7 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T1_RNO_0_2_LC_10_17_7 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.T1_RNO_0_2_LC_10_17_7 .LUT_INIT=16'b0101110100001100;
    LogicCell40 \u1.PIO_control.PIO_access_control.T1_RNO_0_2_LC_10_17_7  (
            .in0(N__27855),
            .in1(N__29252),
            .in2(N__34141),
            .in3(N__29440),
            .lcout(\u1.PIO_control.PIO_access_control.it1_1_iv_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_0_LC_10_18_0 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_0_LC_10_18_0 .SEQ_MODE=4'b1010;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_0_LC_10_18_0 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_0_LC_10_18_0  (
            .in0(N__27460),
            .in1(N__26143),
            .in2(N__52178),
            .in3(N__26468),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.QiZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54161),
            .ce(N__26437),
            .sr(N__53339));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_6_LC_10_18_1 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_6_LC_10_18_1 .SEQ_MODE=4'b1010;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_6_LC_10_18_1 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_6_LC_10_18_1  (
            .in0(N__26472),
            .in1(N__28366),
            .in2(N__27514),
            .in3(N__51987),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.QiZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54161),
            .ce(N__26437),
            .sr(N__53339));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_7_LC_10_18_2 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_7_LC_10_18_2 .SEQ_MODE=4'b1010;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_7_LC_10_18_2 .LUT_INIT=16'b0000110010101010;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_7_LC_10_18_2  (
            .in0(N__29542),
            .in1(N__27502),
            .in2(N__52180),
            .in3(N__26473),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.QiZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54161),
            .ce(N__26437),
            .sr(N__53339));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_1_LC_10_18_3 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_1_LC_10_18_3 .SEQ_MODE=4'b1010;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_1_LC_10_18_3 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_1_LC_10_18_3  (
            .in0(N__26469),
            .in1(N__51982),
            .in2(N__27451),
            .in3(N__28900),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.QiZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54161),
            .ce(N__26437),
            .sr(N__53339));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_3_LC_10_18_4 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_3_LC_10_18_4 .SEQ_MODE=4'b1011;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_3_LC_10_18_4 .LUT_INIT=16'b1111101011001100;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_3_LC_10_18_4  (
            .in0(N__27394),
            .in1(N__28834),
            .in2(N__52179),
            .in3(N__26470),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.QiZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54161),
            .ce(N__26437),
            .sr(N__53339));
    defparam \u1.PIO_control.PIO_access_control.it4_1_iv_i_i_a2_2_2_LC_10_18_5 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.it4_1_iv_i_i_a2_2_2_LC_10_18_5 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.it4_1_iv_i_i_a2_2_2_LC_10_18_5 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \u1.PIO_control.PIO_access_control.it4_1_iv_i_i_a2_2_2_LC_10_18_5  (
            .in0(N__27690),
            .in1(N__26493),
            .in2(N__36251),
            .in3(N__26678),
            .lcout(\u1.PIO_control.PIO_access_control.N_2110 ),
            .ltout(\u1.PIO_control.PIO_access_control.N_2110_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T1_RNO_0_5_LC_10_18_6 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T1_RNO_0_5_LC_10_18_6 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.T1_RNO_0_5_LC_10_18_6 .LUT_INIT=16'b0111001101010000;
    LogicCell40 \u1.PIO_control.PIO_access_control.T1_RNO_0_5_LC_10_18_6  (
            .in0(N__46173),
            .in1(N__31176),
            .in2(N__26482),
            .in3(N__29365),
            .lcout(\u1.PIO_control.PIO_access_control.it1_1_iv_i_i_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_4_LC_10_18_7 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_4_LC_10_18_7 .SEQ_MODE=4'b1011;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_4_LC_10_18_7 .LUT_INIT=16'b1111101011011000;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_4_LC_10_18_7  (
            .in0(N__26471),
            .in1(N__51986),
            .in2(N__28798),
            .in3(N__27352),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.QiZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54161),
            .ce(N__26437),
            .sr(N__53339));
    defparam \u1.DA_0_LC_10_19_0 .C_ON=1'b0;
    defparam \u1.DA_0_LC_10_19_0 .SEQ_MODE=4'b1010;
    defparam \u1.DA_0_LC_10_19_0 .LUT_INIT=16'b0000110000001010;
    LogicCell40 \u1.DA_0_LC_10_19_0  (
            .in0(N__26416),
            .in1(N__26403),
            .in2(N__52297),
            .in3(N__26904),
            .lcout(da_pad_o_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54171),
            .ce(),
            .sr(N__53344));
    defparam \u1.PIO_control.gen_pingpong_rpp_LC_10_19_1 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_rpp_LC_10_19_1 .SEQ_MODE=4'b1010;
    defparam \u1.PIO_control.gen_pingpong_rpp_LC_10_19_1 .LUT_INIT=16'b0000101000000110;
    LogicCell40 \u1.PIO_control.gen_pingpong_rpp_LC_10_19_1  (
            .in0(N__26903),
            .in1(N__26360),
            .in2(N__26326),
            .in3(N__26307),
            .lcout(\u1.rpp ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54171),
            .ce(),
            .sr(N__53344));
    defparam \u1.PIO_control.PIO_access_control.it4_1_iv_i_i_o2_0_x1_2_LC_10_19_2 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.it4_1_iv_i_i_o2_0_x1_2_LC_10_19_2 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.it4_1_iv_i_i_o2_0_x1_2_LC_10_19_2 .LUT_INIT=16'b1111110111111101;
    LogicCell40 \u1.PIO_control.PIO_access_control.it4_1_iv_i_i_o2_0_x1_2_LC_10_19_2  (
            .in0(N__26790),
            .in1(N__26274),
            .in2(N__26226),
            .in3(_gnd_net_),
            .lcout(\u1.PIO_control.PIO_access_control.it4_1_iv_i_i_o2_0_x1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.it4_1_iv_i_i_o2_0_x0_2_LC_10_19_3 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.it4_1_iv_i_i_o2_0_x0_2_LC_10_19_3 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.it4_1_iv_i_i_o2_0_x0_2_LC_10_19_3 .LUT_INIT=16'b1111110010111000;
    LogicCell40 \u1.PIO_control.PIO_access_control.it4_1_iv_i_i_o2_0_x0_2_LC_10_19_3  (
            .in0(N__26275),
            .in1(N__26791),
            .in2(N__26257),
            .in3(N__26219),
            .lcout(),
            .ltout(\u1.PIO_control.PIO_access_control.it4_1_iv_i_i_o2_0_x0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.it4_1_iv_i_i_o2_0_ns_2_LC_10_19_4 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.it4_1_iv_i_i_o2_0_ns_2_LC_10_19_4 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.it4_1_iv_i_i_o2_0_ns_2_LC_10_19_4 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \u1.PIO_control.PIO_access_control.it4_1_iv_i_i_o2_0_ns_2_LC_10_19_4  (
            .in0(_gnd_net_),
            .in1(N__26574),
            .in2(N__26563),
            .in3(N__26560),
            .lcout(\u1.PIO_control.PIO_access_control.it4_1_iv_i_i_o2_0_2 ),
            .ltout(\u1.PIO_control.PIO_access_control.it4_1_iv_i_i_o2_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.it4_1_iv_i_i_o3_x0_2_LC_10_19_5 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.it4_1_iv_i_i_o3_x0_2_LC_10_19_5 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.it4_1_iv_i_i_o3_x0_2_LC_10_19_5 .LUT_INIT=16'b1111001011110111;
    LogicCell40 \u1.PIO_control.PIO_access_control.it4_1_iv_i_i_o3_x0_2_LC_10_19_5  (
            .in0(N__36209),
            .in1(N__40623),
            .in2(N__26554),
            .in3(N__27683),
            .lcout(),
            .ltout(\u1.PIO_control.PIO_access_control.it4_1_iv_i_i_o3_x0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.it4_1_iv_i_i_o3_ns_2_LC_10_19_6 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.it4_1_iv_i_i_o3_ns_2_LC_10_19_6 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.it4_1_iv_i_i_o3_ns_2_LC_10_19_6 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \u1.PIO_control.PIO_access_control.it4_1_iv_i_i_o3_ns_2_LC_10_19_6  (
            .in0(N__28708),
            .in1(_gnd_net_),
            .in2(N__26551),
            .in3(N__26677),
            .lcout(\u1.PIO_control.PIO_access_control.N_1319 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.IORDYen_RNO_0_LC_10_20_0 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.IORDYen_RNO_0_LC_10_20_0 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.IORDYen_RNO_0_LC_10_20_0 .LUT_INIT=16'b0111010100110000;
    LogicCell40 \u1.PIO_control.PIO_access_control.IORDYen_RNO_0_LC_10_20_0  (
            .in0(N__27792),
            .in1(N__39237),
            .in2(N__29439),
            .in3(N__29243),
            .lcout(),
            .ltout(\u1.PIO_control.PIO_access_control.iiordyen_1_iv_i_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.IORDYen_LC_10_20_1 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.IORDYen_LC_10_20_1 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.IORDYen_LC_10_20_1 .LUT_INIT=16'b0000101000001111;
    LogicCell40 \u1.PIO_control.PIO_access_control.IORDYen_LC_10_20_1  (
            .in0(N__27831),
            .in1(_gnd_net_),
            .in2(N__26548),
            .in3(N__29070),
            .lcout(\u1.PIO_control.PIO_access_control.IORDYenZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54183),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T1_RNO_0_1_LC_10_20_3 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T1_RNO_0_1_LC_10_20_3 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.T1_RNO_0_1_LC_10_20_3 .LUT_INIT=16'b0011101100001010;
    LogicCell40 \u1.PIO_control.PIO_access_control.T1_RNO_0_1_LC_10_20_3  (
            .in0(N__29244),
            .in1(N__27651),
            .in2(N__44673),
            .in3(N__29380),
            .lcout(),
            .ltout(\u1.PIO_control.PIO_access_control.it1_1_iv_i_i_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T1_1_LC_10_20_4 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T1_1_LC_10_20_4 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.T1_1_LC_10_20_4 .LUT_INIT=16'b0000111100000101;
    LogicCell40 \u1.PIO_control.PIO_access_control.T1_1_LC_10_20_4  (
            .in0(N__29071),
            .in1(_gnd_net_),
            .in2(N__26530),
            .in3(N__31731),
            .lcout(\u1.PIO_control.PIO_access_control.T1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54183),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_Td_1_LC_10_20_5 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_Td_1_LC_10_20_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.DMA_timing_ctrl_Td_1_LC_10_20_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_Td_1_LC_10_20_5  (
            .in0(N__48384),
            .in1(N__31306),
            .in2(_gnd_net_),
            .in3(N__36170),
            .lcout(\u1.DMA_control.Td_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54183),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.it4_1_iv_i_i_a2_3_2_LC_10_20_6 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.it4_1_iv_i_i_a2_3_2_LC_10_20_6 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.it4_1_iv_i_i_a2_3_2_LC_10_20_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \u1.PIO_control.PIO_access_control.it4_1_iv_i_i_a2_3_2_LC_10_20_6  (
            .in0(N__40619),
            .in1(N__26494),
            .in2(N__36216),
            .in3(N__26679),
            .lcout(\u1.PIO_control.PIO_access_control.N_2112 ),
            .ltout(\u1.PIO_control.PIO_access_control.N_2112_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.Teoc_RNO_0_7_LC_10_20_7 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.Teoc_RNO_0_7_LC_10_20_7 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.Teoc_RNO_0_7_LC_10_20_7 .LUT_INIT=16'b0111001101010000;
    LogicCell40 \u1.PIO_control.PIO_access_control.Teoc_RNO_0_7_LC_10_20_7  (
            .in0(N__40363),
            .in1(N__40341),
            .in2(N__26656),
            .in3(N__29376),
            .lcout(\u1.PIO_control.PIO_access_control.iteoc_1_iv_i_i_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T4_RNO_0_2_LC_10_21_0 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T4_RNO_0_2_LC_10_21_0 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.T4_RNO_0_2_LC_10_21_0 .LUT_INIT=16'b0101110100001100;
    LogicCell40 \u1.PIO_control.PIO_access_control.T4_RNO_0_2_LC_10_21_0  (
            .in0(N__35142),
            .in1(N__29245),
            .in2(N__37017),
            .in3(N__29456),
            .lcout(),
            .ltout(\u1.PIO_control.PIO_access_control.it4_1_iv_i_i_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T4_2_LC_10_21_1 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T4_2_LC_10_21_1 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.T4_2_LC_10_21_1 .LUT_INIT=16'b0000111100000101;
    LogicCell40 \u1.PIO_control.PIO_access_control.T4_2_LC_10_21_1  (
            .in0(N__29068),
            .in1(_gnd_net_),
            .in2(N__26644),
            .in3(N__37546),
            .lcout(\u1.PIO_control.PIO_access_control.T4Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54194),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T4_RNO_0_3_LC_10_21_2 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T4_RNO_0_3_LC_10_21_2 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.T4_RNO_0_3_LC_10_21_2 .LUT_INIT=16'b0101110100001100;
    LogicCell40 \u1.PIO_control.PIO_access_control.T4_RNO_0_3_LC_10_21_2  (
            .in0(N__29595),
            .in1(N__29246),
            .in2(N__34447),
            .in3(N__29457),
            .lcout(),
            .ltout(\u1.PIO_control.PIO_access_control.it4_1_iv_i_i_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T4_3_LC_10_21_3 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T4_3_LC_10_21_3 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.T4_3_LC_10_21_3 .LUT_INIT=16'b0000111100000101;
    LogicCell40 \u1.PIO_control.PIO_access_control.T4_3_LC_10_21_3  (
            .in0(N__29069),
            .in1(_gnd_net_),
            .in2(N__26626),
            .in3(N__34294),
            .lcout(\u1.PIO_control.PIO_access_control.T4Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54194),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T4_RNO_0_4_LC_10_21_4 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T4_RNO_0_4_LC_10_21_4 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.T4_RNO_0_4_LC_10_21_4 .LUT_INIT=16'b0101110100001100;
    LogicCell40 \u1.PIO_control.PIO_access_control.T4_RNO_0_4_LC_10_21_4  (
            .in0(N__29580),
            .in1(N__29066),
            .in2(N__37504),
            .in3(N__29458),
            .lcout(),
            .ltout(\u1.PIO_control.PIO_access_control.it4_1_iv_0_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T4_4_LC_10_21_5 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T4_4_LC_10_21_5 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.T4_4_LC_10_21_5 .LUT_INIT=16'b0000111100000101;
    LogicCell40 \u1.PIO_control.PIO_access_control.T4_4_LC_10_21_5  (
            .in0(N__29247),
            .in1(_gnd_net_),
            .in2(N__26611),
            .in3(N__37524),
            .lcout(\u1.PIO_control.PIO_access_control.T4Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54194),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T4_RNO_0_5_LC_10_21_6 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T4_RNO_0_5_LC_10_21_6 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.T4_RNO_0_5_LC_10_21_6 .LUT_INIT=16'b0101110100001100;
    LogicCell40 \u1.PIO_control.PIO_access_control.T4_RNO_0_5_LC_10_21_6  (
            .in0(N__37911),
            .in1(N__29067),
            .in2(N__37444),
            .in3(N__29459),
            .lcout(),
            .ltout(\u1.PIO_control.PIO_access_control.it4_1_iv_i_i_0_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T4_5_LC_10_21_7 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T4_5_LC_10_21_7 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.T4_5_LC_10_21_7 .LUT_INIT=16'b0000111100000101;
    LogicCell40 \u1.PIO_control.PIO_access_control.T4_5_LC_10_21_7  (
            .in0(N__29248),
            .in1(_gnd_net_),
            .in2(N__26593),
            .in3(N__37468),
            .lcout(\u1.PIO_control.PIO_access_control.T4Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54194),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DDo_0_LC_10_22_0 .C_ON=1'b0;
    defparam \u1.DDo_0_LC_10_22_0 .SEQ_MODE=4'b1010;
    defparam \u1.DDo_0_LC_10_22_0 .LUT_INIT=16'b0000111000000010;
    LogicCell40 \u1.DDo_0_LC_10_22_0  (
            .in0(N__27043),
            .in1(N__36773),
            .in2(N__52422),
            .in3(N__26935),
            .lcout(dd_pad_o_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54204),
            .ce(),
            .sr(N__53363));
    defparam \u1.PIO_control.gen_pingpong_pong_a_RNI35V01_3_LC_10_22_1 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_pong_a_RNI35V01_3_LC_10_22_1 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.gen_pingpong_pong_a_RNI35V01_3_LC_10_22_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.PIO_control.gen_pingpong_pong_a_RNI35V01_3_LC_10_22_1  (
            .in0(N__27010),
            .in1(N__26995),
            .in2(_gnd_net_),
            .in3(N__26876),
            .lcout(\u1.N_1425 ),
            .ltout(\u1.N_1425_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.CS0n_LC_10_22_2 .C_ON=1'b0;
    defparam \u1.CS0n_LC_10_22_2 .SEQ_MODE=4'b1011;
    defparam \u1.CS0n_LC_10_22_2 .LUT_INIT=16'b1111101011111111;
    LogicCell40 \u1.CS0n_LC_10_22_2  (
            .in0(N__52181),
            .in1(_gnd_net_),
            .in2(N__26977),
            .in3(N__36771),
            .lcout(cs0n_pad_o_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54204),
            .ce(),
            .sr(N__53363));
    defparam \u1.PIO_control.gen_pingpong_pong_d_RNI3HHN_0_LC_10_22_3 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_pong_d_RNI3HHN_0_LC_10_22_3 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.gen_pingpong_pong_d_RNI3HHN_0_LC_10_22_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.PIO_control.gen_pingpong_pong_d_RNI3HHN_0_LC_10_22_3  (
            .in0(N__26956),
            .in1(N__26944),
            .in2(_gnd_net_),
            .in3(N__26877),
            .lcout(\u1.N_1426 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.gen_pingpong_pong_d_RNI5JHN_1_LC_10_22_4 .C_ON=1'b0;
    defparam \u1.PIO_control.gen_pingpong_pong_d_RNI5JHN_1_LC_10_22_4 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.gen_pingpong_pong_d_RNI5JHN_1_LC_10_22_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \u1.PIO_control.gen_pingpong_pong_d_RNI5JHN_1_LC_10_22_4  (
            .in0(N__26878),
            .in1(_gnd_net_),
            .in2(N__26755),
            .in3(N__26743),
            .lcout(),
            .ltout(\u1.N_1427_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DDo_1_LC_10_22_5 .C_ON=1'b0;
    defparam \u1.DDo_1_LC_10_22_5 .SEQ_MODE=4'b1010;
    defparam \u1.DDo_1_LC_10_22_5 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \u1.DDo_1_LC_10_22_5  (
            .in0(N__36774),
            .in1(N__52186),
            .in2(N__26731),
            .in3(N__26728),
            .lcout(dd_pad_o_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54204),
            .ce(),
            .sr(N__53363));
    defparam \u1.CS1n_LC_10_22_6 .C_ON=1'b0;
    defparam \u1.CS1n_LC_10_22_6 .SEQ_MODE=4'b1011;
    defparam \u1.CS1n_LC_10_22_6 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \u1.CS1n_LC_10_22_6  (
            .in0(N__52182),
            .in1(N__36772),
            .in2(_gnd_net_),
            .in3(N__26701),
            .lcout(cs1n_pad_o_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54204),
            .ce(),
            .sr(N__53363));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__5_LC_10_23_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__5_LC_10_23_0 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__5_LC_10_23_0 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__5_LC_10_23_0  (
            .in0(N__35557),
            .in1(_gnd_net_),
            .in2(N__35637),
            .in3(N__42727),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54217),
            .ce(N__41269),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__21_LC_10_23_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__21_LC_10_23_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__21_LC_10_23_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__21_LC_10_23_1  (
            .in0(N__42724),
            .in1(N__35605),
            .in2(_gnd_net_),
            .in3(N__35556),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54217),
            .ce(N__41269),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__15_LC_10_23_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__15_LC_10_23_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__15_LC_10_23_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__15_LC_10_23_2  (
            .in0(N__32598),
            .in1(N__32485),
            .in2(_gnd_net_),
            .in3(N__42726),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54217),
            .ce(N__41269),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI61KT_31_LC_10_23_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI61KT_31_LC_10_23_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI61KT_31_LC_10_23_3 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI61KT_31_LC_10_23_3  (
            .in0(N__27091),
            .in1(N__27193),
            .in2(N__45461),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI61KTZ0Z_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI4VG71_31_LC_10_23_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI4VG71_31_LC_10_23_4 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI4VG71_31_LC_10_23_4 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI4VG71_31_LC_10_23_4  (
            .in0(N__27076),
            .in1(_gnd_net_),
            .in2(N__27079),
            .in3(N__50038),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI4VG71Z0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__31_LC_10_23_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__31_LC_10_23_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__31_LC_10_23_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__31_LC_10_23_5  (
            .in0(N__42725),
            .in1(_gnd_net_),
            .in2(N__32496),
            .in3(N__32599),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54217),
            .ce(N__41269),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIIGLM1_2_LC_10_23_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIIGLM1_2_LC_10_23_6 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIIGLM1_2_LC_10_23_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIIGLM1_2_LC_10_23_6  (
            .in0(N__27070),
            .in1(N__28003),
            .in2(_gnd_net_),
            .in3(N__50039),
            .lcout(),
            .ltout(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIIGLM1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI9RD53_3_LC_10_23_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI9RD53_3_LC_10_23_7 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI9RD53_3_LC_10_23_7 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI9RD53_3_LC_10_23_7  (
            .in0(N__27058),
            .in1(_gnd_net_),
            .in2(N__27052),
            .in3(N__48868),
            .lcout(DMAq_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIQ0CM_2_LC_10_24_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIQ0CM_2_LC_10_24_0 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIQ0CM_2_LC_10_24_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIQ0CM_2_LC_10_24_0  (
            .in0(N__45417),
            .in1(N__27049),
            .in2(_gnd_net_),
            .in3(N__27175),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIQ0CMZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__2_LC_10_24_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__2_LC_10_24_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__2_LC_10_24_1 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__2_LC_10_24_1  (
            .in0(N__30362),
            .in1(_gnd_net_),
            .in2(N__30498),
            .in3(N__42723),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54230),
            .ce(N__35890),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__18_LC_10_24_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__18_LC_10_24_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__18_LC_10_24_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__18_LC_10_24_2  (
            .in0(N__42719),
            .in1(N__30487),
            .in2(_gnd_net_),
            .in3(N__30361),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54230),
            .ce(N__35890),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIS2CM_3_LC_10_24_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIS2CM_3_LC_10_24_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIS2CM_3_LC_10_24_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIS2CM_3_LC_10_24_3  (
            .in0(N__27223),
            .in1(N__27157),
            .in2(_gnd_net_),
            .in3(N__45418),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIS2CMZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__3_LC_10_24_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__3_LC_10_24_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__3_LC_10_24_4 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__3_LC_10_24_4  (
            .in0(N__42720),
            .in1(N__36536),
            .in2(N__36438),
            .in3(_gnd_net_),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54230),
            .ce(N__35890),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__19_LC_10_24_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__19_LC_10_24_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__19_LC_10_24_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__19_LC_10_24_5  (
            .in0(N__36535),
            .in1(N__36427),
            .in2(_gnd_net_),
            .in3(N__42722),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54230),
            .ce(N__35890),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNISIUQ_12_LC_10_24_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNISIUQ_12_LC_10_24_6 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNISIUQ_12_LC_10_24_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNISIUQ_12_LC_10_24_6  (
            .in0(N__45419),
            .in1(N__27166),
            .in2(_gnd_net_),
            .in3(N__27145),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNISIUQZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__12_LC_10_24_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__12_LC_10_24_7 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__12_LC_10_24_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__12_LC_10_24_7  (
            .in0(N__32140),
            .in1(N__32049),
            .in2(_gnd_net_),
            .in3(N__42721),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54230),
            .ce(N__35890),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI8VFT_14_LC_10_25_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI8VFT_14_LC_10_25_0 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI8VFT_14_LC_10_25_0 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI8VFT_14_LC_10_25_0  (
            .in0(N__45424),
            .in1(_gnd_net_),
            .in2(N__27130),
            .in3(N__27139),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI8VFTZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__14_LC_10_25_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__14_LC_10_25_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__14_LC_10_25_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__14_LC_10_25_1  (
            .in0(N__33039),
            .in1(N__32959),
            .in2(_gnd_net_),
            .in3(N__42730),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54241),
            .ce(N__41855),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__30_LC_10_25_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__30_LC_10_25_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__30_LC_10_25_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__30_LC_10_25_2  (
            .in0(N__42729),
            .in1(_gnd_net_),
            .in2(N__32977),
            .in3(N__33040),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54241),
            .ce(N__41855),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIA1GT_15_LC_10_25_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIA1GT_15_LC_10_25_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIA1GT_15_LC_10_25_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIA1GT_15_LC_10_25_3  (
            .in0(N__27121),
            .in1(N__27199),
            .in2(_gnd_net_),
            .in3(N__45425),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIA1GTZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__15_LC_10_25_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__15_LC_10_25_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__15_LC_10_25_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__15_LC_10_25_4  (
            .in0(N__42728),
            .in1(N__32585),
            .in2(_gnd_net_),
            .in3(N__32444),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54241),
            .ce(N__41855),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__31_LC_10_25_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__31_LC_10_25_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__31_LC_10_25_5 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__31_LC_10_25_5  (
            .in0(N__32445),
            .in1(_gnd_net_),
            .in2(N__32607),
            .in3(N__42732),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54241),
            .ce(N__41855),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIE5GT_17_LC_10_25_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIE5GT_17_LC_10_25_6 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIE5GT_17_LC_10_25_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIE5GT_17_LC_10_25_6  (
            .in0(N__45426),
            .in1(N__27181),
            .in2(_gnd_net_),
            .in3(N__27235),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIE5GTZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__17_LC_10_25_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__17_LC_10_25_7 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__17_LC_10_25_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__17_LC_10_25_7  (
            .in0(N__41535),
            .in1(N__41417),
            .in2(_gnd_net_),
            .in3(N__42731),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54241),
            .ce(N__41855),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__31_LC_10_26_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__31_LC_10_26_0 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__31_LC_10_26_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__31_LC_10_26_0  (
            .in0(N__32597),
            .in1(N__32477),
            .in2(_gnd_net_),
            .in3(N__42351),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54256),
            .ce(N__33260),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__9_LC_10_26_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__9_LC_10_26_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__9_LC_10_26_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__9_LC_10_26_1  (
            .in0(N__42348),
            .in1(N__35426),
            .in2(_gnd_net_),
            .in3(N__35323),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54256),
            .ce(N__33260),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__2_LC_10_26_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__2_LC_10_26_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__2_LC_10_26_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__2_LC_10_26_2  (
            .in0(N__30486),
            .in1(N__30338),
            .in2(_gnd_net_),
            .in3(N__42350),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54256),
            .ce(N__33260),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__24_LC_10_26_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__24_LC_10_26_3 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__24_LC_10_26_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__24_LC_10_26_3  (
            .in0(N__42346),
            .in1(N__38485),
            .in2(_gnd_net_),
            .in3(N__38609),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54256),
            .ce(N__33260),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__12_LC_10_26_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__12_LC_10_26_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__12_LC_10_26_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__12_LC_10_26_4  (
            .in0(N__32163),
            .in1(N__32059),
            .in2(_gnd_net_),
            .in3(N__42349),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54256),
            .ce(N__33260),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__28_LC_10_26_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__28_LC_10_26_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__28_LC_10_26_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__28_LC_10_26_5  (
            .in0(N__42347),
            .in1(_gnd_net_),
            .in2(N__32083),
            .in3(N__32164),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54256),
            .ce(N__33260),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__3_LC_10_26_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__3_LC_10_26_6 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__3_LC_10_26_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__3_LC_10_26_6  (
            .in0(N__36411),
            .in1(N__36503),
            .in2(_gnd_net_),
            .in3(N__42352),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54256),
            .ce(N__33260),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__19_LC_10_26_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__19_LC_10_26_7 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__19_LC_10_26_7 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__19_LC_10_26_7  (
            .in0(N__42345),
            .in1(_gnd_net_),
            .in2(N__36529),
            .in3(N__36412),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54256),
            .ce(N__33260),
            .sr(_gnd_net_));
    defparam \u0.register_block_gen_ctrl_reg_un6_sel_ctrl_i_LC_10_27_0 .C_ON=1'b0;
    defparam \u0.register_block_gen_ctrl_reg_un6_sel_ctrl_i_LC_10_27_0 .SEQ_MODE=4'b0000;
    defparam \u0.register_block_gen_ctrl_reg_un6_sel_ctrl_i_LC_10_27_0 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \u0.register_block_gen_ctrl_reg_un6_sel_ctrl_i_LC_10_27_0  (
            .in0(N__52425),
            .in1(N__50838),
            .in2(_gnd_net_),
            .in3(N__48337),
            .lcout(\u0.N_286 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.CtrlReg_2_LC_10_27_4 .C_ON=1'b0;
    defparam \u0.CtrlReg_2_LC_10_27_4 .SEQ_MODE=4'b1010;
    defparam \u0.CtrlReg_2_LC_10_27_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.CtrlReg_2_LC_10_27_4  (
            .in0(N__52423),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34242),
            .lcout(PIO_dport0_IORDYen),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54268),
            .ce(N__53549),
            .sr(N__53394));
    defparam \u0.CtrlReg_3_LC_10_27_5 .C_ON=1'b0;
    defparam \u0.CtrlReg_3_LC_10_27_5 .SEQ_MODE=4'b1010;
    defparam \u0.CtrlReg_3_LC_10_27_5 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \u0.CtrlReg_3_LC_10_27_5  (
            .in0(N__37378),
            .in1(N__52424),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(PIO_dport1_IORDYen),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54268),
            .ce(N__53549),
            .sr(N__53394));
    defparam \u1.DMA_control.gen_DMA_sigs_gen_writed_pipe_writeDlw_4_i_m2_0_LC_10_27_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_gen_writed_pipe_writeDlw_4_i_m2_0_LC_10_27_7 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMA_sigs_gen_writed_pipe_writeDlw_4_i_m2_0_LC_10_27_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_gen_writed_pipe_writeDlw_4_i_m2_0_LC_10_27_7  (
            .in0(N__44730),
            .in1(N__54357),
            .in2(_gnd_net_),
            .in3(N__36252),
            .lcout(\u1.DMA_control.N_1313 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__11_LC_10_28_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__11_LC_10_28_0 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__11_LC_10_28_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__11_LC_10_28_0  (
            .in0(N__43137),
            .in1(N__43232),
            .in2(_gnd_net_),
            .in3(N__42357),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54278),
            .ce(N__28138),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__27_LC_10_28_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__27_LC_10_28_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__27_LC_10_28_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__27_LC_10_28_1  (
            .in0(N__42356),
            .in1(_gnd_net_),
            .in2(N__43237),
            .in3(N__43138),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54278),
            .ce(N__28138),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__2_LC_10_28_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__2_LC_10_28_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__2_LC_10_28_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__2_LC_10_28_2  (
            .in0(N__30336),
            .in1(N__30473),
            .in2(_gnd_net_),
            .in3(N__42359),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54278),
            .ce(N__28138),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__18_LC_10_28_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__18_LC_10_28_3 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__18_LC_10_28_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__18_LC_10_28_3  (
            .in0(N__42353),
            .in1(N__30472),
            .in2(_gnd_net_),
            .in3(N__30335),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54278),
            .ce(N__28138),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__12_LC_10_28_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__12_LC_10_28_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__12_LC_10_28_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__12_LC_10_28_4  (
            .in0(N__32185),
            .in1(N__32081),
            .in2(_gnd_net_),
            .in3(N__42358),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54278),
            .ce(N__28138),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__25_LC_10_28_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__25_LC_10_28_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__25_LC_10_28_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__25_LC_10_28_5  (
            .in0(N__42355),
            .in1(_gnd_net_),
            .in2(N__35443),
            .in3(N__35341),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54278),
            .ce(N__28138),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__8_LC_10_28_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__8_LC_10_28_6 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__8_LC_10_28_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__8_LC_10_28_6  (
            .in0(N__38527),
            .in1(N__38619),
            .in2(_gnd_net_),
            .in3(N__42360),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54278),
            .ce(N__28138),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__19_LC_10_28_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__19_LC_10_28_7 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__19_LC_10_28_7 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__19_LC_10_28_7  (
            .in0(N__42354),
            .in1(N__36537),
            .in2(N__36435),
            .in3(_gnd_net_),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54278),
            .ce(N__28138),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__11_LC_10_29_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__11_LC_10_29_0 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__11_LC_10_29_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__11_LC_10_29_0  (
            .in0(N__43139),
            .in1(N__43225),
            .in2(_gnd_net_),
            .in3(N__42479),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54288),
            .ce(N__28293),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__27_LC_10_29_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__27_LC_10_29_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__27_LC_10_29_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__27_LC_10_29_1  (
            .in0(N__42478),
            .in1(_gnd_net_),
            .in2(N__43236),
            .in3(N__43140),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54288),
            .ce(N__28293),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__17_LC_10_29_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__17_LC_10_29_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__17_LC_10_29_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__17_LC_10_29_2  (
            .in0(N__41514),
            .in1(N__41418),
            .in2(_gnd_net_),
            .in3(N__42480),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54288),
            .ce(N__28293),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__25_LC_10_29_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__25_LC_10_29_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__25_LC_10_29_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__25_LC_10_29_4  (
            .in0(N__35438),
            .in1(N__35337),
            .in2(_gnd_net_),
            .in3(N__42481),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54288),
            .ce(N__28293),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__3_LC_10_29_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__3_LC_10_29_6 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__3_LC_10_29_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__3_LC_10_29_6  (
            .in0(_gnd_net_),
            .in1(N__36402),
            .in2(N__36549),
            .in3(N__42482),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54288),
            .ce(N__28293),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__19_LC_10_29_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__19_LC_10_29_7 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__19_LC_10_29_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__19_LC_10_29_7  (
            .in0(N__42477),
            .in1(N__36530),
            .in2(_gnd_net_),
            .in3(N__36403),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54288),
            .ce(N__28293),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__0_LC_10_30_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__0_LC_10_30_0 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__0_LC_10_30_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__0_LC_10_30_0  (
            .in0(N__41738),
            .in1(N__41642),
            .in2(_gnd_net_),
            .in3(N__42487),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54299),
            .ce(N__28146),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__1_LC_10_30_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__1_LC_10_30_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__1_LC_10_30_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__1_LC_10_30_1  (
            .in0(N__42483),
            .in1(_gnd_net_),
            .in2(N__41536),
            .in3(N__41419),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54299),
            .ce(N__28146),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__16_LC_10_30_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__16_LC_10_30_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__16_LC_10_30_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__16_LC_10_30_2  (
            .in0(N__41739),
            .in1(N__41643),
            .in2(_gnd_net_),
            .in3(N__42488),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54299),
            .ce(N__28146),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__22_LC_10_30_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__22_LC_10_30_3 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__22_LC_10_30_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__22_LC_10_30_3  (
            .in0(N__42485),
            .in1(N__32821),
            .in2(_gnd_net_),
            .in3(N__32713),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54299),
            .ce(N__28146),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__7_LC_10_30_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__7_LC_10_30_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__7_LC_10_30_4 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__7_LC_10_30_4  (
            .in0(N__38745),
            .in1(_gnd_net_),
            .in2(N__38857),
            .in3(N__42490),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54299),
            .ce(N__28146),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__23_LC_10_30_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__23_LC_10_30_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__23_LC_10_30_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__23_LC_10_30_5  (
            .in0(N__42486),
            .in1(N__38851),
            .in2(_gnd_net_),
            .in3(N__38744),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54299),
            .ce(N__28146),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__28_LC_10_30_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__28_LC_10_30_6 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__28_LC_10_30_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__28_LC_10_30_6  (
            .in0(N__32206),
            .in1(N__32082),
            .in2(_gnd_net_),
            .in3(N__42489),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54299),
            .ce(N__28146),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__21_LC_10_30_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__21_LC_10_30_7 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__21_LC_10_30_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__21_LC_10_30_7  (
            .in0(N__42484),
            .in1(N__35666),
            .in2(_gnd_net_),
            .in3(N__35560),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54299),
            .ce(N__28146),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI6F9K_24_LC_10_31_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI6F9K_24_LC_10_31_0 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI6F9K_24_LC_10_31_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI6F9K_24_LC_10_31_0  (
            .in0(N__45632),
            .in1(N__27331),
            .in2(_gnd_net_),
            .in3(N__27286),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI6F9KZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__24_LC_10_31_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__24_LC_10_31_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__24_LC_10_31_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__24_LC_10_31_1  (
            .in0(N__38626),
            .in1(N__38531),
            .in2(_gnd_net_),
            .in3(N__43031),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54307),
            .ce(N__30812),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__8_LC_10_31_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__8_LC_10_31_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__8_LC_10_31_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__8_LC_10_31_2  (
            .in0(N__43029),
            .in1(N__38532),
            .in2(_gnd_net_),
            .in3(N__38627),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54307),
            .ce(N__30812),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIAT4N_8_LC_10_31_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIAT4N_8_LC_10_31_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIAT4N_8_LC_10_31_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIAT4N_8_LC_10_31_3  (
            .in0(N__27325),
            .in1(N__27319),
            .in2(_gnd_net_),
            .in3(N__45634),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIAT4NZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI8F7K_16_LC_10_31_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI8F7K_16_LC_10_31_4 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI8F7K_16_LC_10_31_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI8F7K_16_LC_10_31_4  (
            .in0(N__45633),
            .in1(N__27310),
            .in2(_gnd_net_),
            .in3(N__27304),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI8F7KZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__16_LC_10_31_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__16_LC_10_31_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__16_LC_10_31_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__16_LC_10_31_5  (
            .in0(N__41740),
            .in1(N__41644),
            .in2(_gnd_net_),
            .in3(N__43030),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54307),
            .ce(N__30812),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIQC4N_0_LC_10_31_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIQC4N_0_LC_10_31_7 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIQC4N_0_LC_10_31_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIQC4N_0_LC_10_31_7  (
            .in0(N__27295),
            .in1(N__28213),
            .in2(_gnd_net_),
            .in3(N__45635),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIQC4NZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__24_LC_10_32_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__24_LC_10_32_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__24_LC_10_32_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__24_LC_10_32_5  (
            .in0(N__38533),
            .in1(N__38628),
            .in2(_gnd_net_),
            .in3(N__43025),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54316),
            .ce(N__28147),
            .sr(_gnd_net_));
    defparam \u0.PIO_cmdport_T1_4_LC_11_12_3 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_T1_4_LC_11_12_3 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_cmdport_T1_4_LC_11_12_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \u0.PIO_cmdport_T1_4_LC_11_12_3  (
            .in0(_gnd_net_),
            .in1(N__51754),
            .in2(_gnd_net_),
            .in3(N__37190),
            .lcout(PIO_cmdport_T1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54218),
            .ce(N__49691),
            .sr(N__53355));
    defparam \u0.register_block_gen_PIO_dport1_reg_un6_sel_pio_dport1_i_0_LC_11_15_3 .C_ON=1'b0;
    defparam \u0.register_block_gen_PIO_dport1_reg_un6_sel_pio_dport1_i_0_LC_11_15_3 .SEQ_MODE=4'b0000;
    defparam \u0.register_block_gen_PIO_dport1_reg_un6_sel_pio_dport1_i_0_LC_11_15_3 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \u0.register_block_gen_PIO_dport1_reg_un6_sel_pio_dport1_i_0_LC_11_15_3  (
            .in0(N__51947),
            .in1(N__50868),
            .in2(_gnd_net_),
            .in3(N__46938),
            .lcout(\u0.N_446 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev0_Tm_RNIF1HR3_2_LC_11_15_7 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Tm_RNIF1HR3_2_LC_11_15_7 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev0_Tm_RNIF1HR3_2_LC_11_15_7 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \u0.DMA_dev0_Tm_RNIF1HR3_2_LC_11_15_7  (
            .in0(N__48600),
            .in1(N__46937),
            .in2(N__31206),
            .in3(N__34137),
            .lcout(\u0.dat_o_0_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_cmdport_Teoc_4_LC_11_16_2 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_Teoc_4_LC_11_16_2 .SEQ_MODE=4'b1011;
    defparam \u0.PIO_cmdport_Teoc_4_LC_11_16_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \u0.PIO_cmdport_Teoc_4_LC_11_16_2  (
            .in0(N__46105),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51950),
            .lcout(PIO_cmdport_Teoc_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54172),
            .ce(N__49698),
            .sr(N__53330));
    defparam \u0.PIO_cmdport_T1_3_LC_11_16_3 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_T1_3_LC_11_16_3 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_cmdport_T1_3_LC_11_16_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.PIO_cmdport_T1_3_LC_11_16_3  (
            .in0(N__51948),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37368),
            .lcout(PIO_cmdport_T1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54172),
            .ce(N__49698),
            .sr(N__53330));
    defparam \u0.PIO_cmdport_T1_7_LC_11_16_7 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_T1_7_LC_11_16_7 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_cmdport_T1_7_LC_11_16_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.PIO_cmdport_T1_7_LC_11_16_7  (
            .in0(N__51949),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39640),
            .lcout(PIO_cmdport_T1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54172),
            .ce(N__49698),
            .sr(N__53330));
    defparam \u1.PIO_control.PIO_access_control.T1_RNO_0_6_LC_11_17_0 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T1_RNO_0_6_LC_11_17_0 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.T1_RNO_0_6_LC_11_17_0 .LUT_INIT=16'b0101110100001100;
    LogicCell40 \u1.PIO_control.PIO_access_control.T1_RNO_0_6_LC_11_17_0  (
            .in0(N__40578),
            .in1(N__29276),
            .in2(N__40725),
            .in3(N__29460),
            .lcout(),
            .ltout(\u1.PIO_control.PIO_access_control.it1_1_iv_i_i_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T1_6_LC_11_17_1 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T1_6_LC_11_17_1 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.T1_6_LC_11_17_1 .LUT_INIT=16'b0000110000001111;
    LogicCell40 \u1.PIO_control.PIO_access_control.T1_6_LC_11_17_1  (
            .in0(_gnd_net_),
            .in1(N__40561),
            .in2(N__27376),
            .in3(N__29035),
            .lcout(\u1.PIO_control.PIO_access_control.T1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54159),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T2_4_LC_11_17_2 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T2_4_LC_11_17_2 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.T2_4_LC_11_17_2 .LUT_INIT=16'b0000000010111011;
    LogicCell40 \u1.PIO_control.PIO_access_control.T2_4_LC_11_17_2  (
            .in0(N__27363),
            .in1(N__29279),
            .in2(_gnd_net_),
            .in3(N__27388),
            .lcout(\u1.PIO_control.PIO_access_control.T2Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54159),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T1_7_LC_11_17_3 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T1_7_LC_11_17_3 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.T1_7_LC_11_17_3 .LUT_INIT=16'b0000000010111011;
    LogicCell40 \u1.PIO_control.PIO_access_control.T1_7_LC_11_17_3  (
            .in0(N__36613),
            .in1(N__29036),
            .in2(_gnd_net_),
            .in3(N__27382),
            .lcout(\u1.PIO_control.PIO_access_control.T1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54159),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T2_RNO_0_0_LC_11_17_4 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T2_RNO_0_0_LC_11_17_4 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.T2_RNO_0_0_LC_11_17_4 .LUT_INIT=16'b0011101100001010;
    LogicCell40 \u1.PIO_control.PIO_access_control.T2_RNO_0_0_LC_11_17_4  (
            .in0(N__29034),
            .in1(N__33960),
            .in2(N__36043),
            .in3(N__29461),
            .lcout(),
            .ltout(\u1.PIO_control.PIO_access_control.it2_1_iv_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T2_0_LC_11_17_5 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T2_0_LC_11_17_5 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.T2_0_LC_11_17_5 .LUT_INIT=16'b0000111100000101;
    LogicCell40 \u1.PIO_control.PIO_access_control.T2_0_LC_11_17_5  (
            .in0(N__29278),
            .in1(_gnd_net_),
            .in2(N__27463),
            .in3(N__33937),
            .lcout(\u1.PIO_control.PIO_access_control.T2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54159),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T2_RNO_0_1_LC_11_17_6 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T2_RNO_0_1_LC_11_17_6 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.T2_RNO_0_1_LC_11_17_6 .LUT_INIT=16'b0101110100001100;
    LogicCell40 \u1.PIO_control.PIO_access_control.T2_RNO_0_1_LC_11_17_6  (
            .in0(N__33981),
            .in1(N__29277),
            .in2(N__31396),
            .in3(N__29462),
            .lcout(),
            .ltout(\u1.PIO_control.PIO_access_control.it2_1_iv_i_i_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T2_1_LC_11_17_7 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T2_1_LC_11_17_7 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.T2_1_LC_11_17_7 .LUT_INIT=16'b0000110000001111;
    LogicCell40 \u1.PIO_control.PIO_access_control.T2_1_LC_11_17_7  (
            .in0(_gnd_net_),
            .in1(N__46017),
            .in2(N__27454),
            .in3(N__29037),
            .lcout(\u1.PIO_control.PIO_access_control.T2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54159),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T2_RNO_0_2_LC_11_18_0 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T2_RNO_0_2_LC_11_18_0 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.T2_RNO_0_2_LC_11_18_0 .LUT_INIT=16'b0111001101010000;
    LogicCell40 \u1.PIO_control.PIO_access_control.T2_RNO_0_2_LC_11_18_0  (
            .in0(N__39121),
            .in1(N__40197),
            .in2(N__29446),
            .in3(N__29028),
            .lcout(),
            .ltout(\u1.PIO_control.PIO_access_control.it2_1_iv_0_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T2_2_LC_11_18_1 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T2_2_LC_11_18_1 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.T2_2_LC_11_18_1 .LUT_INIT=16'b0000110000001111;
    LogicCell40 \u1.PIO_control.PIO_access_control.T2_2_LC_11_18_1  (
            .in0(_gnd_net_),
            .in1(N__43536),
            .in2(N__27442),
            .in3(N__29270),
            .lcout(\u1.PIO_control.PIO_access_control.T2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54173),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T2_RNO_0_3_LC_11_18_2 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T2_RNO_0_3_LC_11_18_2 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.T2_RNO_0_3_LC_11_18_2 .LUT_INIT=16'b0010001011110010;
    LogicCell40 \u1.PIO_control.PIO_access_control.T2_RNO_0_3_LC_11_18_2  (
            .in0(N__29268),
            .in1(N__43779),
            .in2(N__29447),
            .in3(N__43584),
            .lcout(),
            .ltout(\u1.PIO_control.PIO_access_control.it2_1_iv_i_i_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T2_3_LC_11_18_3 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T2_3_LC_11_18_3 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.T2_3_LC_11_18_3 .LUT_INIT=16'b0000111100000101;
    LogicCell40 \u1.PIO_control.PIO_access_control.T2_3_LC_11_18_3  (
            .in0(N__29029),
            .in1(_gnd_net_),
            .in2(N__27430),
            .in3(N__27423),
            .lcout(\u1.PIO_control.PIO_access_control.T2Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54173),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T2_RNO_0_4_LC_11_18_4 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T2_RNO_0_4_LC_11_18_4 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.T2_RNO_0_4_LC_11_18_4 .LUT_INIT=16'b0111010100110000;
    LogicCell40 \u1.PIO_control.PIO_access_control.T2_RNO_0_4_LC_11_18_4  (
            .in0(N__28344),
            .in1(N__36879),
            .in2(N__29445),
            .in3(N__29027),
            .lcout(\u1.PIO_control.PIO_access_control.it2_1_iv_0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T1_RNO_0_7_LC_11_18_5 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T1_RNO_0_7_LC_11_18_5 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.T1_RNO_0_7_LC_11_18_5 .LUT_INIT=16'b0101110100001100;
    LogicCell40 \u1.PIO_control.PIO_access_control.T1_RNO_0_7_LC_11_18_5  (
            .in0(N__36798),
            .in1(N__29267),
            .in2(N__36090),
            .in3(N__29389),
            .lcout(\u1.PIO_control.PIO_access_control.it1_1_iv_i_i_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T2_RNO_0_5_LC_11_18_6 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T2_RNO_0_5_LC_11_18_6 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.T2_RNO_0_5_LC_11_18_6 .LUT_INIT=16'b0010001011110010;
    LogicCell40 \u1.PIO_control.PIO_access_control.T2_RNO_0_5_LC_11_18_6  (
            .in0(N__29269),
            .in1(N__31506),
            .in2(N__29448),
            .in3(N__29634),
            .lcout(),
            .ltout(\u1.PIO_control.PIO_access_control.it2_1_iv_0_0_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T2_5_LC_11_18_7 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T2_5_LC_11_18_7 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.T2_5_LC_11_18_7 .LUT_INIT=16'b0000111100000101;
    LogicCell40 \u1.PIO_control.PIO_access_control.T2_5_LC_11_18_7  (
            .in0(N__29030),
            .in1(_gnd_net_),
            .in2(N__27529),
            .in3(N__34587),
            .lcout(\u1.PIO_control.PIO_access_control.T2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54173),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T2_RNO_0_6_LC_11_19_0 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T2_RNO_0_6_LC_11_19_0 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.T2_RNO_0_6_LC_11_19_0 .LUT_INIT=16'b0010001011110010;
    LogicCell40 \u1.PIO_control.PIO_access_control.T2_RNO_0_6_LC_11_19_0  (
            .in0(N__29213),
            .in1(N__44094),
            .in2(N__29436),
            .in3(N__43944),
            .lcout(),
            .ltout(\u1.PIO_control.PIO_access_control.it2_1_iv_i_i_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T2_6_LC_11_19_1 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T2_6_LC_11_19_1 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.T2_6_LC_11_19_1 .LUT_INIT=16'b0000111100000101;
    LogicCell40 \u1.PIO_control.PIO_access_control.T2_6_LC_11_19_1  (
            .in0(N__29039),
            .in1(_gnd_net_),
            .in2(N__27517),
            .in3(N__43509),
            .lcout(\u1.PIO_control.PIO_access_control.T2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54184),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T2_RNO_0_7_LC_11_19_2 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T2_RNO_0_7_LC_11_19_2 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.T2_RNO_0_7_LC_11_19_2 .LUT_INIT=16'b0010001011110010;
    LogicCell40 \u1.PIO_control.PIO_access_control.T2_RNO_0_7_LC_11_19_2  (
            .in0(N__29214),
            .in1(N__31483),
            .in2(N__29437),
            .in3(N__29620),
            .lcout(),
            .ltout(\u1.PIO_control.PIO_access_control.it2_1_iv_i_i_0_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T2_7_LC_11_19_3 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T2_7_LC_11_19_3 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.T2_7_LC_11_19_3 .LUT_INIT=16'b0000111100000101;
    LogicCell40 \u1.PIO_control.PIO_access_control.T2_7_LC_11_19_3  (
            .in0(N__29040),
            .in1(_gnd_net_),
            .in2(N__27505),
            .in3(N__34399),
            .lcout(\u1.PIO_control.PIO_access_control.T2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54184),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T4_RNO_0_0_LC_11_19_4 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T4_RNO_0_0_LC_11_19_4 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.T4_RNO_0_0_LC_11_19_4 .LUT_INIT=16'b0111010100110000;
    LogicCell40 \u1.PIO_control.PIO_access_control.T4_RNO_0_0_LC_11_19_4  (
            .in0(N__37059),
            .in1(N__41034),
            .in2(N__29438),
            .in3(N__29038),
            .lcout(),
            .ltout(\u1.PIO_control.PIO_access_control.it4_1_iv_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T4_0_LC_11_19_5 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T4_0_LC_11_19_5 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.T4_0_LC_11_19_5 .LUT_INIT=16'b0000110000001111;
    LogicCell40 \u1.PIO_control.PIO_access_control.T4_0_LC_11_19_5  (
            .in0(_gnd_net_),
            .in1(N__37041),
            .in2(N__27496),
            .in3(N__29215),
            .lcout(\u1.PIO_control.PIO_access_control.T4Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54184),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.Teoc_2_LC_11_19_6 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.Teoc_2_LC_11_19_6 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.Teoc_2_LC_11_19_6 .LUT_INIT=16'b0000000010111011;
    LogicCell40 \u1.PIO_control.PIO_access_control.Teoc_2_LC_11_19_6  (
            .in0(N__44301),
            .in1(N__29041),
            .in2(_gnd_net_),
            .in3(N__27550),
            .lcout(\u1.PIO_control.PIO_access_control.TeocZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54184),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.Teoc_RNO_0_3_LC_11_19_7 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.Teoc_RNO_0_3_LC_11_19_7 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.Teoc_RNO_0_3_LC_11_19_7 .LUT_INIT=16'b0101110100001100;
    LogicCell40 \u1.PIO_control.PIO_access_control.Teoc_RNO_0_3_LC_11_19_7  (
            .in0(N__37800),
            .in1(N__29212),
            .in2(N__37620),
            .in3(N__29366),
            .lcout(\u1.PIO_control.PIO_access_control.iteoc_1_iv_i_i_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T4_RNO_0_6_LC_11_20_0 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T4_RNO_0_6_LC_11_20_0 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.T4_RNO_0_6_LC_11_20_0 .LUT_INIT=16'b0101110100001100;
    LogicCell40 \u1.PIO_control.PIO_access_control.T4_RNO_0_6_LC_11_20_0  (
            .in0(N__38928),
            .in1(N__29206),
            .in2(N__37420),
            .in3(N__29402),
            .lcout(\u1.PIO_control.PIO_access_control.it4_1_iv_i_i_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.Teoc_RNO_0_0_LC_11_20_1 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.Teoc_RNO_0_0_LC_11_20_1 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.Teoc_RNO_0_0_LC_11_20_1 .LUT_INIT=16'b0010001011110010;
    LogicCell40 \u1.PIO_control.PIO_access_control.Teoc_RNO_0_0_LC_11_20_1  (
            .in0(N__29207),
            .in1(N__39993),
            .in2(N__29449),
            .in3(N__39949),
            .lcout(\u1.PIO_control.PIO_access_control.iteoc_1_iv_i_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T4_RNO_0_7_LC_11_20_2 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T4_RNO_0_7_LC_11_20_2 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.T4_RNO_0_7_LC_11_20_2 .LUT_INIT=16'b0101110100001100;
    LogicCell40 \u1.PIO_control.PIO_access_control.T4_RNO_0_7_LC_11_20_2  (
            .in0(N__44949),
            .in1(N__29210),
            .in2(N__49218),
            .in3(N__29410),
            .lcout(),
            .ltout(\u1.PIO_control.PIO_access_control.it4_1_iv_i_i_0_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T4_7_LC_11_20_3 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T4_7_LC_11_20_3 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.T4_7_LC_11_20_3 .LUT_INIT=16'b0000101000001111;
    LogicCell40 \u1.PIO_control.PIO_access_control.T4_7_LC_11_20_3  (
            .in0(N__49242),
            .in1(_gnd_net_),
            .in2(N__27586),
            .in3(N__29097),
            .lcout(\u1.PIO_control.PIO_access_control.T4Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54195),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.Teoc_RNO_0_5_LC_11_20_4 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.Teoc_RNO_0_5_LC_11_20_4 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.Teoc_RNO_0_5_LC_11_20_4 .LUT_INIT=16'b0101110100001100;
    LogicCell40 \u1.PIO_control.PIO_access_control.Teoc_RNO_0_5_LC_11_20_4  (
            .in0(N__49720),
            .in1(N__29211),
            .in2(N__44415),
            .in3(N__29411),
            .lcout(),
            .ltout(\u1.PIO_control.PIO_access_control.iteoc_1_iv_i_i_0_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.Teoc_5_LC_11_20_5 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.Teoc_5_LC_11_20_5 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.Teoc_5_LC_11_20_5 .LUT_INIT=16'b0000101000001111;
    LogicCell40 \u1.PIO_control.PIO_access_control.Teoc_5_LC_11_20_5  (
            .in0(N__43819),
            .in1(_gnd_net_),
            .in2(N__27568),
            .in3(N__29098),
            .lcout(\u1.PIO_control.PIO_access_control.TeocZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54195),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.Teoc_RNO_0_1_LC_11_20_6 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.Teoc_RNO_0_1_LC_11_20_6 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.Teoc_RNO_0_1_LC_11_20_6 .LUT_INIT=16'b0101110100001100;
    LogicCell40 \u1.PIO_control.PIO_access_control.Teoc_RNO_0_1_LC_11_20_6  (
            .in0(N__40275),
            .in1(N__29208),
            .in2(N__40240),
            .in3(N__29406),
            .lcout(\u1.PIO_control.PIO_access_control.iteoc_1_iv_i_i_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.Teoc_RNO_0_2_LC_11_20_7 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.Teoc_RNO_0_2_LC_11_20_7 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.Teoc_RNO_0_2_LC_11_20_7 .LUT_INIT=16'b0010001011110010;
    LogicCell40 \u1.PIO_control.PIO_access_control.Teoc_RNO_0_2_LC_11_20_7  (
            .in0(N__29209),
            .in1(N__44280),
            .in2(N__29450),
            .in3(N__47010),
            .lcout(\u1.PIO_control.PIO_access_control.iteoc_1_iv_i_i_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_Teoc_3_LC_11_21_2 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_Teoc_3_LC_11_21_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.DMA_timing_ctrl_Teoc_3_LC_11_21_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_Teoc_3_LC_11_21_2  (
            .in0(N__37756),
            .in1(N__37582),
            .in2(_gnd_net_),
            .in3(N__36217),
            .lcout(\u1.DMA_control.Teoc_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54205),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_cmdport_T1_RNI1BUP3_2_LC_11_21_3 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_T1_RNI1BUP3_2_LC_11_21_3 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_cmdport_T1_RNI1BUP3_2_LC_11_21_3 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \u0.PIO_cmdport_T1_RNI1BUP3_2_LC_11_21_3  (
            .in0(N__48124),
            .in1(N__48275),
            .in2(N__27862),
            .in3(N__27835),
            .lcout(\u0.dat_o_0_0_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_cmdport_T1_RNI3DUP3_3_LC_11_21_4 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_T1_RNI3DUP3_3_LC_11_21_4 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_cmdport_T1_RNI3DUP3_3_LC_11_21_4 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \u0.PIO_cmdport_T1_RNI3DUP3_3_LC_11_21_4  (
            .in0(N__48276),
            .in1(N__48125),
            .in2(N__27814),
            .in3(N__27796),
            .lcout(\u0.dat_o_0_0_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_cmdport_T1_RNI5FUP3_4_LC_11_21_5 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_T1_RNI5FUP3_4_LC_11_21_5 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_cmdport_T1_RNI5FUP3_4_LC_11_21_5 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \u0.PIO_cmdport_T1_RNI5FUP3_4_LC_11_21_5  (
            .in0(N__48126),
            .in1(N__48277),
            .in2(N__27771),
            .in3(N__27738),
            .lcout(\u0.dat_o_0_0_2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_cmdport_T1_RNI7HUP3_5_LC_11_21_6 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_T1_RNI7HUP3_5_LC_11_21_6 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_cmdport_T1_RNI7HUP3_5_LC_11_21_6 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \u0.PIO_cmdport_T1_RNI7HUP3_5_LC_11_21_6  (
            .in0(N__48278),
            .in1(N__48127),
            .in2(N__27697),
            .in3(N__31180),
            .lcout(\u0.dat_o_0_2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_cmdport_T1_RNIV8UP3_1_LC_11_21_7 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_T1_RNIV8UP3_1_LC_11_21_7 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_cmdport_T1_RNIV8UP3_1_LC_11_21_7 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \u0.PIO_cmdport_T1_RNIV8UP3_1_LC_11_21_7  (
            .in0(N__48128),
            .in1(N__27658),
            .in2(N__39241),
            .in3(N__48279),
            .lcout(\u0.dat_o_0_0_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.CtrlReg_RNI27LU1_20_LC_11_22_0 .C_ON=1'b0;
    defparam \u0.CtrlReg_RNI27LU1_20_LC_11_22_0 .SEQ_MODE=4'b0000;
    defparam \u0.CtrlReg_RNI27LU1_20_LC_11_22_0 .LUT_INIT=16'b0101000011011100;
    LogicCell40 \u0.CtrlReg_RNI27LU1_20_LC_11_22_0  (
            .in0(N__29581),
            .in1(N__45025),
            .in2(N__44911),
            .in3(N__27634),
            .lcout(),
            .ltout(\u0.dat_o_0_a2_i_2_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport0_T4_RNI8IPO9_4_LC_11_22_1 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T4_RNI8IPO9_4_LC_11_22_1 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport0_T4_RNI8IPO9_4_LC_11_22_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \u0.PIO_dport0_T4_RNI8IPO9_4_LC_11_22_1  (
            .in0(N__49644),
            .in1(N__37483),
            .in2(N__27619),
            .in3(N__27934),
            .lcout(N_211_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIQI0R_20_LC_11_22_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIQI0R_20_LC_11_22_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIQI0R_20_LC_11_22_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIQI0R_20_LC_11_22_3  (
            .in0(N__45294),
            .in1(N__30040),
            .in2(_gnd_net_),
            .in3(N__28072),
            .lcout(),
            .ltout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIQI0RZ0Z_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIA4HM1_2_LC_11_22_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIA4HM1_2_LC_11_22_4 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIA4HM1_2_LC_11_22_4 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIA4HM1_2_LC_11_22_4  (
            .in0(N__49853),
            .in1(_gnd_net_),
            .in2(N__27589),
            .in3(N__31033),
            .lcout(iQ_RNIA4HM1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNO_0_1_LC_11_22_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNO_0_1_LC_11_22_5 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNO_0_1_LC_11_22_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNO_0_1_LC_11_22_5  (
            .in0(_gnd_net_),
            .in1(N__49851),
            .in2(_gnd_net_),
            .in3(N__48768),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.N_1386_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIULD71_20_LC_11_22_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIULD71_20_LC_11_22_6 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIULD71_20_LC_11_22_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIULD71_20_LC_11_22_6  (
            .in0(N__49852),
            .in1(N__27955),
            .in2(_gnd_net_),
            .in3(N__28081),
            .lcout(),
            .ltout(mem_mem_ram6__RNIULD71_20_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.dat_o_0_a2_i_a2_20_LC_11_22_7 .C_ON=1'b0;
    defparam \u0.dat_o_0_a2_i_a2_20_LC_11_22_7 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_0_a2_i_a2_20_LC_11_22_7 .LUT_INIT=16'b0000101000100010;
    LogicCell40 \u0.dat_o_0_a2_i_a2_20_LC_11_22_7  (
            .in0(N__50466),
            .in1(N__27943),
            .in2(N__27937),
            .in3(N__48769),
            .lcout(\u0.N_1559 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIEDOD1_2_LC_11_23_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIEDOD1_2_LC_11_23_0 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIEDOD1_2_LC_11_23_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIEDOD1_2_LC_11_23_0  (
            .in0(N__28048),
            .in1(N__30196),
            .in2(_gnd_net_),
            .in3(N__49977),
            .lcout(),
            .ltout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIEDOD1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIBLN93_3_LC_11_23_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIBLN93_3_LC_11_23_1 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIBLN93_3_LC_11_23_1 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIBLN93_3_LC_11_23_1  (
            .in0(N__48830),
            .in1(N__27868),
            .in2(N__27925),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(DMAq_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.dat_o_0_0_1_2_LC_11_23_2 .C_ON=1'b0;
    defparam \u0.dat_o_0_0_1_2_LC_11_23_2 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_0_0_1_2_LC_11_23_2 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \u0.dat_o_0_0_1_2_LC_11_23_2  (
            .in0(N__47487),
            .in1(N__47213),
            .in2(N__27922),
            .in3(N__27880),
            .lcout(),
            .ltout(\u0.dat_o_0_0_1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_cmdport_T1_RNI8AUSG_2_LC_11_23_3 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_T1_RNI8AUSG_2_LC_11_23_3 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_cmdport_T1_RNI8AUSG_2_LC_11_23_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \u0.PIO_cmdport_T1_RNI8AUSG_2_LC_11_23_3  (
            .in0(N__31663),
            .in1(N__27919),
            .in2(N__27907),
            .in3(N__27904),
            .lcout(wb_dat_o_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.q_2_LC_11_23_4 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.q_2_LC_11_23_4 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.q_2_LC_11_23_4 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \u1.PIO_control.PIO_access_control.q_2_LC_11_23_4  (
            .in0(_gnd_net_),
            .in1(N__32355),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(PIOq_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54231),
            .ce(N__45907),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIASNK1_2_LC_11_23_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIASNK1_2_LC_11_23_6 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIASNK1_2_LC_11_23_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIASNK1_2_LC_11_23_6  (
            .in0(N__29947),
            .in1(N__27874),
            .in2(_gnd_net_),
            .in3(N__49978),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIASNK1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI2PUQ_15_LC_11_24_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI2PUQ_15_LC_11_24_0 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI2PUQ_15_LC_11_24_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI2PUQ_15_LC_11_24_0  (
            .in0(N__28063),
            .in1(N__28024),
            .in2(_gnd_net_),
            .in3(N__45420),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI2PUQZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__15_LC_11_24_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__15_LC_11_24_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__15_LC_11_24_1 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__15_LC_11_24_1  (
            .in0(N__32589),
            .in1(N__32473),
            .in2(N__43006),
            .in3(_gnd_net_),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54242),
            .ce(N__35891),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__31_LC_11_24_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__31_LC_11_24_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__31_LC_11_24_2 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__31_LC_11_24_2  (
            .in0(_gnd_net_),
            .in1(N__42834),
            .in2(N__32491),
            .in3(N__32590),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54242),
            .ce(N__35891),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIUO2R_31_LC_11_24_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIUO2R_31_LC_11_24_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIUO2R_31_LC_11_24_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIUO2R_31_LC_11_24_3  (
            .in0(N__45423),
            .in1(N__28018),
            .in2(_gnd_net_),
            .in3(N__28012),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIUO2RZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI2R0R_24_LC_11_24_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI2R0R_24_LC_11_24_4 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI2R0R_24_LC_11_24_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI2R0R_24_LC_11_24_4  (
            .in0(N__27982),
            .in1(N__27991),
            .in2(_gnd_net_),
            .in3(N__45421),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI2R0RZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__24_LC_11_24_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__24_LC_11_24_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__24_LC_11_24_5 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__24_LC_11_24_5  (
            .in0(N__38528),
            .in1(_gnd_net_),
            .in2(N__43007),
            .in3(N__38623),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54242),
            .ce(N__35891),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__8_LC_11_24_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__8_LC_11_24_6 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__8_LC_11_24_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__8_LC_11_24_6  (
            .in0(N__38624),
            .in1(N__42835),
            .in2(_gnd_net_),
            .in3(N__38529),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54242),
            .ce(N__35891),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI6DCM_8_LC_11_24_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI6DCM_8_LC_11_24_7 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI6DCM_8_LC_11_24_7 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI6DCM_8_LC_11_24_7  (
            .in0(N__45422),
            .in1(N__27976),
            .in2(N__28057),
            .in3(_gnd_net_),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI6DCMZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__30_LC_11_25_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__30_LC_11_25_0 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__30_LC_11_25_0 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__30_LC_11_25_0  (
            .in0(N__42579),
            .in1(N__33030),
            .in2(N__32978),
            .in3(_gnd_net_),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54257),
            .ce(N__33262),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__14_LC_11_25_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__14_LC_11_25_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__14_LC_11_25_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__14_LC_11_25_1  (
            .in0(N__33029),
            .in1(N__32963),
            .in2(_gnd_net_),
            .in3(N__42583),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54257),
            .ce(N__33262),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__4_LC_11_25_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__4_LC_11_25_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__4_LC_11_25_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__4_LC_11_25_2  (
            .in0(N__42580),
            .in1(N__31008),
            .in2(_gnd_net_),
            .in3(N__30912),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54257),
            .ce(N__33262),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__20_LC_11_25_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__20_LC_11_25_3 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__20_LC_11_25_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__20_LC_11_25_3  (
            .in0(N__31007),
            .in1(N__30911),
            .in2(_gnd_net_),
            .in3(N__42585),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54257),
            .ce(N__33262),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__5_LC_11_25_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__5_LC_11_25_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__5_LC_11_25_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__5_LC_11_25_4  (
            .in0(N__42581),
            .in1(_gnd_net_),
            .in2(N__35547),
            .in3(N__35668),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54257),
            .ce(N__33262),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__15_LC_11_25_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__15_LC_11_25_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__15_LC_11_25_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__15_LC_11_25_5  (
            .in0(N__32584),
            .in1(N__32443),
            .in2(_gnd_net_),
            .in3(N__42584),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54257),
            .ce(N__33262),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__8_LC_11_25_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__8_LC_11_25_6 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__8_LC_11_25_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__8_LC_11_25_6  (
            .in0(N__42582),
            .in1(N__38508),
            .in2(_gnd_net_),
            .in3(N__38629),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54257),
            .ce(N__33262),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__21_LC_11_25_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__21_LC_11_25_7 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__21_LC_11_25_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__21_LC_11_25_7  (
            .in0(N__35667),
            .in1(N__35517),
            .in2(_gnd_net_),
            .in3(N__42586),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54257),
            .ce(N__33262),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__2_LC_11_26_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__2_LC_11_26_0 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__2_LC_11_26_0 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__2_LC_11_26_0  (
            .in0(N__30360),
            .in1(_gnd_net_),
            .in2(N__30499),
            .in3(N__42397),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54269),
            .ce(N__41268),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__18_LC_11_26_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__18_LC_11_26_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__18_LC_11_26_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__18_LC_11_26_1  (
            .in0(N__42392),
            .in1(N__30494),
            .in2(_gnd_net_),
            .in3(N__30359),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54269),
            .ce(N__41268),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__3_LC_11_26_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__3_LC_11_26_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__3_LC_11_26_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__3_LC_11_26_2  (
            .in0(N__36409),
            .in1(N__36499),
            .in2(_gnd_net_),
            .in3(N__42398),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54269),
            .ce(N__41268),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__19_LC_11_26_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__19_LC_11_26_3 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__19_LC_11_26_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__19_LC_11_26_3  (
            .in0(N__42393),
            .in1(N__36498),
            .in2(_gnd_net_),
            .in3(N__36410),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54269),
            .ce(N__41268),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__4_LC_11_26_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__4_LC_11_26_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__4_LC_11_26_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__4_LC_11_26_4  (
            .in0(N__30914),
            .in1(N__31010),
            .in2(_gnd_net_),
            .in3(N__42399),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54269),
            .ce(N__41268),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__20_LC_11_26_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__20_LC_11_26_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__20_LC_11_26_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__20_LC_11_26_5  (
            .in0(N__42394),
            .in1(N__31009),
            .in2(_gnd_net_),
            .in3(N__30913),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54269),
            .ce(N__41268),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__14_LC_11_26_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__14_LC_11_26_6 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__14_LC_11_26_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__14_LC_11_26_6  (
            .in0(N__33054),
            .in1(N__32940),
            .in2(_gnd_net_),
            .in3(N__42396),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54269),
            .ce(N__41268),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__30_LC_11_26_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__30_LC_11_26_7 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__30_LC_11_26_7 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__30_LC_11_26_7  (
            .in0(N__42395),
            .in1(N__33055),
            .in2(N__32967),
            .in3(_gnd_net_),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54269),
            .ce(N__41268),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__9_LC_11_27_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__9_LC_11_27_0 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__9_LC_11_27_0 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__9_LC_11_27_0  (
            .in0(N__35339),
            .in1(_gnd_net_),
            .in2(N__35441),
            .in3(N__42368),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54279),
            .ce(N__41818),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__25_LC_11_27_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__25_LC_11_27_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__25_LC_11_27_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__25_LC_11_27_1  (
            .in0(N__42363),
            .in1(N__35427),
            .in2(_gnd_net_),
            .in3(N__35338),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54279),
            .ce(N__41818),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__10_LC_11_27_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__10_LC_11_27_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__10_LC_11_27_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__10_LC_11_27_2  (
            .in0(N__33853),
            .in1(N__33737),
            .in2(_gnd_net_),
            .in3(N__42365),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54279),
            .ce(N__41818),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__26_LC_11_27_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__26_LC_11_27_3 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__26_LC_11_27_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__26_LC_11_27_3  (
            .in0(N__42364),
            .in1(_gnd_net_),
            .in2(N__33755),
            .in3(N__33854),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54279),
            .ce(N__41818),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__1_LC_11_27_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__1_LC_11_27_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__1_LC_11_27_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__1_LC_11_27_4  (
            .in0(N__41520),
            .in1(N__41411),
            .in2(_gnd_net_),
            .in3(N__42366),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54279),
            .ce(N__41818),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__12_LC_11_27_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__12_LC_11_27_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__12_LC_11_27_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__12_LC_11_27_5  (
            .in0(N__42361),
            .in1(N__32194),
            .in2(_gnd_net_),
            .in3(N__32088),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54279),
            .ce(N__41818),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__28_LC_11_27_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__28_LC_11_27_6 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__28_LC_11_27_6 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__28_LC_11_27_6  (
            .in0(N__32087),
            .in1(_gnd_net_),
            .in2(N__32211),
            .in3(N__42367),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54279),
            .ce(N__41818),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__13_LC_11_27_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__13_LC_11_27_7 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__13_LC_11_27_7 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__13_LC_11_27_7  (
            .in0(N__42362),
            .in1(N__33571),
            .in2(N__33460),
            .in3(_gnd_net_),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54279),
            .ce(N__41818),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__9_LC_11_28_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__9_LC_11_28_0 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__9_LC_11_28_0 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__9_LC_11_28_0  (
            .in0(N__42387),
            .in1(_gnd_net_),
            .in2(N__35442),
            .in3(N__35340),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54289),
            .ce(N__28289),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__24_LC_11_28_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__24_LC_11_28_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__24_LC_11_28_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__24_LC_11_28_1  (
            .in0(N__38526),
            .in1(N__38618),
            .in2(_gnd_net_),
            .in3(N__42389),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54289),
            .ce(N__28289),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__16_LC_11_28_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__16_LC_11_28_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__16_LC_11_28_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__16_LC_11_28_2  (
            .in0(N__42385),
            .in1(N__41733),
            .in2(_gnd_net_),
            .in3(N__41629),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54289),
            .ce(N__28289),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__0_LC_11_28_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__0_LC_11_28_3 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__0_LC_11_28_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__0_LC_11_28_3  (
            .in0(N__41732),
            .in1(N__41628),
            .in2(_gnd_net_),
            .in3(N__42388),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54289),
            .ce(N__28289),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__10_LC_11_28_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__10_LC_11_28_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__10_LC_11_28_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__10_LC_11_28_4  (
            .in0(N__42384),
            .in1(N__33855),
            .in2(_gnd_net_),
            .in3(N__33735),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54289),
            .ce(N__28289),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__26_LC_11_28_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__26_LC_11_28_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__26_LC_11_28_5 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__26_LC_11_28_5  (
            .in0(N__33736),
            .in1(_gnd_net_),
            .in2(N__33865),
            .in3(N__42390),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54289),
            .ce(N__28289),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__1_LC_11_28_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__1_LC_11_28_6 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__1_LC_11_28_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__1_LC_11_28_6  (
            .in0(N__42386),
            .in1(_gnd_net_),
            .in2(N__41534),
            .in3(N__41412),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54289),
            .ce(N__28289),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__29_LC_11_28_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__29_LC_11_28_7 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__29_LC_11_28_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__29_LC_11_28_7  (
            .in0(N__33600),
            .in1(N__33440),
            .in2(_gnd_net_),
            .in3(N__42391),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54289),
            .ce(N__28289),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__9_LC_11_29_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__9_LC_11_29_0 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__9_LC_11_29_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__9_LC_11_29_0  (
            .in0(N__43012),
            .in1(N__35437),
            .in2(_gnd_net_),
            .in3(N__35336),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54300),
            .ce(N__28145),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__10_LC_11_29_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__10_LC_11_29_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__10_LC_11_29_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__10_LC_11_29_1  (
            .in0(N__33861),
            .in1(N__33757),
            .in2(_gnd_net_),
            .in3(N__43013),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54300),
            .ce(N__28145),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__6_LC_11_29_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__6_LC_11_29_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__6_LC_11_29_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__6_LC_11_29_2  (
            .in0(N__43011),
            .in1(N__32824),
            .in2(_gnd_net_),
            .in3(N__32692),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54300),
            .ce(N__28145),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__15_LC_11_29_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__15_LC_11_29_3 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__15_LC_11_29_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__15_LC_11_29_3  (
            .in0(N__32600),
            .in1(N__32478),
            .in2(_gnd_net_),
            .in3(N__43014),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54300),
            .ce(N__28145),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__13_LC_11_29_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__13_LC_11_29_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__13_LC_11_29_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__13_LC_11_29_4  (
            .in0(N__43009),
            .in1(N__33604),
            .in2(_gnd_net_),
            .in3(N__33457),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54300),
            .ce(N__28145),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__26_LC_11_29_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__26_LC_11_29_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__26_LC_11_29_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__26_LC_11_29_5  (
            .in0(N__33862),
            .in1(N__33758),
            .in2(_gnd_net_),
            .in3(N__43016),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54300),
            .ce(N__28145),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__31_LC_11_29_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__31_LC_11_29_6 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__31_LC_11_29_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__31_LC_11_29_6  (
            .in0(N__43010),
            .in1(N__32601),
            .in2(_gnd_net_),
            .in3(N__32479),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54300),
            .ce(N__28145),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__17_LC_11_29_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__17_LC_11_29_7 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__17_LC_11_29_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__17_LC_11_29_7  (
            .in0(N__41413),
            .in1(N__41521),
            .in2(_gnd_net_),
            .in3(N__43015),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram3_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54300),
            .ce(N__28145),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__10_LC_11_30_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__10_LC_11_30_0 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__10_LC_11_30_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__10_LC_11_30_0  (
            .in0(N__43017),
            .in1(N__33864),
            .in2(_gnd_net_),
            .in3(N__33759),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54308),
            .ce(N__30806),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__26_LC_11_30_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__26_LC_11_30_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__26_LC_11_30_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__26_LC_11_30_1  (
            .in0(N__33760),
            .in1(N__33863),
            .in2(_gnd_net_),
            .in3(N__43022),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54308),
            .ce(N__30806),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__12_LC_11_30_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__12_LC_11_30_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__12_LC_11_30_2 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__12_LC_11_30_2  (
            .in0(N__43018),
            .in1(N__32207),
            .in2(N__32102),
            .in3(_gnd_net_),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54308),
            .ce(N__30806),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__28_LC_11_30_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__28_LC_11_30_3 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__28_LC_11_30_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__28_LC_11_30_3  (
            .in0(_gnd_net_),
            .in1(N__32092),
            .in2(N__32215),
            .in3(N__43023),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54308),
            .ce(N__30806),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__13_LC_11_30_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__13_LC_11_30_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__13_LC_11_30_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__13_LC_11_30_4  (
            .in0(N__43019),
            .in1(N__33598),
            .in2(_gnd_net_),
            .in3(N__33456),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54308),
            .ce(N__30806),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__29_LC_11_30_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__29_LC_11_30_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__29_LC_11_30_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__29_LC_11_30_5  (
            .in0(N__33455),
            .in1(N__33599),
            .in2(_gnd_net_),
            .in3(N__43024),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54308),
            .ce(N__30806),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__4_LC_11_30_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__4_LC_11_30_6 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__4_LC_11_30_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__4_LC_11_30_6  (
            .in0(N__43020),
            .in1(N__31018),
            .in2(_gnd_net_),
            .in3(N__30922),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54308),
            .ce(N__30806),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__0_LC_11_30_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__0_LC_11_30_7 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__0_LC_11_30_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__0_LC_11_30_7  (
            .in0(N__41737),
            .in1(N__41641),
            .in2(_gnd_net_),
            .in3(N__43021),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54308),
            .ce(N__30806),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNISM2R_30_LC_11_31_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNISM2R_30_LC_11_31_0 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNISM2R_30_LC_11_31_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNISM2R_30_LC_11_31_0  (
            .in0(N__45656),
            .in1(N__28300),
            .in2(_gnd_net_),
            .in3(N__28207),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNISM2RZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI4VJT_30_LC_11_31_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI4VJT_30_LC_11_31_1 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI4VJT_30_LC_11_31_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI4VJT_30_LC_11_31_1  (
            .in0(N__28198),
            .in1(N__28186),
            .in2(_gnd_net_),
            .in3(N__45658),
            .lcout(),
            .ltout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI4VJTZ0Z_30_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI1SG71_30_LC_11_31_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI1SG71_30_LC_11_31_2 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI1SG71_30_LC_11_31_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI1SG71_30_LC_11_31_2  (
            .in0(N__50134),
            .in1(_gnd_net_),
            .in2(N__28333),
            .in3(N__28330),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI1SG71Z0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI0BBK_30_LC_11_31_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI0BBK_30_LC_11_31_4 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI0BBK_30_LC_11_31_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI0BBK_30_LC_11_31_4  (
            .in0(N__45657),
            .in1(N__28321),
            .in2(_gnd_net_),
            .in3(N__30592),
            .lcout(),
            .ltout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI0BBKZ0Z_30_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIECLM1_2_LC_11_31_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIECLM1_2_LC_11_31_5 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIECLM1_2_LC_11_31_5 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIECLM1_2_LC_11_31_5  (
            .in0(N__28309),
            .in1(_gnd_net_),
            .in2(N__28303),
            .in3(N__50135),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIECLM1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__30_LC_11_31_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__30_LC_11_31_6 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__30_LC_11_31_6 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__30_LC_11_31_6  (
            .in0(N__43026),
            .in1(N__33073),
            .in2(N__32968),
            .in3(_gnd_net_),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54317),
            .ce(N__35901),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__14_LC_11_31_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__14_LC_11_31_7 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__14_LC_11_31_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__14_LC_11_31_7  (
            .in0(N__33072),
            .in1(N__32945),
            .in2(_gnd_net_),
            .in3(N__43027),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54317),
            .ce(N__35901),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__12_LC_11_32_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__12_LC_11_32_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__12_LC_11_32_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__12_LC_11_32_5  (
            .in0(N__32212),
            .in1(N__32096),
            .in2(_gnd_net_),
            .in3(N__43008),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram5_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54323),
            .ce(N__28290),
            .sr(_gnd_net_));
    defparam \u0.PIO_cmdport_T1_6_LC_12_11_1 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_T1_6_LC_12_11_1 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_cmdport_T1_6_LC_12_11_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.PIO_cmdport_T1_6_LC_12_11_1  (
            .in0(N__39430),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51685),
            .lcout(PIO_cmdport_T1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54243),
            .ce(N__49690),
            .sr(N__53370));
    defparam \u0.DMA_dev0_Tm_1_LC_12_13_7 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Tm_1_LC_12_13_7 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev0_Tm_1_LC_12_13_7 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.DMA_dev0_Tm_1_LC_12_13_7  (
            .in0(N__39295),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50998),
            .lcout(DMA_dev0_Tm_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54219),
            .ce(N__39740),
            .sr(N__53356));
    defparam \u0.dat_o_0_a2_i_a2_7_16_LC_12_15_2 .C_ON=1'b0;
    defparam \u0.dat_o_0_a2_i_a2_7_16_LC_12_15_2 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_0_a2_i_a2_7_16_LC_12_15_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.dat_o_0_a2_i_a2_7_16_LC_12_15_2  (
            .in0(N__50581),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47653),
            .lcout(\u0.N_2142 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport1_T1_4_LC_12_16_0 .C_ON=1'b0;
    defparam \u0.PIO_dport1_T1_4_LC_12_16_0 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport1_T1_4_LC_12_16_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.PIO_dport1_T1_4_LC_12_16_0  (
            .in0(N__51626),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37237),
            .lcout(PIO_dport1_T1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54185),
            .ce(N__39155),
            .sr(N__53337));
    defparam \u0.PIO_dport1_T1_5_LC_12_16_1 .C_ON=1'b0;
    defparam \u0.PIO_dport1_T1_5_LC_12_16_1 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport1_T1_5_LC_12_16_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.PIO_dport1_T1_5_LC_12_16_1  (
            .in0(N__46272),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51627),
            .lcout(PIO_dport1_T1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54185),
            .ce(N__39155),
            .sr(N__53337));
    defparam \u0.PIO_dport1_T1_6_LC_12_16_2 .C_ON=1'b0;
    defparam \u0.PIO_dport1_T1_6_LC_12_16_2 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport1_T1_6_LC_12_16_2 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \u0.PIO_dport1_T1_6_LC_12_16_2  (
            .in0(N__39449),
            .in1(_gnd_net_),
            .in2(N__51867),
            .in3(_gnd_net_),
            .lcout(PIO_dport1_T1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54185),
            .ce(N__39155),
            .sr(N__53337));
    defparam \u0.PIO_dport1_T1_7_LC_12_16_3 .C_ON=1'b0;
    defparam \u0.PIO_dport1_T1_7_LC_12_16_3 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport1_T1_7_LC_12_16_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.PIO_dport1_T1_7_LC_12_16_3  (
            .in0(N__39628),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51631),
            .lcout(PIO_dport1_T1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54185),
            .ce(N__39155),
            .sr(N__53337));
    defparam \u0.PIO_dport1_T2_1_LC_12_16_5 .C_ON=1'b0;
    defparam \u0.PIO_dport1_T2_1_LC_12_16_5 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport1_T2_1_LC_12_16_5 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \u0.PIO_dport1_T2_1_LC_12_16_5  (
            .in0(N__35965),
            .in1(N__51632),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(PIO_dport1_T2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54185),
            .ce(N__39155),
            .sr(N__53337));
    defparam \u0.PIO_dport0_T1_1_LC_12_17_0 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T1_1_LC_12_17_0 .SEQ_MODE=4'b1011;
    defparam \u0.PIO_dport0_T1_1_LC_12_17_0 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \u0.PIO_dport0_T1_1_LC_12_17_0  (
            .in0(N__51633),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39341),
            .lcout(PIO_dport0_T1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54170),
            .ce(N__49380),
            .sr(N__53345));
    defparam \u0.PIO_dport0_T1_3_LC_12_17_2 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T1_3_LC_12_17_2 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport0_T1_3_LC_12_17_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.PIO_dport0_T1_3_LC_12_17_2  (
            .in0(N__51634),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37318),
            .lcout(PIO_dport0_T1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54170),
            .ce(N__49380),
            .sr(N__53345));
    defparam \u0.PIO_dport0_T2_2_LC_12_17_3 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T2_2_LC_12_17_3 .SEQ_MODE=4'b1011;
    defparam \u0.PIO_dport0_T2_2_LC_12_17_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \u0.PIO_dport0_T2_2_LC_12_17_3  (
            .in0(N__40128),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51635),
            .lcout(PIO_dport0_T2_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54170),
            .ce(N__49380),
            .sr(N__53345));
    defparam \u0.PIO_dport0_T2_4_LC_12_17_5 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T2_4_LC_12_17_5 .SEQ_MODE=4'b1011;
    defparam \u0.PIO_dport0_T2_4_LC_12_17_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \u0.PIO_dport0_T2_4_LC_12_17_5  (
            .in0(N__36990),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51636),
            .lcout(PIO_dport0_T2_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54170),
            .ce(N__49380),
            .sr(N__53345));
    defparam \u0.PIO_dport0_T4_1_LC_12_17_6 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T4_1_LC_12_17_6 .SEQ_MODE=4'b1011;
    defparam \u0.PIO_dport0_T4_1_LC_12_17_6 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \u0.PIO_dport0_T4_1_LC_12_17_6  (
            .in0(N__51637),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45134),
            .lcout(PIO_dport0_T4_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54170),
            .ce(N__49380),
            .sr(N__53345));
    defparam \u0.PIO_dport0_Teoc_0_LC_12_17_7 .C_ON=1'b0;
    defparam \u0.PIO_dport0_Teoc_0_LC_12_17_7 .SEQ_MODE=4'b1011;
    defparam \u0.PIO_dport0_Teoc_0_LC_12_17_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \u0.PIO_dport0_Teoc_0_LC_12_17_7  (
            .in0(_gnd_net_),
            .in1(N__39907),
            .in2(_gnd_net_),
            .in3(N__51638),
            .lcout(PIO_dport0_Teoc_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54170),
            .ce(N__49380),
            .sr(N__53345));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_cry_c_0_LC_12_18_0 .C_ON=1'b1;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_cry_c_0_LC_12_18_0 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_cry_c_0_LC_12_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_cry_c_0_LC_12_18_0  (
            .in0(_gnd_net_),
            .in1(N__28942),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_18_0_),
            .carryout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNO_0_1_LC_12_18_1 .C_ON=1'b1;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNO_0_1_LC_12_18_1 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNO_0_1_LC_12_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNO_0_1_LC_12_18_1  (
            .in0(_gnd_net_),
            .in1(N__28921),
            .in2(N__28727),
            .in3(N__28888),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_s_1 ),
            .ltout(),
            .carryin(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_cry_0 ),
            .carryout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNO_0_2_LC_12_18_2 .C_ON=1'b1;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNO_0_2_LC_12_18_2 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNO_0_2_LC_12_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNO_0_2_LC_12_18_2  (
            .in0(_gnd_net_),
            .in1(N__28885),
            .in2(N__28730),
            .in3(N__28861),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_s_2 ),
            .ltout(),
            .carryin(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_cry_1 ),
            .carryout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNO_0_3_LC_12_18_3 .C_ON=1'b1;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNO_0_3_LC_12_18_3 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNO_0_3_LC_12_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNO_0_3_LC_12_18_3  (
            .in0(_gnd_net_),
            .in1(N__28858),
            .in2(N__28728),
            .in3(N__28825),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_s_3 ),
            .ltout(),
            .carryin(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_cry_2 ),
            .carryout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNO_0_4_LC_12_18_4 .C_ON=1'b1;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNO_0_4_LC_12_18_4 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNO_0_4_LC_12_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNO_0_4_LC_12_18_4  (
            .in0(_gnd_net_),
            .in1(N__28822),
            .in2(N__28731),
            .in3(N__28786),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_s_4 ),
            .ltout(),
            .carryin(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_cry_3 ),
            .carryout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNO_0_5_LC_12_18_5 .C_ON=1'b1;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNO_0_5_LC_12_18_5 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNO_0_5_LC_12_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNO_0_5_LC_12_18_5  (
            .in0(_gnd_net_),
            .in1(N__28783),
            .in2(N__28729),
            .in3(N__28750),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_s_5 ),
            .ltout(),
            .carryin(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_cry_4 ),
            .carryout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNO_0_6_LC_12_18_6 .C_ON=1'b1;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNO_0_6_LC_12_18_6 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNO_0_6_LC_12_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNO_0_6_LC_12_18_6  (
            .in0(_gnd_net_),
            .in1(N__28747),
            .in2(N__28732),
            .in3(N__28357),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_s_6 ),
            .ltout(),
            .carryin(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_cry_5 ),
            .carryout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNO_0_7_LC_12_18_7 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNO_0_7_LC_12_18_7 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNO_0_7_LC_12_18_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_RNO_0_7_LC_12_18_7  (
            .in0(_gnd_net_),
            .in1(N__29563),
            .in2(_gnd_net_),
            .in3(N__29545),
            .lcout(\u1.PIO_control.PIO_access_control.PIO_timing_controller.t2_cnt.cnt.Qi_s_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.Teoc_1_LC_12_19_0 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.Teoc_1_LC_12_19_0 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.Teoc_1_LC_12_19_0 .LUT_INIT=16'b0000000011011101;
    LogicCell40 \u1.PIO_control.PIO_access_control.Teoc_1_LC_12_19_0  (
            .in0(N__29094),
            .in1(N__40260),
            .in2(_gnd_net_),
            .in3(N__29533),
            .lcout(\u1.PIO_control.PIO_access_control.TeocZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54196),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T4_RNO_0_1_LC_12_19_1 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T4_RNO_0_1_LC_12_19_1 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.T4_RNO_0_1_LC_12_19_1 .LUT_INIT=16'b0101110100001100;
    LogicCell40 \u1.PIO_control.PIO_access_control.T4_RNO_0_1_LC_12_19_1  (
            .in0(N__45750),
            .in1(N__29091),
            .in2(N__52860),
            .in3(N__29452),
            .lcout(),
            .ltout(\u1.PIO_control.PIO_access_control.it4_1_iv_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T4_1_LC_12_19_2 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T4_1_LC_12_19_2 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.T4_1_LC_12_19_2 .LUT_INIT=16'b0000110000001111;
    LogicCell40 \u1.PIO_control.PIO_access_control.T4_1_LC_12_19_2  (
            .in0(_gnd_net_),
            .in1(N__52827),
            .in2(N__29509),
            .in3(N__29281),
            .lcout(\u1.PIO_control.PIO_access_control.T4Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54196),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.Teoc_3_LC_12_19_3 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.Teoc_3_LC_12_19_3 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.Teoc_3_LC_12_19_3 .LUT_INIT=16'b0000000010111011;
    LogicCell40 \u1.PIO_control.PIO_access_control.Teoc_3_LC_12_19_3  (
            .in0(N__37779),
            .in1(N__29095),
            .in2(_gnd_net_),
            .in3(N__29488),
            .lcout(\u1.PIO_control.PIO_access_control.TeocZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54196),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.Teoc_RNO_0_4_LC_12_19_4 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.Teoc_RNO_0_4_LC_12_19_4 .SEQ_MODE=4'b0000;
    defparam \u1.PIO_control.PIO_access_control.Teoc_RNO_0_4_LC_12_19_4 .LUT_INIT=16'b0111010100110000;
    LogicCell40 \u1.PIO_control.PIO_access_control.Teoc_RNO_0_4_LC_12_19_4  (
            .in0(N__46518),
            .in1(N__36822),
            .in2(N__29464),
            .in3(N__29280),
            .lcout(),
            .ltout(\u1.PIO_control.PIO_access_control.iteoc_1_iv_i_i_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.Teoc_4_LC_12_19_5 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.Teoc_4_LC_12_19_5 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.Teoc_4_LC_12_19_5 .LUT_INIT=16'b0000110000001111;
    LogicCell40 \u1.PIO_control.PIO_access_control.Teoc_4_LC_12_19_5  (
            .in0(_gnd_net_),
            .in1(N__46623),
            .in2(N__29137),
            .in3(N__29096),
            .lcout(\u1.PIO_control.PIO_access_control.TeocZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54196),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.T4_6_LC_12_19_6 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.T4_6_LC_12_19_6 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.T4_6_LC_12_19_6 .LUT_INIT=16'b0000000011011101;
    LogicCell40 \u1.PIO_control.PIO_access_control.T4_6_LC_12_19_6  (
            .in0(N__29092),
            .in1(N__37398),
            .in2(_gnd_net_),
            .in3(N__29122),
            .lcout(\u1.PIO_control.PIO_access_control.T4Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54196),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.Teoc_0_LC_12_19_7 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.Teoc_0_LC_12_19_7 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.Teoc_0_LC_12_19_7 .LUT_INIT=16'b0000000010111011;
    LogicCell40 \u1.PIO_control.PIO_access_control.Teoc_0_LC_12_19_7  (
            .in0(N__39963),
            .in1(N__29093),
            .in2(_gnd_net_),
            .in3(N__28960),
            .lcout(\u1.PIO_control.PIO_access_control.TeocZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54196),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_cmdport_Teoc_1_LC_12_20_0 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_Teoc_1_LC_12_20_0 .SEQ_MODE=4'b1011;
    defparam \u0.PIO_cmdport_Teoc_1_LC_12_20_0 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \u0.PIO_cmdport_Teoc_1_LC_12_20_0  (
            .in0(N__51873),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40867),
            .lcout(PIO_cmdport_Teoc_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54206),
            .ce(N__49701),
            .sr(N__53364));
    defparam \u0.PIO_cmdport_Teoc_2_LC_12_20_1 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_Teoc_2_LC_12_20_1 .SEQ_MODE=4'b1011;
    defparam \u0.PIO_cmdport_Teoc_2_LC_12_20_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \u0.PIO_cmdport_Teoc_2_LC_12_20_1  (
            .in0(_gnd_net_),
            .in1(N__44230),
            .in2(_gnd_net_),
            .in3(N__51874),
            .lcout(PIO_cmdport_Teoc_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54206),
            .ce(N__49701),
            .sr(N__53364));
    defparam \u0.PIO_cmdport_T2_5_LC_12_20_3 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_T2_5_LC_12_20_3 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_cmdport_T2_5_LC_12_20_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \u0.PIO_cmdport_T2_5_LC_12_20_3  (
            .in0(_gnd_net_),
            .in1(N__34688),
            .in2(_gnd_net_),
            .in3(N__51868),
            .lcout(PIO_cmdport_T2_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54206),
            .ce(N__49701),
            .sr(N__53364));
    defparam \u0.PIO_cmdport_T2_6_LC_12_20_4 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_T2_6_LC_12_20_4 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_cmdport_T2_6_LC_12_20_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.PIO_cmdport_T2_6_LC_12_20_4  (
            .in0(N__51869),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44060),
            .lcout(PIO_cmdport_T2_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54206),
            .ce(N__49701),
            .sr(N__53364));
    defparam \u0.PIO_cmdport_T2_7_LC_12_20_5 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_T2_7_LC_12_20_5 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_cmdport_T2_7_LC_12_20_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.PIO_cmdport_T2_7_LC_12_20_5  (
            .in0(N__34542),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51870),
            .lcout(PIO_cmdport_T2_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54206),
            .ce(N__49701),
            .sr(N__53364));
    defparam \u0.PIO_cmdport_T4_0_LC_12_20_6 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_T4_0_LC_12_20_6 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_cmdport_T4_0_LC_12_20_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.PIO_cmdport_T4_0_LC_12_20_6  (
            .in0(N__51871),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41018),
            .lcout(PIO_cmdport_T4_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54206),
            .ce(N__49701),
            .sr(N__53364));
    defparam \u0.PIO_cmdport_T4_2_LC_12_20_7 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_T4_2_LC_12_20_7 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_cmdport_T4_2_LC_12_20_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \u0.PIO_cmdport_T4_2_LC_12_20_7  (
            .in0(_gnd_net_),
            .in1(N__35021),
            .in2(_gnd_net_),
            .in3(N__51872),
            .lcout(PIO_cmdport_T4_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54206),
            .ce(N__49701),
            .sr(N__53364));
    defparam \u0.PIO_cmdport_T4_3_LC_12_21_0 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_T4_3_LC_12_21_0 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_cmdport_T4_3_LC_12_21_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.PIO_cmdport_T4_3_LC_12_21_0  (
            .in0(N__34337),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51875),
            .lcout(PIO_cmdport_T4_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54220),
            .ce(N__49702),
            .sr(N__53371));
    defparam \u0.PIO_cmdport_T4_4_LC_12_21_1 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_T4_4_LC_12_21_1 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_cmdport_T4_4_LC_12_21_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.PIO_cmdport_T4_4_LC_12_21_1  (
            .in0(N__51876),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34803),
            .lcout(PIO_cmdport_T4_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54220),
            .ce(N__49702),
            .sr(N__53371));
    defparam \u0.PIO_cmdport_T4_5_LC_12_21_2 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_T4_5_LC_12_21_2 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_cmdport_T4_5_LC_12_21_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.PIO_cmdport_T4_5_LC_12_21_2  (
            .in0(N__38056),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51877),
            .lcout(PIO_cmdport_T4_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54220),
            .ce(N__49702),
            .sr(N__53371));
    defparam \u0.PIO_cmdport_T4_6_LC_12_21_3 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_T4_6_LC_12_21_3 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_cmdport_T4_6_LC_12_21_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.PIO_cmdport_T4_6_LC_12_21_3  (
            .in0(N__51878),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38183),
            .lcout(PIO_cmdport_T4_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54220),
            .ce(N__49702),
            .sr(N__53371));
    defparam \u0.PIO_cmdport_T4_7_LC_12_21_4 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_T4_7_LC_12_21_4 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_cmdport_T4_7_LC_12_21_4 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.PIO_cmdport_T4_7_LC_12_21_4  (
            .in0(N__44818),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51879),
            .lcout(PIO_cmdport_T4_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54220),
            .ce(N__49702),
            .sr(N__53371));
    defparam \u0.PIO_cmdport_Teoc_3_LC_12_21_5 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_Teoc_3_LC_12_21_5 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_cmdport_Teoc_3_LC_12_21_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.PIO_cmdport_Teoc_3_LC_12_21_5  (
            .in0(N__51880),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37707),
            .lcout(PIO_cmdport_Teoc_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54220),
            .ce(N__49702),
            .sr(N__53371));
    defparam \u0.CtrlReg_RNILK6Q3_12_LC_12_22_0 .C_ON=1'b0;
    defparam \u0.CtrlReg_RNILK6Q3_12_LC_12_22_0 .SEQ_MODE=4'b0000;
    defparam \u0.CtrlReg_RNILK6Q3_12_LC_12_22_0 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \u0.CtrlReg_RNILK6Q3_12_LC_12_22_0  (
            .in0(N__48120),
            .in1(N__48329),
            .in2(N__36883),
            .in3(N__29701),
            .lcout(),
            .ltout(\u0.dat_o_0_0_2_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev1_Td_RNISSFKG_4_LC_12_22_1 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Td_RNISSFKG_4_LC_12_22_1 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev1_Td_RNISSFKG_4_LC_12_22_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \u0.DMA_dev1_Td_RNISSFKG_4_LC_12_22_1  (
            .in0(N__29743),
            .in1(N__29671),
            .in2(N__29728),
            .in3(N__29911),
            .lcout(wb_dat_o_c_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.CtrlReg_12_LC_12_22_2 .C_ON=1'b0;
    defparam \u0.CtrlReg_12_LC_12_22_2 .SEQ_MODE=4'b1010;
    defparam \u0.CtrlReg_12_LC_12_22_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \u0.CtrlReg_12_LC_12_22_2  (
            .in0(_gnd_net_),
            .in1(N__36989),
            .in2(_gnd_net_),
            .in3(N__52059),
            .lcout(\u0.CtrlRegZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54232),
            .ce(N__53645),
            .sr(N__53380));
    defparam \u0.DMA_dev1_Td_RNITPHP3_4_LC_12_22_3 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Td_RNITPHP3_4_LC_12_22_3 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev1_Td_RNITPHP3_4_LC_12_22_3 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \u0.DMA_dev1_Td_RNITPHP3_4_LC_12_22_3  (
            .in0(N__48565),
            .in1(N__54713),
            .in2(N__29695),
            .in3(N__31560),
            .lcout(\u0.dat_o_0_0_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI26V43_3_LC_12_22_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI26V43_3_LC_12_22_4 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI26V43_3_LC_12_22_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI26V43_3_LC_12_22_4  (
            .in0(N__48831),
            .in1(N__30049),
            .in2(_gnd_net_),
            .in3(N__29992),
            .lcout(),
            .ltout(DMAq_12_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.dat_o_0_0_1_12_LC_12_22_5 .C_ON=1'b0;
    defparam \u0.dat_o_0_0_1_12_LC_12_22_5 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_0_0_1_12_LC_12_22_5 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \u0.dat_o_0_0_1_12_LC_12_22_5  (
            .in0(N__47481),
            .in1(N__47168),
            .in2(N__29932),
            .in3(N__29929),
            .lcout(\u0.dat_o_0_0_1Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.dat_o_0_0_1_4_LC_12_23_0 .C_ON=1'b0;
    defparam \u0.dat_o_0_0_1_4_LC_12_23_0 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_0_0_1_4_LC_12_23_0 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \u0.dat_o_0_0_1_4_LC_12_23_0  (
            .in0(N__47482),
            .in1(N__29821),
            .in2(N__47238),
            .in3(N__29779),
            .lcout(),
            .ltout(\u0.dat_o_0_0_1Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_cmdport_T1_RNI47VSG_4_LC_12_23_1 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_T1_RNI47VSG_4_LC_12_23_1 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_cmdport_T1_RNI47VSG_4_LC_12_23_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \u0.PIO_cmdport_T1_RNI47VSG_4_LC_12_23_1  (
            .in0(N__34411),
            .in1(N__29848),
            .in2(N__29905),
            .in3(N__29902),
            .lcout(wb_dat_o_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev0_Tm_RNIJ5HR3_4_LC_12_23_2 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Tm_RNIJ5HR3_4_LC_12_23_2 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev0_Tm_RNIJ5HR3_4_LC_12_23_2 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \u0.DMA_dev0_Tm_RNIJ5HR3_4_LC_12_23_2  (
            .in0(N__29868),
            .in1(N__46978),
            .in2(N__34822),
            .in3(N__48583),
            .lcout(\u0.dat_o_0_0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNII4OK1_2_LC_12_23_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNII4OK1_2_LC_12_23_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNII4OK1_2_LC_12_23_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNII4OK1_2_LC_12_23_3  (
            .in0(N__50059),
            .in1(N__29749),
            .in2(_gnd_net_),
            .in3(N__29839),
            .lcout(),
            .ltout(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNII4OK1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIP3O93_3_LC_12_23_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIP3O93_3_LC_12_23_4 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIP3O93_3_LC_12_23_4 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIP3O93_3_LC_12_23_4  (
            .in0(N__48910),
            .in1(_gnd_net_),
            .in2(N__29824),
            .in3(N__29761),
            .lcout(DMAq_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.q_4_LC_12_23_5 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.q_4_LC_12_23_5 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.q_4_LC_12_23_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \u1.PIO_control.PIO_access_control.q_4_LC_12_23_5  (
            .in0(N__29815),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(PIOq_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54244),
            .ce(N__45881),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIKJOD1_4_LC_12_23_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIKJOD1_4_LC_12_23_6 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIKJOD1_4_LC_12_23_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIKJOD1_4_LC_12_23_6  (
            .in0(N__29770),
            .in1(N__30136),
            .in2(_gnd_net_),
            .in3(N__50058),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIKJOD1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIU4CM_4_LC_12_24_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIU4CM_4_LC_12_24_0 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIU4CM_4_LC_12_24_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIU4CM_4_LC_12_24_0  (
            .in0(N__29755),
            .in1(N__30082),
            .in2(_gnd_net_),
            .in3(N__45464),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIU4CMZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__4_LC_12_24_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__4_LC_12_24_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__4_LC_12_24_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__4_LC_12_24_1  (
            .in0(N__42842),
            .in1(N__31006),
            .in2(_gnd_net_),
            .in3(N__30890),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54258),
            .ce(N__35878),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI4RFT_12_LC_12_24_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI4RFT_12_LC_12_24_2 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI4RFT_12_LC_12_24_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI4RFT_12_LC_12_24_2  (
            .in0(N__30076),
            .in1(N__30061),
            .in2(_gnd_net_),
            .in3(N__45466),
            .lcout(),
            .ltout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI4RFTZ0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI1MA71_12_LC_12_24_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI1MA71_12_LC_12_24_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI1MA71_12_LC_12_24_3 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI1MA71_12_LC_12_24_3  (
            .in0(N__50060),
            .in1(N__31057),
            .in2(N__30052),
            .in3(_gnd_net_),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI1MA71Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__20_LC_12_24_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__20_LC_12_24_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__20_LC_12_24_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__20_LC_12_24_4  (
            .in0(N__31005),
            .in1(N__30889),
            .in2(_gnd_net_),
            .in3(N__42843),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54258),
            .ce(N__35878),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI077K_12_LC_12_24_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI077K_12_LC_12_24_5 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI077K_12_LC_12_24_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI077K_12_LC_12_24_5  (
            .in0(N__45465),
            .in1(N__30031),
            .in2(_gnd_net_),
            .in3(N__30019),
            .lcout(),
            .ltout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI077KZ0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIE4DM1_2_LC_12_24_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIE4DM1_2_LC_12_24_6 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIE4DM1_2_LC_12_24_6 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIE4DM1_2_LC_12_24_6  (
            .in0(_gnd_net_),
            .in1(N__50064),
            .in2(N__30004),
            .in3(N__30001),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIE4DM1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI7SA71_14_LC_12_24_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI7SA71_14_LC_12_24_7 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI7SA71_14_LC_12_24_7 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI7SA71_14_LC_12_24_7  (
            .in0(N__29983),
            .in1(N__29971),
            .in2(N__50136),
            .in3(_gnd_net_),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI7SA71Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIUG4N_2_LC_12_25_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIUG4N_2_LC_12_25_0 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIUG4N_2_LC_12_25_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIUG4N_2_LC_12_25_0  (
            .in0(N__29959),
            .in1(N__29938),
            .in2(_gnd_net_),
            .in3(N__45505),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIUG4NZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__2_LC_12_25_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__2_LC_12_25_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__2_LC_12_25_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__2_LC_12_25_1  (
            .in0(N__42896),
            .in1(_gnd_net_),
            .in2(N__30367),
            .in3(N__30493),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54270),
            .ce(N__30817),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__18_LC_12_25_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__18_LC_12_25_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__18_LC_12_25_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__18_LC_12_25_2  (
            .in0(N__30492),
            .in1(N__30363),
            .in2(_gnd_net_),
            .in3(N__42897),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54270),
            .ce(N__30817),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNI0VSN_1_LC_12_25_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNI0VSN_1_LC_12_25_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNI0VSN_1_LC_12_25_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNI0VSN_1_LC_12_25_3  (
            .in0(N__45506),
            .in1(N__30241),
            .in2(_gnd_net_),
            .in3(N__30229),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNI0VSNZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNI21TN_2_LC_12_25_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNI21TN_2_LC_12_25_4 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNI21TN_2_LC_12_25_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNI21TN_2_LC_12_25_4  (
            .in0(N__30220),
            .in1(N__30205),
            .in2(_gnd_net_),
            .in3(N__45507),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNI21TNZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNI43TN_3_LC_12_25_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNI43TN_3_LC_12_25_5 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNI43TN_3_LC_12_25_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNI43TN_3_LC_12_25_5  (
            .in0(N__45508),
            .in1(N__30187),
            .in2(_gnd_net_),
            .in3(N__30175),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNI43TNZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNI65TN_4_LC_12_25_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNI65TN_4_LC_12_25_6 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNI65TN_4_LC_12_25_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNI65TN_4_LC_12_25_6  (
            .in0(N__30163),
            .in1(N__30145),
            .in2(_gnd_net_),
            .in3(N__45509),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNI65TNZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNI87TN_5_LC_12_25_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNI87TN_5_LC_12_25_7 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNI87TN_5_LC_12_25_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNI87TN_5_LC_12_25_7  (
            .in0(N__45510),
            .in1(N__30127),
            .in2(_gnd_net_),
            .in3(N__30115),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNI87TNZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI8R4N_7_LC_12_26_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI8R4N_7_LC_12_26_0 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI8R4N_7_LC_12_26_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI8R4N_7_LC_12_26_0  (
            .in0(N__45511),
            .in1(N__30088),
            .in2(_gnd_net_),
            .in3(N__30100),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI8R4NZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__7_LC_12_26_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__7_LC_12_26_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__7_LC_12_26_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__7_LC_12_26_1  (
            .in0(N__42968),
            .in1(N__38830),
            .in2(_gnd_net_),
            .in3(N__38693),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54280),
            .ce(N__30807),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__23_LC_12_26_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__23_LC_12_26_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__23_LC_12_26_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__23_LC_12_26_2  (
            .in0(N__38829),
            .in1(N__38692),
            .in2(_gnd_net_),
            .in3(N__42970),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54280),
            .ce(N__30807),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIAH7K_17_LC_12_26_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIAH7K_17_LC_12_26_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIAH7K_17_LC_12_26_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIAH7K_17_LC_12_26_3  (
            .in0(_gnd_net_),
            .in1(N__30547),
            .in2(N__30565),
            .in3(N__45512),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIAH7KZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__17_LC_12_26_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__17_LC_12_26_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__17_LC_12_26_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__17_LC_12_26_4  (
            .in0(N__41509),
            .in1(N__41382),
            .in2(_gnd_net_),
            .in3(N__42969),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54280),
            .ce(N__30807),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__1_LC_12_26_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__1_LC_12_26_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__1_LC_12_26_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__1_LC_12_26_5  (
            .in0(N__42967),
            .in1(N__41510),
            .in2(_gnd_net_),
            .in3(N__41383),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54280),
            .ce(N__30807),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNISE4N_1_LC_12_26_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNISE4N_1_LC_12_26_6 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNISE4N_1_LC_12_26_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNISE4N_1_LC_12_26_6  (
            .in0(N__45514),
            .in1(N__30541),
            .in2(_gnd_net_),
            .in3(N__30526),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNISE4NZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNICJ7K_18_LC_12_26_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNICJ7K_18_LC_12_26_7 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNICJ7K_18_LC_12_26_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNICJ7K_18_LC_12_26_7  (
            .in0(N__30520),
            .in1(N__30514),
            .in2(_gnd_net_),
            .in3(N__45513),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNICJ7KZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__29_LC_12_27_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__29_LC_12_27_0 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__29_LC_12_27_0 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__29_LC_12_27_0  (
            .in0(N__42704),
            .in1(_gnd_net_),
            .in2(N__33593),
            .in3(N__33454),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54290),
            .ce(N__33261),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__18_LC_12_27_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__18_LC_12_27_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__18_LC_12_27_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__18_LC_12_27_1  (
            .in0(N__30491),
            .in1(N__30358),
            .in2(_gnd_net_),
            .in3(N__42708),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54290),
            .ce(N__33261),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__6_LC_12_27_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__6_LC_12_27_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__6_LC_12_27_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__6_LC_12_27_2  (
            .in0(N__42705),
            .in1(N__32806),
            .in2(_gnd_net_),
            .in3(N__32682),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54290),
            .ce(N__33261),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__22_LC_12_27_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__22_LC_12_27_3 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__22_LC_12_27_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__22_LC_12_27_3  (
            .in0(N__32805),
            .in1(N__32681),
            .in2(_gnd_net_),
            .in3(N__42709),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54290),
            .ce(N__33261),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__7_LC_12_27_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__7_LC_12_27_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__7_LC_12_27_4 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__7_LC_12_27_4  (
            .in0(N__42706),
            .in1(_gnd_net_),
            .in2(N__38856),
            .in3(N__38716),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54290),
            .ce(N__33261),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__23_LC_12_27_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__23_LC_12_27_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__23_LC_12_27_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__23_LC_12_27_5  (
            .in0(N__38715),
            .in1(N__38845),
            .in2(_gnd_net_),
            .in3(N__42710),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54290),
            .ce(N__33261),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__11_LC_12_27_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__11_LC_12_27_6 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__11_LC_12_27_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__11_LC_12_27_6  (
            .in0(N__42703),
            .in1(N__43074),
            .in2(_gnd_net_),
            .in3(N__43177),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54290),
            .ce(N__33261),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__10_LC_12_27_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__10_LC_12_27_7 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__10_LC_12_27_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__10_LC_12_27_7  (
            .in0(N__33801),
            .in1(N__33696),
            .in2(_gnd_net_),
            .in3(N__42707),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54290),
            .ce(N__33261),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI4B7K_14_LC_12_28_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI4B7K_14_LC_12_28_0 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI4B7K_14_LC_12_28_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI4B7K_14_LC_12_28_0  (
            .in0(N__30598),
            .in1(N__30610),
            .in2(_gnd_net_),
            .in3(N__45615),
            .lcout(),
            .ltout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI4B7KZ0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIMCDM1_2_LC_12_28_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIMCDM1_2_LC_12_28_1 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIMCDM1_2_LC_12_28_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIMCDM1_2_LC_12_28_1  (
            .in0(N__50138),
            .in1(_gnd_net_),
            .in2(N__30601),
            .in3(N__32227),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIMCDM1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__14_LC_12_28_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__14_LC_12_28_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__14_LC_12_28_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__14_LC_12_28_2  (
            .in0(N__42830),
            .in1(N__33068),
            .in2(_gnd_net_),
            .in3(N__32944),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54301),
            .ce(N__30808),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__30_LC_12_28_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__30_LC_12_28_3 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__30_LC_12_28_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__30_LC_12_28_3  (
            .in0(_gnd_net_),
            .in1(N__32926),
            .in2(N__33076),
            .in3(N__42831),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54301),
            .ce(N__30808),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIE7IT_26_LC_12_28_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIE7IT_26_LC_12_28_4 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIE7IT_26_LC_12_28_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIE7IT_26_LC_12_28_4  (
            .in0(N__30580),
            .in1(N__30571),
            .in2(_gnd_net_),
            .in3(N__45617),
            .lcout(),
            .ltout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIE7ITZ0Z_26_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIG8E71_26_LC_12_28_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIG8E71_26_LC_12_28_5 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIG8E71_26_LC_12_28_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIG8E71_26_LC_12_28_5  (
            .in0(N__50137),
            .in1(_gnd_net_),
            .in2(N__30673),
            .in3(N__33658),
            .lcout(),
            .ltout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIG8E71Z0Z_26_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI5H753_3_LC_12_28_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI5H753_3_LC_12_28_6 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI5H753_3_LC_12_28_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI5H753_3_LC_12_28_6  (
            .in0(N__48929),
            .in1(_gnd_net_),
            .in2(N__30670),
            .in3(N__30682),
            .lcout(DMAq_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI4D9K_23_LC_12_28_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI4D9K_23_LC_12_28_7 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI4D9K_23_LC_12_28_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI4D9K_23_LC_12_28_7  (
            .in0(N__45616),
            .in1(N__30667),
            .in2(_gnd_net_),
            .in3(N__30652),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI4D9KZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNICV4N_9_LC_12_29_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNICV4N_9_LC_12_29_0 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNICV4N_9_LC_12_29_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNICV4N_9_LC_12_29_0  (
            .in0(N__45650),
            .in1(N__30634),
            .in2(_gnd_net_),
            .in3(N__30640),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNICV4NZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__9_LC_12_29_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__9_LC_12_29_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__9_LC_12_29_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__9_LC_12_29_1  (
            .in0(N__42758),
            .in1(_gnd_net_),
            .in2(N__35335),
            .in3(N__35440),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54309),
            .ce(N__30813),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__25_LC_12_29_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__25_LC_12_29_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__25_LC_12_29_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__25_LC_12_29_2  (
            .in0(N__35439),
            .in1(N__35313),
            .in2(_gnd_net_),
            .in3(N__42760),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54309),
            .ce(N__30813),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIU47K_11_LC_12_29_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIU47K_11_LC_12_29_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIU47K_11_LC_12_29_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIU47K_11_LC_12_29_3  (
            .in0(N__30628),
            .in1(N__30616),
            .in2(_gnd_net_),
            .in3(N__45651),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIU47KZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__11_LC_12_29_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__11_LC_12_29_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__11_LC_12_29_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__11_LC_12_29_4  (
            .in0(N__43205),
            .in1(N__43117),
            .in2(_gnd_net_),
            .in3(N__42759),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54309),
            .ce(N__30813),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__27_LC_12_29_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__27_LC_12_29_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__27_LC_12_29_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__27_LC_12_29_5  (
            .in0(N__42757),
            .in1(_gnd_net_),
            .in2(N__43136),
            .in3(N__43206),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54309),
            .ce(N__30813),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIU69K_20_LC_12_29_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIU69K_20_LC_12_29_6 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIU69K_20_LC_12_29_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIU69K_20_LC_12_29_6  (
            .in0(N__45652),
            .in1(N__31045),
            .in2(_gnd_net_),
            .in3(N__30823),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIU69KZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__20_LC_12_29_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__20_LC_12_29_7 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__20_LC_12_29_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram2__20_LC_12_29_7  (
            .in0(N__42756),
            .in1(N__31017),
            .in2(_gnd_net_),
            .in3(N__30921),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram2_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54309),
            .ce(N__30813),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI4BCM_7_LC_12_30_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI4BCM_7_LC_12_30_0 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI4BCM_7_LC_12_30_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI4BCM_7_LC_12_30_0  (
            .in0(N__45653),
            .in1(N__30715),
            .in2(_gnd_net_),
            .in3(N__30724),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI4BCMZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__7_LC_12_30_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__7_LC_12_30_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__7_LC_12_30_1 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__7_LC_12_30_1  (
            .in0(N__38740),
            .in1(_gnd_net_),
            .in2(N__38855),
            .in3(N__42905),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54318),
            .ce(N__35905),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__23_LC_12_30_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__23_LC_12_30_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__23_LC_12_30_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__23_LC_12_30_2  (
            .in0(N__42902),
            .in1(N__38841),
            .in2(_gnd_net_),
            .in3(N__38739),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54318),
            .ce(N__35905),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIAJ9K_26_LC_12_30_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIAJ9K_26_LC_12_30_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIAJ9K_26_LC_12_30_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIAJ9K_26_LC_12_30_3  (
            .in0(N__30709),
            .in1(N__30703),
            .in2(_gnd_net_),
            .in3(N__45655),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIAJ9KZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__26_LC_12_30_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__26_LC_12_30_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__26_LC_12_30_4 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__26_LC_12_30_4  (
            .in0(N__42903),
            .in1(_gnd_net_),
            .in2(N__33756),
            .in3(N__33860),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54318),
            .ce(N__35905),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI6V0R_26_LC_12_30_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI6V0R_26_LC_12_30_5 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI6V0R_26_LC_12_30_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI6V0R_26_LC_12_30_5  (
            .in0(N__30697),
            .in1(N__33085),
            .in2(_gnd_net_),
            .in3(N__45654),
            .lcout(),
            .ltout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI6V0RZ0Z_26_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI2THM1_2_LC_12_30_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI2THM1_2_LC_12_30_6 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI2THM1_2_LC_12_30_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI2THM1_2_LC_12_30_6  (
            .in0(_gnd_net_),
            .in1(N__30691),
            .in2(N__30685),
            .in3(N__50141),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI2THM1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__10_LC_12_30_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__10_LC_12_30_7 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__10_LC_12_30_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__10_LC_12_30_7  (
            .in0(N__33859),
            .in1(N__33741),
            .in2(_gnd_net_),
            .in3(N__42904),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54318),
            .ce(N__35905),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIA31R_28_LC_12_31_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIA31R_28_LC_12_31_0 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIA31R_28_LC_12_31_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIA31R_28_LC_12_31_0  (
            .in0(N__31990),
            .in1(N__45618),
            .in2(_gnd_net_),
            .in3(N__31141),
            .lcout(),
            .ltout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIA31RZ0Z_28_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIA5IM1_2_LC_12_31_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIA5IM1_2_LC_12_31_1 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIA5IM1_2_LC_12_31_1 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIA5IM1_2_LC_12_31_1  (
            .in0(_gnd_net_),
            .in1(N__31069),
            .in2(N__31126),
            .in3(N__50140),
            .lcout(u1_DMA_control_gen_DMAbuf_Rxbuf_mem_N_1165),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIIBIT_28_LC_12_31_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIIBIT_28_LC_12_31_2 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIIBIT_28_LC_12_31_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIIBIT_28_LC_12_31_2  (
            .in0(N__45659),
            .in1(N__31123),
            .in2(_gnd_net_),
            .in3(N__31111),
            .lcout(),
            .ltout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_N_1197_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIMEE71_28_LC_12_31_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIMEE71_28_LC_12_31_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIMEE71_28_LC_12_31_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIMEE71_28_LC_12_31_3  (
            .in0(_gnd_net_),
            .in1(N__31063),
            .in2(N__31099),
            .in3(N__50139),
            .lcout(),
            .ltout(u1_DMA_control_gen_DMAbuf_Rxbuf_mem_N_1229_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.dat_o_i_i_a2_2_28_LC_12_31_4 .C_ON=1'b0;
    defparam \u0.dat_o_i_i_a2_2_28_LC_12_31_4 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_i_i_a2_2_28_LC_12_31_4 .LUT_INIT=16'b1100010010000000;
    LogicCell40 \u0.dat_o_i_i_a2_2_28_LC_12_31_4  (
            .in0(N__48970),
            .in1(N__47254),
            .in2(N__31096),
            .in3(N__31093),
            .lcout(\u0.N_1689 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIEN9K_28_LC_12_31_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIEN9K_28_LC_12_31_5 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIEN9K_28_LC_12_31_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIEN9K_28_LC_12_31_5  (
            .in0(N__45619),
            .in1(N__31087),
            .in2(_gnd_net_),
            .in3(N__31081),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIEN9KZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__28_LC_12_31_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__28_LC_12_31_6 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__28_LC_12_31_6 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__28_LC_12_31_6  (
            .in0(N__42908),
            .in1(N__32214),
            .in2(N__32107),
            .in3(_gnd_net_),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54324),
            .ce(N__41299),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__12_LC_12_31_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__12_LC_12_31_7 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__12_LC_12_31_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__12_LC_12_31_7  (
            .in0(N__32213),
            .in1(N__32103),
            .in2(_gnd_net_),
            .in3(N__42909),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54324),
            .ce(N__41299),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI6P4N_6_LC_12_32_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI6P4N_6_LC_12_32_0 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI6P4N_6_LC_12_32_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI6P4N_6_LC_12_32_0  (
            .in0(N__45692),
            .in1(N__31261),
            .in2(_gnd_net_),
            .in3(N__31252),
            .lcout(),
            .ltout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI6P4NZ0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIQCOK1_2_LC_12_32_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIQCOK1_2_LC_12_32_1 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIQCOK1_2_LC_12_32_1 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIQCOK1_2_LC_12_32_1  (
            .in0(_gnd_net_),
            .in1(N__50205),
            .in2(N__31240),
            .in3(N__31216),
            .lcout(iQ_RNIQCOK1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI29CM_6_LC_12_32_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI29CM_6_LC_12_32_6 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI29CM_6_LC_12_32_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI29CM_6_LC_12_32_6  (
            .in0(N__45691),
            .in1(N__31966),
            .in2(_gnd_net_),
            .in3(N__31225),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI29CMZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev0_Tm_2_LC_13_15_1 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Tm_2_LC_13_15_1 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev0_Tm_2_LC_13_15_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.DMA_dev0_Tm_2_LC_13_15_1  (
            .in0(N__34236),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51696),
            .lcout(DMA_dev0_Tm_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54207),
            .ce(N__39736),
            .sr(N__53351));
    defparam \u0.PIO_cmdport_T1_0_LC_13_16_0 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_T1_0_LC_13_16_0 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_cmdport_T1_0_LC_13_16_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.PIO_cmdport_T1_0_LC_13_16_0  (
            .in0(N__49493),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51549),
            .lcout(PIO_cmdport_T1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54197),
            .ce(N__49694),
            .sr(N__53343));
    defparam \u0.PIO_cmdport_Teoc_6_LC_13_17_0 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_Teoc_6_LC_13_17_0 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_cmdport_Teoc_6_LC_13_17_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.PIO_cmdport_Teoc_6_LC_13_17_0  (
            .in0(N__47838),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51551),
            .lcout(PIO_cmdport_Teoc_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54181),
            .ce(N__49697),
            .sr(N__53352));
    defparam \u0.PIO_cmdport_Teoc_7_LC_13_17_1 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_Teoc_7_LC_13_17_1 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_cmdport_Teoc_7_LC_13_17_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.PIO_cmdport_Teoc_7_LC_13_17_1  (
            .in0(N__51552),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40527),
            .lcout(PIO_cmdport_Teoc_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54181),
            .ce(N__49697),
            .sr(N__53352));
    defparam \u0.PIO_cmdport_T1_5_LC_13_17_3 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_T1_5_LC_13_17_3 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_cmdport_T1_5_LC_13_17_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.PIO_cmdport_T1_5_LC_13_17_3  (
            .in0(N__51550),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46271),
            .lcout(PIO_cmdport_T1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54181),
            .ce(N__49697),
            .sr(N__53352));
    defparam \u0.DMA_dev1_Td_RNI4B7N3_0_LC_13_18_0 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Td_RNI4B7N3_0_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev1_Td_RNI4B7N3_0_LC_13_18_0 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \u0.DMA_dev1_Td_RNI4B7N3_0_LC_13_18_0  (
            .in0(N__31326),
            .in1(N__46960),
            .in2(N__33936),
            .in3(N__54708),
            .lcout(\u0.dat_o_0_0_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_cmdport_T2_RNIGRQJ3_0_LC_13_18_2 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_T2_RNIGRQJ3_0_LC_13_18_2 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_cmdport_T2_RNIGRQJ3_0_LC_13_18_2 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \u0.PIO_cmdport_T2_RNIGRQJ3_0_LC_13_18_2  (
            .in0(N__50757),
            .in1(N__48134),
            .in2(N__33961),
            .in3(N__36042),
            .lcout(\u0.dat_o_0_0_3_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_cmdport_T2_RNI2D6I3_1_LC_13_18_3 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_T2_RNI2D6I3_1_LC_13_18_3 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_cmdport_T2_RNI2D6I3_1_LC_13_18_3 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \u0.PIO_cmdport_T2_RNI2D6I3_1_LC_13_18_3  (
            .in0(N__48133),
            .in1(N__46589),
            .in2(N__33985),
            .in3(N__31447),
            .lcout(\u0.dat_o_0_0_3_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev1_Td_RNI6D7N3_1_LC_13_18_5 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Td_RNI6D7N3_1_LC_13_18_5 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev1_Td_RNI6D7N3_1_LC_13_18_5 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \u0.DMA_dev1_Td_RNI6D7N3_1_LC_13_18_5  (
            .in0(N__46961),
            .in1(N__31302),
            .in2(N__54718),
            .in3(N__31395),
            .lcout(\u0.dat_o_0_0_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev1_Td_RNIIP7N3_7_LC_13_18_6 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Td_RNIIP7N3_7_LC_13_18_6 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev1_Td_RNIIP7N3_7_LC_13_18_6 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \u0.DMA_dev1_Td_RNIIP7N3_7_LC_13_18_6  (
            .in0(N__31482),
            .in1(N__46962),
            .in2(N__31375),
            .in3(N__54712),
            .lcout(\u0.dat_o_0_0_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.register_block_gen_DMA_dev1_reg_un6_sel_dma_dev1_i_0_LC_13_19_0 .C_ON=1'b0;
    defparam \u0.register_block_gen_DMA_dev1_reg_un6_sel_dma_dev1_i_0_LC_13_19_0 .SEQ_MODE=4'b0000;
    defparam \u0.register_block_gen_DMA_dev1_reg_un6_sel_dma_dev1_i_0_LC_13_19_0 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \u0.register_block_gen_DMA_dev1_reg_un6_sel_dma_dev1_i_0_LC_13_19_0  (
            .in0(N__51541),
            .in1(N__50850),
            .in2(_gnd_net_),
            .in3(N__54707),
            .lcout(\u0.N_442 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev1_Td_0_LC_13_19_1 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Td_0_LC_13_19_1 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev1_Td_0_LC_13_19_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.DMA_dev1_Td_0_LC_13_19_1  (
            .in0(N__51917),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54465),
            .lcout(DMA_dev1_Td_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54208),
            .ce(N__39532),
            .sr(N__53365));
    defparam \u0.DMA_dev1_Td_1_LC_13_19_2 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Td_1_LC_13_19_2 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev1_Td_1_LC_13_19_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \u0.DMA_dev1_Td_1_LC_13_19_2  (
            .in0(_gnd_net_),
            .in1(N__35985),
            .in2(_gnd_net_),
            .in3(N__51918),
            .lcout(DMA_dev1_Td_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54208),
            .ce(N__39532),
            .sr(N__53365));
    defparam \u0.DMA_dev1_Td_2_LC_13_19_3 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Td_2_LC_13_19_3 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev1_Td_2_LC_13_19_3 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \u0.DMA_dev1_Td_2_LC_13_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__52110),
            .in3(N__40185),
            .lcout(DMA_dev1_Td_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54208),
            .ce(N__39532),
            .sr(N__53365));
    defparam \u0.DMA_dev1_Td_3_LC_13_19_4 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Td_3_LC_13_19_4 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev1_Td_3_LC_13_19_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \u0.DMA_dev1_Td_3_LC_13_19_4  (
            .in0(_gnd_net_),
            .in1(N__51922),
            .in2(_gnd_net_),
            .in3(N__43701),
            .lcout(DMA_dev1_Td_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54208),
            .ce(N__39532),
            .sr(N__53365));
    defparam \u0.DMA_dev1_Td_4_LC_13_19_5 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Td_4_LC_13_19_5 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev1_Td_4_LC_13_19_5 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \u0.DMA_dev1_Td_4_LC_13_19_5  (
            .in0(N__51923),
            .in1(N__36971),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(DMA_dev1_Td_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54208),
            .ce(N__39532),
            .sr(N__53365));
    defparam \u0.DMA_dev1_Td_5_LC_13_19_6 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Td_5_LC_13_19_6 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev1_Td_5_LC_13_19_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.DMA_dev1_Td_5_LC_13_19_6  (
            .in0(N__34666),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51924),
            .lcout(DMA_dev1_Td_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54208),
            .ce(N__39532),
            .sr(N__53365));
    defparam \u0.DMA_dev1_Td_6_LC_13_19_7 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Td_6_LC_13_19_7 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev1_Td_6_LC_13_19_7 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \u0.DMA_dev1_Td_6_LC_13_19_7  (
            .in0(N__44058),
            .in1(_gnd_net_),
            .in2(N__52111),
            .in3(_gnd_net_),
            .lcout(DMA_dev1_Td_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54208),
            .ce(N__39532),
            .sr(N__53365));
    defparam \u0.PIO_dport1_T2_5_LC_13_20_1 .C_ON=1'b0;
    defparam \u0.PIO_dport1_T2_5_LC_13_20_1 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport1_T2_5_LC_13_20_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \u0.PIO_dport1_T2_5_LC_13_20_1  (
            .in0(_gnd_net_),
            .in1(N__34687),
            .in2(_gnd_net_),
            .in3(N__51542),
            .lcout(PIO_dport1_T2_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54221),
            .ce(N__39206),
            .sr(N__53372));
    defparam \u0.PIO_dport1_T2_6_LC_13_20_2 .C_ON=1'b0;
    defparam \u0.PIO_dport1_T2_6_LC_13_20_2 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport1_T2_6_LC_13_20_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.PIO_dport1_T2_6_LC_13_20_2  (
            .in0(N__51543),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44061),
            .lcout(PIO_dport1_T2_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54221),
            .ce(N__39206),
            .sr(N__53372));
    defparam \u0.PIO_dport1_T2_7_LC_13_20_3 .C_ON=1'b0;
    defparam \u0.PIO_dport1_T2_7_LC_13_20_3 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport1_T2_7_LC_13_20_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.PIO_dport1_T2_7_LC_13_20_3  (
            .in0(N__34541),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51544),
            .lcout(PIO_dport1_T2_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54221),
            .ce(N__39206),
            .sr(N__53372));
    defparam \u0.PIO_dport1_T4_0_LC_13_20_4 .C_ON=1'b0;
    defparam \u0.PIO_dport1_T4_0_LC_13_20_4 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport1_T4_0_LC_13_20_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.PIO_dport1_T4_0_LC_13_20_4  (
            .in0(N__51545),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41019),
            .lcout(PIO_dport1_T4_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54221),
            .ce(N__39206),
            .sr(N__53372));
    defparam \u0.PIO_dport1_T4_2_LC_13_20_5 .C_ON=1'b0;
    defparam \u0.PIO_dport1_T4_2_LC_13_20_5 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport1_T4_2_LC_13_20_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.PIO_dport1_T4_2_LC_13_20_5  (
            .in0(N__35036),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51546),
            .lcout(PIO_dport1_T4_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54221),
            .ce(N__39206),
            .sr(N__53372));
    defparam \u0.PIO_dport1_T4_3_LC_13_20_6 .C_ON=1'b0;
    defparam \u0.PIO_dport1_T4_3_LC_13_20_6 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport1_T4_3_LC_13_20_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.PIO_dport1_T4_3_LC_13_20_6  (
            .in0(N__51547),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34369),
            .lcout(PIO_dport1_T4_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54221),
            .ce(N__39206),
            .sr(N__53372));
    defparam \u0.PIO_dport1_T4_4_LC_13_20_7 .C_ON=1'b0;
    defparam \u0.PIO_dport1_T4_4_LC_13_20_7 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport1_T4_4_LC_13_20_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \u0.PIO_dport1_T4_4_LC_13_20_7  (
            .in0(_gnd_net_),
            .in1(N__34804),
            .in2(_gnd_net_),
            .in3(N__51548),
            .lcout(PIO_dport1_T4_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54221),
            .ce(N__39206),
            .sr(N__53372));
    defparam \u0.PIO_dport0_T1_RNIDVGR3_1_LC_13_21_1 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T1_RNIDVGR3_1_LC_13_21_1 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport0_T1_RNIDVGR3_1_LC_13_21_1 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \u0.PIO_dport0_T1_RNIDVGR3_1_LC_13_21_1  (
            .in0(N__50748),
            .in1(N__54686),
            .in2(N__31761),
            .in3(N__31735),
            .lcout(\u0.dat_o_0_0_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport0_T1_RNIF1HR3_2_LC_13_21_2 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T1_RNIF1HR3_2_LC_13_21_2 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport0_T1_RNIF1HR3_2_LC_13_21_2 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \u0.PIO_dport0_T1_RNIF1HR3_2_LC_13_21_2  (
            .in0(N__54687),
            .in1(N__50749),
            .in2(N__31714),
            .in3(N__31683),
            .lcout(\u0.dat_o_0_0_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport0_T1_RNIH3HR3_3_LC_13_21_3 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T1_RNIH3HR3_3_LC_13_21_3 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport0_T1_RNIH3HR3_3_LC_13_21_3 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \u0.PIO_dport0_T1_RNIH3HR3_3_LC_13_21_3  (
            .in0(N__50750),
            .in1(N__54688),
            .in2(N__37273),
            .in3(N__31651),
            .lcout(\u0.dat_o_0_0_3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport0_T1_RNIL7HR3_5_LC_13_21_5 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T1_RNIL7HR3_5_LC_13_21_5 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport0_T1_RNIL7HR3_5_LC_13_21_5 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \u0.PIO_dport0_T1_RNIL7HR3_5_LC_13_21_5  (
            .in0(N__50751),
            .in1(N__54689),
            .in2(N__46177),
            .in3(N__37828),
            .lcout(\u0.dat_o_0_3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_Td_6_LC_13_21_6 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_Td_6_LC_13_21_6 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.DMA_timing_ctrl_Td_6_LC_13_21_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_Td_6_LC_13_21_6  (
            .in0(N__43485),
            .in1(N__44122),
            .in2(_gnd_net_),
            .in3(N__36241),
            .lcout(\u1.DMA_control.Td_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54233),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNINMOD1_5_LC_13_22_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNINMOD1_5_LC_13_22_0 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNINMOD1_5_LC_13_22_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNINMOD1_5_LC_13_22_0  (
            .in0(N__49937),
            .in1(N__31615),
            .in2(_gnd_net_),
            .in3(N__31603),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNINMOD1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIM8OK1_2_LC_13_22_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIM8OK1_2_LC_13_22_1 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIM8OK1_2_LC_13_22_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIM8OK1_2_LC_13_22_1  (
            .in0(N__31591),
            .in1(N__31768),
            .in2(_gnd_net_),
            .in3(N__49938),
            .lcout(),
            .ltout(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIM8OK1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI0BO93_3_LC_13_22_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI0BO93_3_LC_13_22_2 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI0BO93_3_LC_13_22_2 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI0BO93_3_LC_13_22_2  (
            .in0(_gnd_net_),
            .in1(N__31573),
            .in2(N__31567),
            .in3(N__48832),
            .lcout(),
            .ltout(DMAq_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.dat_o_0_1_5_LC_13_22_3 .C_ON=1'b0;
    defparam \u0.dat_o_0_1_5_LC_13_22_3 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_0_1_5_LC_13_22_3 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \u0.dat_o_0_1_5_LC_13_22_3  (
            .in0(N__31840),
            .in1(N__47183),
            .in2(N__31564),
            .in3(N__47435),
            .lcout(),
            .ltout(\u0.dat_o_0_1Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_cmdport_T1_RNIILVSG_5_LC_13_22_4 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_T1_RNIILVSG_5_LC_13_22_4 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_cmdport_T1_RNIILVSG_5_LC_13_22_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \u0.PIO_cmdport_T1_RNIILVSG_5_LC_13_22_4  (
            .in0(N__31876),
            .in1(N__31951),
            .in2(N__31939),
            .in3(N__31936),
            .lcout(wb_dat_o_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev0_Tm_RNIL7HR3_5_LC_13_22_5 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Tm_RNIL7HR3_5_LC_13_22_5 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev0_Tm_RNIL7HR3_5_LC_13_22_5 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \u0.DMA_dev0_Tm_RNIL7HR3_5_LC_13_22_5  (
            .in0(N__46940),
            .in1(N__35161),
            .in2(N__31906),
            .in3(N__48582),
            .lcout(\u0.dat_o_0_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.q_5_LC_13_22_6 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.q_5_LC_13_22_6 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.q_5_LC_13_22_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \u1.PIO_control.PIO_access_control.q_5_LC_13_22_6  (
            .in0(N__31870),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(PIOq_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54245),
            .ce(N__45899),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_Tm_3_LC_13_23_1 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_Tm_3_LC_13_23_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.DMA_timing_ctrl_Tm_3_LC_13_23_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_Tm_3_LC_13_23_1  (
            .in0(N__37269),
            .in1(N__34833),
            .in2(_gnd_net_),
            .in3(N__36253),
            .lcout(\u1.DMA_control.Tm_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54259),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_Tm_4_LC_13_23_2 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_Tm_4_LC_13_23_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.DMA_timing_ctrl_Tm_4_LC_13_23_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_Tm_4_LC_13_23_2  (
            .in0(N__36254),
            .in1(_gnd_net_),
            .in2(N__37855),
            .in3(N__34815),
            .lcout(\u1.DMA_control.Tm_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54259),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_Tm_5_LC_13_23_3 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_Tm_5_LC_13_23_3 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.DMA_timing_ctrl_Tm_5_LC_13_23_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_Tm_5_LC_13_23_3  (
            .in0(N__37827),
            .in1(N__35157),
            .in2(_gnd_net_),
            .in3(N__36255),
            .lcout(\u1.DMA_control.Tm_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54259),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.DMA_timing_ctrl_Tm_6_LC_13_23_4 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_Tm_6_LC_13_23_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.DMA_timing_ctrl_Tm_6_LC_13_23_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_Tm_6_LC_13_23_4  (
            .in0(N__36256),
            .in1(N__40705),
            .in2(_gnd_net_),
            .in3(N__40746),
            .lcout(\u1.DMA_control.Tm_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54259),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI07CM_5_LC_13_23_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI07CM_5_LC_13_23_6 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI07CM_5_LC_13_23_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI07CM_5_LC_13_23_6  (
            .in0(N__31780),
            .in1(N__45462),
            .in2(_gnd_net_),
            .in3(N__31972),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI07CMZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI0NUQ_14_LC_13_23_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI0NUQ_14_LC_13_23_7 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI0NUQ_14_LC_13_23_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI0NUQ_14_LC_13_23_7  (
            .in0(N__32257),
            .in1(N__32245),
            .in2(_gnd_net_),
            .in3(N__45463),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI0NUQZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__17_LC_13_24_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__17_LC_13_24_0 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__17_LC_13_24_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__17_LC_13_24_0  (
            .in0(N__41402),
            .in1(N__41513),
            .in2(_gnd_net_),
            .in3(N__42849),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54271),
            .ce(N__35892),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__28_LC_13_24_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__28_LC_13_24_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__28_LC_13_24_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__28_LC_13_24_1  (
            .in0(N__42846),
            .in1(N__32173),
            .in2(_gnd_net_),
            .in3(N__32075),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54271),
            .ce(N__35892),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__13_LC_13_24_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__13_LC_13_24_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__13_LC_13_24_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__13_LC_13_24_2  (
            .in0(N__33560),
            .in1(N__33450),
            .in2(_gnd_net_),
            .in3(N__42848),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54271),
            .ce(N__35892),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__29_LC_13_24_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__29_LC_13_24_3 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__29_LC_13_24_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__29_LC_13_24_3  (
            .in0(N__42847),
            .in1(_gnd_net_),
            .in2(N__33463),
            .in3(N__33561),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54271),
            .ce(N__35892),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__5_LC_13_24_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__5_LC_13_24_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__5_LC_13_24_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__5_LC_13_24_4  (
            .in0(N__35495),
            .in1(N__35654),
            .in2(_gnd_net_),
            .in3(N__42850),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54271),
            .ce(N__35892),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__21_LC_13_24_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__21_LC_13_24_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__21_LC_13_24_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__21_LC_13_24_5  (
            .in0(N__42844),
            .in1(N__35653),
            .in2(_gnd_net_),
            .in3(N__35494),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54271),
            .ce(N__35892),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__6_LC_13_24_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__6_LC_13_24_6 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__6_LC_13_24_6 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__6_LC_13_24_6  (
            .in0(N__32634),
            .in1(_gnd_net_),
            .in2(N__32795),
            .in3(N__42851),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54271),
            .ce(N__35892),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__22_LC_13_24_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__22_LC_13_24_7 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__22_LC_13_24_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__22_LC_13_24_7  (
            .in0(N__42845),
            .in1(N__32763),
            .in2(_gnd_net_),
            .in3(N__32633),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54271),
            .ce(N__35892),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_14_LC_13_25_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_14_LC_13_25_0 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_14_LC_13_25_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_readDlw_14_LC_13_25_0  (
            .in0(N__32865),
            .in1(N__40682),
            .in2(_gnd_net_),
            .in3(N__42898),
            .lcout(\u1.DMA_control.readDlw_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54281),
            .ce(N__36324),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_14_LC_13_25_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_14_LC_13_25_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_14_LC_13_25_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_readDfw_14_LC_13_25_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33028),
            .lcout(\u1.DMA_control.readDfw_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54281),
            .ce(N__36324),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_6_LC_13_25_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_6_LC_13_25_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_6_LC_13_25_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_readDlw_6_LC_13_25_2  (
            .in0(N__32866),
            .in1(N__40683),
            .in2(_gnd_net_),
            .in3(N__42900),
            .lcout(\u1.DMA_control.readDlw_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54281),
            .ce(N__36324),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_6_LC_13_25_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_6_LC_13_25_3 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_6_LC_13_25_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_readDfw_6_LC_13_25_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32762),
            .lcout(\u1.DMA_control.readDfw_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54281),
            .ce(N__36324),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_15_LC_13_25_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_15_LC_13_25_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_15_LC_13_25_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_readDlw_15_LC_13_25_4  (
            .in0(N__32391),
            .in1(N__38390),
            .in2(_gnd_net_),
            .in3(N__42899),
            .lcout(\u1.DMA_control.readDlw_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54281),
            .ce(N__36324),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_15_LC_13_25_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_15_LC_13_25_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_15_LC_13_25_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_readDfw_15_LC_13_25_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32549),
            .lcout(\u1.DMA_control.readDfw_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54281),
            .ce(N__36324),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_7_LC_13_25_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_7_LC_13_25_6 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_7_LC_13_25_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_readDlw_7_LC_13_25_6  (
            .in0(N__32392),
            .in1(N__38391),
            .in2(_gnd_net_),
            .in3(N__42901),
            .lcout(\u1.DMA_control.readDlw_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54281),
            .ce(N__36324),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_7_LC_13_25_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_7_LC_13_25_7 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_7_LC_13_25_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_readDfw_7_LC_13_25_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38804),
            .lcout(\u1.DMA_control.readDfw_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54281),
            .ce(N__36324),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_10_LC_13_26_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_10_LC_13_26_0 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_10_LC_13_26_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_readDlw_10_LC_13_26_0  (
            .in0(N__32356),
            .in1(N__32302),
            .in2(_gnd_net_),
            .in3(N__42971),
            .lcout(\u1.DMA_control.readDlw_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54291),
            .ce(N__36323),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_10_LC_13_26_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_10_LC_13_26_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_10_LC_13_26_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_readDfw_10_LC_13_26_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33824),
            .lcout(\u1.DMA_control.readDfw_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54291),
            .ce(N__36323),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_11_LC_13_26_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_11_LC_13_26_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_11_LC_13_26_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_readDlw_11_LC_13_26_4  (
            .in0(N__33123),
            .in1(N__34911),
            .in2(_gnd_net_),
            .in3(N__42972),
            .lcout(\u1.DMA_control.readDlw_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54291),
            .ce(N__36323),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_11_LC_13_26_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_11_LC_13_26_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_11_LC_13_26_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_readDfw_11_LC_13_26_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43094),
            .lcout(\u1.DMA_control.readDfw_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54291),
            .ce(N__36323),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_3_LC_13_26_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_3_LC_13_26_6 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_3_LC_13_26_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_readDlw_3_LC_13_26_6  (
            .in0(N__33124),
            .in1(N__34912),
            .in2(_gnd_net_),
            .in3(N__42973),
            .lcout(\u1.DMA_control.readDlw_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54291),
            .ce(N__36323),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_9_LC_13_26_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_9_LC_13_26_7 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_9_LC_13_26_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_readDfw_9_LC_13_26_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35398),
            .lcout(\u1.DMA_control.readDfw_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54291),
            .ce(N__36323),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__27_LC_13_27_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__27_LC_13_27_0 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__27_LC_13_27_0 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__27_LC_13_27_0  (
            .in0(N__42928),
            .in1(_gnd_net_),
            .in2(N__43095),
            .in3(N__43176),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54302),
            .ce(N__33256),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__25_LC_13_27_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__25_LC_13_27_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__25_LC_13_27_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__25_LC_13_27_1  (
            .in0(N__35375),
            .in1(N__35310),
            .in2(_gnd_net_),
            .in3(N__42931),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54302),
            .ce(N__33256),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__16_LC_13_27_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__16_LC_13_27_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__16_LC_13_27_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__16_LC_13_27_2  (
            .in0(N__42926),
            .in1(N__41584),
            .in2(_gnd_net_),
            .in3(N__41684),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54302),
            .ce(N__33256),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__0_LC_13_27_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__0_LC_13_27_3 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__0_LC_13_27_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__0_LC_13_27_3  (
            .in0(N__41683),
            .in1(N__41583),
            .in2(_gnd_net_),
            .in3(N__42929),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54302),
            .ce(N__33256),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__13_LC_13_27_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__13_LC_13_27_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__13_LC_13_27_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__13_LC_13_27_4  (
            .in0(N__42925),
            .in1(N__33575),
            .in2(_gnd_net_),
            .in3(N__33462),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54302),
            .ce(N__33256),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__26_LC_13_27_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__26_LC_13_27_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__26_LC_13_27_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__26_LC_13_27_5  (
            .in0(N__33712),
            .in1(N__33800),
            .in2(_gnd_net_),
            .in3(N__42932),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54302),
            .ce(N__33256),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__1_LC_13_27_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__1_LC_13_27_6 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__1_LC_13_27_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__1_LC_13_27_6  (
            .in0(N__42927),
            .in1(N__41512),
            .in2(_gnd_net_),
            .in3(N__41372),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54302),
            .ce(N__33256),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__17_LC_13_27_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__17_LC_13_27_7 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__17_LC_13_27_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram1__17_LC_13_27_7  (
            .in0(N__41511),
            .in1(N__41371),
            .in2(_gnd_net_),
            .in3(N__42930),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram1_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54302),
            .ce(N__33256),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIGP9K_29_LC_13_28_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIGP9K_29_LC_13_28_0 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIGP9K_29_LC_13_28_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIGP9K_29_LC_13_28_0  (
            .in0(N__45661),
            .in1(N__33217),
            .in2(_gnd_net_),
            .in3(N__33205),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIGP9KZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIKDIT_29_LC_13_28_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIKDIT_29_LC_13_28_1 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIKDIT_29_LC_13_28_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIKDIT_29_LC_13_28_1  (
            .in0(N__33193),
            .in1(N__33184),
            .in2(_gnd_net_),
            .in3(N__45662),
            .lcout(),
            .ltout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIKDITZ0Z_29_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIPHE71_29_LC_13_28_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIPHE71_29_LC_13_28_2 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIPHE71_29_LC_13_28_2 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIPHE71_29_LC_13_28_2  (
            .in0(_gnd_net_),
            .in1(N__33130),
            .in2(N__33169),
            .in3(N__50152),
            .lcout(),
            .ltout(mem_mem_ram6__RNIPHE71_29_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.dat_o_i_i_a2_2_29_LC_13_28_3 .C_ON=1'b0;
    defparam \u0.dat_o_i_i_a2_2_29_LC_13_28_3 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_i_i_a2_2_29_LC_13_28_3 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \u0.dat_o_i_i_a2_2_29_LC_13_28_3  (
            .in0(N__33136),
            .in1(N__47249),
            .in2(N__33166),
            .in3(N__48930),
            .lcout(\u0.N_1696 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIC51R_29_LC_13_28_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIC51R_29_LC_13_28_4 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIC51R_29_LC_13_28_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIC51R_29_LC_13_28_4  (
            .in0(N__45660),
            .in1(N__33163),
            .in2(_gnd_net_),
            .in3(N__33151),
            .lcout(),
            .ltout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIC51RZ0Z_29_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIE9IM1_2_LC_13_28_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIE9IM1_2_LC_13_28_5 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIE9IM1_2_LC_13_28_5 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIE9IM1_2_LC_13_28_5  (
            .in0(N__50153),
            .in1(N__33145),
            .in2(N__33139),
            .in3(_gnd_net_),
            .lcout(iQ_RNIE9IM1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__29_LC_13_28_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__29_LC_13_28_6 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__29_LC_13_28_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__29_LC_13_28_6  (
            .in0(N__42832),
            .in1(N__33459),
            .in2(_gnd_net_),
            .in3(N__33592),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54310),
            .ce(N__41288),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__13_LC_13_28_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__13_LC_13_28_7 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__13_LC_13_28_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__13_LC_13_28_7  (
            .in0(N__33591),
            .in1(N__33458),
            .in2(_gnd_net_),
            .in3(N__42833),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54310),
            .ce(N__41288),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__9_LC_13_29_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__9_LC_13_29_0 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__9_LC_13_29_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__9_LC_13_29_0  (
            .in0(N__42761),
            .in1(N__35420),
            .in2(_gnd_net_),
            .in3(N__35312),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54319),
            .ce(N__41296),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__25_LC_13_29_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__25_LC_13_29_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__25_LC_13_29_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__25_LC_13_29_1  (
            .in0(N__35419),
            .in1(N__35311),
            .in2(_gnd_net_),
            .in3(N__42762),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54319),
            .ce(N__41296),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI4T0R_25_LC_13_29_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI4T0R_25_LC_13_29_2 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI4T0R_25_LC_13_29_2 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI4T0R_25_LC_13_29_2  (
            .in0(N__35236),
            .in1(_gnd_net_),
            .in2(N__33343),
            .in3(N__45676),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI4T0RZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI8H9K_25_LC_13_29_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI8H9K_25_LC_13_29_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI8H9K_25_LC_13_29_3 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI8H9K_25_LC_13_29_3  (
            .in0(N__33331),
            .in1(N__33319),
            .in2(N__45703),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI8H9KZ0Z_25_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIUOHM1_2_LC_13_29_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIUOHM1_2_LC_13_29_4 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIUOHM1_2_LC_13_29_4 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIUOHM1_2_LC_13_29_4  (
            .in0(N__50208),
            .in1(N__33313),
            .in2(N__33307),
            .in3(_gnd_net_),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIUOHM1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIOEUQ_10_LC_13_30_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIOEUQ_10_LC_13_30_0 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIOEUQ_10_LC_13_30_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIOEUQ_10_LC_13_30_0  (
            .in0(N__45673),
            .in1(N__33304),
            .in2(_gnd_net_),
            .in3(N__33289),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIOEUQZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIS27K_10_LC_13_30_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIS27K_10_LC_13_30_1 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIS27K_10_LC_13_30_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIS27K_10_LC_13_30_1  (
            .in0(N__33283),
            .in1(N__33274),
            .in2(_gnd_net_),
            .in3(N__45674),
            .lcout(),
            .ltout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNIS27KZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI6SCM1_2_LC_13_30_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI6SCM1_2_LC_13_30_2 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI6SCM1_2_LC_13_30_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI6SCM1_2_LC_13_30_2  (
            .in0(_gnd_net_),
            .in1(N__33916),
            .in2(N__33910),
            .in3(N__50170),
            .lcout(iQ_RNI6SCM1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI0NFT_10_LC_13_30_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI0NFT_10_LC_13_30_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI0NFT_10_LC_13_30_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI0NFT_10_LC_13_30_3  (
            .in0(N__33907),
            .in1(N__33895),
            .in2(_gnd_net_),
            .in3(N__45675),
            .lcout(),
            .ltout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI0NFTZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIRFA71_10_LC_13_30_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIRFA71_10_LC_13_30_4 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIRFA71_10_LC_13_30_4 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIRFA71_10_LC_13_30_4  (
            .in0(N__33871),
            .in1(_gnd_net_),
            .in2(N__33883),
            .in3(N__50169),
            .lcout(),
            .ltout(mem_mem_ram6__RNIRFA71_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.dat_o_i_i_a2_1_10_LC_13_30_5 .C_ON=1'b0;
    defparam \u0.dat_o_i_i_a2_1_10_LC_13_30_5 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_i_i_a2_1_10_LC_13_30_5 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \u0.dat_o_i_i_a2_1_10_LC_13_30_5  (
            .in0(N__33880),
            .in1(N__48969),
            .in2(N__33874),
            .in3(N__47253),
            .lcout(\u0.N_1989 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__10_LC_13_30_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__10_LC_13_30_6 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__10_LC_13_30_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__10_LC_13_30_6  (
            .in0(N__33830),
            .in1(N__33728),
            .in2(_gnd_net_),
            .in3(N__42907),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54325),
            .ce(N__41295),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__26_LC_13_30_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__26_LC_13_30_7 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__26_LC_13_30_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__26_LC_13_30_7  (
            .in0(N__42906),
            .in1(N__33831),
            .in2(_gnd_net_),
            .in3(N__33729),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54325),
            .ce(N__41295),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI6TFT_13_LC_13_31_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI6TFT_13_LC_13_31_0 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI6TFT_13_LC_13_31_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI6TFT_13_LC_13_31_0  (
            .in0(N__33646),
            .in1(N__33631),
            .in2(_gnd_net_),
            .in3(N__45695),
            .lcout(),
            .ltout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI6TFTZ0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI4PA71_13_LC_13_31_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI4PA71_13_LC_13_31_1 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI4PA71_13_LC_13_31_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI4PA71_13_LC_13_31_1  (
            .in0(N__50188),
            .in1(_gnd_net_),
            .in2(N__33619),
            .in3(N__33616),
            .lcout(),
            .ltout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI4PA71Z0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI9DV43_3_LC_13_31_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI9DV43_3_LC_13_31_2 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI9DV43_3_LC_13_31_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI9DV43_3_LC_13_31_2  (
            .in0(N__48971),
            .in1(_gnd_net_),
            .in2(N__33607),
            .in3(N__34081),
            .lcout(DMAq_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI297K_13_LC_13_31_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI297K_13_LC_13_31_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI297K_13_LC_13_31_3 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI297K_13_LC_13_31_3  (
            .in0(N__45694),
            .in1(N__34111),
            .in2(N__34099),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNI297KZ0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNII8DM1_2_LC_13_31_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNII8DM1_2_LC_13_31_4 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNII8DM1_2_LC_13_31_4 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNII8DM1_2_LC_13_31_4  (
            .in0(N__34036),
            .in1(_gnd_net_),
            .in2(N__34084),
            .in3(N__50189),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNII8DM1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.dat_o_0_0_1_13_LC_13_31_5 .C_ON=1'b0;
    defparam \u0.dat_o_0_0_1_13_LC_13_31_5 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_0_0_1_13_LC_13_31_5 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \u0.dat_o_0_0_1_13_LC_13_31_5  (
            .in0(N__34075),
            .in1(N__33991),
            .in2(N__47263),
            .in3(N__47467),
            .lcout(\u0.dat_o_0_0_1Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIUKUQ_13_LC_13_31_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIUKUQ_13_LC_13_31_6 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIUKUQ_13_LC_13_31_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIUKUQ_13_LC_13_31_6  (
            .in0(N__34057),
            .in1(N__34048),
            .in2(_gnd_net_),
            .in3(N__45693),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIUKUQZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.q_13_LC_13_31_7 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.q_13_LC_13_31_7 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.q_13_LC_13_31_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.PIO_control.PIO_access_control.q_13_LC_13_31_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34030),
            .lcout(PIOq_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54329),
            .ce(N__45932),
            .sr(_gnd_net_));
    defparam \u0.PIO_cmdport_T2_1_LC_14_15_0 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_T2_1_LC_14_15_0 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_cmdport_T2_1_LC_14_15_0 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \u0.PIO_cmdport_T2_1_LC_14_15_0  (
            .in0(N__51458),
            .in1(N__35952),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(PIO_cmdport_T2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54222),
            .ce(N__49692),
            .sr(N__53357));
    defparam \u0.PIO_cmdport_T2_0_LC_14_16_3 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_T2_0_LC_14_16_3 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_cmdport_T2_0_LC_14_16_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.PIO_cmdport_T2_0_LC_14_16_3  (
            .in0(N__54459),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51264),
            .lcout(PIO_cmdport_T2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54209),
            .ce(N__49693),
            .sr(N__53350));
    defparam \u0.PIO_dport1_T2_0_LC_14_17_1 .C_ON=1'b0;
    defparam \u0.PIO_dport1_T2_0_LC_14_17_1 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport1_T2_0_LC_14_17_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.PIO_dport1_T2_0_LC_14_17_1  (
            .in0(N__51500),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54461),
            .lcout(PIO_dport1_T2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54193),
            .ce(N__39188),
            .sr(N__53358));
    defparam \u0.PIO_dport1_T1_1_LC_14_18_0 .C_ON=1'b0;
    defparam \u0.PIO_dport1_T1_1_LC_14_18_0 .SEQ_MODE=4'b1011;
    defparam \u0.PIO_dport1_T1_1_LC_14_18_0 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \u0.PIO_dport1_T1_1_LC_14_18_0  (
            .in0(N__39352),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51265),
            .lcout(PIO_dport1_T1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54210),
            .ce(N__39205),
            .sr(N__53366));
    defparam \u0.PIO_dport1_T1_2_LC_14_18_1 .C_ON=1'b0;
    defparam \u0.PIO_dport1_T1_2_LC_14_18_1 .SEQ_MODE=4'b1011;
    defparam \u0.PIO_dport1_T1_2_LC_14_18_1 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \u0.PIO_dport1_T1_2_LC_14_18_1  (
            .in0(N__51266),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34237),
            .lcout(PIO_dport1_T1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54210),
            .ce(N__39205),
            .sr(N__53366));
    defparam \u0.PIO_dport1_T2_2_LC_14_18_2 .C_ON=1'b0;
    defparam \u0.PIO_dport1_T2_2_LC_14_18_2 .SEQ_MODE=4'b1011;
    defparam \u0.PIO_dport1_T2_2_LC_14_18_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \u0.PIO_dport1_T2_2_LC_14_18_2  (
            .in0(N__40186),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51267),
            .lcout(PIO_dport1_T2_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54210),
            .ce(N__39205),
            .sr(N__53366));
    defparam \u0.PIO_dport1_T2_3_LC_14_18_3 .C_ON=1'b0;
    defparam \u0.PIO_dport1_T2_3_LC_14_18_3 .SEQ_MODE=4'b1011;
    defparam \u0.PIO_dport1_T2_3_LC_14_18_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \u0.PIO_dport1_T2_3_LC_14_18_3  (
            .in0(N__43702),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51271),
            .lcout(PIO_dport1_T2_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54210),
            .ce(N__39205),
            .sr(N__53366));
    defparam \u0.PIO_dport1_T4_1_LC_14_18_4 .C_ON=1'b0;
    defparam \u0.PIO_dport1_T4_1_LC_14_18_4 .SEQ_MODE=4'b1011;
    defparam \u0.PIO_dport1_T4_1_LC_14_18_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \u0.PIO_dport1_T4_1_LC_14_18_4  (
            .in0(N__45145),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51268),
            .lcout(PIO_dport1_T4_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54210),
            .ce(N__39205),
            .sr(N__53366));
    defparam \u0.PIO_dport1_Teoc_0_LC_14_18_5 .C_ON=1'b0;
    defparam \u0.PIO_dport1_Teoc_0_LC_14_18_5 .SEQ_MODE=4'b1011;
    defparam \u0.PIO_dport1_Teoc_0_LC_14_18_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \u0.PIO_dport1_Teoc_0_LC_14_18_5  (
            .in0(N__39922),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51272),
            .lcout(PIO_dport1_Teoc_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54210),
            .ce(N__39205),
            .sr(N__53366));
    defparam \u0.PIO_dport1_Teoc_1_LC_14_18_6 .C_ON=1'b0;
    defparam \u0.PIO_dport1_Teoc_1_LC_14_18_6 .SEQ_MODE=4'b1011;
    defparam \u0.PIO_dport1_Teoc_1_LC_14_18_6 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \u0.PIO_dport1_Teoc_1_LC_14_18_6  (
            .in0(N__40873),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51269),
            .lcout(PIO_dport1_Teoc_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54210),
            .ce(N__39205),
            .sr(N__53366));
    defparam \u0.PIO_dport1_T1_3_LC_14_18_7 .C_ON=1'b0;
    defparam \u0.PIO_dport1_T1_3_LC_14_18_7 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport1_T1_3_LC_14_18_7 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.PIO_dport1_T1_3_LC_14_18_7  (
            .in0(N__37341),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51270),
            .lcout(PIO_dport1_T1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54210),
            .ce(N__39205),
            .sr(N__53366));
    defparam \u0.PIO_dport0_Teoc_1_LC_14_19_0 .C_ON=1'b0;
    defparam \u0.PIO_dport0_Teoc_1_LC_14_19_0 .SEQ_MODE=4'b1011;
    defparam \u0.PIO_dport0_Teoc_1_LC_14_19_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \u0.PIO_dport0_Teoc_1_LC_14_19_0  (
            .in0(_gnd_net_),
            .in1(N__40872),
            .in2(_gnd_net_),
            .in3(N__51278),
            .lcout(PIO_dport0_Teoc_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54223),
            .ce(N__49381),
            .sr(N__53373));
    defparam \u0.PIO_dport0_Teoc_2_LC_14_19_1 .C_ON=1'b0;
    defparam \u0.PIO_dport0_Teoc_2_LC_14_19_1 .SEQ_MODE=4'b1011;
    defparam \u0.PIO_dport0_Teoc_2_LC_14_19_1 .LUT_INIT=16'b1110111011101110;
    LogicCell40 \u0.PIO_dport0_Teoc_2_LC_14_19_1  (
            .in0(N__44238),
            .in1(N__51717),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(PIO_dport0_Teoc_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54223),
            .ce(N__49381),
            .sr(N__53373));
    defparam \u0.PIO_dport0_Teoc_4_LC_14_19_2 .C_ON=1'b0;
    defparam \u0.PIO_dport0_Teoc_4_LC_14_19_2 .SEQ_MODE=4'b1011;
    defparam \u0.PIO_dport0_Teoc_4_LC_14_19_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \u0.PIO_dport0_Teoc_4_LC_14_19_2  (
            .in0(N__46124),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51279),
            .lcout(PIO_dport0_Teoc_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54223),
            .ce(N__49381),
            .sr(N__53373));
    defparam \u0.PIO_dport0_T2_5_LC_14_19_3 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T2_5_LC_14_19_3 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport0_T2_5_LC_14_19_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.PIO_dport0_T2_5_LC_14_19_3  (
            .in0(N__51273),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34646),
            .lcout(PIO_dport0_T2_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54223),
            .ce(N__49381),
            .sr(N__53373));
    defparam \u0.PIO_dport0_T2_6_LC_14_19_4 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T2_6_LC_14_19_4 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport0_T2_6_LC_14_19_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \u0.PIO_dport0_T2_6_LC_14_19_4  (
            .in0(_gnd_net_),
            .in1(N__44059),
            .in2(_gnd_net_),
            .in3(N__51274),
            .lcout(PIO_dport0_T2_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54223),
            .ce(N__49381),
            .sr(N__53373));
    defparam \u0.PIO_dport0_T2_7_LC_14_19_5 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T2_7_LC_14_19_5 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport0_T2_7_LC_14_19_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.PIO_dport0_T2_7_LC_14_19_5  (
            .in0(N__51275),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34522),
            .lcout(PIO_dport0_T2_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54223),
            .ce(N__49381),
            .sr(N__53373));
    defparam \u0.PIO_dport0_T4_0_LC_14_19_6 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T4_0_LC_14_19_6 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport0_T4_0_LC_14_19_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.PIO_dport0_T4_0_LC_14_19_6  (
            .in0(N__41000),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51276),
            .lcout(PIO_dport0_T4_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54223),
            .ce(N__49381),
            .sr(N__53373));
    defparam \u0.PIO_dport0_T4_5_LC_14_19_7 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T4_5_LC_14_19_7 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport0_T4_5_LC_14_19_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.PIO_dport0_T4_5_LC_14_19_7  (
            .in0(N__51277),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38077),
            .lcout(PIO_dport0_T4_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54223),
            .ce(N__49381),
            .sr(N__53373));
    defparam \u0.PIO_dport0_T4_RNIBRI22_3_LC_14_20_0 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T4_RNIBRI22_3_LC_14_20_0 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport0_T4_RNIBRI22_3_LC_14_20_0 .LUT_INIT=16'b0100010011110100;
    LogicCell40 \u0.PIO_dport0_T4_RNIBRI22_3_LC_14_20_0  (
            .in0(N__34440),
            .in1(N__52912),
            .in2(N__50293),
            .in3(N__34290),
            .lcout(\u0.dat_o_i_0_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport0_T1_RNIJ5HR3_4_LC_14_20_4 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T1_RNIJ5HR3_4_LC_14_20_4 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport0_T1_RNIJ5HR3_4_LC_14_20_4 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \u0.PIO_dport0_T1_RNIJ5HR3_4_LC_14_20_4  (
            .in0(N__36063),
            .in1(N__54675),
            .in2(N__37854),
            .in3(N__50725),
            .lcout(\u0.dat_o_0_0_3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport0_T2_RNIF0OR1_7_LC_14_20_7 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T2_RNIF0OR1_7_LC_14_20_7 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport0_T2_RNIF0OR1_7_LC_14_20_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \u0.PIO_dport0_T2_RNIF0OR1_7_LC_14_20_7  (
            .in0(N__46741),
            .in1(N__53006),
            .in2(N__47736),
            .in3(N__34398),
            .lcout(\u0.N_2033 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport0_T4_3_LC_14_21_0 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T4_3_LC_14_21_0 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport0_T4_3_LC_14_21_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.PIO_dport0_T4_3_LC_14_21_0  (
            .in0(N__34368),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51299),
            .lcout(PIO_dport0_T4_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54246),
            .ce(N__49382),
            .sr(N__53385));
    defparam \u0.PIO_dport0_T4_4_LC_14_21_1 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T4_4_LC_14_21_1 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport0_T4_4_LC_14_21_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.PIO_dport0_T4_4_LC_14_21_1  (
            .in0(N__51300),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34787),
            .lcout(PIO_dport0_T4_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54246),
            .ce(N__49382),
            .sr(N__53385));
    defparam \u0.PIO_dport0_T4_2_LC_14_21_2 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T4_2_LC_14_21_2 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport0_T4_2_LC_14_21_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \u0.PIO_dport0_T4_2_LC_14_21_2  (
            .in0(_gnd_net_),
            .in1(N__35043),
            .in2(_gnd_net_),
            .in3(N__51298),
            .lcout(PIO_dport0_T4_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54246),
            .ce(N__49382),
            .sr(N__53385));
    defparam \u0.PIO_dport0_T4_6_LC_14_21_3 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T4_6_LC_14_21_3 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport0_T4_6_LC_14_21_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.PIO_dport0_T4_6_LC_14_21_3  (
            .in0(N__51301),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38184),
            .lcout(PIO_dport0_T4_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54246),
            .ce(N__49382),
            .sr(N__53385));
    defparam \u0.PIO_dport0_T4_7_LC_14_21_4 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T4_7_LC_14_21_4 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport0_T4_7_LC_14_21_4 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.PIO_dport0_T4_7_LC_14_21_4  (
            .in0(N__44838),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51302),
            .lcout(PIO_dport0_T4_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54246),
            .ce(N__49382),
            .sr(N__53385));
    defparam \u0.PIO_dport0_Teoc_3_LC_14_21_5 .C_ON=1'b0;
    defparam \u0.PIO_dport0_Teoc_3_LC_14_21_5 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport0_Teoc_3_LC_14_21_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.PIO_dport0_Teoc_3_LC_14_21_5  (
            .in0(N__37715),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51304),
            .lcout(PIO_dport0_Teoc_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54246),
            .ce(N__49382),
            .sr(N__53385));
    defparam \u0.PIO_dport0_Teoc_5_LC_14_21_6 .C_ON=1'b0;
    defparam \u0.PIO_dport0_Teoc_5_LC_14_21_6 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport0_Teoc_5_LC_14_21_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \u0.PIO_dport0_Teoc_5_LC_14_21_6  (
            .in0(_gnd_net_),
            .in1(N__49335),
            .in2(_gnd_net_),
            .in3(N__51303),
            .lcout(PIO_dport0_Teoc_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54246),
            .ce(N__49382),
            .sr(N__53385));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIE0OK1_2_LC_14_22_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIE0OK1_2_LC_14_22_0 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIE0OK1_2_LC_14_22_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIE0OK1_2_LC_14_22_0  (
            .in0(N__34744),
            .in1(N__34732),
            .in2(_gnd_net_),
            .in3(N__49918),
            .lcout(),
            .ltout(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIE0OK1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIISN93_3_LC_14_22_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIISN93_3_LC_14_22_1 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIISN93_3_LC_14_22_1 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIISN93_3_LC_14_22_1  (
            .in0(_gnd_net_),
            .in1(N__34840),
            .in2(N__34714),
            .in3(N__48833),
            .lcout(),
            .ltout(DMAq_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.dat_o_0_0_1_3_LC_14_22_2 .C_ON=1'b0;
    defparam \u0.dat_o_0_0_1_3_LC_14_22_2 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_0_0_1_3_LC_14_22_2 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \u0.dat_o_0_0_1_3_LC_14_22_2  (
            .in0(N__34876),
            .in1(N__47167),
            .in2(N__34711),
            .in3(N__47398),
            .lcout(\u0.dat_o_0_0_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev0_Tm_RNIH3HR3_3_LC_14_22_3 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Tm_RNIH3HR3_3_LC_14_22_3 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev0_Tm_RNIH3HR3_3_LC_14_22_3 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \u0.DMA_dev0_Tm_RNIH3HR3_3_LC_14_22_3  (
            .in0(N__46939),
            .in1(N__34834),
            .in2(N__48597),
            .in3(N__34971),
            .lcout(),
            .ltout(\u0.dat_o_0_0_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_cmdport_T1_RNIMOUSG_3_LC_14_22_4 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_T1_RNIMOUSG_3_LC_14_22_4 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_cmdport_T1_RNIMOUSG_3_LC_14_22_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \u0.PIO_cmdport_T1_RNIMOUSG_3_LC_14_22_4  (
            .in0(N__34951),
            .in1(N__34939),
            .in2(N__34933),
            .in3(N__34930),
            .lcout(wb_dat_o_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.q_3_LC_14_22_5 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.q_3_LC_14_22_5 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.q_3_LC_14_22_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \u1.PIO_control.PIO_access_control.q_3_LC_14_22_5  (
            .in0(N__34910),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(PIOq_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54260),
            .ce(N__45903),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIHGOD1_3_LC_14_22_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIHGOD1_3_LC_14_22_6 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIHGOD1_3_LC_14_22_6 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIHGOD1_3_LC_14_22_6  (
            .in0(N__34870),
            .in1(_gnd_net_),
            .in2(N__34858),
            .in3(N__49917),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIHGOD1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev0_Teoc_4_LC_14_23_0 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Teoc_4_LC_14_23_0 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev0_Teoc_4_LC_14_23_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \u0.DMA_dev0_Teoc_4_LC_14_23_0  (
            .in0(_gnd_net_),
            .in1(N__46131),
            .in2(_gnd_net_),
            .in3(N__51306),
            .lcout(DMA_dev0_Teoc_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54272),
            .ce(N__39741),
            .sr(N__53395));
    defparam \u0.DMA_dev0_Teoc_5_LC_14_23_1 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Teoc_5_LC_14_23_1 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev0_Teoc_5_LC_14_23_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.DMA_dev0_Teoc_5_LC_14_23_1  (
            .in0(N__51307),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49344),
            .lcout(DMA_dev0_Teoc_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54272),
            .ce(N__39741),
            .sr(N__53395));
    defparam \u0.DMA_dev0_Tm_3_LC_14_23_2 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Tm_3_LC_14_23_2 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev0_Tm_3_LC_14_23_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.DMA_dev0_Tm_3_LC_14_23_2  (
            .in0(N__37364),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51308),
            .lcout(DMA_dev0_Tm_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54272),
            .ce(N__39741),
            .sr(N__53395));
    defparam \u0.DMA_dev0_Teoc_3_LC_14_23_3 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Teoc_3_LC_14_23_3 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev0_Teoc_3_LC_14_23_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.DMA_dev0_Teoc_3_LC_14_23_3  (
            .in0(N__51305),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37714),
            .lcout(DMA_dev0_Teoc_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54272),
            .ce(N__39741),
            .sr(N__53395));
    defparam \u0.DMA_dev0_Tm_4_LC_14_23_5 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Tm_4_LC_14_23_5 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev0_Tm_4_LC_14_23_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.DMA_dev0_Tm_4_LC_14_23_5  (
            .in0(N__51309),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37241),
            .lcout(DMA_dev0_Tm_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54272),
            .ce(N__39741),
            .sr(N__53395));
    defparam \u0.DMA_dev0_Tm_5_LC_14_23_6 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Tm_5_LC_14_23_6 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev0_Tm_5_LC_14_23_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.DMA_dev0_Tm_5_LC_14_23_6  (
            .in0(N__46290),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51310),
            .lcout(DMA_dev0_Tm_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54272),
            .ce(N__39741),
            .sr(N__53395));
    defparam \u0.DMA_dev0_Tm_6_LC_14_23_7 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Tm_6_LC_14_23_7 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev0_Tm_6_LC_14_23_7 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \u0.DMA_dev0_Tm_6_LC_14_23_7  (
            .in0(N__39475),
            .in1(N__51942),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(DMA_dev0_Tm_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54272),
            .ce(N__39741),
            .sr(N__53395));
    defparam \u0.CtrlReg_RNI7BKU1_18_LC_14_24_0 .C_ON=1'b0;
    defparam \u0.CtrlReg_RNI7BKU1_18_LC_14_24_0 .SEQ_MODE=4'b0000;
    defparam \u0.CtrlReg_RNI7BKU1_18_LC_14_24_0 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \u0.CtrlReg_RNI7BKU1_18_LC_14_24_0  (
            .in0(N__44928),
            .in1(N__45029),
            .in2(N__35146),
            .in3(N__34981),
            .lcout(\u0.dat_o_i_0_2_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIJ8B71_18_LC_14_24_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIJ8B71_18_LC_14_24_2 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIJ8B71_18_LC_14_24_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIJ8B71_18_LC_14_24_2  (
            .in0(N__50019),
            .in1(N__35119),
            .in2(_gnd_net_),
            .in3(N__35104),
            .lcout(),
            .ltout(mem_mem_ram6__RNIJ8B71_18_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.dat_o_i_0_a2_18_LC_14_24_3 .C_ON=1'b0;
    defparam \u0.dat_o_i_0_a2_18_LC_14_24_3 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_i_0_a2_18_LC_14_24_3 .LUT_INIT=16'b0001101100000000;
    LogicCell40 \u0.dat_o_i_0_a2_18_LC_14_24_3  (
            .in0(N__48889),
            .in1(N__35050),
            .in2(N__35092),
            .in3(N__50465),
            .lcout(\u0.N_1729 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI8VUQ_18_LC_14_24_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI8VUQ_18_LC_14_24_4 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI8VUQ_18_LC_14_24_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI8VUQ_18_LC_14_24_4  (
            .in0(N__35089),
            .in1(N__35077),
            .in2(_gnd_net_),
            .in3(N__45551),
            .lcout(),
            .ltout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI8VUQZ0Z_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI6TDM1_2_LC_14_24_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI6TDM1_2_LC_14_24_5 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI6TDM1_2_LC_14_24_5 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI6TDM1_2_LC_14_24_5  (
            .in0(N__35065),
            .in1(_gnd_net_),
            .in2(N__35053),
            .in3(N__50020),
            .lcout(iQ_RNI6TDM1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.CtrlReg_18_LC_14_24_6 .C_ON=1'b0;
    defparam \u0.CtrlReg_18_LC_14_24_6 .SEQ_MODE=4'b1010;
    defparam \u0.CtrlReg_18_LC_14_24_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.CtrlReg_18_LC_14_24_6  (
            .in0(N__35044),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51311),
            .lcout(\u0.CtrlRegZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54282),
            .ce(N__53530),
            .sr(N__53400));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__7_LC_14_25_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__7_LC_14_25_0 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__7_LC_14_25_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__7_LC_14_25_0  (
            .in0(N__43032),
            .in1(N__38803),
            .in2(_gnd_net_),
            .in3(N__38691),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54292),
            .ce(N__41297),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__23_LC_14_25_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__23_LC_14_25_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__23_LC_14_25_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__23_LC_14_25_1  (
            .in0(N__38802),
            .in1(N__38690),
            .in2(_gnd_net_),
            .in3(N__43034),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54292),
            .ce(N__41297),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__8_LC_14_25_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__8_LC_14_25_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__8_LC_14_25_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__8_LC_14_25_2  (
            .in0(N__43033),
            .in1(N__38460),
            .in2(_gnd_net_),
            .in3(N__38584),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54292),
            .ce(N__41297),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__24_LC_14_25_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__24_LC_14_25_3 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__24_LC_14_25_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__24_LC_14_25_3  (
            .in0(N__38583),
            .in1(N__38459),
            .in2(_gnd_net_),
            .in3(N__43035),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54292),
            .ce(N__41297),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIQKHM1_2_LC_14_25_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIQKHM1_2_LC_14_25_4 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIQKHM1_2_LC_14_25_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIQKHM1_2_LC_14_25_4  (
            .in0(N__35221),
            .in1(N__35206),
            .in2(_gnd_net_),
            .in3(N__50015),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIQKHM1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIA3IT_24_LC_14_25_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIA3IT_24_LC_14_25_5 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIA3IT_24_LC_14_25_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIA3IT_24_LC_14_25_5  (
            .in0(N__38419),
            .in1(N__35191),
            .in2(_gnd_net_),
            .in3(N__45552),
            .lcout(),
            .ltout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIA3ITZ0Z_24_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIA2E71_24_LC_14_25_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIA2E71_24_LC_14_25_6 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIA2E71_24_LC_14_25_6 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIA2E71_24_LC_14_25_6  (
            .in0(_gnd_net_),
            .in1(N__50014),
            .in2(N__35179),
            .in3(N__35176),
            .lcout(),
            .ltout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIA2E71Z0Z_24_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIN2753_3_LC_14_25_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIN2753_3_LC_14_25_7 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIN2753_3_LC_14_25_7 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIN2753_3_LC_14_25_7  (
            .in0(N__35170),
            .in1(_gnd_net_),
            .in2(N__35164),
            .in3(N__48891),
            .lcout(DMAq_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_0_LC_14_26_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_0_LC_14_26_0 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_0_LC_14_26_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_readDlw_0_LC_14_26_0  (
            .in0(N__44480),
            .in1(N__43379),
            .in2(_gnd_net_),
            .in3(N__43036),
            .lcout(\u1.DMA_control.readDlw_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54303),
            .ce(N__36322),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_0_LC_14_26_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_0_LC_14_26_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_0_LC_14_26_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_readDfw_0_LC_14_26_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41701),
            .lcout(\u1.DMA_control.readDfw_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54303),
            .ce(N__36322),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_8_LC_14_26_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_8_LC_14_26_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_8_LC_14_26_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_readDlw_8_LC_14_26_2  (
            .in0(N__44481),
            .in1(N__43380),
            .in2(_gnd_net_),
            .in3(N__43038),
            .lcout(\u1.DMA_control.readDlw_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54303),
            .ce(N__36322),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_8_LC_14_26_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_8_LC_14_26_3 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_8_LC_14_26_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_readDfw_8_LC_14_26_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38483),
            .lcout(\u1.DMA_control.readDfw_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54303),
            .ce(N__36322),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_1_LC_14_26_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_1_LC_14_26_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_1_LC_14_26_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_readDlw_1_LC_14_26_4  (
            .in0(N__44570),
            .in1(N__45974),
            .in2(_gnd_net_),
            .in3(N__43037),
            .lcout(\u1.DMA_control.readDlw_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54303),
            .ce(N__36322),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_5_LC_14_26_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_5_LC_14_26_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_5_LC_14_26_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_readDfw_5_LC_14_26_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35674),
            .lcout(\u1.DMA_control.readDfw_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54303),
            .ce(N__36322),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_9_LC_14_26_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_9_LC_14_26_6 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_readDlw_9_LC_14_26_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_readDlw_9_LC_14_26_6  (
            .in0(N__44571),
            .in1(N__45975),
            .in2(_gnd_net_),
            .in3(N__43039),
            .lcout(\u1.DMA_control.readDlw_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54303),
            .ce(N__36322),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_1_LC_14_26_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_1_LC_14_26_7 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_1_LC_14_26_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_readDfw_1_LC_14_26_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41485),
            .lcout(\u1.DMA_control.readDfw_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54303),
            .ce(N__36322),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI8FCM_9_LC_14_27_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI8FCM_9_LC_14_27_0 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI8FCM_9_LC_14_27_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI8FCM_9_LC_14_27_0  (
            .in0(N__35461),
            .in1(N__35449),
            .in2(_gnd_net_),
            .in3(N__45636),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI8FCMZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__9_LC_14_27_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__9_LC_14_27_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__9_LC_14_27_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__9_LC_14_27_1  (
            .in0(N__42935),
            .in1(N__35374),
            .in2(_gnd_net_),
            .in3(N__35297),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54311),
            .ce(N__35899),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__25_LC_14_27_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__25_LC_14_27_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__25_LC_14_27_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__25_LC_14_27_2  (
            .in0(N__35373),
            .in1(N__35296),
            .in2(_gnd_net_),
            .in3(N__42937),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54311),
            .ce(N__35899),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIMSBM_0_LC_14_27_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIMSBM_0_LC_14_27_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIMSBM_0_LC_14_27_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIMSBM_0_LC_14_27_3  (
            .in0(N__35227),
            .in1(N__45663),
            .in2(_gnd_net_),
            .in3(N__35740),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIMSBMZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__0_LC_14_27_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__0_LC_14_27_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__0_LC_14_27_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__0_LC_14_27_4  (
            .in0(N__41681),
            .in1(N__41581),
            .in2(_gnd_net_),
            .in3(N__42936),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54311),
            .ce(N__35899),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__16_LC_14_27_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__16_LC_14_27_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__16_LC_14_27_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__16_LC_14_27_5  (
            .in0(N__42933),
            .in1(N__41682),
            .in2(_gnd_net_),
            .in3(N__41582),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54311),
            .ce(N__35899),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIOUBM_1_LC_14_27_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIOUBM_1_LC_14_27_6 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIOUBM_1_LC_14_27_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIOUBM_1_LC_14_27_6  (
            .in0(N__35734),
            .in1(N__35725),
            .in2(_gnd_net_),
            .in3(N__45637),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIOUBMZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__1_LC_14_27_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__1_LC_14_27_7 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__1_LC_14_27_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__1_LC_14_27_7  (
            .in0(N__42934),
            .in1(N__41484),
            .in2(_gnd_net_),
            .in3(N__41350),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54311),
            .ce(N__35899),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI811R_27_LC_14_28_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI811R_27_LC_14_28_0 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI811R_27_LC_14_28_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI811R_27_LC_14_28_0  (
            .in0(N__45667),
            .in1(N__35680),
            .in2(_gnd_net_),
            .in3(N__35719),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI811RZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNICL9K_27_LC_14_28_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNICL9K_27_LC_14_28_1 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNICL9K_27_LC_14_28_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNICL9K_27_LC_14_28_1  (
            .in0(N__35713),
            .in1(N__35704),
            .in2(_gnd_net_),
            .in3(N__45669),
            .lcout(),
            .ltout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram3__RNICL9KZ0Z_27_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI61IM1_2_LC_14_28_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI61IM1_2_LC_14_28_2 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI61IM1_2_LC_14_28_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI61IM1_2_LC_14_28_2  (
            .in0(_gnd_net_),
            .in1(N__35692),
            .in2(N__35686),
            .in3(N__50165),
            .lcout(),
            .ltout(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI61IM1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNICO753_3_LC_14_28_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNICO753_3_LC_14_28_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNICO753_3_LC_14_28_3 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNICO753_3_LC_14_28_3  (
            .in0(N__41185),
            .in1(_gnd_net_),
            .in2(N__35683),
            .in3(N__48937),
            .lcout(DMAq_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__27_LC_14_28_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__27_LC_14_28_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__27_LC_14_28_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__27_LC_14_28_4  (
            .in0(N__42816),
            .in1(N__43097),
            .in2(_gnd_net_),
            .in3(N__43203),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54320),
            .ce(N__35900),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__11_LC_14_28_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__11_LC_14_28_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__11_LC_14_28_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__11_LC_14_28_5  (
            .in0(N__43202),
            .in1(N__43096),
            .in2(_gnd_net_),
            .in3(N__42817),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54320),
            .ce(N__35900),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIQGUQ_11_LC_14_28_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIQGUQ_11_LC_14_28_6 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIQGUQ_11_LC_14_28_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIQGUQ_11_LC_14_28_6  (
            .in0(N__45668),
            .in1(N__35815),
            .in2(_gnd_net_),
            .in3(N__35803),
            .lcout(),
            .ltout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIQGUQZ0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIA0DM1_2_LC_14_28_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIA0DM1_2_LC_14_28_7 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIA0DM1_2_LC_14_28_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIA0DM1_2_LC_14_28_7  (
            .in0(N__50166),
            .in1(_gnd_net_),
            .in2(N__35797),
            .in3(N__35794),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIA0DM1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__0_LC_14_29_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__0_LC_14_29_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__0_LC_14_29_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__0_LC_14_29_1  (
            .in0(N__41702),
            .in1(N__41602),
            .in2(_gnd_net_),
            .in3(N__42986),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54326),
            .ce(N__41860),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__16_LC_14_29_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__16_LC_14_29_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__16_LC_14_29_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__16_LC_14_29_2  (
            .in0(N__42985),
            .in1(_gnd_net_),
            .in2(N__41625),
            .in3(N__41703),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54326),
            .ce(N__41860),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIC3GT_16_LC_14_29_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIC3GT_16_LC_14_29_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIC3GT_16_LC_14_29_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIC3GT_16_LC_14_29_3  (
            .in0(N__35782),
            .in1(N__35770),
            .in2(_gnd_net_),
            .in3(N__45681),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIC3GTZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI2PFT_11_LC_14_29_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI2PFT_11_LC_14_29_4 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI2PFT_11_LC_14_29_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI2PFT_11_LC_14_29_4  (
            .in0(N__45680),
            .in1(N__35764),
            .in2(_gnd_net_),
            .in3(N__35755),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI2PFTZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__11_LC_14_29_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__11_LC_14_29_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__11_LC_14_29_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__11_LC_14_29_5  (
            .in0(N__43204),
            .in1(N__43108),
            .in2(_gnd_net_),
            .in3(N__42987),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54326),
            .ce(N__41860),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIG9IT_27_LC_14_29_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIG9IT_27_LC_14_29_7 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIG9IT_27_LC_14_29_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIG9IT_27_LC_14_29_7  (
            .in0(N__41869),
            .in1(N__35749),
            .in2(_gnd_net_),
            .in3(N__45682),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIG9ITZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_3_LC_14_30_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_3_LC_14_30_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMA_sigs_readDfw_3_LC_14_30_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.DMA_control.gen_DMA_sigs_readDfw_3_LC_14_30_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36534),
            .lcout(\u1.DMA_control.readDfw_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54330),
            .ce(N__36321),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport0_T1_7_LC_15_14_1 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T1_7_LC_15_14_1 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport0_T1_7_LC_15_14_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.PIO_dport0_T1_7_LC_15_14_1  (
            .in0(N__51457),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39614),
            .lcout(PIO_dport0_T1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54247),
            .ce(N__49379),
            .sr(N__53374));
    defparam \u1.DMA_control.DMA_timing_ctrl_Tm_7_LC_15_15_5 .C_ON=1'b0;
    defparam \u1.DMA_control.DMA_timing_ctrl_Tm_7_LC_15_15_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.DMA_timing_ctrl_Tm_7_LC_15_15_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.DMA_timing_ctrl_Tm_7_LC_15_15_5  (
            .in0(N__39552),
            .in1(N__39753),
            .in2(_gnd_net_),
            .in3(N__36295),
            .lcout(\u1.DMA_control.Tm_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54234),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport1_T1_RNIQH004_7_LC_15_15_6 .C_ON=1'b0;
    defparam \u0.PIO_dport1_T1_RNIQH004_7_LC_15_15_6 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport1_T1_RNIQH004_7_LC_15_15_6 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \u0.PIO_dport1_T1_RNIQH004_7_LC_15_15_6  (
            .in0(N__54717),
            .in1(N__46936),
            .in2(N__36091),
            .in3(N__39553),
            .lcout(\u0.dat_o_0_0_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport0_Teoc_6_LC_15_17_0 .C_ON=1'b0;
    defparam \u0.PIO_dport0_Teoc_6_LC_15_17_0 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport0_Teoc_6_LC_15_17_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \u0.PIO_dport0_Teoc_6_LC_15_17_0  (
            .in0(_gnd_net_),
            .in1(N__51808),
            .in2(_gnd_net_),
            .in3(N__47839),
            .lcout(PIO_dport0_Teoc_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54203),
            .ce(N__49378),
            .sr(N__53367));
    defparam \u0.PIO_dport0_Teoc_7_LC_15_17_1 .C_ON=1'b0;
    defparam \u0.PIO_dport0_Teoc_7_LC_15_17_1 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport0_Teoc_7_LC_15_17_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.PIO_dport0_Teoc_7_LC_15_17_1  (
            .in0(N__51809),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40531),
            .lcout(PIO_dport0_Teoc_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54203),
            .ce(N__49378),
            .sr(N__53367));
    defparam \u0.PIO_dport0_T1_4_LC_15_17_2 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T1_4_LC_15_17_2 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport0_T1_4_LC_15_17_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.PIO_dport0_T1_4_LC_15_17_2  (
            .in0(N__37221),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51806),
            .lcout(PIO_dport0_T1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54203),
            .ce(N__49378),
            .sr(N__53367));
    defparam \u0.PIO_dport0_T2_0_LC_15_17_6 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T2_0_LC_15_17_6 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport0_T2_0_LC_15_17_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.PIO_dport0_T2_0_LC_15_17_6  (
            .in0(N__54460),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51807),
            .lcout(PIO_dport0_T2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54203),
            .ce(N__49378),
            .sr(N__53367));
    defparam \u0.PIO_dport0_T2_1_LC_15_17_7 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T2_1_LC_15_17_7 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport0_T2_1_LC_15_17_7 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.PIO_dport0_T2_1_LC_15_17_7  (
            .in0(N__35953),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51459),
            .lcout(PIO_dport0_T2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54203),
            .ce(N__49378),
            .sr(N__53367));
    defparam \u0.PIO_cmdport_T2_2_LC_15_18_3 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_T2_2_LC_15_18_3 .SEQ_MODE=4'b1011;
    defparam \u0.PIO_cmdport_T2_2_LC_15_18_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \u0.PIO_cmdport_T2_2_LC_15_18_3  (
            .in0(_gnd_net_),
            .in1(N__40166),
            .in2(_gnd_net_),
            .in3(N__51712),
            .lcout(PIO_cmdport_T2_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54224),
            .ce(N__49695),
            .sr(N__53375));
    defparam \u0.PIO_cmdport_T2_3_LC_15_18_4 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_T2_3_LC_15_18_4 .SEQ_MODE=4'b1011;
    defparam \u0.PIO_cmdport_T2_3_LC_15_18_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \u0.PIO_cmdport_T2_3_LC_15_18_4  (
            .in0(N__51713),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43699),
            .lcout(PIO_cmdport_T2_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54224),
            .ce(N__49695),
            .sr(N__53375));
    defparam \u0.PIO_cmdport_T2_4_LC_15_18_5 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_T2_4_LC_15_18_5 .SEQ_MODE=4'b1011;
    defparam \u0.PIO_cmdport_T2_4_LC_15_18_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \u0.PIO_cmdport_T2_4_LC_15_18_5  (
            .in0(N__36991),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51714),
            .lcout(PIO_cmdport_T2_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54224),
            .ce(N__49695),
            .sr(N__53375));
    defparam \u0.PIO_cmdport_T4_1_LC_15_18_6 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_T4_1_LC_15_18_6 .SEQ_MODE=4'b1011;
    defparam \u0.PIO_cmdport_T4_1_LC_15_18_6 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \u0.PIO_cmdport_T4_1_LC_15_18_6  (
            .in0(N__51715),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45141),
            .lcout(PIO_cmdport_T4_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54224),
            .ce(N__49695),
            .sr(N__53375));
    defparam \u0.PIO_cmdport_Teoc_0_LC_15_18_7 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_Teoc_0_LC_15_18_7 .SEQ_MODE=4'b1011;
    defparam \u0.PIO_cmdport_Teoc_0_LC_15_18_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \u0.PIO_cmdport_Teoc_0_LC_15_18_7  (
            .in0(N__39920),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51716),
            .lcout(PIO_cmdport_Teoc_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54224),
            .ce(N__49695),
            .sr(N__53375));
    defparam \u0.DMA_dev1_Teoc_RNI3P9J3_4_LC_15_19_0 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Teoc_RNI3P9J3_4_LC_15_19_0 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev1_Teoc_RNI3P9J3_4_LC_15_19_0 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \u0.DMA_dev1_Teoc_RNI3P9J3_4_LC_15_19_0  (
            .in0(N__48112),
            .in1(N__36856),
            .in2(N__54716),
            .in3(N__36826),
            .lcout(\u0.dat_o_i_i_1_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_cmdport_T1_RNIV52H3_7_LC_15_19_2 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_T1_RNIV52H3_7_LC_15_19_2 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_cmdport_T1_RNIV52H3_7_LC_15_19_2 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \u0.PIO_cmdport_T1_RNIV52H3_7_LC_15_19_2  (
            .in0(N__48114),
            .in1(N__46566),
            .in2(N__36808),
            .in3(N__36784),
            .lcout(),
            .ltout(\u0.dat_o_0_0_3_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport0_T1_RNI7LNB9_7_LC_15_19_3 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T1_RNI7LNB9_7_LC_15_19_3 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport0_T1_RNI7LNB9_7_LC_15_19_3 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \u0.PIO_dport0_T1_RNI7LNB9_7_LC_15_19_3  (
            .in0(N__36609),
            .in1(N__36589),
            .in2(N__36580),
            .in3(N__50718),
            .lcout(\u0.dat_o_0_0_6_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_cmdport_T1_RNIELKH3_0_LC_15_19_5 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_T1_RNIELKH3_0_LC_15_19_5 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_cmdport_T1_RNIELKH3_0_LC_15_19_5 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \u0.PIO_cmdport_T1_RNIELKH3_0_LC_15_19_5  (
            .in0(N__49416),
            .in1(N__48113),
            .in2(N__36577),
            .in3(N__50717),
            .lcout(),
            .ltout(\u0.dat_o_0_0_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.register_block_gen_stat_reg_int_RNITGPG9_LC_15_19_6 .C_ON=1'b0;
    defparam \u0.register_block_gen_stat_reg_int_RNITGPG9_LC_15_19_6 .SEQ_MODE=4'b0000;
    defparam \u0.register_block_gen_stat_reg_int_RNITGPG9_LC_15_19_6 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \u0.register_block_gen_stat_reg_int_RNITGPG9_LC_15_19_6  (
            .in0(N__37123),
            .in1(N__46567),
            .in2(N__37102),
            .in3(N__37099),
            .lcout(\u0.dat_o_0_0_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport1_T4_5_LC_15_20_0 .C_ON=1'b0;
    defparam \u0.PIO_dport1_T4_5_LC_15_20_0 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport1_T4_5_LC_15_20_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.PIO_dport1_T4_5_LC_15_20_0  (
            .in0(N__38076),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51718),
            .lcout(PIO_dport1_T4_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54248),
            .ce(N__39207),
            .sr(N__53386));
    defparam \u0.PIO_dport1_T4_6_LC_15_20_1 .C_ON=1'b0;
    defparam \u0.PIO_dport1_T4_6_LC_15_20_1 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport1_T4_6_LC_15_20_1 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \u0.PIO_dport1_T4_6_LC_15_20_1  (
            .in0(N__51719),
            .in1(_gnd_net_),
            .in2(N__38188),
            .in3(_gnd_net_),
            .lcout(PIO_dport1_T4_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54248),
            .ce(N__39207),
            .sr(N__53386));
    defparam \u0.PIO_dport1_T4_7_LC_15_20_2 .C_ON=1'b0;
    defparam \u0.PIO_dport1_T4_7_LC_15_20_2 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport1_T4_7_LC_15_20_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.PIO_dport1_T4_7_LC_15_20_2  (
            .in0(N__44842),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51720),
            .lcout(PIO_dport1_T4_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54248),
            .ce(N__39207),
            .sr(N__53386));
    defparam \u0.PIO_dport1_Teoc_5_LC_15_20_4 .C_ON=1'b0;
    defparam \u0.PIO_dport1_Teoc_5_LC_15_20_4 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport1_Teoc_5_LC_15_20_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \u0.PIO_dport1_Teoc_5_LC_15_20_4  (
            .in0(_gnd_net_),
            .in1(N__49342),
            .in2(_gnd_net_),
            .in3(N__51722),
            .lcout(PIO_dport1_Teoc_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54248),
            .ce(N__39207),
            .sr(N__53386));
    defparam \u0.PIO_dport1_Teoc_2_LC_15_20_5 .C_ON=1'b0;
    defparam \u0.PIO_dport1_Teoc_2_LC_15_20_5 .SEQ_MODE=4'b1011;
    defparam \u0.PIO_dport1_Teoc_2_LC_15_20_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \u0.PIO_dport1_Teoc_2_LC_15_20_5  (
            .in0(N__51721),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44239),
            .lcout(PIO_dport1_Teoc_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54248),
            .ce(N__39207),
            .sr(N__53386));
    defparam \u0.PIO_dport1_Teoc_6_LC_15_20_6 .C_ON=1'b0;
    defparam \u0.PIO_dport1_Teoc_6_LC_15_20_6 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport1_Teoc_6_LC_15_20_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \u0.PIO_dport1_Teoc_6_LC_15_20_6  (
            .in0(_gnd_net_),
            .in1(N__47831),
            .in2(_gnd_net_),
            .in3(N__51723),
            .lcout(PIO_dport1_Teoc_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54248),
            .ce(N__39207),
            .sr(N__53386));
    defparam \u0.PIO_dport1_Teoc_7_LC_15_20_7 .C_ON=1'b0;
    defparam \u0.PIO_dport1_Teoc_7_LC_15_20_7 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport1_Teoc_7_LC_15_20_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.PIO_dport1_Teoc_7_LC_15_20_7  (
            .in0(N__51724),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40519),
            .lcout(PIO_dport1_Teoc_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54248),
            .ce(N__39207),
            .sr(N__53386));
    defparam \u0.PIO_dport0_T4_RNI5LI22_0_LC_15_21_0 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T4_RNI5LI22_0_LC_15_21_0 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport0_T4_RNI5LI22_0_LC_15_21_0 .LUT_INIT=16'b0000110010101110;
    LogicCell40 \u0.PIO_dport0_T4_RNI5LI22_0_LC_15_21_0  (
            .in0(N__52907),
            .in1(N__50288),
            .in2(N__37063),
            .in3(N__37042),
            .lcout(\u0.dat_o_0_a2_i_0_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport0_T4_RNI9PI22_2_LC_15_21_2 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T4_RNI9PI22_2_LC_15_21_2 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport0_T4_RNI9PI22_2_LC_15_21_2 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \u0.PIO_dport0_T4_RNI9PI22_2_LC_15_21_2  (
            .in0(N__52908),
            .in1(N__50289),
            .in2(N__37018),
            .in3(N__37542),
            .lcout(\u0.dat_o_i_0_0_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport0_T4_RNIDTI22_4_LC_15_21_4 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T4_RNIDTI22_4_LC_15_21_4 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport0_T4_RNIDTI22_4_LC_15_21_4 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \u0.PIO_dport0_T4_RNIDTI22_4_LC_15_21_4  (
            .in0(N__52909),
            .in1(N__50290),
            .in2(N__37528),
            .in3(N__37500),
            .lcout(\u0.dat_o_0_a2_i_0_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport0_T4_RNIFVI22_5_LC_15_21_5 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T4_RNIFVI22_5_LC_15_21_5 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport0_T4_RNIFVI22_5_LC_15_21_5 .LUT_INIT=16'b0000110010101110;
    LogicCell40 \u0.PIO_dport0_T4_RNIFVI22_5_LC_15_21_5  (
            .in0(N__50291),
            .in1(N__52910),
            .in2(N__37464),
            .in3(N__37440),
            .lcout(\u0.dat_o_i_0_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport0_T4_RNIH1J22_6_LC_15_21_6 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T4_RNIH1J22_6_LC_15_21_6 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport0_T4_RNIH1J22_6_LC_15_21_6 .LUT_INIT=16'b0010111100100010;
    LogicCell40 \u0.PIO_dport0_T4_RNIH1J22_6_LC_15_21_6  (
            .in0(N__52911),
            .in1(N__37413),
            .in2(N__37399),
            .in3(N__50292),
            .lcout(\u0.dat_o_i_0_0_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev1_Teoc_3_LC_15_22_0 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Teoc_3_LC_15_22_0 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev1_Teoc_3_LC_15_22_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \u0.DMA_dev1_Teoc_3_LC_15_22_0  (
            .in0(_gnd_net_),
            .in1(N__37717),
            .in2(_gnd_net_),
            .in3(N__51928),
            .lcout(DMA_dev1_Teoc_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54273),
            .ce(N__39542),
            .sr(N__53396));
    defparam \u0.DMA_dev1_Teoc_5_LC_15_22_1 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Teoc_5_LC_15_22_1 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev1_Teoc_5_LC_15_22_1 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \u0.DMA_dev1_Teoc_5_LC_15_22_1  (
            .in0(N__49343),
            .in1(_gnd_net_),
            .in2(N__52112),
            .in3(_gnd_net_),
            .lcout(DMA_dev1_Teoc_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54273),
            .ce(N__39542),
            .sr(N__53396));
    defparam \u0.DMA_dev1_Tm_3_LC_15_22_2 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Tm_3_LC_15_22_2 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev1_Tm_3_LC_15_22_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \u0.DMA_dev1_Tm_3_LC_15_22_2  (
            .in0(_gnd_net_),
            .in1(N__51934),
            .in2(_gnd_net_),
            .in3(N__37363),
            .lcout(DMA_dev1_Tm_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54273),
            .ce(N__39542),
            .sr(N__53396));
    defparam \u0.DMA_dev1_Teoc_6_LC_15_22_3 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Teoc_6_LC_15_22_3 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev1_Teoc_6_LC_15_22_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.DMA_dev1_Teoc_6_LC_15_22_3  (
            .in0(N__51932),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47822),
            .lcout(DMA_dev1_Teoc_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54273),
            .ce(N__39542),
            .sr(N__53396));
    defparam \u0.DMA_dev1_Teoc_7_LC_15_22_4 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Teoc_7_LC_15_22_4 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev1_Teoc_7_LC_15_22_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \u0.DMA_dev1_Teoc_7_LC_15_22_4  (
            .in0(_gnd_net_),
            .in1(N__51933),
            .in2(_gnd_net_),
            .in3(N__40504),
            .lcout(DMA_dev1_Teoc_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54273),
            .ce(N__39542),
            .sr(N__53396));
    defparam \u0.DMA_dev1_Tm_4_LC_15_22_5 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Tm_4_LC_15_22_5 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev1_Tm_4_LC_15_22_5 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \u0.DMA_dev1_Tm_4_LC_15_22_5  (
            .in0(N__37225),
            .in1(_gnd_net_),
            .in2(N__52113),
            .in3(_gnd_net_),
            .lcout(DMA_dev1_Tm_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54273),
            .ce(N__39542),
            .sr(N__53396));
    defparam \u0.DMA_dev1_Tm_5_LC_15_22_6 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Tm_5_LC_15_22_6 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev1_Tm_5_LC_15_22_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.DMA_dev1_Tm_5_LC_15_22_6  (
            .in0(N__46289),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51938),
            .lcout(DMA_dev1_Tm_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54273),
            .ce(N__39542),
            .sr(N__53396));
    defparam \u0.DMA_dev1_Tm_6_LC_15_22_7 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Tm_6_LC_15_22_7 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev1_Tm_6_LC_15_22_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.DMA_dev1_Tm_6_LC_15_22_7  (
            .in0(N__51939),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39421),
            .lcout(DMA_dev1_Tm_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54273),
            .ce(N__39542),
            .sr(N__53396));
    defparam \u0.CtrlReg_RNIVM5S3_27_LC_15_23_0 .C_ON=1'b0;
    defparam \u0.CtrlReg_RNIVM5S3_27_LC_15_23_0 .SEQ_MODE=4'b0000;
    defparam \u0.CtrlReg_RNIVM5S3_27_LC_15_23_0 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \u0.CtrlReg_RNIVM5S3_27_LC_15_23_0  (
            .in0(N__37804),
            .in1(N__48111),
            .in2(N__37633),
            .in3(N__48327),
            .lcout(),
            .ltout(\u0.dat_o_i_i_1_27_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport0_Teoc_RNI0G9H7_3_LC_15_23_1 .C_ON=1'b0;
    defparam \u0.PIO_dport0_Teoc_RNI0G9H7_3_LC_15_23_1 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport0_Teoc_RNI0G9H7_3_LC_15_23_1 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \u0.PIO_dport0_Teoc_RNI0G9H7_3_LC_15_23_1  (
            .in0(N__37588),
            .in1(N__50724),
            .in2(N__37783),
            .in3(N__37780),
            .lcout(),
            .ltout(\u0.dat_o_i_i_4_27_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev1_Teoc_RNILDL3G_3_LC_15_23_2 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Teoc_RNILDL3G_3_LC_15_23_2 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev1_Teoc_RNILDL3G_3_LC_15_23_2 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \u0.DMA_dev1_Teoc_RNILDL3G_3_LC_15_23_2  (
            .in0(N__54704),
            .in1(N__37552),
            .in2(N__37759),
            .in3(N__37749),
            .lcout(N_269),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.CtrlReg_27_LC_15_23_3 .C_ON=1'b0;
    defparam \u0.CtrlReg_27_LC_15_23_3 .SEQ_MODE=4'b1010;
    defparam \u0.CtrlReg_27_LC_15_23_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.CtrlReg_27_LC_15_23_3  (
            .in0(N__51940),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37716),
            .lcout(\u0.CtrlRegZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54283),
            .ce(N__53651),
            .sr(N__53401));
    defparam \u0.PIO_dport1_Teoc_RNIH00N1_3_LC_15_23_4 .C_ON=1'b0;
    defparam \u0.PIO_dport1_Teoc_RNIH00N1_3_LC_15_23_4 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport1_Teoc_RNIH00N1_3_LC_15_23_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \u0.PIO_dport1_Teoc_RNIH00N1_3_LC_15_23_4  (
            .in0(N__37621),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46951),
            .lcout(\u0.N_1682 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev0_Teoc_RNI483P6_3_LC_15_23_5 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Teoc_RNI483P6_3_LC_15_23_5 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev0_Teoc_RNI483P6_3_LC_15_23_5 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \u0.DMA_dev0_Teoc_RNI483P6_3_LC_15_23_5  (
            .in0(N__37578),
            .in1(N__37564),
            .in2(N__48577),
            .in3(N__47181),
            .lcout(\u0.dat_o_i_i_0_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.dat_o_i_a2_21_LC_15_24_0 .C_ON=1'b0;
    defparam \u0.dat_o_i_a2_21_LC_15_24_0 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_i_a2_21_LC_15_24_0 .LUT_INIT=16'b0000110001000100;
    LogicCell40 \u0.dat_o_i_a2_21_LC_15_24_0  (
            .in0(N__37966),
            .in1(N__50464),
            .in2(N__37933),
            .in3(N__48890),
            .lcout(),
            .ltout(\u0.N_1636_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport0_T4_RNIJTPO9_5_LC_15_24_1 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T4_RNIJTPO9_5_LC_15_24_1 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport0_T4_RNIJTPO9_5_LC_15_24_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \u0.PIO_dport0_T4_RNIJTPO9_5_LC_15_24_1  (
            .in0(N__49624),
            .in1(N__37894),
            .in2(N__38113),
            .in3(N__38110),
            .lcout(N_259_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.CtrlReg_21_LC_15_24_2 .C_ON=1'b0;
    defparam \u0.CtrlReg_21_LC_15_24_2 .SEQ_MODE=4'b1010;
    defparam \u0.CtrlReg_21_LC_15_24_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.CtrlReg_21_LC_15_24_2  (
            .in0(N__51941),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38069),
            .lcout(\u0.CtrlRegZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54293),
            .ce(N__53561),
            .sr(N__53404));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNISK0R_21_LC_15_24_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNISK0R_21_LC_15_24_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNISK0R_21_LC_15_24_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNISK0R_21_LC_15_24_3  (
            .in0(N__38008),
            .in1(N__37993),
            .in2(_gnd_net_),
            .in3(N__45687),
            .lcout(),
            .ltout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNISK0RZ0Z_21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIE8HM1_2_LC_15_24_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIE8HM1_2_LC_15_24_4 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIE8HM1_2_LC_15_24_4 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIE8HM1_2_LC_15_24_4  (
            .in0(N__50013),
            .in1(_gnd_net_),
            .in2(N__37981),
            .in3(N__37978),
            .lcout(iQ_RNIE8HM1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI1PD71_21_LC_15_24_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI1PD71_21_LC_15_24_5 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI1PD71_21_LC_15_24_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI1PD71_21_LC_15_24_5  (
            .in0(N__37960),
            .in1(N__37945),
            .in2(_gnd_net_),
            .in3(N__50012),
            .lcout(mem_mem_ram6__RNI1PD71_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.CtrlReg_RNI49LU1_21_LC_15_24_6 .C_ON=1'b0;
    defparam \u0.CtrlReg_RNI49LU1_21_LC_15_24_6 .SEQ_MODE=4'b0000;
    defparam \u0.CtrlReg_RNI49LU1_21_LC_15_24_6 .LUT_INIT=16'b0100010011110100;
    LogicCell40 \u0.CtrlReg_RNI49LU1_21_LC_15_24_6  (
            .in0(N__37924),
            .in1(N__45030),
            .in2(N__44937),
            .in3(N__37915),
            .lcout(\u0.dat_o_i_2_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.dat_o_0_0_a2_0_7_LC_15_25_0 .C_ON=1'b0;
    defparam \u0.dat_o_0_0_a2_0_7_LC_15_25_0 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_0_0_a2_0_7_LC_15_25_0 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \u0.dat_o_0_0_a2_0_7_LC_15_25_0  (
            .in0(N__47182),
            .in1(N__38248),
            .in2(N__48938),
            .in3(N__38266),
            .lcout(),
            .ltout(\u0.N_1979_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport0_T1_RNIVH2NI_7_LC_15_25_1 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T1_RNIVH2NI_7_LC_15_25_1 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport0_T1_RNIVH2NI_7_LC_15_25_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \u0.PIO_dport0_T1_RNIVH2NI_7_LC_15_25_1  (
            .in0(N__37888),
            .in1(N__38260),
            .in2(N__37879),
            .in3(N__38299),
            .lcout(wb_dat_o_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.q_7_LC_15_25_2 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.q_7_LC_15_25_2 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.q_7_LC_15_25_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \u1.PIO_control.PIO_access_control.q_7_LC_15_25_2  (
            .in0(N__38395),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(PIOq_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54304),
            .ce(N__45931),
            .sr(_gnd_net_));
    defparam \u0.CtrlReg_RNIOOLH2_7_LC_15_25_3 .C_ON=1'b0;
    defparam \u0.CtrlReg_RNIOOLH2_7_LC_15_25_3 .SEQ_MODE=4'b0000;
    defparam \u0.CtrlReg_RNIOOLH2_7_LC_15_25_3 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \u0.CtrlReg_RNIOOLH2_7_LC_15_25_3  (
            .in0(N__47454),
            .in1(N__38353),
            .in2(N__38347),
            .in3(N__48328),
            .lcout(\u0.dat_o_0_0_2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIUGOK1_2_LC_15_25_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIUGOK1_2_LC_15_25_4 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIUGOK1_2_LC_15_25_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIUGOK1_2_LC_15_25_4  (
            .in0(N__50017),
            .in1(N__38293),
            .in2(_gnd_net_),
            .in3(N__38281),
            .lcout(iQ_RNIUGOK1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev0_Tm_RNIA8DS1_7_LC_15_25_5 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Tm_RNIA8DS1_7_LC_15_25_5 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev0_Tm_RNIA8DS1_7_LC_15_25_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \u0.DMA_dev0_Tm_RNIA8DS1_7_LC_15_25_5  (
            .in0(N__48544),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39763),
            .lcout(\u0.N_1980 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNITSOD1_7_LC_15_25_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNITSOD1_7_LC_15_25_6 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNITSOD1_7_LC_15_25_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNITSOD1_7_LC_15_25_6  (
            .in0(N__50016),
            .in1(N__38872),
            .in2(_gnd_net_),
            .in3(N__38254),
            .lcout(mem_mem_ram6__RNITSOD1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI4SD71_22_LC_15_26_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI4SD71_22_LC_15_26_0 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI4SD71_22_LC_15_26_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI4SD71_22_LC_15_26_0  (
            .in0(N__38242),
            .in1(N__38227),
            .in2(_gnd_net_),
            .in3(N__50018),
            .lcout(mem_mem_ram6__RNI4SD71_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIUM0R_22_LC_15_26_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIUM0R_22_LC_15_26_1 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIUM0R_22_LC_15_26_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIUM0R_22_LC_15_26_1  (
            .in0(N__38212),
            .in1(N__45701),
            .in2(_gnd_net_),
            .in3(N__38200),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNIUM0RZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.CtrlReg_22_LC_15_26_4 .C_ON=1'b0;
    defparam \u0.CtrlReg_22_LC_15_26_4 .SEQ_MODE=4'b1010;
    defparam \u0.CtrlReg_22_LC_15_26_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \u0.CtrlReg_22_LC_15_26_4  (
            .in0(_gnd_net_),
            .in1(N__38182),
            .in2(_gnd_net_),
            .in3(N__52114),
            .lcout(\u0.CtrlRegZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54312),
            .ce(N__53560),
            .sr(N__53408));
    defparam \u0.CtrlReg_RNI6BLU1_22_LC_15_26_5 .C_ON=1'b0;
    defparam \u0.CtrlReg_RNI6BLU1_22_LC_15_26_5 .SEQ_MODE=4'b0000;
    defparam \u0.CtrlReg_RNI6BLU1_22_LC_15_26_5 .LUT_INIT=16'b0010001011110010;
    LogicCell40 \u0.CtrlReg_RNI6BLU1_22_LC_15_26_5  (
            .in0(N__45048),
            .in1(N__38944),
            .in2(N__44938),
            .in3(N__38938),
            .lcout(),
            .ltout(\u0.dat_o_i_0_2_22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport0_T4_RNIU8QO9_6_LC_15_26_6 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T4_RNIU8QO9_6_LC_15_26_6 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport0_T4_RNIU8QO9_6_LC_15_26_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \u0.PIO_dport0_T4_RNIU8QO9_6_LC_15_26_6  (
            .in0(N__40897),
            .in1(N__49637),
            .in2(N__38917),
            .in3(N__38914),
            .lcout(N_330_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNICBTN_7_LC_15_27_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNICBTN_7_LC_15_27_0 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNICBTN_7_LC_15_27_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNICBTN_7_LC_15_27_0  (
            .in0(N__38887),
            .in1(N__38863),
            .in2(_gnd_net_),
            .in3(N__45689),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNICBTNZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__7_LC_15_27_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__7_LC_15_27_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__7_LC_15_27_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__7_LC_15_27_1  (
            .in0(N__42938),
            .in1(N__38840),
            .in2(_gnd_net_),
            .in3(N__38742),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54321),
            .ce(N__41849),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__23_LC_15_27_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__23_LC_15_27_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__23_LC_15_27_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__23_LC_15_27_2  (
            .in0(N__38839),
            .in1(N__38741),
            .in2(_gnd_net_),
            .in3(N__42940),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54321),
            .ce(N__41849),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNIEDTN_8_LC_15_27_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNIEDTN_8_LC_15_27_4 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNIEDTN_8_LC_15_27_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNIEDTN_8_LC_15_27_4  (
            .in0(N__38635),
            .in1(N__38650),
            .in2(_gnd_net_),
            .in3(N__45690),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNIEDTNZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__8_LC_15_27_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__8_LC_15_27_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__8_LC_15_27_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__8_LC_15_27_5  (
            .in0(N__42939),
            .in1(_gnd_net_),
            .in2(N__38484),
            .in3(N__38586),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54321),
            .ce(N__41849),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__24_LC_15_27_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__24_LC_15_27_6 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__24_LC_15_27_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__24_LC_15_27_6  (
            .in0(N__38585),
            .in1(N__38461),
            .in2(_gnd_net_),
            .in3(N__42941),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54321),
            .ce(N__41849),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI7VD71_23_LC_15_28_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI7VD71_23_LC_15_28_0 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI7VD71_23_LC_15_28_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI7VD71_23_LC_15_28_0  (
            .in0(N__38407),
            .in1(N__39085),
            .in2(_gnd_net_),
            .in3(N__50168),
            .lcout(u1_DMA_control_gen_DMAbuf_Rxbuf_mem_N_1224),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI81IT_23_LC_15_28_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI81IT_23_LC_15_28_1 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI81IT_23_LC_15_28_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI81IT_23_LC_15_28_1  (
            .in0(N__45698),
            .in1(N__39106),
            .in2(_gnd_net_),
            .in3(N__39100),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNI81ITZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNIGFTN_9_LC_15_28_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNIGFTN_9_LC_15_28_2 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNIGFTN_9_LC_15_28_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNIGFTN_9_LC_15_28_2  (
            .in0(N__39079),
            .in1(N__39070),
            .in2(_gnd_net_),
            .in3(N__45696),
            .lcout(),
            .ltout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNIGFTNZ0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI33PD1_9_LC_15_28_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI33PD1_9_LC_15_28_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI33PD1_9_LC_15_28_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI33PD1_9_LC_15_28_3  (
            .in0(N__50167),
            .in1(_gnd_net_),
            .in2(N__39058),
            .in3(N__39055),
            .lcout(mem_mem_ram6__RNI33PD1_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNIUSSN_0_LC_15_28_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNIUSSN_0_LC_15_28_5 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNIUSSN_0_LC_15_28_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNIUSSN_0_LC_15_28_5  (
            .in0(N__45697),
            .in1(N__39043),
            .in2(_gnd_net_),
            .in3(N__39031),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__RNIUSSNZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIU9753_3_LC_15_28_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIU9753_3_LC_15_28_7 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIU9753_3_LC_15_28_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIU9753_3_LC_15_28_7  (
            .in0(N__48944),
            .in1(N__39787),
            .in2(_gnd_net_),
            .in3(N__39019),
            .lcout(DMAq_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIMGHM1_2_LC_15_29_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIMGHM1_2_LC_15_29_0 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIMGHM1_2_LC_15_29_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIMGHM1_2_LC_15_29_0  (
            .in0(N__50112),
            .in1(N__39007),
            .in2(_gnd_net_),
            .in3(N__38971),
            .lcout(u1_DMA_control_gen_DMAbuf_Rxbuf_mem_N_1160),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI0P0R_23_LC_15_29_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI0P0R_23_LC_15_29_2 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI0P0R_23_LC_15_29_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI0P0R_23_LC_15_29_2  (
            .in0(N__45699),
            .in1(N__38995),
            .in2(_gnd_net_),
            .in3(N__38983),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI0P0RZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIC5IT_25_LC_15_29_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIC5IT_25_LC_15_29_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIC5IT_25_LC_15_29_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIC5IT_25_LC_15_29_3  (
            .in0(N__38965),
            .in1(N__45700),
            .in2(_gnd_net_),
            .in3(N__38956),
            .lcout(),
            .ltout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram5__RNIC5ITZ0Z_25_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNID5E71_25_LC_15_29_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNID5E71_25_LC_15_29_4 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNID5E71_25_LC_15_29_4 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNID5E71_25_LC_15_29_4  (
            .in0(_gnd_net_),
            .in1(N__50111),
            .in2(N__39799),
            .in3(N__39796),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNID5E71Z0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIUIA71_11_LC_15_30_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIUIA71_11_LC_15_30_2 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIUIA71_11_LC_15_30_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIUIA71_11_LC_15_30_2  (
            .in0(N__41311),
            .in1(N__39781),
            .in2(_gnd_net_),
            .in3(N__50113),
            .lcout(),
            .ltout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIUIA71Z0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIRUU43_3_LC_15_30_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIRUU43_3_LC_15_30_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIRUU43_3_LC_15_30_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIRUU43_3_LC_15_30_3  (
            .in0(N__48945),
            .in1(_gnd_net_),
            .in2(N__39775),
            .in3(N__39772),
            .lcout(DMAq_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev0_Tm_7_LC_16_14_0 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Tm_7_LC_16_14_0 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev0_Tm_7_LC_16_14_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \u0.DMA_dev0_Tm_7_LC_16_14_0  (
            .in0(_gnd_net_),
            .in1(N__51363),
            .in2(_gnd_net_),
            .in3(N__39607),
            .lcout(DMA_dev0_Tm_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54261),
            .ce(N__39742),
            .sr(N__53381));
    defparam \u0.DMA_dev1_Tm_7_LC_16_15_0 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Tm_7_LC_16_15_0 .SEQ_MODE=4'b1010;
    defparam \u0.DMA_dev1_Tm_7_LC_16_15_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \u0.DMA_dev1_Tm_7_LC_16_15_0  (
            .in0(_gnd_net_),
            .in1(N__51364),
            .in2(_gnd_net_),
            .in3(N__39624),
            .lcout(DMA_dev1_Tm_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54249),
            .ce(N__39543),
            .sr(N__53376));
    defparam \u0.PIO_dport0_T1_6_LC_16_16_7 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T1_6_LC_16_16_7 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport0_T1_6_LC_16_16_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.PIO_dport0_T1_6_LC_16_16_7  (
            .in0(N__51366),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39455),
            .lcout(PIO_dport0_T1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54235),
            .ce(N__49377),
            .sr(N__53362));
    defparam \u0.CtrlReg_1_LC_16_17_5 .C_ON=1'b0;
    defparam \u0.CtrlReg_1_LC_16_17_5 .SEQ_MODE=4'b1010;
    defparam \u0.CtrlReg_1_LC_16_17_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.CtrlReg_1_LC_16_17_5  (
            .in0(N__39308),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51373),
            .lcout(PIO_cmdport_IORDYen),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54216),
            .ce(N__53653),
            .sr(N__53377));
    defparam \u0.PIO_dport1_Teoc_4_LC_16_18_7 .C_ON=1'b0;
    defparam \u0.PIO_dport1_Teoc_4_LC_16_18_7 .SEQ_MODE=4'b1011;
    defparam \u0.PIO_dport1_Teoc_4_LC_16_18_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \u0.PIO_dport1_Teoc_4_LC_16_18_7  (
            .in0(N__51611),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46123),
            .lcout(PIO_dport1_Teoc_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54236),
            .ce(N__39201),
            .sr(N__53382));
    defparam \u0.CtrlReg_RNIHG6Q3_10_LC_16_19_0 .C_ON=1'b0;
    defparam \u0.CtrlReg_RNIHG6Q3_10_LC_16_19_0 .SEQ_MODE=4'b0000;
    defparam \u0.CtrlReg_RNIHG6Q3_10_LC_16_19_0 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \u0.CtrlReg_RNIHG6Q3_10_LC_16_19_0  (
            .in0(N__39120),
            .in1(N__48065),
            .in2(N__48330),
            .in3(N__40069),
            .lcout(),
            .ltout(\u0.dat_o_i_i_3_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport0_T2_RNI3R5D9_2_LC_16_19_1 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T2_RNI3R5D9_2_LC_16_19_1 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport0_T2_RNI3R5D9_2_LC_16_19_1 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \u0.PIO_dport0_T2_RNI3R5D9_2_LC_16_19_1  (
            .in0(N__50716),
            .in1(N__43519),
            .in2(N__40207),
            .in3(N__40204),
            .lcout(\u0.dat_o_i_i_6_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.CtrlReg_10_LC_16_19_3 .C_ON=1'b0;
    defparam \u0.CtrlReg_10_LC_16_19_3 .SEQ_MODE=4'b1010;
    defparam \u0.CtrlReg_10_LC_16_19_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \u0.CtrlReg_10_LC_16_19_3  (
            .in0(_gnd_net_),
            .in1(N__40173),
            .in2(_gnd_net_),
            .in3(N__51612),
            .lcout(\u0.CtrlRegZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54250),
            .ce(N__53610),
            .sr(N__53387));
    defparam \u0.DMA_dev0_Td_RNIS7H22_2_LC_16_19_4 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Td_RNIS7H22_2_LC_16_19_4 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev0_Td_RNIS7H22_2_LC_16_19_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \u0.DMA_dev0_Td_RNIS7H22_2_LC_16_19_4  (
            .in0(N__40063),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48570),
            .lcout(),
            .ltout(\u0.N_1990_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport0_T2_RNI7C9HJ_2_LC_16_19_5 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T2_RNI7C9HJ_2_LC_16_19_5 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport0_T2_RNI7C9HJ_2_LC_16_19_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \u0.PIO_dport0_T2_RNI7C9HJ_2_LC_16_19_5  (
            .in0(N__40045),
            .in1(N__40033),
            .in2(N__40021),
            .in3(N__40018),
            .lcout(N_1097),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport1_Teoc_RNIETVM1_0_LC_16_20_0 .C_ON=1'b0;
    defparam \u0.PIO_dport1_Teoc_RNIETVM1_0_LC_16_20_0 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport1_Teoc_RNIETVM1_0_LC_16_20_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \u0.PIO_dport1_Teoc_RNIETVM1_0_LC_16_20_0  (
            .in0(N__46905),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39994),
            .lcout(),
            .ltout(\u0.N_1661_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport0_Teoc_RNIK39H7_0_LC_16_20_1 .C_ON=1'b0;
    defparam \u0.PIO_dport0_Teoc_RNIK39H7_0_LC_16_20_1 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport0_Teoc_RNIK39H7_0_LC_16_20_1 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \u0.PIO_dport0_Teoc_RNIK39H7_0_LC_16_20_1  (
            .in0(N__39928),
            .in1(N__50678),
            .in2(N__39973),
            .in3(N__39970),
            .lcout(\u0.dat_o_i_i_4_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.CtrlReg_RNIPG5S3_24_LC_16_20_3 .C_ON=1'b0;
    defparam \u0.CtrlReg_RNIPG5S3_24_LC_16_20_3 .SEQ_MODE=4'b0000;
    defparam \u0.CtrlReg_RNIPG5S3_24_LC_16_20_3 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \u0.CtrlReg_RNIPG5S3_24_LC_16_20_3  (
            .in0(N__39805),
            .in1(N__48283),
            .in2(N__48061),
            .in3(N__39948),
            .lcout(\u0.dat_o_i_i_1_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.CtrlReg_24_LC_16_20_4 .C_ON=1'b0;
    defparam \u0.CtrlReg_24_LC_16_20_4 .SEQ_MODE=4'b1010;
    defparam \u0.CtrlReg_24_LC_16_20_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.CtrlReg_24_LC_16_20_4  (
            .in0(N__51614),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39921),
            .lcout(\u0.CtrlRegZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54262),
            .ce(N__53647),
            .sr(N__53391));
    defparam \u0.CtrlReg_31_LC_16_21_0 .C_ON=1'b0;
    defparam \u0.CtrlReg_31_LC_16_21_0 .SEQ_MODE=4'b1010;
    defparam \u0.CtrlReg_31_LC_16_21_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \u0.CtrlReg_31_LC_16_21_0  (
            .in0(_gnd_net_),
            .in1(N__40526),
            .in2(_gnd_net_),
            .in3(N__52003),
            .lcout(\u0.CtrlRegZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54274),
            .ce(N__53652),
            .sr(N__53397));
    defparam \u0.DMA_dev0_Teoc_RNI5F9P6_7_LC_16_21_1 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Teoc_RNI5F9P6_7_LC_16_21_1 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev0_Teoc_RNI5F9P6_7_LC_16_21_1 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \u0.DMA_dev0_Teoc_RNI5F9P6_7_LC_16_21_1  (
            .in0(N__40453),
            .in1(N__48480),
            .in2(N__47209),
            .in3(N__40438),
            .lcout(),
            .ltout(\u0.dat_o_i_i_0_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev1_Teoc_RNI11T3G_7_LC_16_21_2 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Teoc_RNI11T3G_7_LC_16_21_2 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev1_Teoc_RNI11T3G_7_LC_16_21_2 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \u0.DMA_dev1_Teoc_RNI11T3G_7_LC_16_21_2  (
            .in0(N__40288),
            .in1(N__54588),
            .in2(N__40411),
            .in3(N__40398),
            .lcout(N_277),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport1_Teoc_RNIL40N1_7_LC_16_21_3 .C_ON=1'b0;
    defparam \u0.PIO_dport1_Teoc_RNIL40N1_7_LC_16_21_3 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport1_Teoc_RNIL40N1_7_LC_16_21_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \u0.PIO_dport1_Teoc_RNIL40N1_7_LC_16_21_3  (
            .in0(_gnd_net_),
            .in1(N__46867),
            .in2(_gnd_net_),
            .in3(N__40362),
            .lcout(\u0.N_1710 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.CtrlReg_RNIUM6S3_31_LC_16_21_4 .C_ON=1'b0;
    defparam \u0.CtrlReg_RNIUM6S3_31_LC_16_21_4 .SEQ_MODE=4'b0000;
    defparam \u0.CtrlReg_RNIUM6S3_31_LC_16_21_4 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \u0.CtrlReg_RNIUM6S3_31_LC_16_21_4  (
            .in0(N__40348),
            .in1(N__48253),
            .in2(N__48060),
            .in3(N__40342),
            .lcout(),
            .ltout(\u0.dat_o_i_i_1_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport0_Teoc_RNI7OAH7_7_LC_16_21_5 .C_ON=1'b0;
    defparam \u0.PIO_dport0_Teoc_RNI7OAH7_7_LC_16_21_5 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport0_Teoc_RNI7OAH7_7_LC_16_21_5 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \u0.PIO_dport0_Teoc_RNI7OAH7_7_LC_16_21_5  (
            .in0(N__50719),
            .in1(N__40318),
            .in2(N__40312),
            .in3(N__40309),
            .lcout(\u0.dat_o_i_i_4_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.CtrlReg_RNIRI5S3_25_LC_16_22_0 .C_ON=1'b0;
    defparam \u0.CtrlReg_RNIRI5S3_25_LC_16_22_0 .SEQ_MODE=4'b0000;
    defparam \u0.CtrlReg_RNIRI5S3_25_LC_16_22_0 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \u0.CtrlReg_RNIRI5S3_25_LC_16_22_0  (
            .in0(N__40792),
            .in1(N__48027),
            .in2(N__48326),
            .in3(N__40282),
            .lcout(),
            .ltout(\u0.dat_o_i_i_1_25_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport0_Teoc_RNIO79H7_1_LC_16_22_1 .C_ON=1'b0;
    defparam \u0.PIO_dport0_Teoc_RNIO79H7_1_LC_16_22_1 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport0_Teoc_RNIO79H7_1_LC_16_22_1 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \u0.PIO_dport0_Teoc_RNIO79H7_1_LC_16_22_1  (
            .in0(N__40213),
            .in1(N__50720),
            .in2(N__40264),
            .in3(N__40261),
            .lcout(\u0.dat_o_i_i_4_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport1_Teoc_RNIFUVM1_1_LC_16_22_3 .C_ON=1'b0;
    defparam \u0.PIO_dport1_Teoc_RNIFUVM1_1_LC_16_22_3 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport1_Teoc_RNIFUVM1_1_LC_16_22_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \u0.PIO_dport1_Teoc_RNIFUVM1_1_LC_16_22_3  (
            .in0(_gnd_net_),
            .in1(N__46888),
            .in2(_gnd_net_),
            .in3(N__40239),
            .lcout(\u0.N_1668 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.CtrlReg_25_LC_16_22_4 .C_ON=1'b0;
    defparam \u0.CtrlReg_25_LC_16_22_4 .SEQ_MODE=4'b1010;
    defparam \u0.CtrlReg_25_LC_16_22_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \u0.CtrlReg_25_LC_16_22_4  (
            .in0(_gnd_net_),
            .in1(N__40871),
            .in2(_gnd_net_),
            .in3(N__51862),
            .lcout(\u0.CtrlRegZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54284),
            .ce(N__53646),
            .sr(N__53402));
    defparam \u0.DMA_dev0_Teoc_RNIKN2P6_1_LC_16_22_5 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Teoc_RNIKN2P6_1_LC_16_22_5 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev0_Teoc_RNIKN2P6_1_LC_16_22_5 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \u0.DMA_dev0_Teoc_RNIKN2P6_1_LC_16_22_5  (
            .in0(N__47111),
            .in1(N__40786),
            .in2(N__40774),
            .in3(N__48531),
            .lcout(\u0.dat_o_i_i_0_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev0_Tm_RNIN9HR3_6_LC_16_23_0 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Tm_RNIN9HR3_6_LC_16_23_0 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev0_Tm_RNIN9HR3_6_LC_16_23_0 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \u0.DMA_dev0_Tm_RNIN9HR3_6_LC_16_23_0  (
            .in0(N__40750),
            .in1(N__46906),
            .in2(N__40735),
            .in3(N__48540),
            .lcout(),
            .ltout(\u0.dat_o_0_0_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev1_Tm_RNIRO2E9_6_LC_16_23_1 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Tm_RNIRO2E9_6_LC_16_23_1 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev1_Tm_RNIRO2E9_6_LC_16_23_1 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \u0.DMA_dev1_Tm_RNIRO2E9_6_LC_16_23_1  (
            .in0(N__54674),
            .in1(N__40537),
            .in2(N__40708),
            .in3(N__40701),
            .lcout(\u0.dat_o_0_0_6_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.dat_o_0_0_a2_0_6_LC_16_23_3 .C_ON=1'b0;
    defparam \u0.dat_o_0_0_a2_0_6_LC_16_23_3 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_0_0_a2_0_6_LC_16_23_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \u0.dat_o_0_0_a2_0_6_LC_16_23_3  (
            .in0(N__47468),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40648),
            .lcout(\u0.N_1970 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.q_6_LC_16_23_4 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.q_6_LC_16_23_4 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.q_6_LC_16_23_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \u1.PIO_control.PIO_access_control.q_6_LC_16_23_4  (
            .in0(N__40687),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(PIOq_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54294),
            .ce(N__45936),
            .sr(_gnd_net_));
    defparam \u0.CtrlReg_RNISQLO4_6_LC_16_23_5 .C_ON=1'b0;
    defparam \u0.CtrlReg_RNISQLO4_6_LC_16_23_5 .SEQ_MODE=4'b0000;
    defparam \u0.CtrlReg_RNISQLO4_6_LC_16_23_5 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \u0.CtrlReg_RNISQLO4_6_LC_16_23_5  (
            .in0(N__40642),
            .in1(N__48331),
            .in2(_gnd_net_),
            .in3(N__40624),
            .lcout(\u0.dat_o_0_0_2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_cmdport_T1_RNIQ1LH3_6_LC_16_23_6 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_T1_RNIQ1LH3_6_LC_16_23_6 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_cmdport_T1_RNIQ1LH3_6_LC_16_23_6 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \u0.PIO_cmdport_T1_RNIQ1LH3_6_LC_16_23_6  (
            .in0(N__40588),
            .in1(N__48110),
            .in2(N__50747),
            .in3(N__40557),
            .lcout(\u0.dat_o_0_0_3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI00PD1_8_LC_16_24_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI00PD1_8_LC_16_24_0 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI00PD1_8_LC_16_24_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI00PD1_8_LC_16_24_0  (
            .in0(N__50171),
            .in1(N__41140),
            .in2(_gnd_net_),
            .in3(N__41128),
            .lcout(mem_mem_ram6__RNI00PD1_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIBAOD1_1_LC_16_24_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIBAOD1_1_LC_16_24_1 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIBAOD1_1_LC_16_24_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIBAOD1_1_LC_16_24_1  (
            .in0(N__41116),
            .in1(N__41545),
            .in2(_gnd_net_),
            .in3(N__50172),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIBAOD1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev1_Tm_RNI0HNIJ_6_LC_16_24_7 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Tm_RNI0HNIJ_6_LC_16_24_7 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev1_Tm_RNI0HNIJ_6_LC_16_24_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \u0.DMA_dev1_Tm_RNI0HNIJ_6_LC_16_24_7  (
            .in0(N__41104),
            .in1(N__41083),
            .in2(N__41077),
            .in3(N__41068),
            .lcout(wb_dat_o_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.CtrlReg_RNI37KU1_16_LC_16_25_0 .C_ON=1'b0;
    defparam \u0.CtrlReg_RNI37KU1_16_LC_16_25_0 .SEQ_MODE=4'b0000;
    defparam \u0.CtrlReg_RNI37KU1_16_LC_16_25_0 .LUT_INIT=16'b0101000011011100;
    LogicCell40 \u0.CtrlReg_RNI37KU1_16_LC_16_25_0  (
            .in0(N__41044),
            .in1(N__45049),
            .in2(N__44904),
            .in3(N__40960),
            .lcout(\u0.dat_o_0_a2_i_2_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.CtrlReg_16_LC_16_25_2 .C_ON=1'b0;
    defparam \u0.CtrlReg_16_LC_16_25_2 .SEQ_MODE=4'b1010;
    defparam \u0.CtrlReg_16_LC_16_25_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \u0.CtrlReg_16_LC_16_25_2  (
            .in0(_gnd_net_),
            .in1(N__41023),
            .in2(_gnd_net_),
            .in3(N__51863),
            .lcout(\u0.CtrlRegZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54313),
            .ce(N__53634),
            .sr(N__53409));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI4RUQ_16_LC_16_25_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI4RUQ_16_LC_16_25_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI4RUQ_16_LC_16_25_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI4RUQ_16_LC_16_25_3  (
            .in0(N__40954),
            .in1(N__40942),
            .in2(_gnd_net_),
            .in3(N__45688),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI4RUQZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIICHM1_2_LC_16_26_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIICHM1_2_LC_16_26_4 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIICHM1_2_LC_16_26_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIICHM1_2_LC_16_26_4  (
            .in0(N__40930),
            .in1(N__40924),
            .in2(_gnd_net_),
            .in3(N__50173),
            .lcout(),
            .ltout(iQ_RNIICHM1_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.dat_o_i_0_a2_22_LC_16_26_5 .C_ON=1'b0;
    defparam \u0.dat_o_i_0_a2_22_LC_16_26_5 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_i_0_a2_22_LC_16_26_5 .LUT_INIT=16'b0010001000001010;
    LogicCell40 \u0.dat_o_i_0_a2_22_LC_16_26_5  (
            .in0(N__50369),
            .in1(N__40906),
            .in2(N__40900),
            .in3(N__48939),
            .lcout(\u0.N_1719 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIUKDM1_2_LC_16_26_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIUKDM1_2_LC_16_26_6 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIUKDM1_2_LC_16_26_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIUKDM1_2_LC_16_26_6  (
            .in0(N__40891),
            .in1(N__41746),
            .in2(_gnd_net_),
            .in3(N__50174),
            .lcout(iQ_RNIUKDM1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__16_LC_16_27_0 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__16_LC_16_27_0 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__16_LC_16_27_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__16_LC_16_27_0  (
            .in0(N__42943),
            .in1(N__41731),
            .in2(_gnd_net_),
            .in3(N__41627),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54327),
            .ce(N__41298),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__0_LC_16_27_1 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__0_LC_16_27_1 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__0_LC_16_27_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__0_LC_16_27_1  (
            .in0(N__41730),
            .in1(N__41626),
            .in2(_gnd_net_),
            .in3(N__42945),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54327),
            .ce(N__41298),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__1_LC_16_27_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__1_LC_16_27_2 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__1_LC_16_27_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__1_LC_16_27_2  (
            .in0(N__42944),
            .in1(N__41519),
            .in2(_gnd_net_),
            .in3(N__41410),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54327),
            .ce(N__41298),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__17_LC_16_27_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__17_LC_16_27_3 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__17_LC_16_27_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__17_LC_16_27_3  (
            .in0(N__41518),
            .in1(N__41409),
            .in2(_gnd_net_),
            .in3(N__42946),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54327),
            .ce(N__41298),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__11_LC_16_27_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__11_LC_16_27_4 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__11_LC_16_27_4 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__11_LC_16_27_4  (
            .in0(N__42942),
            .in1(_gnd_net_),
            .in2(N__43141),
            .in3(N__43229),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54327),
            .ce(N__41298),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__27_LC_16_27_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__27_LC_16_27_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__27_LC_16_27_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__27_LC_16_27_5  (
            .in0(N__43230),
            .in1(N__43134),
            .in2(_gnd_net_),
            .in3(N__42947),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram6_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54327),
            .ce(N__41298),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIJBE71_27_LC_16_27_7 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIJBE71_27_LC_16_27_7 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIJBE71_27_LC_16_27_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIJBE71_27_LC_16_27_7  (
            .in0(N__41203),
            .in1(N__41191),
            .in2(_gnd_net_),
            .in3(N__50175),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIJBE71Z0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev0_Tm_RNI31DS1_0_LC_16_28_0 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Tm_RNI31DS1_0_LC_16_28_0 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev0_Tm_RNI31DS1_0_LC_16_28_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \u0.DMA_dev0_Tm_RNI31DS1_0_LC_16_28_0  (
            .in0(N__48578),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41173),
            .lcout(),
            .ltout(\u0.N_1938_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev0_Tm_RNIF52SI_0_LC_16_28_1 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Tm_RNIF52SI_0_LC_16_28_1 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev0_Tm_RNIF52SI_0_LC_16_28_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \u0.DMA_dev0_Tm_RNIF52SI_0_LC_16_28_1  (
            .in0(N__43312),
            .in1(N__43423),
            .in2(N__43408),
            .in3(N__43261),
            .lcout(wb_dat_o_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.q_0_LC_16_28_2 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.q_0_LC_16_28_2 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.q_0_LC_16_28_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.PIO_control.PIO_access_control.q_0_LC_16_28_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43387),
            .lcout(PIOq_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54331),
            .ce(N__45927),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI2KNK1_2_LC_16_28_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI2KNK1_2_LC_16_28_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI2KNK1_2_LC_16_28_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI2KNK1_2_LC_16_28_3  (
            .in0(N__43342),
            .in1(N__50194),
            .in2(_gnd_net_),
            .in3(N__43330),
            .lcout(),
            .ltout(iQ_RNI2KNK1_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.dat_o_0_0_a2_0_0_LC_16_28_4 .C_ON=1'b0;
    defparam \u0.dat_o_0_0_a2_0_0_LC_16_28_4 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_0_0_a2_0_0_LC_16_28_4 .LUT_INIT=16'b1100100001000000;
    LogicCell40 \u0.dat_o_0_0_a2_0_0_LC_16_28_4  (
            .in0(N__48967),
            .in1(N__47228),
            .in2(N__43315),
            .in3(N__43243),
            .lcout(\u0.N_1937 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.CtrlReg_RNIAALH2_0_LC_16_28_5 .C_ON=1'b0;
    defparam \u0.CtrlReg_RNIAALH2_0_LC_16_28_5 .SEQ_MODE=4'b0000;
    defparam \u0.CtrlReg_RNIAALH2_0_LC_16_28_5 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \u0.CtrlReg_RNIAALH2_0_LC_16_28_5  (
            .in0(N__48325),
            .in1(N__43306),
            .in2(N__47497),
            .in3(N__43300),
            .lcout(\u0.dat_o_0_0_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI87OD1_0_LC_16_28_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI87OD1_0_LC_16_28_6 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI87OD1_0_LC_16_28_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNI87OD1_0_LC_16_28_6  (
            .in0(N__50193),
            .in1(N__43255),
            .in2(_gnd_net_),
            .in3(N__43249),
            .lcout(mem_mem_ram6__RNI87OD1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__27_LC_16_29_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__27_LC_16_29_5 .SEQ_MODE=4'b1000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__27_LC_16_29_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram4__27_LC_16_29_5  (
            .in0(N__43231),
            .in1(N__43135),
            .in2(_gnd_net_),
            .in3(N__42965),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_ram4_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54333),
            .ce(N__41859),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI2KD53_3_LC_16_31_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI2KD53_3_LC_16_31_6 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI2KD53_3_LC_16_31_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI2KD53_3_LC_16_31_6  (
            .in0(N__48985),
            .in1(N__41764),
            .in2(_gnd_net_),
            .in3(N__41755),
            .lcout(DMAq_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.register_block_gen_PIO_cmdport_reg_un6_sel_pio_cmdport_i_0_LC_17_16_2 .C_ON=1'b0;
    defparam \u0.register_block_gen_PIO_cmdport_reg_un6_sel_pio_cmdport_i_0_LC_17_16_2 .SEQ_MODE=4'b0000;
    defparam \u0.register_block_gen_PIO_cmdport_reg_un6_sel_pio_cmdport_i_0_LC_17_16_2 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \u0.register_block_gen_PIO_cmdport_reg_un6_sel_pio_cmdport_i_0_LC_17_16_2  (
            .in0(N__51365),
            .in1(N__50864),
            .in2(_gnd_net_),
            .in3(N__48085),
            .lcout(N_448),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport1_T2_RNI9BO24_3_LC_17_18_0 .C_ON=1'b0;
    defparam \u0.PIO_dport1_T2_RNI9BO24_3_LC_17_18_0 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport1_T2_RNI9BO24_3_LC_17_18_0 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \u0.PIO_dport1_T2_RNI9BO24_3_LC_17_18_0  (
            .in0(N__43780),
            .in1(N__46908),
            .in2(N__48587),
            .in3(N__43765),
            .lcout(),
            .ltout(\u0.dat_o_0_0_0_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev1_Td_RNIEEFKG_3_LC_17_18_1 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Td_RNIEEFKG_3_LC_17_18_1 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev1_Td_RNIEEFKG_3_LC_17_18_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \u0.DMA_dev1_Td_RNIEEFKG_3_LC_17_18_1  (
            .in0(N__43567),
            .in1(N__46354),
            .in2(N__43741),
            .in3(N__43738),
            .lcout(wb_dat_o_c_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.CtrlReg_11_LC_17_18_2 .C_ON=1'b0;
    defparam \u0.CtrlReg_11_LC_17_18_2 .SEQ_MODE=4'b1010;
    defparam \u0.CtrlReg_11_LC_17_18_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.CtrlReg_11_LC_17_18_2  (
            .in0(N__51610),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43700),
            .lcout(\u0.CtrlRegZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54251),
            .ce(N__53643),
            .sr(N__53388));
    defparam \u0.CtrlReg_RNIJI6Q3_11_LC_17_18_5 .C_ON=1'b0;
    defparam \u0.CtrlReg_RNIJI6Q3_11_LC_17_18_5 .SEQ_MODE=4'b0000;
    defparam \u0.CtrlReg_RNIJI6Q3_11_LC_17_18_5 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \u0.CtrlReg_RNIJI6Q3_11_LC_17_18_5  (
            .in0(N__48311),
            .in1(N__43591),
            .in2(N__48106),
            .in3(N__43585),
            .lcout(\u0.dat_o_0_0_2_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev1_Td_RNI8F7N3_2_LC_17_19_1 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Td_RNI8F7N3_2_LC_17_19_1 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev1_Td_RNI8F7N3_2_LC_17_19_1 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \u0.DMA_dev1_Td_RNI8F7N3_2_LC_17_19_1  (
            .in0(N__46907),
            .in1(N__54629),
            .in2(N__43561),
            .in3(N__43540),
            .lcout(\u0.dat_o_i_i_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev1_Td_RNIFHOI3_6_LC_17_19_3 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Td_RNIFHOI3_6_LC_17_19_3 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev1_Td_RNIFHOI3_6_LC_17_19_3 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \u0.DMA_dev1_Td_RNIFHOI3_6_LC_17_19_3  (
            .in0(N__50663),
            .in1(N__54630),
            .in2(N__43510),
            .in3(N__43486),
            .lcout(),
            .ltout(\u0.dat_o_0_0_3_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev1_Td_RNIOPGKG_6_LC_17_19_4 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Td_RNIOPGKG_6_LC_17_19_4 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev1_Td_RNIOPGKG_6_LC_17_19_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \u0.DMA_dev1_Td_RNIOPGKG_6_LC_17_19_4  (
            .in0(N__43933),
            .in1(N__44071),
            .in2(N__43468),
            .in3(N__43429),
            .lcout(wb_dat_o_c_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.dat_o_0_0_1_14_LC_17_19_5 .C_ON=1'b0;
    defparam \u0.dat_o_0_0_1_14_LC_17_19_5 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_0_0_1_14_LC_17_19_5 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \u0.dat_o_0_0_1_14_LC_17_19_5  (
            .in0(N__47405),
            .in1(N__43894),
            .in2(N__47224),
            .in3(N__43450),
            .lcout(\u0.dat_o_0_0_1Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport1_T2_RNIFHO24_6_LC_17_20_0 .C_ON=1'b0;
    defparam \u0.PIO_dport1_T2_RNIFHO24_6_LC_17_20_0 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport1_T2_RNIFHO24_6_LC_17_20_0 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \u0.PIO_dport1_T2_RNIFHO24_6_LC_17_20_0  (
            .in0(N__44121),
            .in1(N__46865),
            .in2(N__44095),
            .in3(N__48469),
            .lcout(\u0.dat_o_0_0_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.CtrlReg_14_LC_17_20_2 .C_ON=1'b0;
    defparam \u0.CtrlReg_14_LC_17_20_2 .SEQ_MODE=4'b1010;
    defparam \u0.CtrlReg_14_LC_17_20_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.CtrlReg_14_LC_17_20_2  (
            .in0(N__51613),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44065),
            .lcout(\u0.CtrlRegZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54275),
            .ce(N__53615),
            .sr(N__53398));
    defparam \u0.CtrlReg_RNIPO6Q3_14_LC_17_20_3 .C_ON=1'b0;
    defparam \u0.CtrlReg_RNIPO6Q3_14_LC_17_20_3 .SEQ_MODE=4'b0000;
    defparam \u0.CtrlReg_RNIPO6Q3_14_LC_17_20_3 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \u0.CtrlReg_RNIPO6Q3_14_LC_17_20_3  (
            .in0(N__43954),
            .in1(N__48018),
            .in2(N__48254),
            .in3(N__43948),
            .lcout(\u0.dat_o_0_0_2_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIGKV43_3_LC_17_20_5 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIGKV43_3_LC_17_20_5 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIGKV43_3_LC_17_20_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNIGKV43_3_LC_17_20_5  (
            .in0(N__43927),
            .in1(N__43912),
            .in2(_gnd_net_),
            .in3(N__48958),
            .lcout(DMAq_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev1_Teoc_RNINVRS6_5_LC_17_21_0 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Teoc_RNINVRS6_5_LC_17_21_0 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev1_Teoc_RNINVRS6_5_LC_17_21_0 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \u0.DMA_dev1_Teoc_RNINVRS6_5_LC_17_21_0  (
            .in0(N__54587),
            .in1(N__46535),
            .in2(N__43887),
            .in3(N__43825),
            .lcout(\u0.dat_o_i_i_4_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.register_block_gen_PIO_cmdport_reg_un6_sel_pio_cmdport_i_0_a2_0_LC_17_21_1 .C_ON=1'b0;
    defparam \u0.register_block_gen_PIO_cmdport_reg_un6_sel_pio_cmdport_i_0_a2_0_LC_17_21_1 .SEQ_MODE=4'b0000;
    defparam \u0.register_block_gen_PIO_cmdport_reg_un6_sel_pio_cmdport_i_0_a2_0_LC_17_21_1 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \u0.register_block_gen_PIO_cmdport_reg_un6_sel_pio_cmdport_i_0_a2_0_LC_17_21_1  (
            .in0(N__46416),
            .in1(N__47720),
            .in2(N__53080),
            .in3(N__50577),
            .lcout(\u0.N_2123 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev0_Teoc_RNIS54G3_5_LC_17_21_2 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Teoc_RNIS54G3_5_LC_17_21_2 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev0_Teoc_RNIS54G3_5_LC_17_21_2 .LUT_INIT=16'b1101110011001100;
    LogicCell40 \u0.DMA_dev0_Teoc_RNIS54G3_5_LC_17_21_2  (
            .in0(N__47715),
            .in1(N__46429),
            .in2(N__43855),
            .in3(N__46730),
            .lcout(\u0.dat_o_i_i_0_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport0_Teoc_RNII5UK_5_LC_17_21_3 .C_ON=1'b0;
    defparam \u0.PIO_dport0_Teoc_RNII5UK_5_LC_17_21_3 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport0_Teoc_RNII5UK_5_LC_17_21_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.PIO_dport0_Teoc_RNII5UK_5_LC_17_21_3  (
            .in0(N__53069),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43818),
            .lcout(),
            .ltout(\u0.dat_o_i_i_a2_0_0_29_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport1_Teoc_RNIUGQA3_5_LC_17_21_4 .C_ON=1'b0;
    defparam \u0.PIO_dport1_Teoc_RNIUGQA3_5_LC_17_21_4 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport1_Teoc_RNIUGQA3_5_LC_17_21_4 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \u0.PIO_dport1_Teoc_RNIUGQA3_5_LC_17_21_4  (
            .in0(N__46864),
            .in1(N__46731),
            .in2(N__44419),
            .in3(N__44416),
            .lcout(),
            .ltout(\u0.dat_o_i_i_2_29_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport1_Teoc_RNI269OG_5_LC_17_21_5 .C_ON=1'b0;
    defparam \u0.PIO_dport1_Teoc_RNI269OG_5_LC_17_21_5 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport1_Teoc_RNI269OG_5_LC_17_21_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \u0.PIO_dport1_Teoc_RNI269OG_5_LC_17_21_5  (
            .in0(N__44386),
            .in1(N__44371),
            .in2(N__44365),
            .in3(N__46060),
            .lcout(N_273),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.dat_o_0_0_a2_7_1_LC_17_21_6 .C_ON=1'b0;
    defparam \u0.dat_o_0_0_a2_7_1_LC_17_21_6 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_0_0_a2_7_1_LC_17_21_6 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \u0.dat_o_0_0_a2_7_1_LC_17_21_6  (
            .in0(N__50575),
            .in1(N__46414),
            .in2(N__47731),
            .in3(N__53070),
            .lcout(\u0.N_2122 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.dat_o_0_0_a2_8_1_LC_17_21_7 .C_ON=1'b0;
    defparam \u0.dat_o_0_0_a2_8_1_LC_17_21_7 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_0_0_a2_8_1_LC_17_21_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \u0.dat_o_0_0_a2_8_1_LC_17_21_7  (
            .in0(N__46415),
            .in1(N__47719),
            .in2(N__53079),
            .in3(N__50576),
            .lcout(\u0.N_2124 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev1_Teoc_RNIGK8P1_2_LC_17_22_0 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Teoc_RNIGK8P1_2_LC_17_22_0 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev1_Teoc_RNIGK8P1_2_LC_17_22_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \u0.DMA_dev1_Teoc_RNIGK8P1_2_LC_17_22_0  (
            .in0(_gnd_net_),
            .in1(N__54589),
            .in2(_gnd_net_),
            .in3(N__44341),
            .lcout(),
            .ltout(\u0.N_1675_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport0_Teoc_RNIS0IJ7_2_LC_17_22_1 .C_ON=1'b0;
    defparam \u0.PIO_dport0_Teoc_RNIS0IJ7_2_LC_17_22_1 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport0_Teoc_RNIS0IJ7_2_LC_17_22_1 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \u0.PIO_dport0_Teoc_RNIS0IJ7_2_LC_17_22_1  (
            .in0(N__50702),
            .in1(N__46990),
            .in2(N__44308),
            .in3(N__44305),
            .lcout(),
            .ltout(\u0.dat_o_i_i_4_26_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport1_Teoc_RNI80L3G_2_LC_17_22_2 .C_ON=1'b0;
    defparam \u0.PIO_dport1_Teoc_RNI80L3G_2_LC_17_22_2 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport1_Teoc_RNI80L3G_2_LC_17_22_2 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \u0.PIO_dport1_Teoc_RNI80L3G_2_LC_17_22_2  (
            .in0(N__46866),
            .in1(N__44128),
            .in2(N__44284),
            .in3(N__44281),
            .lcout(N_267),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.CtrlReg_26_LC_17_22_3 .C_ON=1'b0;
    defparam \u0.CtrlReg_26_LC_17_22_3 .SEQ_MODE=4'b1010;
    defparam \u0.CtrlReg_26_LC_17_22_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.CtrlReg_26_LC_17_22_3  (
            .in0(N__51436),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44237),
            .lcout(\u0.CtrlRegZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54295),
            .ce(N__53614),
            .sr(N__53405));
    defparam \u0.DMA_dev0_Teoc_RNISV2P6_2_LC_17_22_5 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Teoc_RNISV2P6_2_LC_17_22_5 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev0_Teoc_RNISV2P6_2_LC_17_22_5 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \u0.DMA_dev0_Teoc_RNISV2P6_2_LC_17_22_5  (
            .in0(N__48468),
            .in1(N__44161),
            .in2(N__44149),
            .in3(N__47070),
            .lcout(\u0.dat_o_i_i_0_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev0_Tm_RNIDVGR3_1_LC_17_23_0 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Tm_RNIDVGR3_1_LC_17_23_0 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev0_Tm_RNIDVGR3_1_LC_17_23_0 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \u0.DMA_dev0_Tm_RNIDVGR3_1_LC_17_23_0  (
            .in0(N__48549),
            .in1(N__46904),
            .in2(N__44704),
            .in3(N__44674),
            .lcout(),
            .ltout(\u0.dat_o_0_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_cmdport_T1_RNIQRTSG_1_LC_17_23_1 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_T1_RNIQRTSG_1_LC_17_23_1 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_cmdport_T1_RNIQRTSG_1_LC_17_23_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \u0.PIO_cmdport_T1_RNIQRTSG_1_LC_17_23_1  (
            .in0(N__44647),
            .in1(N__44632),
            .in2(N__44620),
            .in3(N__47026),
            .lcout(wb_dat_o_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI6ONK1_2_LC_17_23_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI6ONK1_2_LC_17_23_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI6ONK1_2_LC_17_23_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI6ONK1_2_LC_17_23_3  (
            .in0(N__50179),
            .in1(N__44602),
            .in2(_gnd_net_),
            .in3(N__44587),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI6ONK1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.q_1_LC_17_23_5 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.q_1_LC_17_23_5 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.q_1_LC_17_23_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \u1.PIO_control.PIO_access_control.q_1_LC_17_23_5  (
            .in0(N__44572),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(PIOq_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54305),
            .ce(N__45925),
            .sr(_gnd_net_));
    defparam \u0.CtrlReg_RNIQQLH2_8_LC_17_24_0 .C_ON=1'b0;
    defparam \u0.CtrlReg_RNIQQLH2_8_LC_17_24_0 .SEQ_MODE=4'b0000;
    defparam \u0.CtrlReg_RNIQQLH2_8_LC_17_24_0 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \u0.CtrlReg_RNIQQLH2_8_LC_17_24_0  (
            .in0(N__44452),
            .in1(N__48289),
            .in2(N__47453),
            .in3(N__54358),
            .lcout(),
            .ltout(\u0.dat_o_0_0_2_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev0_Td_RNI9VQMI_0_LC_17_24_1 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Td_RNI9VQMI_0_LC_17_24_1 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev0_Td_RNI9VQMI_0_LC_17_24_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \u0.DMA_dev0_Td_RNI9VQMI_0_LC_17_24_1  (
            .in0(N__44533),
            .in1(N__44521),
            .in2(N__44506),
            .in3(N__45982),
            .lcout(wb_dat_o_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.q_8_LC_17_24_2 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.q_8_LC_17_24_2 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.q_8_LC_17_24_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \u1.PIO_control.PIO_access_control.q_8_LC_17_24_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44482),
            .lcout(PIOq_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54314),
            .ce(N__45937),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI2LOK1_2_LC_17_24_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI2LOK1_2_LC_17_24_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI2LOK1_2_LC_17_24_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI2LOK1_2_LC_17_24_3  (
            .in0(N__44446),
            .in1(N__44437),
            .in2(_gnd_net_),
            .in3(N__50206),
            .lcout(),
            .ltout(iQ_RNI2LOK1_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.dat_o_0_0_a2_0_8_LC_17_24_4 .C_ON=1'b0;
    defparam \u0.dat_o_0_0_a2_0_8_LC_17_24_4 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_0_0_a2_0_8_LC_17_24_4 .LUT_INIT=16'b1101100000000000;
    LogicCell40 \u0.dat_o_0_0_a2_0_8_LC_17_24_4  (
            .in0(N__48986),
            .in1(N__45991),
            .in2(N__45985),
            .in3(N__47145),
            .lcout(\u0.N_1735 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.PIO_control.PIO_access_control.q_9_LC_17_25_2 .C_ON=1'b0;
    defparam \u1.PIO_control.PIO_access_control.q_9_LC_17_25_2 .SEQ_MODE=4'b1000;
    defparam \u1.PIO_control.PIO_access_control.q_9_LC_17_25_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \u1.PIO_control.PIO_access_control.q_9_LC_17_25_2  (
            .in0(N__45976),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(PIOq_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54322),
            .ce(N__45909),
            .sr(_gnd_net_));
    defparam \u0.CtrlReg_RNI59KU1_17_LC_17_26_0 .C_ON=1'b0;
    defparam \u0.CtrlReg_RNI59KU1_17_LC_17_26_0 .SEQ_MODE=4'b0000;
    defparam \u0.CtrlReg_RNI59KU1_17_LC_17_26_0 .LUT_INIT=16'b0100010011110100;
    LogicCell40 \u0.CtrlReg_RNI59KU1_17_LC_17_26_0  (
            .in0(N__45055),
            .in1(N__45046),
            .in2(N__44936),
            .in3(N__45754),
            .lcout(\u0.dat_o_0_a2_i_2_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI6TUQ_17_LC_17_26_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI6TUQ_17_LC_17_26_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI6TUQ_17_LC_17_26_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI6TUQ_17_LC_17_26_3  (
            .in0(N__45727),
            .in1(N__45715),
            .in2(_gnd_net_),
            .in3(N__45702),
            .lcout(\u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram0__RNI6TUQZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.CtrlReg_17_LC_17_26_5 .C_ON=1'b0;
    defparam \u0.CtrlReg_17_LC_17_26_5 .SEQ_MODE=4'b1010;
    defparam \u0.CtrlReg_17_LC_17_26_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.CtrlReg_17_LC_17_26_5  (
            .in0(N__51683),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45133),
            .lcout(\u0.CtrlRegZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54328),
            .ce(N__53575),
            .sr(N__53411));
    defparam \u0.CtrlReg_RNI8DLU1_23_LC_17_27_0 .C_ON=1'b0;
    defparam \u0.CtrlReg_RNI8DLU1_23_LC_17_27_0 .SEQ_MODE=4'b0000;
    defparam \u0.CtrlReg_RNI8DLU1_23_LC_17_27_0 .LUT_INIT=16'b0010111100100010;
    LogicCell40 \u0.CtrlReg_RNI8DLU1_23_LC_17_27_0  (
            .in0(N__45047),
            .in1(N__44773),
            .in2(N__44965),
            .in3(N__44927),
            .lcout(\u0.dat_o_i_0_0_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.CtrlReg_23_LC_17_27_3 .C_ON=1'b0;
    defparam \u0.CtrlReg_23_LC_17_27_3 .SEQ_MODE=4'b1010;
    defparam \u0.CtrlReg_23_LC_17_27_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \u0.CtrlReg_23_LC_17_27_3  (
            .in0(_gnd_net_),
            .in1(N__44831),
            .in2(_gnd_net_),
            .in3(N__51684),
            .lcout(\u0.CtrlRegZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54332),
            .ce(N__53565),
            .sr(N__53412));
    defparam \u0.dat_o_i_0_a2_23_LC_17_27_6 .C_ON=1'b0;
    defparam \u0.dat_o_i_0_a2_23_LC_17_27_6 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_i_0_a2_23_LC_17_27_6 .LUT_INIT=16'b0100010000001100;
    LogicCell40 \u0.dat_o_i_0_a2_23_LC_17_27_6  (
            .in0(N__44767),
            .in1(N__50457),
            .in2(N__44755),
            .in3(N__48975),
            .lcout(\u0.N_1714 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.CtrlReg_RNISSLH2_9_LC_17_28_0 .C_ON=1'b0;
    defparam \u0.CtrlReg_RNISSLH2_9_LC_17_28_0 .SEQ_MODE=4'b0000;
    defparam \u0.CtrlReg_RNISSLH2_9_LC_17_28_0 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \u0.CtrlReg_RNISSLH2_9_LC_17_28_0  (
            .in0(N__44740),
            .in1(N__44713),
            .in2(N__48324),
            .in3(N__47423),
            .lcout(\u0.dat_o_0_0_2_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.dat_o_0_0_1_11_LC_17_28_2 .C_ON=1'b0;
    defparam \u0.dat_o_0_0_1_11_LC_17_28_2 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_0_0_1_11_LC_17_28_2 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \u0.dat_o_0_0_1_11_LC_17_28_2  (
            .in0(N__47483),
            .in1(N__47196),
            .in2(N__46384),
            .in3(N__46369),
            .lcout(\u0.dat_o_0_0_1Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI6POK1_2_LC_17_28_3 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI6POK1_2_LC_17_28_3 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI6POK1_2_LC_17_28_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI6POK1_2_LC_17_28_3  (
            .in0(N__46342),
            .in1(N__46327),
            .in2(_gnd_net_),
            .in3(N__50207),
            .lcout(),
            .ltout(iQ_RNI6POK1_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.dat_o_0_0_a2_0_9_LC_17_28_4 .C_ON=1'b0;
    defparam \u0.dat_o_0_0_a2_0_9_LC_17_28_4 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_0_0_a2_0_9_LC_17_28_4 .LUT_INIT=16'b1000100011000000;
    LogicCell40 \u0.dat_o_0_0_a2_0_9_LC_17_28_4  (
            .in0(N__46315),
            .in1(N__47197),
            .in2(N__46306),
            .in3(N__48968),
            .lcout(\u0.N_1650 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport0_T1_5_LC_18_16_5 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T1_5_LC_18_16_5 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport0_T1_5_LC_18_16_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \u0.PIO_dport0_T1_5_LC_18_16_5  (
            .in0(_gnd_net_),
            .in1(N__51202),
            .in2(_gnd_net_),
            .in3(N__46265),
            .lcout(PIO_dport0_T1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54263),
            .ce(N__49375),
            .sr(N__53379));
    defparam \u0.CtrlReg_28_LC_18_18_6 .C_ON=1'b0;
    defparam \u0.CtrlReg_28_LC_18_18_6 .SEQ_MODE=4'b1010;
    defparam \u0.CtrlReg_28_LC_18_18_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \u0.CtrlReg_28_LC_18_18_6  (
            .in0(N__51203),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46111),
            .lcout(\u0.CtrlRegZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54264),
            .ce(N__53644),
            .sr(N__53392));
    defparam \u0.CtrlReg_RNIBCRN1_29_LC_18_19_0 .C_ON=1'b0;
    defparam \u0.CtrlReg_RNIBCRN1_29_LC_18_19_0 .SEQ_MODE=4'b0000;
    defparam \u0.CtrlReg_RNIBCRN1_29_LC_18_19_0 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \u0.CtrlReg_RNIBCRN1_29_LC_18_19_0  (
            .in0(N__53019),
            .in1(N__49255),
            .in2(N__46423),
            .in3(N__47634),
            .lcout(\u0.N_1695 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport0_T2_RNIHK559_1_LC_18_19_3 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T2_RNIHK559_1_LC_18_19_3 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport0_T2_RNIHK559_1_LC_18_19_3 .LUT_INIT=16'b1111111011101110;
    LogicCell40 \u0.PIO_dport0_T2_RNIHK559_1_LC_18_19_3  (
            .in0(N__46051),
            .in1(N__46036),
            .in2(N__50676),
            .in3(N__46021),
            .lcout(\u0.dat_o_0_0_6_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.CtrlReg_RNIABRN1_28_LC_18_20_0 .C_ON=1'b0;
    defparam \u0.CtrlReg_RNIABRN1_28_LC_18_20_0 .SEQ_MODE=4'b0000;
    defparam \u0.CtrlReg_RNIABRN1_28_LC_18_20_0 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \u0.CtrlReg_RNIABRN1_28_LC_18_20_0  (
            .in0(N__46413),
            .in1(N__46000),
            .in2(N__53056),
            .in3(N__47701),
            .lcout(),
            .ltout(\u0.N_1688_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport0_Teoc_RNIKOLB3_4_LC_18_20_1 .C_ON=1'b0;
    defparam \u0.PIO_dport0_Teoc_RNIKOLB3_4_LC_18_20_1 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport0_Teoc_RNIKOLB3_4_LC_18_20_1 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \u0.PIO_dport0_Teoc_RNIKOLB3_4_LC_18_20_1  (
            .in0(N__46627),
            .in1(N__46732),
            .in2(N__46606),
            .in3(N__53023),
            .lcout(\u0.dat_o_i_i_2_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.dat_o_i_i_a3_28_LC_18_20_4 .C_ON=1'b0;
    defparam \u0.dat_o_i_i_a3_28_LC_18_20_4 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_i_i_a3_28_LC_18_20_4 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \u0.dat_o_i_i_a3_28_LC_18_20_4  (
            .in0(N__46734),
            .in1(_gnd_net_),
            .in2(N__53057),
            .in3(N__47703),
            .lcout(\u0.N_2137 ),
            .ltout(\u0.N_2137_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport1_Teoc_RNITSOT6_4_LC_18_20_5 .C_ON=1'b0;
    defparam \u0.PIO_dport1_Teoc_RNITSOT6_4_LC_18_20_5 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport1_Teoc_RNITSOT6_4_LC_18_20_5 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \u0.PIO_dport1_Teoc_RNITSOT6_4_LC_18_20_5  (
            .in0(N__46519),
            .in1(N__46495),
            .in2(N__46480),
            .in3(N__46890),
            .lcout(),
            .ltout(\u0.dat_o_i_i_4_28_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport1_Teoc_RNILO8OG_4_LC_18_20_6 .C_ON=1'b0;
    defparam \u0.PIO_dport1_Teoc_RNILO8OG_4_LC_18_20_6 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport1_Teoc_RNILO8OG_4_LC_18_20_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \u0.PIO_dport1_Teoc_RNILO8OG_4_LC_18_20_6  (
            .in0(N__46675),
            .in1(N__46477),
            .in2(N__46471),
            .in3(N__46468),
            .lcout(N_271),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.dat_o_0_0_a2_10_1_LC_18_20_7 .C_ON=1'b0;
    defparam \u0.dat_o_0_0_a2_10_1_LC_18_20_7 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_0_0_a2_10_1_LC_18_20_7 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \u0.dat_o_0_0_a2_10_1_LC_18_20_7  (
            .in0(N__47702),
            .in1(N__46733),
            .in2(_gnd_net_),
            .in3(N__53024),
            .lcout(\u0.N_2129 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_cmdport_Teoc_RNII31Q1_5_LC_18_21_0 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_Teoc_RNII31Q1_5_LC_18_21_0 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_cmdport_Teoc_RNII31Q1_5_LC_18_21_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \u0.PIO_cmdport_Teoc_RNII31Q1_5_LC_18_21_0  (
            .in0(_gnd_net_),
            .in1(N__48020),
            .in2(_gnd_net_),
            .in3(N__49716),
            .lcout(\u0.N_1699 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.dat_o_0_0_a2_9_1_LC_18_21_1 .C_ON=1'b0;
    defparam \u0.dat_o_0_0_a2_9_1_LC_18_21_1 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_0_0_a2_9_1_LC_18_21_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \u0.dat_o_0_0_a2_9_1_LC_18_21_1  (
            .in0(N__47705),
            .in1(N__46412),
            .in2(N__53077),
            .in3(N__50558),
            .lcout(\u0.N_2128 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.dat_o_i_i_a2_6_28_LC_18_21_2 .C_ON=1'b0;
    defparam \u0.dat_o_i_i_a2_6_28_LC_18_21_2 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_i_i_a2_6_28_LC_18_21_2 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \u0.dat_o_i_i_a2_6_28_LC_18_21_2  (
            .in0(N__50409),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47373),
            .lcout(\u0.N_2095 ),
            .ltout(\u0.N_2095_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.dat_o_0_0_a2_11_1_LC_18_21_3 .C_ON=1'b0;
    defparam \u0.dat_o_0_0_a2_11_1_LC_18_21_3 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_0_0_a2_11_1_LC_18_21_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \u0.dat_o_0_0_a2_11_1_LC_18_21_3  (
            .in0(N__47704),
            .in1(N__53058),
            .in2(N__46387),
            .in3(N__50557),
            .lcout(\u0.N_2130 ),
            .ltout(\u0.N_2130_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.CtrlReg_RNITK5S3_26_LC_18_21_4 .C_ON=1'b0;
    defparam \u0.CtrlReg_RNITK5S3_26_LC_18_21_4 .SEQ_MODE=4'b0000;
    defparam \u0.CtrlReg_RNITK5S3_26_LC_18_21_4 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \u0.CtrlReg_RNITK5S3_26_LC_18_21_4  (
            .in0(N__47020),
            .in1(N__48019),
            .in2(N__46999),
            .in3(N__46996),
            .lcout(\u0.dat_o_i_i_1_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.dat_o_0_a2_i_o2_0_16_LC_18_21_5 .C_ON=1'b0;
    defparam \u0.dat_o_0_a2_i_o2_0_16_LC_18_21_5 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_0_a2_i_o2_0_16_LC_18_21_5 .LUT_INIT=16'b0010110011101100;
    LogicCell40 \u0.dat_o_0_a2_i_o2_0_16_LC_18_21_5  (
            .in0(N__47706),
            .in1(N__50408),
            .in2(N__53078),
            .in3(N__50559),
            .lcout(\u0.dat_o_0_a2_i_o2_0Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.dat_o_i_i_a2_7_28_LC_18_21_6 .C_ON=1'b0;
    defparam \u0.dat_o_i_i_a2_7_28_LC_18_21_6 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_i_i_a2_7_28_LC_18_21_6 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \u0.dat_o_i_i_a2_7_28_LC_18_21_6  (
            .in0(N__50561),
            .in1(_gnd_net_),
            .in2(N__50442),
            .in3(N__47374),
            .lcout(\u0.N_2104 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.dat_o_0_a2_i_o2_1_16_LC_18_21_7 .C_ON=1'b0;
    defparam \u0.dat_o_0_a2_i_o2_1_16_LC_18_21_7 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_0_a2_i_o2_1_16_LC_18_21_7 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \u0.dat_o_0_a2_i_o2_1_16_LC_18_21_7  (
            .in0(N__53065),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50560),
            .lcout(N_1321),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport1_Teoc_RNIK30N1_6_LC_18_22_2 .C_ON=1'b0;
    defparam \u0.PIO_dport1_Teoc_RNIK30N1_6_LC_18_22_2 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport1_Teoc_RNIK30N1_6_LC_18_22_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \u0.PIO_dport1_Teoc_RNIK30N1_6_LC_18_22_2  (
            .in0(N__46889),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46797),
            .lcout(),
            .ltout(\u0.N_1703_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport0_Teoc_RNI3KAH7_6_LC_18_22_3 .C_ON=1'b0;
    defparam \u0.PIO_dport0_Teoc_RNI3KAH7_6_LC_18_22_3 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport0_Teoc_RNI3KAH7_6_LC_18_22_3 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \u0.PIO_dport0_Teoc_RNI3KAH7_6_LC_18_22_3  (
            .in0(N__46771),
            .in1(N__47938),
            .in2(N__46744),
            .in3(N__50677),
            .lcout(\u0.dat_o_i_i_4_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev0_Teoc_RNI913M1_4_LC_18_22_5 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Teoc_RNI913M1_4_LC_18_22_5 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev0_Teoc_RNI913M1_4_LC_18_22_5 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \u0.DMA_dev0_Teoc_RNI913M1_4_LC_18_22_5  (
            .in0(N__47707),
            .in1(N__46729),
            .in2(_gnd_net_),
            .in3(N__46701),
            .lcout(\u0.N_1686 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.valid_3_0_0_a2_1_LC_18_22_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.valid_3_0_0_a2_1_LC_18_22_6 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Txbuf.valid_3_0_0_a2_1_LC_18_22_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Txbuf.valid_3_0_0_a2_1_LC_18_22_6  (
            .in0(N__46666),
            .in1(N__47375),
            .in2(N__50443),
            .in3(N__47708),
            .lcout(N_2119),
            .ltout(N_2119_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev0_Teoc_RNICF2P6_0_LC_18_22_7 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Teoc_RNICF2P6_0_LC_18_22_7 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev0_Teoc_RNICF2P6_0_LC_18_22_7 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \u0.DMA_dev0_Teoc_RNICF2P6_0_LC_18_22_7  (
            .in0(N__48436),
            .in1(N__46660),
            .in2(N__46648),
            .in3(N__46645),
            .lcout(\u0.dat_o_i_i_0_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.CtrlReg_RNISK6S3_30_LC_18_23_0 .C_ON=1'b0;
    defparam \u0.CtrlReg_RNISK6S3_30_LC_18_23_0 .SEQ_MODE=4'b0000;
    defparam \u0.CtrlReg_RNISK6S3_30_LC_18_23_0 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \u0.CtrlReg_RNISK6S3_30_LC_18_23_0  (
            .in0(N__47752),
            .in1(N__48237),
            .in2(N__48132),
            .in3(N__47962),
            .lcout(\u0.dat_o_i_i_1_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev0_Teoc_RNIT69P6_6_LC_18_23_1 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Teoc_RNIT69P6_6_LC_18_23_1 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev0_Teoc_RNIT69P6_6_LC_18_23_1 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \u0.DMA_dev0_Teoc_RNIT69P6_6_LC_18_23_1  (
            .in0(N__47932),
            .in1(N__47908),
            .in2(N__48548),
            .in3(N__47071),
            .lcout(),
            .ltout(\u0.dat_o_i_i_0_30_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev1_Teoc_RNIKJS3G_6_LC_18_23_2 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Teoc_RNIKJS3G_6_LC_18_23_2 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev1_Teoc_RNIKJS3G_6_LC_18_23_2 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \u0.DMA_dev1_Teoc_RNIKJS3G_6_LC_18_23_2  (
            .in0(N__47896),
            .in1(N__54634),
            .in2(N__47887),
            .in3(N__47883),
            .lcout(N_275),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.CtrlReg_30_LC_18_23_4 .C_ON=1'b0;
    defparam \u0.CtrlReg_30_LC_18_23_4 .SEQ_MODE=4'b1010;
    defparam \u0.CtrlReg_30_LC_18_23_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \u0.CtrlReg_30_LC_18_23_4  (
            .in0(_gnd_net_),
            .in1(N__47821),
            .in2(_gnd_net_),
            .in3(N__51212),
            .lcout(\u0.CtrlRegZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54315),
            .ce(N__53606),
            .sr(N__53410));
    defparam \u0.dat_o_0_a2_i_o2_16_LC_18_24_1 .C_ON=1'b0;
    defparam \u0.dat_o_0_a2_i_o2_16_LC_18_24_1 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_0_a2_i_o2_16_LC_18_24_1 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \u0.dat_o_0_a2_i_o2_16_LC_18_24_1  (
            .in0(N__50562),
            .in1(N__47746),
            .in2(N__47416),
            .in3(N__47727),
            .lcout(\u0.N_1374 ),
            .ltout(\u0.N_1374_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport0_T4_RNI9KQO9_7_LC_18_24_2 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T4_RNI9KQO9_7_LC_18_24_2 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport0_T4_RNI9KQO9_7_LC_18_24_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \u0.PIO_dport0_T4_RNI9KQO9_7_LC_18_24_2  (
            .in0(N__47581),
            .in1(N__47569),
            .in2(N__47557),
            .in3(N__49195),
            .lcout(N_332_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI4EN93_3_LC_18_24_4 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI4EN93_3_LC_18_24_4 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI4EN93_3_LC_18_24_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI4EN93_3_LC_18_24_4  (
            .in0(N__47533),
            .in1(N__48987),
            .in2(_gnd_net_),
            .in3(N__47527),
            .lcout(),
            .ltout(DMAq_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.dat_o_0_0_1_1_LC_18_24_5 .C_ON=1'b0;
    defparam \u0.dat_o_0_0_1_1_LC_18_24_5 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_0_0_1_1_LC_18_24_5 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \u0.dat_o_0_0_1_1_LC_18_24_5  (
            .in0(N__47376),
            .in1(N__47144),
            .in2(N__47035),
            .in3(N__47032),
            .lcout(\u0.dat_o_0_0_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport0_T4_RNIQTIO9_2_LC_18_24_6 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T4_RNIQTIO9_2_LC_18_24_6 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport0_T4_RNIQTIO9_2_LC_18_24_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \u0.PIO_dport0_T4_RNIQTIO9_2_LC_18_24_6  (
            .in0(N__49111),
            .in1(N__49102),
            .in2(N__49087),
            .in3(N__49606),
            .lcout(N_325_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.dat_o_0_a2_i_a2_16_LC_18_26_5 .C_ON=1'b0;
    defparam \u0.dat_o_0_a2_i_a2_16_LC_18_26_5 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_0_a2_i_a2_16_LC_18_26_5 .LUT_INIT=16'b0010001000001010;
    LogicCell40 \u0.dat_o_0_a2_i_a2_16_LC_18_26_5  (
            .in0(N__50444),
            .in1(N__49729),
            .in2(N__49054),
            .in3(N__48940),
            .lcout(\u0.N_1549 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI2PDM1_2_LC_18_26_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI2PDM1_2_LC_18_26_6 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI2PDM1_2_LC_18_26_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.rd_ptr_lfsr.iQ_RNI2PDM1_2_LC_18_26_6  (
            .in0(N__50114),
            .in1(N__49042),
            .in2(_gnd_net_),
            .in3(N__49030),
            .lcout(iQ_RNI2PDM1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIG5B71_17_LC_18_27_2 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIG5B71_17_LC_18_27_2 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIG5B71_17_LC_18_27_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNIG5B71_17_LC_18_27_2  (
            .in0(N__50198),
            .in1(N__49024),
            .in2(_gnd_net_),
            .in3(N__49006),
            .lcout(),
            .ltout(mem_mem_ram6__RNIG5B71_17_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.dat_o_0_a2_i_a2_17_LC_18_27_3 .C_ON=1'b0;
    defparam \u0.dat_o_0_a2_i_a2_17_LC_18_27_3 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_0_a2_i_a2_17_LC_18_27_3 .LUT_INIT=16'b0000101000100010;
    LogicCell40 \u0.dat_o_0_a2_i_a2_17_LC_18_27_3  (
            .in0(N__50463),
            .in1(N__48997),
            .in2(N__48991),
            .in3(N__48988),
            .lcout(\u0.N_1554 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport0_T4_RNI47IO9_0_LC_18_27_7 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T4_RNI47IO9_0_LC_18_27_7 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport0_T4_RNI47IO9_0_LC_18_27_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \u0.PIO_dport0_T4_RNI47IO9_0_LC_18_27_7  (
            .in0(N__48655),
            .in1(N__48649),
            .in2(N__48634),
            .in3(N__49623),
            .lcout(N_207_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev0_Td_RNIR6H22_1_LC_18_28_6 .C_ON=1'b0;
    defparam \u0.DMA_dev0_Td_RNIR6H22_1_LC_18_28_6 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev0_Td_RNIR6H22_1_LC_18_28_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \u0.DMA_dev0_Td_RNIR6H22_1_LC_18_28_6  (
            .in0(_gnd_net_),
            .in1(N__48521),
            .in2(_gnd_net_),
            .in3(N__48394),
            .lcout(),
            .ltout(\u0.N_1651_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport0_T2_RNIC2LMI_1_LC_18_28_7 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T2_RNIC2LMI_1_LC_18_28_7 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport0_T2_RNIC2LMI_1_LC_18_28_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \u0.PIO_dport0_T2_RNIC2LMI_1_LC_18_28_7  (
            .in0(N__48367),
            .in1(N__48361),
            .in2(N__48346),
            .in3(N__48343),
            .lcout(wb_dat_o_c_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNID2B71_16_LC_18_29_6 .C_ON=1'b0;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNID2B71_16_LC_18_29_6 .SEQ_MODE=4'b0000;
    defparam \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNID2B71_16_LC_18_29_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \u1.DMA_control.gen_DMAbuf_Rxbuf.mem_mem_ram6__RNID2B71_16_LC_18_29_6  (
            .in0(N__50212),
            .in1(N__49750),
            .in2(_gnd_net_),
            .in3(N__49738),
            .lcout(mem_mem_ram6__RNID2B71_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_cmdport_Teoc_5_LC_19_20_0 .C_ON=1'b0;
    defparam \u0.PIO_cmdport_Teoc_5_LC_19_20_0 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_cmdport_Teoc_5_LC_19_20_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.PIO_cmdport_Teoc_5_LC_19_20_0  (
            .in0(N__49314),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51802),
            .lcout(PIO_cmdport_Teoc_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54296),
            .ce(N__49700),
            .sr(N__53406));
    defparam \u0.PIO_dport0_T4_RNIFIIO9_1_LC_19_25_6 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T4_RNIFIIO9_1_LC_19_25_6 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport0_T4_RNIFIIO9_1_LC_19_25_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \u0.PIO_dport0_T4_RNIFIIO9_1_LC_19_25_6  (
            .in0(N__49657),
            .in1(N__49607),
            .in2(N__52804),
            .in3(N__49576),
            .lcout(N_209_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport0_T1_0_LC_20_18_3 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T1_0_LC_20_18_3 .SEQ_MODE=4'b1010;
    defparam \u0.PIO_dport0_T1_0_LC_20_18_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \u0.PIO_dport0_T1_0_LC_20_18_3  (
            .in0(_gnd_net_),
            .in1(N__51621),
            .in2(_gnd_net_),
            .in3(N__49465),
            .lcout(PIO_dport0_T1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54285),
            .ce(N__49376),
            .sr(N__53403));
    defparam \u0.CtrlReg_29_LC_20_19_7 .C_ON=1'b0;
    defparam \u0.CtrlReg_29_LC_20_19_7 .SEQ_MODE=4'b1010;
    defparam \u0.CtrlReg_29_LC_20_19_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \u0.CtrlReg_29_LC_20_19_7  (
            .in0(_gnd_net_),
            .in1(N__49288),
            .in2(_gnd_net_),
            .in3(N__51622),
            .lcout(\u0.CtrlRegZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54297),
            .ce(N__53642),
            .sr(N__53407));
    defparam \u0.PIO_dport0_T4_RNIJ3J22_7_LC_20_22_3 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T4_RNIJ3J22_7_LC_20_22_3 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport0_T4_RNIJ3J22_7_LC_20_22_3 .LUT_INIT=16'b0101000011011100;
    LogicCell40 \u0.PIO_dport0_T4_RNIJ3J22_7_LC_20_22_3  (
            .in0(N__49246),
            .in1(N__52887),
            .in2(N__50284),
            .in3(N__49219),
            .lcout(\u0.dat_o_i_0_1_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev1_Teoc_RNIRIK3G_1_LC_20_22_5 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Teoc_RNIRIK3G_1_LC_20_22_5 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev1_Teoc_RNIRIK3G_1_LC_20_22_5 .LUT_INIT=16'b1111111011101110;
    LogicCell40 \u0.DMA_dev1_Teoc_RNIRIK3G_1_LC_20_22_5  (
            .in0(N__49183),
            .in1(N__49174),
            .in2(N__49165),
            .in3(N__54705),
            .lcout(N_265),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.DMA_dev1_Teoc_RNIE5K3G_0_LC_20_23_7 .C_ON=1'b0;
    defparam \u0.DMA_dev1_Teoc_RNIE5K3G_0_LC_20_23_7 .SEQ_MODE=4'b0000;
    defparam \u0.DMA_dev1_Teoc_RNIE5K3G_0_LC_20_23_7 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \u0.DMA_dev1_Teoc_RNIE5K3G_0_LC_20_23_7  (
            .in0(N__54730),
            .in1(N__54706),
            .in2(N__54541),
            .in3(N__54526),
            .lcout(N_263),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.CtrlReg_8_LC_20_27_3 .C_ON=1'b0;
    defparam \u0.CtrlReg_8_LC_20_27_3 .SEQ_MODE=4'b1010;
    defparam \u0.CtrlReg_8_LC_20_27_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.CtrlReg_8_LC_20_27_3  (
            .in0(N__54455),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52058),
            .lcout(DMActrl_BeLeC0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54334),
            .ce(N__53587),
            .sr(N__53413));
    defparam \u0.dat_o_0_a2_i_a2_6_16_LC_21_19_4 .C_ON=1'b0;
    defparam \u0.dat_o_0_a2_i_a2_6_16_LC_21_19_4 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_0_a2_i_a2_6_16_LC_21_19_4 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.dat_o_0_a2_i_a2_6_16_LC_21_19_4  (
            .in0(N__53015),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50370),
            .lcout(\u0.N_2139 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.PIO_dport0_T4_RNI7NI22_1_LC_21_22_6 .C_ON=1'b0;
    defparam \u0.PIO_dport0_T4_RNI7NI22_1_LC_21_22_6 .SEQ_MODE=4'b0000;
    defparam \u0.PIO_dport0_T4_RNI7NI22_1_LC_21_22_6 .LUT_INIT=16'b0000110010101110;
    LogicCell40 \u0.PIO_dport0_T4_RNI7NI22_1_LC_21_22_6  (
            .in0(N__52886),
            .in1(N__50257),
            .in2(N__52864),
            .in3(N__52831),
            .lcout(\u0.dat_o_0_a2_i_0_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.register_block_gen_PIO_dport0_reg_un6_sel_pio_dport0_i_0_LC_22_16_2 .C_ON=1'b0;
    defparam \u0.register_block_gen_PIO_dport0_reg_un6_sel_pio_dport0_i_0_LC_22_16_2 .SEQ_MODE=4'b0000;
    defparam \u0.register_block_gen_PIO_dport0_reg_un6_sel_pio_dport0_i_0_LC_22_16_2 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \u0.register_block_gen_PIO_dport0_reg_un6_sel_pio_dport0_i_0_LC_22_16_2  (
            .in0(N__50997),
            .in1(N__50872),
            .in2(_gnd_net_),
            .in3(N__50761),
            .lcout(N_77),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \u0.dat_o_0_a2_i_a2_8_16_LC_22_20_6 .C_ON=1'b0;
    defparam \u0.dat_o_0_a2_i_a2_8_16_LC_22_20_6 .SEQ_MODE=4'b0000;
    defparam \u0.dat_o_0_a2_i_a2_8_16_LC_22_20_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \u0.dat_o_0_a2_i_a2_8_16_LC_22_20_6  (
            .in0(N__50525),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50377),
            .lcout(\u0.N_2143 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // atahost
