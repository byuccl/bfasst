/*
Random input logic for DLA
*/

`include "../../random_number_generator.sv"

module dla_random(
    input logic clk,
    input logic rst,
    input logic i_ddr_wen_0_0,
    output logic o_dummy_out_0_0,
    input logic i_ddr_wen_0_1,
    output logic o_dummy_out_0_1,
    input logic i_ddr_wen_0_2,
    output logic o_dummy_out_0_2,
    input logic i_ddr_wen_0_3,
    output logic o_dummy_out_0_3,
    input logic i_ddr_wen_0_4,
    output logic o_dummy_out_0_4,
    input logic i_ddr_wen_0_5,
    output logic o_dummy_out_0_5,
	input logic i_ddr_wen_0_6,
    output logic o_dummy_out_0_6,
	input logic i_ddr_wen_0_7,
    output logic o_dummy_out_0_7,
	input logic i_ddr_wen_1_0,
    output logic o_dummy_out_1_0,
	input logic i_ddr_wen_1_1,
    output logic o_dummy_out_1_1,
	input logic i_ddr_wen_1_2,
    output logic o_dummy_out_1_2,
	input logic i_ddr_wen_1_3,
    output logic o_dummy_out_1_3,
	input logic i_ddr_wen_1_4,
    output logic o_dummy_out_1_4,
	input logic i_ddr_wen_1_5,
    output logic o_dummy_out_1_5,
	input logic i_ddr_wen_1_6,
    output logic o_dummy_out_1_6,
	input logic i_ddr_wen_1_7,
    output logic o_dummy_out_1_7,
	input logic i_ddr_wen_2_0,
    output logic o_dummy_out_2_0,
	input logic i_ddr_wen_2_1,
    output logic o_dummy_out_2_1,
	input logic i_ddr_wen_2_2,
    output logic o_dummy_out_2_2,
	input logic i_ddr_wen_2_3,
    output logic o_dummy_out_2_3,
	input logic i_ddr_wen_2_4,
    output logic o_dummy_out_2_4,
    input logic i_ddr_wen_2_5,
    output logic o_dummy_out_2_5,
    input logic i_ddr_wen_2_6,
    output logic o_dummy_out_2_6,
    input logic i_ddr_wen_2_7,
    output logic o_dummy_out_2_7,
    input logic i_ddr_wen_3_0,
    output logic o_dummy_out_3_0,
    input logic i_ddr_wen_3_1,
    output logic o_dummy_out_3_1,
    input logic i_ddr_wen_3_2,
    output logic o_dummy_out_3_2,
    input logic i_ddr_wen_3_3,
    output logic o_dummy_out_3_3,
    input logic i_ddr_wen_3_4,
    output logic o_dummy_out_3_4,
    input logic i_ddr_wen_3_5,
    output logic o_dummy_out_3_5,
    input logic i_ddr_wen_3_6,
    output logic o_dummy_out_3_6,
    input logic i_ddr_wen_3_7,
    output logic o_dummy_out_3_7,
    input logic i_ddr_wen_4_0,
    output logic o_dummy_out_4_0,
    input logic i_ddr_wen_4_1,
    output logic o_dummy_out_4_1,
    input logic i_ddr_wen_4_2,
    output logic o_dummy_out_4_2,
    input logic i_ddr_wen_4_3,
    output logic o_dummy_out_4_3,
    input logic i_ddr_wen_4_4,
    output logic o_dummy_out_4_4,
    input logic i_ddr_wen_4_5,
    output logic o_dummy_out_4_5,
    input logic i_ddr_wen_4_6,
    output logic o_dummy_out_4_6,
    input logic i_ddr_wen_4_7,
    output logic o_dummy_out_4_7,
    input logic i_ddr_wen_5_0,
    output logic o_dummy_out_5_0,
    input logic i_ddr_wen_5_1,
    output logic o_dummy_out_5_1,
    input logic i_ddr_wen_5_2,
    output logic o_dummy_out_5_2,
    input logic i_ddr_wen_5_3,
    output logic o_dummy_out_5_3,
    input logic i_ddr_wen_5_4,
    output logic o_dummy_out_5_4,
    input logic i_ddr_wen_5_5,
    output logic o_dummy_out_5_5,
    input logic i_ddr_wen_5_6,
    output logic o_dummy_out_5_6,
    input logic i_ddr_wen_5_7,
    output logic o_dummy_out_5_7,
    output logic o_valid
);

logic [15:0] i_ddr[5:0][7:0];
generate // generate block for random number generator
genvar i;
genvar j;
for(i=0; i<6; i=i+1) begin
    for(j=0; j<8; j=j+1) begin
        RandomNumberGenerator #(16, i+j) random_number_generator_0(
            .clk(clk),
            .reset(rst),
            .random_number(i_ddr[i][j])
        );
    end
end
endgenerate


DLA dla0(
	clk,
	rst,
	i_ddr_wen_0_0,
	i_ddr[0][0],
	o_dummy_out_0_0,
	i_ddr_wen_0_1,
	i_ddr[0][1],
	o_dummy_out_0_1,
	i_ddr_wen_0_2,
	i_ddr[0][2],
	o_dummy_out_0_2,
	i_ddr_wen_0_3,
	i_ddr[0][3],
	o_dummy_out_0_3,
	i_ddr_wen_0_4,
	i_ddr[0][4],
	o_dummy_out_0_4,
	i_ddr_wen_0_5,
	i_ddr[0][5],
	o_dummy_out_0_5,
	i_ddr_wen_0_6,
	i_ddr[0][6],
	o_dummy_out_0_6,
	i_ddr_wen_0_7,
	i_ddr[0][7],
	o_dummy_out_0_7,
	i_ddr_wen_1_0,
	i_ddr[1][0],
	o_dummy_out_1_0,
	i_ddr_wen_1_1,
	i_ddr[1][1],
	o_dummy_out_1_1,
	i_ddr_wen_1_2,
	i_ddr[1][2],
	o_dummy_out_1_2,
	i_ddr_wen_1_3,
	i_ddr[1][3],
	o_dummy_out_1_3,
	i_ddr_wen_1_4,
	i_ddr[1][4],
	o_dummy_out_1_4,
	i_ddr_wen_1_5,
	i_ddr[1][5],
	o_dummy_out_1_5,
	i_ddr_wen_1_6,
	i_ddr[1][6],
	o_dummy_out_1_6,
	i_ddr_wen_1_7,
	i_ddr[1][7],
	o_dummy_out_1_7,
	i_ddr_wen_2_0,
	i_ddr[2][0],
	o_dummy_out_2_0,
	i_ddr_wen_2_1,
	i_ddr[2][1],
	o_dummy_out_2_1,
	i_ddr_wen_2_2,
	i_ddr[2][2],
	o_dummy_out_2_2,
	i_ddr_wen_2_3,
	i_ddr[2][3],
	o_dummy_out_2_3,
	i_ddr_wen_2_4,
	i_ddr[2][4],
	o_dummy_out_2_4,
	i_ddr_wen_2_5,
	i_ddr[2][5],
	o_dummy_out_2_5,
	i_ddr_wen_2_6,
	i_ddr[2][6],
	o_dummy_out_2_6,
	i_ddr_wen_2_7,
	i_ddr[2][7],
	o_dummy_out_2_7,
	i_ddr_wen_3_0,
	i_ddr[3][0],
	o_dummy_out_3_0,
	i_ddr_wen_3_1,
	i_ddr[3][1],
	o_dummy_out_3_1,
	i_ddr_wen_3_2,
	i_ddr[3][2],
	o_dummy_out_3_2,
	i_ddr_wen_3_3,
	i_ddr[3][3],
	o_dummy_out_3_3,
	i_ddr_wen_3_4,
	i_ddr[3][4],
	o_dummy_out_3_4,
	i_ddr_wen_3_5,
	i_ddr[3][5],
	o_dummy_out_3_5,
	i_ddr_wen_3_6,
	i_ddr[3][6],
	o_dummy_out_3_6,
	i_ddr_wen_3_7,
	i_ddr[3][7],
	o_dummy_out_3_7,
	i_ddr_wen_4_0,
	i_ddr[4][0],
	o_dummy_out_4_0,
	i_ddr_wen_4_1,
	i_ddr[4][1],
	o_dummy_out_4_1,
	i_ddr_wen_4_2,
	i_ddr[4][2],
	o_dummy_out_4_2,
	i_ddr_wen_4_3,
	i_ddr[4][3],
	o_dummy_out_4_3,
	i_ddr_wen_4_4,
	i_ddr[4][4],
	o_dummy_out_4_4,
	i_ddr_wen_4_5,
	i_ddr[4][5],
	o_dummy_out_4_5,
	i_ddr_wen_4_6,
	i_ddr[4][6],
	o_dummy_out_4_6,
	i_ddr_wen_4_7,
	i_ddr[4][7],
	o_dummy_out_4_7,
	i_ddr_wen_5_0,
	i_ddr[5][0],
	o_dummy_out_5_0,
	i_ddr_wen_5_1,
	i_ddr[5][1],
	o_dummy_out_5_1,
	i_ddr_wen_5_2,
	i_ddr[5][2],
	o_dummy_out_5_2,
	i_ddr_wen_5_3,
	i_ddr[5][3],
	o_dummy_out_5_3,
	i_ddr_wen_5_4,
	i_ddr[5][4],
	o_dummy_out_5_4,
	i_ddr_wen_5_5,
	i_ddr[5][5],
	o_dummy_out_5_5,
	i_ddr_wen_5_6,
	i_ddr[5][6],
	o_dummy_out_5_6,
	i_ddr_wen_5_7,
	i_ddr[5][7],
	o_dummy_out_5_7,
	o_valid
);


endmodule