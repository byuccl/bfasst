
module uart (input clk, input rst, output rx_overrun_error, output rx_busy, output tx_busy, input output_axis_tready, input input_axis_tvalid, output input_axis_tready, output output_axis_tvalid, input \input_axis_tdata[3] , input \input_axis_tdata[4] , output \output_axis_tdata[0] , output \output_axis_tdata[3] , input \input_axis_tdata[0] , input \input_axis_tdata[5] , output rx_frame_error, output \output_axis_tdata[6] , output \output_axis_tdata[2] , output \output_axis_tdata[7] , output \output_axis_tdata[4] , output \output_axis_tdata[5] , output \output_axis_tdata[1] , input rxd, input \input_axis_tdata[2] , input \input_axis_tdata[6] , input \input_axis_tdata[7] , input \input_axis_tdata[1] , output txd);

wire clk, n2, rst, n5, output_axis_tready, n10, input_axis_tvalid, n13, n15, n16;
wire n17, n18, n19, n20, n21, n24, n25, n26, n27, n29;
wire n30, n34, n38, n39, n40, n41, n43, n44, n45, n46;
wire n47, n48, n49, n50, n51, n54, n55, n56, n58, n59;
wire n60, n61, n62, n63, n64, n65, n66, n67, \input_axis_tdata[3] , \input_axis_tdata[4] ;
wire n71, n80, n81, n82, n83, n84, n85, n86, n87, n88;
wire n89, n95, n97, n98, n99, n100, n101, n102, n103, n104;
wire n105, n106, n107, n108, n109, n110, n112, n113, n114, n115;
wire n116, n117, n119, n120, n126, n127, n128, n130, n135, n137;
wire n138, n139, n140, n141, n143, n144, n145, n146, n147, n148;
wire n149, \input_axis_tdata[0] , n151, \input_axis_tdata[5] , n153, n154, n156, n157, n158, n159;
wire n160, n161, n162, n163, n164, n165, n166, n167, n168, n169;
wire n170, n171, n172, n173, n174, n175, n176, n177, n178, n179;
wire n180, n181, n182, n183, n184, n185, n186, n187, n188, n189;
wire n190, n191, n192, n193, n194, n195, n196, n204, rxd, \input_axis_tdata[2] ;
wire \input_axis_tdata[6] , n214, n215, n216, n217, n218, n219, \input_axis_tdata[7] , n221, n222;
wire n223, n224, n225, n226, n227, n228, n229, n230, n231, n232;
wire n233, n234, n235, n236, n237, n238, n239, n240, n241, n242;
wire n243, n244, n245, n246, n247, n248, n249, n250, n251, n252;
wire n253, n256, n260, n261, n262, n263, n264, n265, n269, \input_axis_tdata[1] ;
wire n271, n272, n273, n282, n283, n284, n285, n286, n287, n288;
wire n289, n290, n292, n293, n294, n295, n296, n297, n298, n299;
wire n300, n301, n302, n303, n304, n305, n306, n307, n308, n309;
wire n310, n311, n312, n313, n314, n315, n316, n317, n318, n319;
wire n320, n321, n322, n323, n324, n325, n326, n327, n328, n329;
wire n330, n331, n332, n333, n334, n335, n336, n337, n338, n339;
wire n340, n341, n342, n343, n344, n345, n346, n347, n348, n349;
wire n350, n351, n352, n353, n354, n355, n356, n357, n358, n359;
wire n360, n361, n362, n363, n364, n365, n366, n367, n368, n369;
wire n370, n371, n372, n373, n374, n375, n376, n377, n378, n379;
wire n380, n381, n382, n383, n384, n385, n386, n387, n388, n389;
wire n390, n391, n392, n393, n394, n395, n396, n397, n398, n399;
wire n400, n401, n402, n403, n404, n405, n406, n407, n408, n409;
wire n410, n411, n412, n413, n414, n415, n416, n417, n418, n419;
wire n420, n421, n422, n423, n424, n425, n426, n427, n428, n429;
wire n430, n431, n432, n433, n434, n435, n436, n437, n438, n439;
wire n440, n441, n442, n443, n444, n445, n446, n447, n448, n449;
wire n450, n451, n452, n453, n454, n455, n456, n457, n458, n459;
wire n460, n461, n462, n463, n464, n465, n466, n467, n468, n469;
wire n470, n471, n472, n473, n474, n475, n476, n477, n478, n479;
wire n480, n481, n482, n483, n484, n485, n486, n487, n488, n489;
wire n490, n491, n492, n493, n494, n495, n496, n497, n498, n499;
wire n500, n501, n502, n503, n504, n505, n506, n507, n508, n509;
wire n510, n511, n512, n513, n514, n515, n516, n517, n518, n519;
wire n520, n521, n522, n523, n524, n525, n526, n527, n528, n529;
wire n530, n531, n532, n533, n534, n535, n536, n537, n538, n539;
wire n540, n541, n542, n543, n544, n545, n546, n547, n548, n549;
wire n550, n551, n552, n553, n554, n555, n556, n557, n558, n559;
wire n560;
reg n4 = 0, rx_overrun_error = 0, rx_busy = 0, tx_busy = 0, input_axis_tready = 0, n14 = 0, n22 = 0, n23 = 0, n28 = 0, n31 = 0;
reg output_axis_tvalid = 0, n33 = 0, n35 = 0, n36 = 0, n37 = 0, n42 = 0, n52 = 0, n53 = 0, n57 = 0, n70 = 0;
reg n72 = 0, n73 = 0, n74 = 0, n75 = 0, n76 = 0, n77 = 0, n78 = 0, n79 = 0, n90 = 0, n91 = 0;
reg n92 = 0, n93 = 0, n94 = 0, n96 = 0, n111 = 0, n118 = 0, \output_axis_tdata[0]  = 0, \output_axis_tdata[3]  = 0, n123 = 0, n124 = 0;
reg n125 = 0, n129 = 0, n131 = 0, n132 = 0, n133 = 0, n134 = 0, n136 = 0, n142 = 0, n155 = 0, n197 = 0;
reg n198 = 0, n199 = 0, n200 = 0, n201 = 0, n202 = 0, rx_frame_error = 0, \output_axis_tdata[6]  = 0, \output_axis_tdata[2]  = 0, \output_axis_tdata[7]  = 0, \output_axis_tdata[4]  = 0;
reg \output_axis_tdata[5]  = 0, \output_axis_tdata[1]  = 0, n254 = 0, n255 = 0, n257 = 0, n258 = 0, n259 = 0, n266 = 0, n267 = 0, n268 = 0;
reg n274 = 0, n275 = 0, n276 = 0, n277 = 0, n278 = 0, n279 = 0, n280 = 0, n281 = 0, txd = 0;
assign n282 = 1;
assign n322 = 1;
assign n302 = 1;
assign n232 = 1;

assign n343 = /* LUT    6  7  2 */ 1'b1;
assign n177 = /* LUT    8  6  6 */ (n50 ? !n176 : (n176 ? 1'b0 : (n4 ? 1'b1 : n14)));
assign n338 = /* LUT    8  9  0 */ (n53 ? n111 : (n111 ? n14 : !n14));
assign n66  = /* LUT    7  2  3 */ (n33 ? 1'b1 : (n31 ? 1'b1 : (n28 ? 1'b1 : n23)));
assign n339 = /* LUT   11  3  4 */ (n295 ? (n5 ? n254 : !n254) : (n5 ? !n254 : n254));
assign n340 = /* LUT   11  6  7 */ (n317 ? (\input_axis_tdata[7]  ? n5 : !n5) : (\input_axis_tdata[7]  ? !n5 : n5));
assign n341 = /* LUT   12  5  1 */ (n323 ? (\input_axis_tdata[1]  ? n5 : !n5) : (\input_axis_tdata[1]  ? !n5 : n5));
assign n342 = /* LUT    9  8  3 */ (n215 ? n100 : 1'b0);
assign n344 = /* LUT    8  6  0 */ (n86 ? 1'b1 : (n50 ? 1'b1 : n14));
assign n345 = /* LUT    9 13  3 */ n200;
assign n346 = /* LUT    7  1  1 */ (n23 ? n31 : !n31);
assign n347 = /* LUT    9  6  5 */ (n245 ? (n90 ? (n87 ? 1'b1 : n183) : (n87 ? 1'b0 : n183)) : (n90 ? (n87 ? 1'b0 : n183) : (n87 ? 1'b1 : n183)));
assign n65  = /* LUT    7  2  1 */ (n24 ? rst : (n64 ? rst : (n27 ? 1'b1 : rst)));
assign n348 = /* LUT    8 12  4 */ (n119 ? 1'b1 : rst);
assign n349 = /* LUT   11  3  6 */ (n297 ? (n5 ? n133 : !n133) : (n5 ? !n133 : n133));
assign n350 = /* LUT   11  6  5 */ (n315 ? (\input_axis_tdata[5]  ? n5 : !n5) : (\input_axis_tdata[5]  ? !n5 : n5));
assign n351 = /* LUT    8  3  0 */ (n119 ? rst : 1'b1);
assign n352 = /* LUT   12  5  3 */ (n325 ? (\input_axis_tdata[3]  ? n5 : !n5) : (\input_axis_tdata[3]  ? !n5 : n5));
assign n353 = /* LUT    9  8  1 */ (n147 ? n100 : 1'b0);
assign n174 = /* LUT    8  6  2 */ (n79 ? 1'b1 : (n76 ? 1'b1 : (n72 ? 1'b1 : n73)));
assign n355 = /* LUT    9  6  7 */ (n247 ? (n91 ? (n87 ? 1'b1 : n181) : (n87 ? 1'b0 : n181)) : (n91 ? (n87 ? 1'b0 : n181) : (n87 ? 1'b1 : n181)));
assign n356 = /* LUT   11  5  3 */ (n305 ? (\input_axis_tdata[3]  ? n5 : !n5) : (\input_axis_tdata[3]  ? !n5 : n5));
assign n357 = /* LUT   11  6  3 */ (n313 ? (\input_axis_tdata[3]  ? n5 : !n5) : (\input_axis_tdata[3]  ? !n5 : n5));
assign n358 = /* LUT    8  3  6 */ (n24 ? rst : (n61 ? 1'b1 : rst));
assign n359 = /* LUT   12  5  5 */ (n327 ? (\input_axis_tdata[5]  ? n5 : !n5) : (\input_axis_tdata[5]  ? !n5 : n5));
assign n360 = /* LUT    9  8  7 */ (n40 ? n100 : 1'b0);
assign n361 = /* LUT   12  2  4 */ (n2 ? n279 : (n279 ? (\input_axis_tdata[4]  ? 1'b1 : !input_axis_tvalid) : (\input_axis_tdata[4]  ? input_axis_tvalid : 1'b0)));
assign n362 = /* LUT    9  1  1 */ (n24 ? n216 : (n216 ? (\input_axis_tdata[2]  ? 1'b1 : n60) : (\input_axis_tdata[2]  ? !n60 : 1'b0)));
assign n363 = /* LUT    8  8  7 */ (n54 ? 1'b0 : n103);
assign n364 = /* LUT    9  6  1 */ (n241 ? (n77 ? (n87 ? 1'b1 : n180) : (n87 ? 1'b0 : n180)) : (n77 ? (n87 ? 1'b0 : n180) : (n87 ? 1'b1 : n180)));
assign n365 = /* LUT   11  5  1 */ (n303 ? (\input_axis_tdata[1]  ? n5 : !n5) : (\input_axis_tdata[1]  ? !n5 : n5));
assign n366 = /* LUT   11  6  1 */ (n311 ? (\input_axis_tdata[1]  ? n5 : !n5) : (\input_axis_tdata[1]  ? !n5 : n5));
assign n367 = /* LUT   12  5  7 */ (n329 ? (\input_axis_tdata[7]  ? n5 : !n5) : (\input_axis_tdata[7]  ? !n5 : n5));
assign n368 = /* LUT    9  8  5 */ (n229 ? n100 : 1'b0);
assign n369 = /* LUT   12  2  6 */ (n2 ? n281 : (\input_axis_tdata[6]  ? (n281 ? 1'b1 : input_axis_tvalid) : (n281 ? !input_axis_tvalid : 1'b0)));
assign n370 = /* LUT    8  8  5 */ (n54 ? (n196 ? 1'b1 : n4) : n196);
assign n371 = /* LUT    9  1  3 */ (n24 ? n217 : (n217 ? (\input_axis_tdata[4]  ? 1'b1 : n60) : (\input_axis_tdata[4]  ? !n60 : 1'b0)));
assign n372 = /* LUT    9  6  3 */ (n243 ? (n75 ? (n87 ? 1'b1 : n184) : (n87 ? 1'b0 : n184)) : (n75 ? (n87 ? 1'b0 : n184) : (n87 ? 1'b1 : n184)));
assign n373 = /* LUT   11  5  7 */ (n309 ? (\input_axis_tdata[7]  ? n5 : !n5) : (\input_axis_tdata[7]  ? !n5 : n5));
assign n374 = /* LUT    7  2  5 */ (n26 ? 1'b0 : (n30 ? n28 : (n28 ? !n25 : n25)));
assign n375 = /* LUT   12  2  0 */ (n2 ? n275 : (\input_axis_tdata[0]  ? (n275 ? 1'b1 : input_axis_tvalid) : (n275 ? !input_axis_tvalid : 1'b0)));
assign n376 = /* LUT    9  1  5 */ (n24 ? n218 : (n218 ? (\input_axis_tdata[6]  ? 1'b1 : n60) : (\input_axis_tdata[6]  ? !n60 : 1'b0)));
assign n195 = /* LUT    8  8  3 */ (n53 ? 1'b1 : (n111 ? 1'b1 : n52));
assign n377 = /* LUT   11  5  5 */ (n307 ? (\input_axis_tdata[5]  ? n5 : !n5) : (\input_axis_tdata[5]  ? !n5 : n5));
assign n378 = /* LUT    7  5  6 */ (n80 ? (n83 ? 1'b1 : (rst ? 1'b1 : !n84)) : (rst ? 1'b1 : !n84));
assign n379 = /* LUT    8  5  5 */ (n166 ? (n164 ? 1'b1 : n83) : (n164 ? !n83 : 1'b0));
assign n380 = /* LUT   12  2  2 */ (n2 ? n277 : (\input_axis_tdata[2]  ? (n277 ? 1'b1 : input_axis_tvalid) : (n277 ? !input_axis_tvalid : 1'b0)));
assign n381 = /* LUT    9  1  7 */ (n24 ? 1'b1 : (n60 ? 1'b1 : (rst ? 1'b1 : n10)));
assign n194 = /* LUT    8  8  1 */ (n50 ? (n193 ? 1'b1 : n105) : (n193 ? 1'b1 : (n14 ? n105 : 1'b0)));
assign n382 = /* LUT    9  4  4 */ (n160 ? (n230 ? 1'b1 : !n10) : (n230 ? n10 : 1'b0));
assign n383 = /* LUT    8  5  7 */ (n158 ? (n163 ? 1'b1 : n83) : (n163 ? !n83 : 1'b0));
assign n384 = /* LUT    9  9  0 */ (n101 ? (n197 ? n102 : 1'b0) : (n199 ? n102 : 1'b0));
assign n385 = /* LUT    8  2  1 */ (n2 ? (n144 ? 1'b0 : n57) : (n144 ? input_axis_tvalid : n57));
assign n386 = /* LUT    7  5  2 */ (n82 ? (n18 ? 1'b1 : n83) : (n18 ? !n83 : 1'b0));
assign n387 = /* LUT    8  5  1 */ (n162 ? (n161 ? 1'b1 : n83) : (n161 ? !n83 : 1'b0));
assign n388 = /* LUT   11  1  6 */ (n60 ? n273 : (n273 ? (\input_axis_tdata[0]  ? 1'b1 : n24) : (\input_axis_tdata[0]  ? !n24 : 1'b0)));
assign n389 = /* LUT    9  7  2 */ (n253 ? (n188 ? (n73 ? 1'b1 : !n87) : (n73 ? n87 : 1'b0)) : (n188 ? (n73 ? !n87 : 1'b1) : (n73 ? 1'b0 : n87)));
assign n390 = /* LUT    9  9  2 */ (n101 ? (n199 ? n102 : 1'b0) : (n202 ? n102 : 1'b0));
assign n391 = /* LUT    7  8  6 */ (n14 ? 1'b1 : n114);
assign n145 = /* LUT    8  2  3 */ (n33 ? 1'b0 : (n28 ? 1'b0 : !n23));
assign n392 = /* LUT    8  5  3 */ (n168 ? (n154 ? 1'b1 : n83) : (n154 ? !n83 : 1'b0));
assign n393 = /* LUT    7  6  6 */ (rst ? 1'b1 : !n83);
assign n394 = /* LUT    9  7  0 */ (n248 ? (n87 ? n93 : n190) : (n87 ? !n93 : n190));
assign n395 = /* LUT   11  1  4 */ (n254 ? 1'b1 : (n255 ? 1'b1 : (n259 ? 1'b1 : n258)));
assign n396 = /* LUT   11  2  2 */ (n284 ? (n5 ? (n259 ? 1'b1 : n10) : (n259 ? n10 : 1'b1)) : (n5 ? (n259 ? n10 : 1'b1) : (n259 ? 1'b1 : n10)));
assign n397 = /* LUT   11  7  0 */ (n318 ? !n5 : n5);
assign n112 = /* LUT    7  8  0 */ (n86 ? rst : (n49 ? rst : 1'b1));
assign n146 = /* LUT    8  2  5 */ (n33 ? 1'b1 : n28);
assign n399 = /* LUT   12  1  5 */ (n60 ? n320 : (n320 ? (\input_axis_tdata[2]  ? 1'b1 : n24) : (\input_axis_tdata[2]  ? !n24 : 1'b0)));
assign n400 = /* LUT    9  2  0 */ (n24 ? n55 : (\input_axis_tdata[3]  ? (n55 ? 1'b1 : !n60) : (n55 ? n60 : 1'b0)));
assign n401 = /* LUT    8  7  6 */ (n96 ? 1'b1 : (n77 ? 1'b1 : (n42 ? 1'b1 : n94)));
assign n272 = /* LUT   11  1  2 */ (n264 ? (n250 ? 1'b1 : !n10) : (n250 ? n10 : 1'b0));
assign n403 = /* LUT    9  7  6 */ (n100 ? n140 : 1'b0);
assign n404 = /* LUT   11  2  0 */ (n282 ? (n257 ? n10 : 1'b1) : (n257 ? 1'b1 : n10));
assign n405 = /* LUT    9  9  6 */ (n101 ? (n201 ? n102 : 1'b0) : (n22 ? n102 : 1'b0));
assign n406 = /* LUT    7  8  2 */ (n45 ? (n113 ? 1'b0 : !n14) : (n113 ? 1'b0 : n14));
assign n407 = /* LUT   12  1  7 */ (n60 ? n321 : (n321 ? (\input_axis_tdata[5]  ? 1'b1 : n24) : (\input_axis_tdata[5]  ? !n24 : 1'b0)));
assign n408 = /* LUT    9  2  2 */ (n24 ? n224 : (n224 ? (n60 ? 1'b1 : \input_axis_tdata[3] ) : (n60 ? 1'b0 : \input_axis_tdata[3] )));
assign n409 = /* LUT    8  7  4 */ (n178 ? (n107 ? 1'b1 : n83) : (n107 ? !n83 : 1'b0));
assign n410 = /* LUT    9 12  5 */ n198;
assign n271 = /* LUT   11  1  0 */ (n263 ? (n269 ? 1'b1 : !n10) : (n269 ? n10 : 1'b0));
assign n412 = /* LUT    9  7  4 */ (n100 ? n214 : 1'b0);
assign n413 = /* LUT   11  2  6 */ (n288 ? (n134 ? n5 : !n5) : (n134 ? !n5 : n5));
assign n414 = /* LUT   12  6  1 */ (n331 ? (\input_axis_tdata[1]  ? n5 : !n5) : (\input_axis_tdata[1]  ? !n5 : n5));
assign n319 = /* LUT   12  1  1 */ (n40 ? (n10 ? 1'b1 : n261) : (n10 ? 1'b0 : n261));
assign n416 = /* LUT    9 12  3 */ n22;
assign n417 = /* LUT    9  2  4 */ (n24 ? n225 : (n225 ? (n60 ? 1'b1 : \input_axis_tdata[4] ) : (n60 ? 1'b0 : \input_axis_tdata[4] )));
assign n418 = /* LUT    8  7  2 */ (n172 ? (n108 ? 1'b1 : n83) : (n108 ? !n83 : 1'b0));
assign n419 = /* LUT    9  5  5 */ (n237 ? (n87 ? n35 : n43) : (n87 ? !n35 : n43));
assign n420 = /* LUT   11  2  4 */ (n286 ? (n266 ? n5 : !n5) : (n266 ? !n5 : n5));
assign n421 = /* LUT    6  1  0 */ (n24 ? 1'b1 : (n2 ? rst : 1'b1));
assign n422 = /* LUT   12  6  3 */ (n333 ? (\input_axis_tdata[3]  ? n5 : !n5) : (\input_axis_tdata[3]  ? !n5 : n5));
assign n423 = /* LUT    9 12  1 */ n201;
assign n424 = /* LUT    9  2  6 */ (n24 ? n226 : (n226 ? (n60 ? 1'b1 : \input_axis_tdata[7] ) : (n60 ? 1'b0 : \input_axis_tdata[7] )));
assign n425 = /* LUT    8  7  0 */ (n90 ? 1'b1 : (n93 ? 1'b1 : (n91 ? 1'b1 : n92)));
assign n204 = /* LUT    8 10  2 */ (n54 ? 1'b0 : (n103 ? 1'b0 : (n50 ? 1'b0 : n14)));
assign n426 = /* LUT    9  5  7 */ (n239 ? (n87 ? n78 : n191) : (n87 ? !n78 : n191));
assign n427 = /* LUT    6  2  0 */ (input_axis_tready ? !input_axis_tvalid : 1'b1);
assign n428 = /* LUT   12  6  5 */ (n335 ? (\input_axis_tdata[5]  ? n5 : !n5) : (\input_axis_tdata[5]  ? !n5 : n5));
assign n228 = /* LUT    9  3  5 */ (n10 ? n227 : n151);
assign n430 = /* LUT    7  7  1 */ (n98 ? (n83 ? 1'b1 : n99) : (n83 ? 1'b0 : n99));
assign n431 = /* LUT    9  5  1 */ (n233 ? (n87 ? n94 : n100) : (n87 ? !n94 : n100));
assign n432 = /* LUT    7  9  3 */ (n4 ? (n116 ? 1'b0 : (n100 ? n51 : 1'b0)) : (n116 ? !n51 : (n100 ? 1'b1 : !n51)));
assign n137 = /* LUT    8  1  0 */ (n24 ? 1'b0 : (n58 ? n60 : (n27 ? 1'b1 : n60)));
assign n433 = /* LUT    6  1  4 */ (n24 ? 1'b1 : rst);
assign n434 = /* LUT   12  6  7 */ (n337 ? (n5 ? \input_axis_tdata[7]  : !\input_axis_tdata[7] ) : (n5 ? !\input_axis_tdata[7]  : \input_axis_tdata[7] ));
assign n435 = /* LUT    8 10  6 */ (n102 ? (n200 ? (n101 ? n118 : 1'b1) : (n101 ? n118 : 1'b0)) : 1'b0);
assign n436 = /* LUT    9  5  3 */ (n235 ? (n87 ? n72 : n173) : (n87 ? !n72 : n173));
assign n437 = /* LUT    9 10  3 */ !n4;
assign n438 = /* LUT    7  9  1 */ (n4 ? (n115 ? 1'b0 : (n100 ? n51 : 1'b0)) : (n115 ? !n51 : (n100 ? 1'b1 : !n51)));
assign n439 = /* LUT   11  3  1 */ (n292 ? (n255 ? n5 : !n5) : (n255 ? !n5 : n5));
assign n440 = /* LUT    7  2  6 */ (n31 ? !n33 : (n28 ? !n33 : (n23 ? !n33 : n33)));
assign n441 = /* LUT   11  4  1 */ (n300 ? (n125 ? n5 : !n5) : (n125 ? !n5 : n5));
assign n139 = /* LUT    8  1  4 */ (n133 ? 1'b1 : (n138 ? 1'b1 : (n136 ? 1'b1 : n131)));
assign n176 = /* LUT    8  6  5 */ (n85 ? 1'b1 : (n175 ? 1'b1 : (n89 ? 1'b1 : n95)));
assign n443 = /* LUT   12  3  0 */ (n59 ? n2 : (n2 ? n274 : 1'b0));
assign n444 = /* LUT    7  7  7 */ (n47 ? n100 : 1'b0);
assign n445 = /* LUT   11  3  3 */ (n294 ? (n131 ? n5 : !n5) : (n131 ? !n5 : n5));
assign n446 = /* LUT    7  2  4 */ (input_axis_tvalid ? 1'b1 : n66);
assign n447 = /* LUT    8  6  7 */ !n177;
assign n448 = /* LUT    7  2  2 */ (n59 ? n65 : (n65 ? (rst ? 1'b1 : !n2) : 1'b0));
assign n449 = /* LUT   11  3  5 */ (n296 ? (n123 ? n5 : !n5) : (n123 ? !n5 : n5));
assign n450 = /* LUT   11  6  6 */ (n316 ? (\input_axis_tdata[6]  ? n5 : !n5) : (\input_axis_tdata[6]  ? !n5 : n5));
assign n451 = /* LUT    9  8  2 */ (n100 ? n230 : 1'b0);
assign n452 = /* LUT   12  5  0 */ (n322 ? !\input_axis_tdata[0]  : \input_axis_tdata[0] );
assign n453 = /* LUT    9  6  4 */ (n244 ? (n87 ? n96 : n97) : (n87 ? !n96 : n97));
assign n454 = /* LUT   11  3  7 */ (n298 ? (n124 ? n5 : !n5) : (n124 ? !n5 : n5));
assign n64  = /* LUT    7  2  0 */ (n59 ? (n28 ? 1'b1 : (n23 ? 1'b1 : n33)) : 1'b0);
assign n456 = /* LUT   11  6  4 */ (n314 ? (\input_axis_tdata[4]  ? n5 : !n5) : (\input_axis_tdata[4]  ? !n5 : n5));
assign n457 = /* LUT   12  5  2 */ (n324 ? (\input_axis_tdata[2]  ? n5 : !n5) : (\input_axis_tdata[2]  ? !n5 : n5));
assign n458 = /* LUT   11  8  1 */ (n100 ? n269 : 1'b0);
assign n459 = /* LUT    9  8  0 */ (n100 ? n135 : 1'b0);
assign n460 = /* LUT    8  6  3 */ (n74 ? 1'b1 : (n174 ? 1'b1 : (n78 ? 1'b1 : n75)));
assign n461 = /* LUT    9  6  6 */ (n246 ? (n87 ? n74 : n185) : (n87 ? !n74 : n185));
assign n462 = /* LUT   11  6  2 */ (n312 ? (\input_axis_tdata[2]  ? n5 : !n5) : (\input_axis_tdata[2]  ? !n5 : n5));
assign n463 = /* LUT   12  5  4 */ (n326 ? (\input_axis_tdata[4]  ? n5 : !n5) : (\input_axis_tdata[4]  ? !n5 : n5));
assign n464 = /* LUT    9  8  6 */ (n100 ? n223 : 1'b0);
assign n465 = /* LUT   12  2  5 */ (n280 ? (\input_axis_tdata[5]  ? 1'b1 : (input_axis_tvalid ? n2 : 1'b1)) : (\input_axis_tdata[5]  ? (input_axis_tvalid ? !n2 : 1'b0) : 1'b0));
assign n466 = /* LUT    7  4  0 */ output_axis_tvalid;
assign n467 = /* LUT    9  6  0 */ (n240 ? (n87 ? n37 : n182) : (n87 ? !n37 : n182));
assign n468 = /* LUT    8 14  4 */ rxd;
assign n469 = /* LUT   11  5  2 */ (n304 ? (\input_axis_tdata[2]  ? n5 : !n5) : (\input_axis_tdata[2]  ? !n5 : n5));
assign n470 = /* LUT   11  6  0 */ (n310 ? (\input_axis_tdata[0]  ? n5 : !n5) : (\input_axis_tdata[0]  ? !n5 : n5));
assign n471 = /* LUT   12  5  6 */ (n328 ? (\input_axis_tdata[6]  ? n5 : !n5) : (\input_axis_tdata[6]  ? !n5 : n5));
assign n472 = /* LUT    9  8  4 */ (n100 ? n249 : 1'b0);
assign n473 = /* LUT   12  2  7 */ (n57 ? (\input_axis_tdata[7]  ? 1'b1 : (input_axis_tvalid ? n2 : 1'b1)) : (\input_axis_tdata[7]  ? (input_axis_tvalid ? !n2 : 1'b0) : 1'b0));
assign n474 = /* LUT    8  8  6 */ (n86 ? 1'b1 : rst);
assign n216 = /* LUT    9  1  0 */ (n10 ? n140 : n141);
assign n476 = /* LUT    9  6  2 */ (n242 ? (n87 ? n76 : n44) : (n87 ? !n76 : n44));
assign n477 = /* LUT   11  5  0 */ (n302 ? !\input_axis_tdata[0]  : \input_axis_tdata[0] );
assign n478 = /* LUT   12  2  1 */ (n276 ? (\input_axis_tdata[1]  ? 1'b1 : (input_axis_tvalid ? n2 : 1'b1)) : (\input_axis_tdata[1]  ? (input_axis_tvalid ? !n2 : 1'b0) : 1'b0));
assign n196 = /* LUT    8  8  4 */ (n4 ? (n195 ? !n54 : 1'b0) : (n195 ? 1'b1 : n54));
assign n217 = /* LUT    9  1  2 */ (n10 ? n214 : n143);
assign n480 = /* LUT   11  5  6 */ (n308 ? (\input_axis_tdata[6]  ? n5 : !n5) : (\input_axis_tdata[6]  ? !n5 : n5));
assign n481 = /* LUT    7  5  7 */ (n84 ? rst : (n83 ? rst : 1'b1));
assign n482 = /* LUT    8  5  4 */ (n167 ? (n83 ? 1'b1 : n153) : (n83 ? 1'b0 : n153));
assign n483 = /* LUT   12  2  3 */ (n278 ? (\input_axis_tdata[3]  ? 1'b1 : (input_axis_tvalid ? n2 : 1'b1)) : (\input_axis_tdata[3]  ? (input_axis_tvalid ? !n2 : 1'b0) : 1'b0));
assign n484 = /* LUT    8  8  2 */ (n4 ? (n194 ? (n101 ? n22 : 1'b1) : 1'b0) : (n194 ? (n101 ? n22 : 1'b0) : 1'b0));
assign n218 = /* LUT    9  1  4 */ (n10 ? n215 : n62);
assign n486 = /* LUT   11  5  4 */ (n306 ? (\input_axis_tdata[4]  ? n5 : !n5) : (\input_axis_tdata[4]  ? !n5 : n5));
assign n487 = /* LUT    8  5  6 */ (n159 ? (n83 ? 1'b1 : n165) : (n83 ? 1'b0 : n165));
assign n193 = /* LUT    8  8  0 */ (n104 ? 1'b1 : (n51 ? !n105 : n4));
assign n488 = /* LUT    9  1  6 */ (n123 ? 1'b1 : (n142 ? 1'b1 : (n124 ? 1'b1 : n125)));
assign n489 = /* LUT    7  3  1 */ (n2 ? (n29 ? 1'b0 : !n59) : input_axis_tvalid);
assign n490 = /* LUT    8 11  6 */ (n86 ? 1'b0 : (n4 ? n117 : 1'b0));
assign n491 = /* LUT    9  9  1 */ (n102 ? (n201 ? (n101 ? n198 : 1'b1) : (n101 ? n198 : 1'b0)) : 1'b0);
assign n492 = /* LUT    6  6  6 */ !n4;
assign n493 = /* LUT    7  5  3 */ (n71 ? (n83 ? 1'b1 : n41) : (n83 ? 1'b0 : n41));
assign n494 = /* LUT    8  5  0 */ (n157 ? (n83 ? 1'b1 : n39) : (n83 ? 1'b0 : n39));
assign n495 = /* LUT    7  6  3 */ (n84 ? (rst ? 1'b1 : (n83 ? n80 : 1'b0)) : 1'b1);
assign n496 = /* LUT   11  1  7 */ (n24 ? rst : (rst ? 1'b1 : (n10 ? !n60 : 1'b0)));
assign n497 = /* LUT    9  7  3 */ (n250 ? n100 : 1'b0);
assign n498 = /* LUT    7  3  3 */ (n31 ? (input_axis_tvalid ? !n2 : 1'b0) : (input_axis_tvalid ? (n2 ? !n59 : 1'b1) : (n2 ? !n59 : 1'b0)));
assign n144 = /* LUT    8  2  0 */ (n24 ? 1'b0 : (n60 ? !rst : 1'b0));
assign n114 = /* LUT    7  8  5 */ (n53 ? 1'b1 : (n111 ? 1'b1 : n52));
assign n499 = /* LUT    7  5  1 */ (n81 ? (n83 ? 1'b1 : n13) : (n83 ? 1'b0 : n13));
assign n500 = /* LUT    8  5  2 */ (n169 ? (n83 ? 1'b1 : n88) : (n83 ? 1'b0 : n88));
assign n273 = /* LUT   11  1  5 */ (n10 ? n249 : n260);
assign n502 = /* LUT    9  7  1 */ (n252 ? (n92 ? (n87 ? 1'b1 : n189) : (n87 ? 1'b0 : n189)) : (n92 ? (n87 ? 1'b0 : n189) : (n87 ? 1'b1 : n189)));
assign n503 = /* LUT    9  4  1 */ (n10 ? n229 : n231);
assign n504 = /* LUT    9  9  5 */ (n102 ? (n197 ? (n101 ? n200 : 1'b1) : (n101 ? n200 : 1'b0)) : 1'b0);
assign n505 = /* LUT    8  2  2 */ (n23 ? 1'b1 : (n28 ? 1'b1 : (n31 ? n33 : 1'b1)));
assign n320 = /* LUT   12  1  4 */ (n48 ? (n262 ? 1'b1 : n10) : (n262 ? !n10 : 1'b0));
assign n507 = /* LUT   11  1  3 */ (n24 ? n272 : (n272 ? (\input_axis_tdata[6]  ? 1'b1 : n60) : (\input_axis_tdata[6]  ? !n60 : 1'b0)));
assign n508 = /* LUT    9  7  7 */ (n227 ? n100 : 1'b0);
assign n509 = /* LUT   11  2  3 */ (n285 ? (n5 ? n129 : !n129) : (n5 ? !n129 : n129));
assign n510 = /* LUT    9  9  7 */ (n102 ? (n198 ? (n101 ? n202 : 1'b1) : (n101 ? n202 : 1'b0)) : 1'b0);
assign n511 = /* LUT    8  2  4 */ (input_axis_tvalid ? (n145 ? !n2 : 1'b1) : (n145 ? 1'b0 : n2));
assign n113 = /* LUT    7  8  1 */ (n100 ? (n112 ? (n51 ? rst : 1'b1) : 1'b0) : n112);
assign n321 = /* LUT   12  1  6 */ (n265 ? (n10 ? n251 : 1'b1) : (n10 ? n251 : 1'b0));
assign n224 = /* LUT    9  2  1 */ (n10 ? n147 : n221);
assign n514 = /* LUT    8  7  7 */ (n106 ? (n170 ? 1'b1 : !n83) : (n170 ? n83 : 1'b0));
assign n515 = /* LUT    9 12  4 */ n202;
assign n516 = /* LUT   11  1  1 */ (n24 ? n271 : (n271 ? (\input_axis_tdata[1]  ? 1'b1 : n60) : (\input_axis_tdata[1]  ? !n60 : 1'b0)));
assign n517 = /* LUT    9  7  5 */ (n251 ? n100 : 1'b0);
assign n518 = /* LUT   11  2  1 */ (n283 ? (n5 ? (n258 ? 1'b1 : n10) : (n258 ? n10 : 1'b1)) : (n5 ? (n258 ? n10 : 1'b1) : (n258 ? 1'b1 : n10)));
assign n519 = /* LUT    8  2  6 */ (n59 ? (n146 ? (input_axis_tvalid ? !n2 : 1'b0) : (input_axis_tvalid ? 1'b1 : n2)) : (input_axis_tvalid ? 1'b1 : n2));
assign n520 = /* LUT    7  8  3 */ (n80 ? (n14 ? 1'b0 : (n50 ? 1'b0 : n4)) : (n14 ? n50 : (n50 ? 1'b1 : n4)));
assign n521 = /* LUT   12  1  0 */ (n267 ? 1'b1 : (n268 ? 1'b1 : (n257 ? 1'b1 : n266)));
assign n225 = /* LUT    9  2  3 */ (n10 ? n223 : n222);
assign n523 = /* LUT    8  7  5 */ (n156 ? 1'b1 : !n83);
assign n524 = /* LUT    9 12  2 */ n197;
assign n525 = /* LUT   11  2  7 */ (n289 ? (n5 ? n136 : !n136) : (n5 ? !n136 : n136));
assign n526 = /* LUT   12  6  0 */ (n330 ? (\input_axis_tdata[0]  ? n5 : !n5) : (\input_axis_tdata[0]  ? !n5 : n5));
assign n527 = /* LUT    8  4  3 */ (n119 ? 1'b1 : (output_axis_tvalid ? !output_axis_tready : 1'b0));
assign n528 = /* LUT   12  1  2 */ (n24 ? n319 : (n319 ? (n60 ? 1'b1 : \input_axis_tdata[1] ) : (n60 ? 1'b0 : \input_axis_tdata[1] )));
assign n529 = /* LUT    5  1  0 */ input_axis_tvalid;
assign n226 = /* LUT    9  2  5 */ (n10 ? n47 : n219);
assign n531 = /* LUT    8  7  3 */ (n179 ? (n83 ? 1'b1 : n186) : (n83 ? 1'b0 : n186));
assign n532 = /* LUT    8 10  3 */ (n86 ? 1'b1 : (n204 ? rst : 1'b1));
assign n533 = /* LUT    9  5  4 */ (n236 ? (n36 ? (n87 ? 1'b1 : n192) : (n87 ? 1'b0 : n192)) : (n36 ? (n87 ? 1'b0 : n192) : (n87 ? 1'b1 : n192)));
assign n534 = /* LUT   11  2  5 */ (n287 ? (n5 ? n267 : !n267) : (n5 ? !n267 : n267));
assign n535 = /* LUT    8 13  3 */ n118;
assign n536 = /* LUT    6  1  1 */ (n2 ? rst : (rst ? 1'b1 : !n24));
assign n537 = /* LUT   12  6  2 */ (n332 ? (\input_axis_tdata[2]  ? n5 : !n5) : (\input_axis_tdata[2]  ? !n5 : n5));
assign n538 = /* LUT    9  3  6 */ (n24 ? n228 : (n228 ? (n60 ? 1'b1 : \input_axis_tdata[0] ) : (n60 ? 1'b0 : \input_axis_tdata[0] )));
assign n539 = /* LUT    8  7  1 */ (n171 ? (n83 ? 1'b1 : n109) : (n83 ? 1'b0 : n109));
assign n540 = /* LUT    9  5  6 */ (n238 ? (n79 ? (n87 ? 1'b1 : n187) : (n87 ? 1'b0 : n187)) : (n79 ? (n87 ? 1'b0 : n187) : (n87 ? 1'b1 : n187)));
assign n541 = /* LUT   12  6  4 */ (n334 ? (\input_axis_tdata[4]  ? n5 : !n5) : (\input_axis_tdata[4]  ? !n5 : n5));
assign n542 = /* LUT    9  3  4 */ (n24 ? n149 : (\input_axis_tdata[7]  ? (n149 ? 1'b1 : !n60) : (n149 ? n60 : 1'b0)));
assign n543 = /* LUT    9  5  0 */ (n232 ? (n155 ? (n84 ? n100 : 1'b0) : (n84 ? n100 : 1'b1)) : (n155 ? (n84 ? n100 : 1'b1) : (n84 ? n100 : 1'b0)));
assign n116 = /* LUT    7  9  2 */ (n53 ? !n14 : n14);
assign n545 = /* LUT    8  1  1 */ (n63 ? (n137 ? n135 : 1'b1) : (n137 ? n135 : 1'b0));
assign n546 = /* LUT   12  6  6 */ (n336 ? (\input_axis_tdata[6]  ? n5 : !n5) : (\input_axis_tdata[6]  ? !n5 : n5));
assign n547 = /* LUT    9  3  2 */ (n24 ? n148 : (\input_axis_tdata[5]  ? (n148 ? 1'b1 : !n60) : (n148 ? n60 : 1'b0)));
assign n548 = /* LUT    9  5  2 */ (n234 ? (n42 ? (n87 ? 1'b1 : n100) : (n87 ? 1'b0 : n100)) : (n42 ? (n87 ? 1'b0 : n100) : (n87 ? 1'b1 : n100)));
assign n549 = /* LUT   11  4  0 */ (n299 ? (n5 ? n142 : !n142) : (n5 ? !n142 : n142));
assign n115 = /* LUT    7  9  0 */ (n14 ? !n52 : (n53 ? !n52 : (n111 ? !n52 : n52)));
assign n138 = /* LUT    8  1  3 */ (n129 ? 1'b1 : (n70 ? 1'b1 : (n132 ? 1'b1 : n134)));
assign n552 = /* LUT    7  7  4 */ (n100 ? n48 : 1'b0);
assign n553 = /* LUT   11  3  0 */ (n290 ? (n5 ? n268 : !n268) : (n5 ? !n268 : n268));
assign n554 = /* LUT    7  2  7 */ (n31 ? 1'b1 : n23);
assign n555 = /* LUT   11  4  2 */ (n301 ? (n70 ? n5 : !n5) : (n70 ? !n5 : n5));
assign n556 = /* LUT    8  1  5 */ (n130 ? 1'b1 : (n139 ? 1'b1 : (n128 ? 1'b1 : n126)));
assign n557 = /* LUT    7  9  6 */ (n53 ? n52 : (n111 ? n52 : 1'b0));
assign n558 = /* LUT    9 13  7 */ n199;
assign n175 = /* LUT    8  6  4 */ (n35 ? 1'b1 : (n37 ? 1'b1 : (n36 ? 1'b1 : n155)));
assign n560 = /* LUT   11  3  2 */ (n293 ? (n5 ? n132 : !n132) : (n5 ? !n132 : n132));
assign n296 = /* CARRY 11  3  4 */ (n254 & n5) | ((n254 | n5) & n295);
assign n318 = /* CARRY 11  6  7 */ (n5 & \input_axis_tdata[7] ) | ((n5 | \input_axis_tdata[7] ) & n317);
assign n324 = /* CARRY 12  5  1 */ (n5 & \input_axis_tdata[1] ) | ((n5 | \input_axis_tdata[1] ) & n323);
assign n246 = /* CARRY  9  6  5 */ (n87 & n90) | ((n87 | n90) & n245);
assign n298 = /* CARRY 11  3  6 */ (n133 & n5) | ((n133 | n5) & n297);
assign n316 = /* CARRY 11  6  5 */ (n5 & \input_axis_tdata[5] ) | ((n5 | \input_axis_tdata[5] ) & n315);
assign n326 = /* CARRY 12  5  3 */ (n5 & \input_axis_tdata[3] ) | ((n5 | \input_axis_tdata[3] ) & n325);
assign n248 = /* CARRY  9  6  7 */ (n87 & n91) | ((n87 | n91) & n247);
assign n306 = /* CARRY 11  5  3 */ (n5 & \input_axis_tdata[3] ) | ((n5 | \input_axis_tdata[3] ) & n305);
assign n314 = /* CARRY 11  6  3 */ (n5 & \input_axis_tdata[3] ) | ((n5 | \input_axis_tdata[3] ) & n313);
assign n328 = /* CARRY 12  5  5 */ (n5 & \input_axis_tdata[5] ) | ((n5 | \input_axis_tdata[5] ) & n327);
assign n242 = /* CARRY  9  6  1 */ (n87 & n77) | ((n87 | n77) & n241);
assign n304 = /* CARRY 11  5  1 */ (n5 & \input_axis_tdata[1] ) | ((n5 | \input_axis_tdata[1] ) & n303);
assign n312 = /* CARRY 11  6  1 */ (n5 & \input_axis_tdata[1] ) | ((n5 | \input_axis_tdata[1] ) & n311);
assign n330 = /* CARRY 12  5  7 */ (n5 & \input_axis_tdata[7] ) | ((n5 | \input_axis_tdata[7] ) & n329);
assign n244 = /* CARRY  9  6  3 */ (n87 & n75) | ((n87 | n75) & n243);
assign n310 = /* CARRY 11  5  7 */ (n5 & \input_axis_tdata[7] ) | ((n5 | \input_axis_tdata[7] ) & n309);
assign n308 = /* CARRY 11  5  5 */ (n5 & \input_axis_tdata[5] ) | ((n5 | \input_axis_tdata[5] ) & n307);
assign n252 = /* CARRY  9  7  0 */ (n93 & n87) | ((n93 | n87) & n248);
assign n285 = /* CARRY 11  2  2 */ (n259 & n5) | ((n259 | n5) & n284);
assign n283 = /* CARRY 11  2  0 */ (n257 & 1'b0) | ((n257 | 1'b0) & n282);
assign n289 = /* CARRY 11  2  6 */ (n5 & n134) | ((n5 | n134) & n288);
assign n332 = /* CARRY 12  6  1 */ (n5 & \input_axis_tdata[1] ) | ((n5 | \input_axis_tdata[1] ) & n331);
assign n238 = /* CARRY  9  5  5 */ (n35 & n87) | ((n35 | n87) & n237);
assign n287 = /* CARRY 11  2  4 */ (n5 & n266) | ((n5 | n266) & n286);
assign n334 = /* CARRY 12  6  3 */ (n5 & \input_axis_tdata[3] ) | ((n5 | \input_axis_tdata[3] ) & n333);
assign n240 = /* CARRY  9  5  7 */ (n78 & n87) | ((n78 | n87) & n239);
assign n336 = /* CARRY 12  6  5 */ (n5 & \input_axis_tdata[5] ) | ((n5 | \input_axis_tdata[5] ) & n335);
assign n234 = /* CARRY  9  5  1 */ (n94 & n87) | ((n94 | n87) & n233);
assign n236 = /* CARRY  9  5  3 */ (n72 & n87) | ((n72 | n87) & n235);
assign n293 = /* CARRY 11  3  1 */ (n5 & n255) | ((n5 | n255) & n292);
assign n301 = /* CARRY 11  4  1 */ (n5 & n125) | ((n5 | n125) & n300);
assign n295 = /* CARRY 11  3  3 */ (n5 & n131) | ((n5 | n131) & n294);
assign n297 = /* CARRY 11  3  5 */ (n5 & n123) | ((n5 | n123) & n296);
assign n317 = /* CARRY 11  6  6 */ (n5 & \input_axis_tdata[6] ) | ((n5 | \input_axis_tdata[6] ) & n316);
assign n323 = /* CARRY 12  5  0 */ (\input_axis_tdata[0]  & 1'b0) | ((\input_axis_tdata[0]  | 1'b0) & n322);
assign n245 = /* CARRY  9  6  4 */ (n96 & n87) | ((n96 | n87) & n244);
assign n299 = /* CARRY 11  3  7 */ (n5 & n124) | ((n5 | n124) & n298);
assign n315 = /* CARRY 11  6  4 */ (n5 & \input_axis_tdata[4] ) | ((n5 | \input_axis_tdata[4] ) & n314);
assign n325 = /* CARRY 12  5  2 */ (n5 & \input_axis_tdata[2] ) | ((n5 | \input_axis_tdata[2] ) & n324);
assign n247 = /* CARRY  9  6  6 */ (n74 & n87) | ((n74 | n87) & n246);
assign n313 = /* CARRY 11  6  2 */ (n5 & \input_axis_tdata[2] ) | ((n5 | \input_axis_tdata[2] ) & n312);
assign n327 = /* CARRY 12  5  4 */ (n5 & \input_axis_tdata[4] ) | ((n5 | \input_axis_tdata[4] ) & n326);
assign n241 = /* CARRY  9  6  0 */ (n37 & n87) | ((n37 | n87) & n240);
assign n305 = /* CARRY 11  5  2 */ (n5 & \input_axis_tdata[2] ) | ((n5 | \input_axis_tdata[2] ) & n304);
assign n311 = /* CARRY 11  6  0 */ (n5 & \input_axis_tdata[0] ) | ((n5 | \input_axis_tdata[0] ) & n310);
assign n329 = /* CARRY 12  5  6 */ (n5 & \input_axis_tdata[6] ) | ((n5 | \input_axis_tdata[6] ) & n328);
assign n243 = /* CARRY  9  6  2 */ (n76 & n87) | ((n76 | n87) & n242);
assign n303 = /* CARRY 11  5  0 */ (\input_axis_tdata[0]  & 1'b0) | ((\input_axis_tdata[0]  | 1'b0) & n302);
assign n309 = /* CARRY 11  5  6 */ (n5 & \input_axis_tdata[6] ) | ((n5 | \input_axis_tdata[6] ) & n308);
assign n307 = /* CARRY 11  5  4 */ (n5 & \input_axis_tdata[4] ) | ((n5 | \input_axis_tdata[4] ) & n306);
assign n253 = /* CARRY  9  7  1 */ (n87 & n92) | ((n87 | n92) & n252);
assign n286 = /* CARRY 11  2  3 */ (n129 & n5) | ((n129 | n5) & n285);
assign n284 = /* CARRY 11  2  1 */ (n258 & n5) | ((n258 | n5) & n283);
assign n290 = /* CARRY 11  2  7 */ (n136 & n5) | ((n136 | n5) & n289);
assign n331 = /* CARRY 12  6  0 */ (n5 & \input_axis_tdata[0] ) | ((n5 | \input_axis_tdata[0] ) & n330);
assign n237 = /* CARRY  9  5  4 */ (n87 & n36) | ((n87 | n36) & n236);
assign n288 = /* CARRY 11  2  5 */ (n267 & n5) | ((n267 | n5) & n287);
assign n333 = /* CARRY 12  6  2 */ (n5 & \input_axis_tdata[2] ) | ((n5 | \input_axis_tdata[2] ) & n332);
assign n239 = /* CARRY  9  5  6 */ (n87 & n79) | ((n87 | n79) & n238);
assign n335 = /* CARRY 12  6  4 */ (n5 & \input_axis_tdata[4] ) | ((n5 | \input_axis_tdata[4] ) & n334);
assign n233 = /* CARRY  9  5  0 */ (n84 & n155) | ((n84 | n155) & n232);
assign n337 = /* CARRY 12  6  6 */ (n5 & \input_axis_tdata[6] ) | ((n5 | \input_axis_tdata[6] ) & n336);
assign n235 = /* CARRY  9  5  2 */ (n87 & n42) | ((n87 | n42) & n234);
assign n300 = /* CARRY 11  4  0 */ (n142 & n5) | ((n142 | n5) & n299);
assign n292 = /* CARRY 11  3  0 */ (n268 & n5) | ((n268 | n5) & n290);
assign n294 = /* CARRY 11  3  2 */ (n132 & n5) | ((n132 | n5) & n293);
/* FF  8  6  6 */ assign n84 = n177;
/* FF  8  9  0 */ always @(posedge clk) if (n45) n111 <= n46 ? 1'b0 : n338;
/* FF  7  2  3 */ assign n2 = n66;
/* FF 11  3  4 */ assign n263 = n339;
/* FF 11  6  7 */ assign n186 = n340;
/* FF 12  5  1 */ assign n40 = n341;
/* FF  9  8  3 */ assign n189 = n342;
/* FF  6  7  2 */ assign n5 = n343;
/* FF  8  6  0 */ assign n83 = n344;
/* FF  9 13  3 */ always @(posedge clk) if (n120) \output_axis_tdata[1]  <= rst ? 1'b0 : n345;
/* FF  7  1  1 */ always @(posedge clk) if (n25) n23 <= n26 ? 1'b0 : n346;
/* FF  9  6  5 */ assign n171 = n347;
/* FF  7  2  1 */ assign n25 = n65;
/* FF  8 12  4 */ assign n120 = n348;
/* FF 11  3  6 */ assign n63 = n349;
/* FF 11  6  5 */ assign n108 = n350;
/* FF  8  3  0 */ assign n67 = n351;
/* FF 12  5  3 */ assign n147 = n352;
/* FF  9  8  1 */ assign n187 = n353;
/* FF  8  6  2 */ assign n354 = n174;
/* FF  9  6  7 */ assign n172 = n355;
/* FF 11  5  3 */ assign n13 = n356;
/* FF 11  6  3 */ assign n109 = n357;
/* FF  8  3  6 */ assign n34 = n358;
/* FF 12  5  5 */ assign n251 = n359;
/* FF  9  8  7 */ assign n192 = n360;
/* FF 12  2  4 */ always @(posedge clk) if (n56) n278 <= 1'b0 ? 1'b0 : n361;
/* FF  9  1  1 */ always @(posedge clk) if (n127) n123 <= rst ? 1'b0 : n362;
/* FF  8  8  7 */ assign n105 = n363;
/* FF  9  6  1 */ assign n166 = n364;
/* FF 11  5  1 */ assign n39 = n365;
/* FF 11  6  1 */ assign n154 = n366;
/* FF 12  5  7 */ assign n47 = n367;
/* FF  9  8  5 */ assign n190 = n368;
/* FF 12  2  6 */ always @(posedge clk) if (n56) n280 <= 1'b0 ? 1'b0 : n369;
/* FF  8  8  5 */ assign n80 = n370;
/* FF  9  1  3 */ always @(posedge clk) if (n127) n124 <= rst ? 1'b0 : n371;
/* FF  9  6  3 */ assign n168 = n372;
/* FF 11  5  7 */ assign n164 = n373;
/* FF  7  2  5 */ always @(posedge clk) if (1'b1) n28 <= 1'b0 ? 1'b0 : n374;
/* FF 12  2  0 */ always @(posedge clk) if (n56) n274 <= 1'b0 ? 1'b0 : n375;
/* FF  9  1  5 */ always @(posedge clk) if (n127) n125 <= rst ? 1'b0 : n376;
/* FF  8  8  3 */ assign n103 = n195;
/* FF 11  5  5 */ assign n165 = n377;
/* FF  7  5  6 */ assign n19 = n378;
/* FF  8  5  5 */ always @(posedge clk) if (n38) n77 <= rst ? 1'b0 : n379;
/* FF 12  2  2 */ always @(posedge clk) if (n56) n276 <= 1'b0 ? 1'b0 : n380;
/* FF  9  1  7 */ assign n127 = n381;
/* FF  8  8  1 */ assign n102 = n194;
/* FF  9  4  4 */ assign n149 = n382;
/* FF  8  5  7 */ always @(posedge clk) if (n38) n79 <= rst ? 1'b0 : n383;
/* FF  9  9  0 */ always @(posedge clk) if (1'b1) n197 <= 1'b0 ? 1'b0 : n384;
/* FF  8  2  1 */ always @(posedge clk) if (1'b1) n57 <= 1'b0 ? 1'b0 : n385;
/* FF  7  5  2 */ always @(posedge clk) if (n38) n36 <= rst ? 1'b0 : n386;
/* FF  8  5  1 */ always @(posedge clk) if (n38) n73 <= rst ? 1'b0 : n387;
/* FF 11  1  6 */ always @(posedge clk) if (n127) n129 <= rst ? 1'b0 : n388;
/* FF  9  7  2 */ assign n162 = n389;
/* FF  9  9  2 */ always @(posedge clk) if (1'b1) n199 <= 1'b0 ? 1'b0 : n390;
/* FF  7  8  6 */ assign n51 = n391;
/* FF  8  2  3 */ assign n59 = n145;
/* FF  8  5  3 */ always @(posedge clk) if (n38) n75 <= rst ? 1'b0 : n392;
/* FF  7  6  6 */ assign n21 = n393;
/* FF  9  7  0 */ assign n178 = n394;
/* FF 11  1  4 */ assign n130 = n395;
/* FF 11  2  2 */ always @(posedge clk) if (n127) n259 <= n256 ? 1'b0 : n396;
/* FF 11  7  0 */ assign n161 = n397;
/* FF  7  8  0 */ assign n45 = n112;
/* FF  8  2  5 */ assign n398 = n146;
/* FF 12  1  5 */ always @(posedge clk) if (n127) n267 <= rst ? 1'b0 : n399;
/* FF  9  2  0 */ always @(posedge clk) if (n127) n133 <= rst ? 1'b0 : n400;
/* FF  8  7  6 */ assign n95 = n401;
/* FF 11  1  2 */ assign n402 = n272;
/* FF  9  7  6 */ assign n183 = n403;
/* FF 11  2  0 */ always @(posedge clk) if (n127) n257 <= n256 ? 1'b0 : n404;
/* FF  9  9  6 */ always @(posedge clk) if (1'b1) n201 <= 1'b0 ? 1'b0 : n405;
/* FF  7  8  2 */ always @(posedge clk) if (1'b1) n14 <= 1'b0 ? 1'b0 : n406;
/* FF 12  1  7 */ always @(posedge clk) if (n127) n268 <= rst ? 1'b0 : n407;
/* FF  9  2  2 */ always @(posedge clk) if (n127) n134 <= rst ? 1'b0 : n408;
/* FF  8  7  4 */ always @(posedge clk) if (n38) n93 <= rst ? 1'b0 : n409;
/* FF  9 12  5 */ always @(posedge clk) if (n120) \output_axis_tdata[5]  <= rst ? 1'b0 : n410;
/* FF 11  1  0 */ assign n411 = n271;
/* FF  9  7  4 */ assign n181 = n412;
/* FF 11  2  6 */ assign n221 = n413;
/* FF 12  6  1 */ assign n269 = n414;
/* FF 12  1  1 */ assign n415 = n319;
/* FF  9 12  3 */ always @(posedge clk) if (n120) \output_axis_tdata[7]  <= rst ? 1'b0 : n416;
/* FF  9  2  4 */ always @(posedge clk) if (n127) n136 <= rst ? 1'b0 : n417;
/* FF  8  7  2 */ always @(posedge clk) if (n38) n91 <= rst ? 1'b0 : n418;
/* FF  9  5  5 */ assign n81 = n419;
/* FF 11  2  4 */ assign n261 = n420;
/* FF  6  1  0 */ assign n15 = n421;
/* FF 12  6  3 */ assign n135 = n422;
/* FF  9 12  1 */ always @(posedge clk) if (n120) \output_axis_tdata[6]  <= rst ? 1'b0 : n423;
/* FF  9  2  6 */ always @(posedge clk) if (n127) n132 <= rst ? 1'b0 : n424;
/* FF  8  7  0 */ assign n89 = n425;
/* FF  8 10  2 */ assign n117 = n204;
/* FF  9  5  7 */ assign n159 = n426;
/* FF  6  2  0 */ always @(posedge clk) if (n15) input_axis_tready <= n17 ? 1'b0 : n427;
/* FF 12  6  5 */ assign n229 = n428;
/* FF  9  3  5 */ assign n429 = n228;
/* FF  7  7  1 */ always @(posedge clk) if (n38) n42 <= rst ? 1'b0 : n430;
/* FF  9  5  1 */ assign n156 = n431;
/* FF  7  9  3 */ always @(posedge clk) if (n45) n53 <= rst ? 1'b0 : n432;
/* FF  8  1  0 */ assign n10 = n137;
/* FF  6  1  4 */ assign n17 = n433;
/* FF 12  6  7 */ assign n230 = n434;
/* FF  8 10  6 */ always @(posedge clk) if (1'b1) n118 <= 1'b0 ? 1'b0 : n435;
/* FF  9  5  3 */ assign n157 = n436;
/* FF  9 10  3 */ always @(posedge clk) if (1'b1) rx_frame_error <= n110 ? 1'b0 : n437;
/* FF  7  9  1 */ always @(posedge clk) if (n45) n52 <= rst ? 1'b0 : n438;
/* FF 11  3  1 */ assign n264 = n439;
/* FF  7  2  6 */ assign n29 = n440;
/* FF 11  4  1 */ assign n62 = n441;
/* FF  8  1  4 */ assign n442 = n139;
/* FF  8  6  5 */ assign n86 = n176;
/* FF 12  3  0 */ always @(posedge clk) if (n34) txd <= rst ? 1'b1 : n443;
/* FF  7  7  7 */ assign n44 = n444;
/* FF 11  3  3 */ assign n151 = n445;
/* FF  7  2  4 */ assign n27 = n446;
/* FF  8  6  7 */ assign n87 = n447;
/* FF  7  2  2 */ assign n26 = n448;
/* FF 11  3  5 */ assign n141 = n449;
/* FF 11  6  6 */ assign n107 = n450;
/* FF  9  8  2 */ assign n188 = n451;
/* FF 12  5  0 */ assign n249 = n452;
/* FF  9  6  4 */ assign n170 = n453;
/* FF 11  3  7 */ assign n143 = n454;
/* FF  7  2  0 */ assign n455 = n64;
/* FF 11  6  4 */ assign n88 = n456;
/* FF 12  5  2 */ assign n48 = n457;
/* FF 11  8  1 */ assign n97 = n458;
/* FF  9  8  0 */ assign n185 = n459;
/* FF  8  6  3 */ assign n85 = n460;
/* FF  9  6  6 */ assign n169 = n461;
/* FF 11  6  2 */ assign n106 = n462;
/* FF 12  5  4 */ assign n223 = n463;
/* FF  9  8  6 */ assign n191 = n464;
/* FF 12  2  5 */ always @(posedge clk) if (n56) n279 <= 1'b0 ? 1'b0 : n465;
/* FF  7  4  0 */ always @(posedge clk) if (1'b1) rx_overrun_error <= n67 ? 1'b0 : n466;
/* FF  9  6  0 */ assign n71 = n467;
/* FF  8 14  4 */ always @(posedge clk) if (1'b1) n4 <= rst ? 1'b1 : n468;
/* FF 11  5  2 */ assign n18 = n469;
/* FF 11  6  0 */ assign n153 = n470;
/* FF 12  5  6 */ assign n250 = n471;
/* FF  9  8  4 */ assign n173 = n472;
/* FF 12  2  7 */ always @(posedge clk) if (n56) n281 <= 1'b0 ? 1'b0 : n473;
/* FF  8  8  6 */ assign n104 = n474;
/* FF  9  1  0 */ assign n475 = n216;
/* FF  9  6  2 */ assign n167 = n476;
/* FF 11  5  0 */ assign n99 = n477;
/* FF 12  2  1 */ always @(posedge clk) if (n56) n275 <= 1'b0 ? 1'b0 : n478;
/* FF  8  8  4 */ assign n100 = n196;
/* FF  9  1  2 */ assign n479 = n217;
/* FF 11  5  6 */ assign n41 = n480;
/* FF  7  5  7 */ assign n20 = n481;
/* FF  8  5  4 */ always @(posedge clk) if (n38) n76 <= rst ? 1'b0 : n482;
/* FF 12  2  3 */ always @(posedge clk) if (n56) n277 <= 1'b0 ? 1'b0 : n483;
/* FF  8  8  2 */ always @(posedge clk) if (1'b1) n22 <= 1'b0 ? 1'b0 : n484;
/* FF  9  1  4 */ assign n485 = n218;
/* FF 11  5  4 */ assign n163 = n486;
/* FF  8  5  6 */ always @(posedge clk) if (n38) n78 <= rst ? 1'b0 : n487;
/* FF  8  8  0 */ assign n101 = n193;
/* FF  9  1  6 */ assign n126 = n488;
/* FF  7  3  1 */ always @(posedge clk) if (n25) n33 <= rst ? 1'b0 : n489;
/* FF  8 11  6 */ assign n119 = n490;
/* FF  9  9  1 */ always @(posedge clk) if (1'b1) n198 <= 1'b0 ? 1'b0 : n491;
/* FF  6  6  6 */ always @(posedge clk) if (n21) rx_busy <= rst ? 1'b0 : n492;
/* FF  7  5  3 */ always @(posedge clk) if (n38) n37 <= rst ? 1'b0 : n493;
/* FF  8  5  0 */ always @(posedge clk) if (n38) n72 <= rst ? 1'b0 : n494;
/* FF  7  6  3 */ assign n38 = n495;
/* FF 11  1  7 */ assign n256 = n496;
/* FF  9  7  3 */ assign n180 = n497;
/* FF  7  3  3 */ always @(posedge clk) if (n25) n31 <= rst ? 1'b0 : n498;
/* FF  8  2  0 */ assign n56 = n144;
/* FF  7  8  5 */ assign n50 = n114;
/* FF  7  5  1 */ always @(posedge clk) if (n38) n35 <= rst ? 1'b0 : n499;
/* FF  8  5  2 */ always @(posedge clk) if (n38) n74 <= rst ? 1'b0 : n500;
/* FF 11  1  5 */ assign n501 = n273;
/* FF  9  7  1 */ assign n179 = n502;
/* FF  9  4  1 */ assign n148 = n503;
/* FF  9  9  5 */ always @(posedge clk) if (1'b1) n200 <= 1'b0 ? 1'b0 : n504;
/* FF  8  2  2 */ assign n58 = n505;
/* FF 12  1  4 */ assign n506 = n320;
/* FF 11  1  3 */ always @(posedge clk) if (n127) n255 <= rst ? 1'b0 : n507;
/* FF  9  7  7 */ assign n184 = n508;
/* FF 11  2  3 */ assign n260 = n509;
/* FF  9  9  7 */ always @(posedge clk) if (1'b1) n202 <= 1'b0 ? 1'b0 : n510;
/* FF  8  2  4 */ assign n60 = n511;
/* FF  7  8  1 */ assign n46 = n113;
/* FF 12  1  6 */ assign n512 = n321;
/* FF  9  2  1 */ assign n513 = n224;
/* FF  8  7  7 */ always @(posedge clk) if (n38) n96 <= rst ? 1'b0 : n514;
/* FF  9 12  4 */ always @(posedge clk) if (n120) \output_axis_tdata[4]  <= rst ? 1'b0 : n515;
/* FF 11  1  1 */ always @(posedge clk) if (n127) n254 <= rst ? 1'b0 : n516;
/* FF  9  7  5 */ assign n182 = n517;
/* FF 11  2  1 */ always @(posedge clk) if (n127) n258 <= n256 ? 1'b0 : n518;
/* FF  8  2  6 */ assign n61 = n519;
/* FF  7  8  3 */ assign n49 = n520;
/* FF 12  1  0 */ assign n128 = n521;
/* FF  9  2  3 */ assign n522 = n225;
/* FF  8  7  5 */ always @(posedge clk) if (n38) n94 <= rst ? 1'b0 : n523;
/* FF  9 12  2 */ always @(posedge clk) if (n120) \output_axis_tdata[2]  <= rst ? 1'b0 : n524;
/* FF 11  2  7 */ assign n222 = n525;
/* FF 12  6  0 */ assign n227 = n526;
/* FF  8  4  3 */ always @(posedge clk) if (1'b1) output_axis_tvalid <= rst ? 1'b0 : n527;
/* FF 12  1  2 */ always @(posedge clk) if (n127) n266 <= rst ? 1'b0 : n528;
/* FF  5  1  0 */ always @(posedge clk) if (n16) tx_busy <= rst ? 1'b0 : n529;
/* FF  9  2  5 */ assign n530 = n226;
/* FF  8  7  3 */ always @(posedge clk) if (n38) n92 <= rst ? 1'b0 : n531;
/* FF  8 10  3 */ assign n110 = n532;
/* FF  9  5  4 */ assign n82 = n533;
/* FF 11  2  5 */ assign n262 = n534;
/* FF  8 13  3 */ always @(posedge clk) if (n120) \output_axis_tdata[0]  <= rst ? 1'b0 : n535;
/* FF  6  1  1 */ assign n16 = n536;
/* FF 12  6  2 */ assign n140 = n537;
/* FF  9  3  6 */ always @(posedge clk) if (n127) n131 <= rst ? 1'b0 : n538;
/* FF  8  7  1 */ always @(posedge clk) if (n38) n90 <= rst ? 1'b0 : n539;
/* FF  9  5  6 */ assign n158 = n540;
/* FF 12  6  4 */ assign n214 = n541;
/* FF  9  3  4 */ always @(posedge clk) if (n127) n70 <= rst ? 1'b0 : n542;
/* FF  9  5  0 */ always @(posedge clk) if (n19) n155 <= n20 ? 1'b0 : n543;
/* FF  7  9  2 */ assign n544 = n116;
/* FF  8  1  1 */ assign n55 = n545;
/* FF 12  6  6 */ assign n215 = n546;
/* FF  9  3  2 */ always @(posedge clk) if (n127) n142 <= rst ? 1'b0 : n547;
/* FF  9  5  2 */ assign n98 = n548;
/* FF 11  4  0 */ assign n231 = n549;
/* FF  7  9  0 */ assign n550 = n115;
/* FF  8  1  3 */ assign n551 = n138;
/* FF  7  7  4 */ assign n43 = n552;
/* FF 11  3  0 */ assign n265 = n553;
/* FF  7  2  7 */ assign n30 = n554;
/* FF 11  4  2 */ assign n160 = n555;
/* FF  8  1  5 */ assign n24 = n556;
/* FF  7  9  6 */ assign n54 = n557;
/* FF  9 13  7 */ always @(posedge clk) if (n120) \output_axis_tdata[3]  <= rst ? 1'b0 : n558;
/* FF  8  6  4 */ assign n559 = n175;
/* FF 11  3  2 */ assign n219 = n560;

endmodule

