module top(
  input [3:0] alu_op,
  input [31:0] op1,
  input [31:0] op2,
  output [31:0] result,
  output zero
  );
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_A;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_A1;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_A2;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_A3;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_A4;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_A5;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_A6;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_AO5;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_AO6;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_A_CY;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_A_XOR;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_B;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_B1;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_B2;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_B3;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_B4;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_B5;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_B6;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_BO5;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_BO6;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_B_CY;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_B_XOR;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_C;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_C1;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_C2;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_C3;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_C4;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_C5;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_C6;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_CO5;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_CO6;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_C_CY;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_C_XOR;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_D;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_D1;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_D2;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_D3;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_D4;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_D5;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_D6;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_DO5;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_DO6;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_D_CY;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X50Y114_D_XOR;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_A;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_A1;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_A2;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_A3;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_A4;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_A5;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_A6;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_AO5;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_AO6;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_A_CY;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_A_XOR;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_B;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_B1;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_B2;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_B3;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_B4;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_B5;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_B6;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_BO5;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_BO6;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_B_CY;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_B_XOR;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_C;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_C1;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_C2;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_C3;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_C4;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_C5;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_C6;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_CO5;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_CO6;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_C_CY;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_C_XOR;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_D;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_D1;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_D2;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_D3;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_D4;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_D5;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_D6;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_DO5;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_DO6;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_D_CY;
  wire [0:0] CLBLL_L_X34Y114_SLICE_X51Y114_D_XOR;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_A;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_A1;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_A2;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_A3;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_A4;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_A5;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_A6;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_AMUX;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_AO5;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_AO6;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_A_CY;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_A_XOR;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_B;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_B1;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_B2;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_B3;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_B4;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_B5;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_B6;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_BO5;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_BO6;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_B_CY;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_B_XOR;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_C;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_C1;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_C2;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_C3;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_C4;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_C5;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_C6;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_CO5;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_CO6;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_C_CY;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_C_XOR;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_D;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_D1;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_D2;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_D3;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_D4;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_D5;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_D6;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_DO5;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_DO6;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_D_CY;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X50Y115_D_XOR;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_A;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_A1;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_A2;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_A3;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_A4;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_A5;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_A6;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_AO5;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_AO6;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_A_CY;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_A_XOR;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_B;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_B1;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_B2;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_B3;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_B4;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_B5;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_B6;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_BO5;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_BO6;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_B_CY;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_B_XOR;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_C;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_C1;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_C2;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_C3;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_C4;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_C5;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_C6;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_CO5;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_CO6;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_C_CY;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_C_XOR;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_D;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_D1;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_D2;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_D3;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_D4;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_D5;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_D6;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_DO5;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_DO6;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_D_CY;
  wire [0:0] CLBLL_L_X34Y115_SLICE_X51Y115_D_XOR;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_A;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_A1;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_A2;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_A3;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_A4;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_A5;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_A6;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_AMUX;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_AO5;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_AO6;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_A_CY;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_A_XOR;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_B;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_B1;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_B2;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_B3;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_B4;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_B5;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_B6;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_BO5;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_BO6;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_B_CY;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_B_XOR;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_C;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_C1;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_C2;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_C3;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_C4;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_C5;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_C6;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_CO5;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_CO6;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_C_CY;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_C_XOR;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_D;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_D1;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_D2;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_D3;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_D4;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_D5;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_D6;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_DO5;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_DO6;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_D_CY;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X50Y116_D_XOR;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_A;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_A1;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_A2;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_A3;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_A4;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_A5;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_A6;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_AMUX;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_AO5;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_AO6;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_A_CY;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_A_XOR;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_B;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_B1;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_B2;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_B3;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_B4;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_B5;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_B6;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_BO5;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_BO6;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_B_CY;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_B_XOR;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_C;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_C1;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_C2;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_C3;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_C4;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_C5;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_C6;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_CO5;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_CO6;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_C_CY;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_C_XOR;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_D;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_D1;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_D2;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_D3;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_D4;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_D5;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_D6;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_DO5;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_DO6;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_D_CY;
  wire [0:0] CLBLL_L_X34Y116_SLICE_X51Y116_D_XOR;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_A;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_A1;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_A2;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_A3;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_A4;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_A5;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_A6;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_AO5;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_AO6;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_A_CY;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_A_XOR;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_B;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_B1;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_B2;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_B3;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_B4;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_B5;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_B6;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_BO5;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_BO6;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_B_CY;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_B_XOR;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_C;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_C1;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_C2;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_C3;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_C4;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_C5;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_C6;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_CO5;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_CO6;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_C_CY;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_C_XOR;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_D;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_D1;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_D2;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_D3;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_D4;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_D5;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_D6;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_DO5;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_DO6;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_D_CY;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X50Y117_D_XOR;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_A;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_A1;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_A2;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_A3;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_A4;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_A5;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_A6;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_AO5;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_AO6;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_A_CY;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_A_XOR;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_B;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_B1;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_B2;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_B3;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_B4;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_B5;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_B6;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_BMUX;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_BO5;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_BO6;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_B_CY;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_B_XOR;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_C;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_C1;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_C2;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_C3;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_C4;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_C5;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_C6;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_CO5;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_CO6;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_C_CY;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_C_XOR;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_D;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_D1;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_D2;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_D3;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_D4;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_D5;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_D6;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_DO5;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_DO6;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_D_CY;
  wire [0:0] CLBLL_L_X34Y117_SLICE_X51Y117_D_XOR;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_A;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_A1;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_A2;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_A3;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_A4;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_A5;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_A6;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_AO5;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_AO6;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_A_CY;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_A_XOR;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_B;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_B1;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_B2;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_B3;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_B4;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_B5;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_B6;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_BO5;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_BO6;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_B_CY;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_B_XOR;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_C;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_C1;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_C2;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_C3;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_C4;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_C5;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_C6;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_CO5;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_CO6;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_C_CY;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_C_XOR;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_D;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_D1;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_D2;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_D3;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_D4;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_D5;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_D6;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_DO5;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_DO6;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_D_CY;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X50Y118_D_XOR;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_A;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_A1;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_A2;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_A3;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_A4;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_A5;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_A6;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_AO5;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_AO6;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_A_CY;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_A_XOR;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_B;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_B1;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_B2;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_B3;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_B4;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_B5;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_B6;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_BO5;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_BO6;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_B_CY;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_B_XOR;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_C;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_C1;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_C2;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_C3;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_C4;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_C5;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_C6;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_CO5;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_CO6;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_C_CY;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_C_XOR;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_D;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_D1;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_D2;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_D3;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_D4;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_D5;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_D6;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_DO5;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_DO6;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_D_CY;
  wire [0:0] CLBLL_L_X34Y118_SLICE_X51Y118_D_XOR;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_A;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_A1;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_A2;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_A3;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_A4;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_A5;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_A6;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_AO5;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_AO6;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_A_CY;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_A_XOR;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_B;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_B1;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_B2;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_B3;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_B4;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_B5;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_B6;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_BO5;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_BO6;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_B_CY;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_B_XOR;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_C;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_C1;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_C2;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_C3;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_C4;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_C5;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_C6;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_CO5;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_CO6;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_C_CY;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_C_XOR;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_D;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_D1;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_D2;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_D3;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_D4;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_D5;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_D6;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_DO5;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_DO6;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_D_CY;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X50Y119_D_XOR;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_A;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_A1;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_A2;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_A3;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_A4;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_A5;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_A6;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_AMUX;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_AO5;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_AO6;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_A_CY;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_A_XOR;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_B;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_B1;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_B2;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_B3;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_B4;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_B5;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_B6;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_BO5;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_BO6;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_B_CY;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_B_XOR;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_C;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_C1;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_C2;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_C3;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_C4;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_C5;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_C6;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_CMUX;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_CO5;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_CO6;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_C_CY;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_C_XOR;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_D;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_D1;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_D2;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_D3;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_D4;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_D5;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_D6;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_DO5;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_DO6;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_D_CY;
  wire [0:0] CLBLL_L_X34Y119_SLICE_X51Y119_D_XOR;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_A;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_A1;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_A2;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_A3;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_A4;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_A5;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_A6;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_AO5;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_AO6;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_A_CY;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_A_XOR;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_B;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_B1;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_B2;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_B3;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_B4;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_B5;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_B6;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_BO5;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_BO6;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_B_CY;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_B_XOR;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_C;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_C1;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_C2;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_C3;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_C4;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_C5;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_C6;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_CO5;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_CO6;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_C_CY;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_C_XOR;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_D;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_D1;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_D2;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_D3;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_D4;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_D5;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_D6;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_DO5;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_DO6;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_D_CY;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X50Y120_D_XOR;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_A;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_A1;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_A2;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_A3;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_A4;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_A5;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_A6;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_AO5;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_AO6;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_A_CY;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_A_XOR;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_B;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_B1;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_B2;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_B3;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_B4;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_B5;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_B6;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_BO5;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_BO6;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_B_CY;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_B_XOR;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_C;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_C1;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_C2;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_C3;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_C4;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_C5;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_C6;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_CO5;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_CO6;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_C_CY;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_C_XOR;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_D;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_D1;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_D2;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_D3;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_D4;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_D5;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_D6;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_DO5;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_DO6;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_D_CY;
  wire [0:0] CLBLL_L_X34Y120_SLICE_X51Y120_D_XOR;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_A;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_A1;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_A2;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_A3;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_A4;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_A5;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_A6;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_AO5;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_AO6;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_A_CY;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_A_XOR;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_B;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_B1;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_B2;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_B3;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_B4;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_B5;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_B6;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_BO5;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_BO6;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_B_CY;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_B_XOR;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_C;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_C1;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_C2;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_C3;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_C4;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_C5;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_C6;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_CO5;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_CO6;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_C_CY;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_C_XOR;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_D;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_D1;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_D2;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_D3;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_D4;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_D5;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_D6;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_DO5;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_DO6;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_D_CY;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X50Y121_D_XOR;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_A;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_A1;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_A2;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_A3;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_A4;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_A5;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_A6;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_AO5;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_AO6;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_A_CY;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_A_XOR;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_B;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_B1;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_B2;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_B3;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_B4;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_B5;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_B6;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_BO5;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_BO6;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_B_CY;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_B_XOR;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_C;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_C1;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_C2;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_C3;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_C4;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_C5;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_C6;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_CO5;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_CO6;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_C_CY;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_C_XOR;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_D;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_D1;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_D2;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_D3;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_D4;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_D5;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_D6;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_DO5;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_DO6;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_D_CY;
  wire [0:0] CLBLL_L_X34Y121_SLICE_X51Y121_D_XOR;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_A;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_A1;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_A2;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_A3;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_A4;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_A5;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_A6;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_AO5;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_AO6;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_A_CY;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_A_XOR;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_B;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_B1;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_B2;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_B3;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_B4;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_B5;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_B6;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_BO5;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_BO6;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_B_CY;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_B_XOR;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_C;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_C1;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_C2;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_C3;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_C4;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_C5;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_C6;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_CO5;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_CO6;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_C_CY;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_C_XOR;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_D;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_D1;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_D2;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_D3;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_D4;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_D5;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_D6;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_DO5;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_DO6;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_D_CY;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X50Y122_D_XOR;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_A;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_A1;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_A2;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_A3;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_A4;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_A5;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_A6;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_AO5;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_AO6;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_A_CY;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_A_XOR;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_B;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_B1;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_B2;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_B3;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_B4;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_B5;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_B6;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_BO5;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_BO6;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_B_CY;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_B_XOR;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_C;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_C1;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_C2;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_C3;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_C4;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_C5;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_C6;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_CO5;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_CO6;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_C_CY;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_C_XOR;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_D;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_D1;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_D2;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_D3;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_D4;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_D5;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_D6;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_DO5;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_DO6;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_D_CY;
  wire [0:0] CLBLL_L_X34Y122_SLICE_X51Y122_D_XOR;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_A;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_A1;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_A2;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_A3;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_A4;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_A5;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_A6;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_AMUX;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_AO5;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_AO6;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_A_CY;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_A_XOR;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_B;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_B1;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_B2;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_B3;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_B4;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_B5;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_B6;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_BMUX;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_BO5;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_BO6;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_B_CY;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_B_XOR;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_C;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_C1;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_C2;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_C3;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_C4;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_C5;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_C6;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_CO5;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_CO6;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_C_CY;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_C_XOR;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_D;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_D1;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_D2;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_D3;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_D4;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_D5;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_D6;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_DO5;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_DO6;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_D_CY;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X50Y123_D_XOR;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_A;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_A1;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_A2;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_A3;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_A4;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_A5;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_A6;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_AO5;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_AO6;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_A_CY;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_A_XOR;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_B;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_B1;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_B2;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_B3;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_B4;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_B5;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_B6;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_BO5;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_BO6;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_B_CY;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_B_XOR;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_C;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_C1;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_C2;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_C3;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_C4;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_C5;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_C6;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_CO5;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_CO6;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_COUT;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_C_CY;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_C_XOR;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_D;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_D1;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_D2;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_D3;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_D4;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_D5;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_D6;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_DO5;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_DO6;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_D_CY;
  wire [0:0] CLBLL_L_X34Y123_SLICE_X51Y123_D_XOR;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_A;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_A1;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_A2;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_A3;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_A4;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_A5;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_A6;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_AO5;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_AO6;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_A_CY;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_A_XOR;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_B;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_B1;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_B2;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_B3;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_B4;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_B5;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_B6;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_BO5;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_BO6;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_B_CY;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_B_XOR;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_C;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_C1;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_C2;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_C3;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_C4;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_C5;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_C6;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_CMUX;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_CO5;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_CO6;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_C_CY;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_C_XOR;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_D;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_D1;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_D2;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_D3;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_D4;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_D5;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_D6;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_DO5;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_DO6;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_D_CY;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X50Y124_D_XOR;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_A;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_A1;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_A2;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_A3;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_A4;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_A5;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_A6;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_AO5;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_AO6;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_A_CY;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_A_XOR;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_B;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_B1;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_B2;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_B3;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_B4;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_B5;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_B6;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_BO5;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_BO6;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_B_CY;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_B_XOR;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_C;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_C1;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_C2;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_C3;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_C4;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_C5;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_C6;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_CIN;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_CO5;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_CO6;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_COUT;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_C_CY;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_C_XOR;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_D;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_D1;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_D2;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_D3;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_D4;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_D5;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_D6;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_DO5;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_DO6;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_D_CY;
  wire [0:0] CLBLL_L_X34Y124_SLICE_X51Y124_D_XOR;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_A;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_A1;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_A2;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_A3;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_A4;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_A5;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_A6;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_AO5;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_AO6;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_A_CY;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_A_XOR;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_B;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_B1;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_B2;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_B3;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_B4;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_B5;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_B6;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_BO5;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_BO6;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_B_CY;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_B_XOR;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_C;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_C1;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_C2;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_C3;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_C4;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_C5;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_C6;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_CO5;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_CO6;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_C_CY;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_C_XOR;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_D;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_D1;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_D2;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_D3;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_D4;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_D5;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_D6;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_DO5;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_DO6;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_D_CY;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X50Y125_D_XOR;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_A;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_A1;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_A2;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_A3;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_A4;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_A5;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_A6;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_AO5;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_AO6;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_A_CY;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_A_XOR;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_B;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_B1;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_B2;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_B3;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_B4;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_B5;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_B6;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_BO5;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_BO6;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_B_CY;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_B_XOR;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_C;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_C1;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_C2;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_C3;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_C4;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_C5;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_C6;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_CIN;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_CO5;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_CO6;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_COUT;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_C_CY;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_C_XOR;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_D;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_D1;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_D2;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_D3;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_D4;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_D5;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_D6;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_DO5;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_DO6;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_D_CY;
  wire [0:0] CLBLL_L_X34Y125_SLICE_X51Y125_D_XOR;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_A;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_A1;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_A2;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_A3;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_A4;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_A5;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_A6;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_AO5;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_AO6;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_A_CY;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_A_XOR;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_B;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_B1;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_B2;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_B3;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_B4;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_B5;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_B6;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_BO5;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_BO6;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_B_CY;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_B_XOR;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_C;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_C1;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_C2;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_C3;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_C4;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_C5;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_C6;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_CO5;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_CO6;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_C_CY;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_C_XOR;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_D;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_D1;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_D2;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_D3;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_D4;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_D5;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_D6;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_DO5;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_DO6;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_D_CY;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X50Y126_D_XOR;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_A;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_A1;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_A2;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_A3;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_A4;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_A5;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_A6;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_AO5;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_AO6;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_A_CY;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_A_XOR;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_B;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_B1;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_B2;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_B3;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_B4;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_B5;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_B6;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_BO5;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_BO6;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_B_CY;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_B_XOR;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_C;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_C1;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_C2;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_C3;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_C4;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_C5;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_C6;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_CIN;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_CO5;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_CO6;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_COUT;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_C_CY;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_C_XOR;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_D;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_D1;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_D2;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_D3;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_D4;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_D5;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_D6;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_DMUX;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_DO5;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_DO6;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_D_CY;
  wire [0:0] CLBLL_L_X34Y126_SLICE_X51Y126_D_XOR;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_A;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_A1;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_A2;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_A3;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_A4;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_A5;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_A6;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_AO5;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_AO6;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_A_CY;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_A_XOR;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_B;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_B1;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_B2;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_B3;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_B4;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_B5;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_B6;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_BO5;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_BO6;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_B_CY;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_B_XOR;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_C;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_C1;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_C2;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_C3;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_C4;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_C5;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_C6;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_CO5;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_CO6;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_C_CY;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_C_XOR;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_D;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_D1;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_D2;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_D3;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_D4;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_D5;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_D6;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_DO5;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_D_CY;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X50Y127_D_XOR;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_A;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_A1;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_A2;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_A3;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_A4;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_A5;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_A6;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_AO5;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_AO6;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_A_CY;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_A_XOR;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_B;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_B1;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_B2;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_B3;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_B4;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_B5;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_B6;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_BO5;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_BO6;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_B_CY;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_B_XOR;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_C;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_C1;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_C2;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_C3;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_C4;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_C5;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_C6;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_CO5;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_CO6;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_C_CY;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_C_XOR;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_D;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_D1;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_D2;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_D3;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_D4;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_D5;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_D6;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_DO5;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_DO6;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_D_CY;
  wire [0:0] CLBLL_L_X34Y127_SLICE_X51Y127_D_XOR;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_A;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_A1;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_A2;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_A3;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_A4;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_A5;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_A6;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_AO5;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_AO6;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_A_CY;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_A_XOR;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_B;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_B1;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_B2;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_B3;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_B4;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_B5;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_B6;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_BO5;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_BO6;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_B_CY;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_B_XOR;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_C;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_C1;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_C2;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_C3;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_C4;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_C5;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_C6;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_CO5;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_CO6;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_C_CY;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_C_XOR;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_D;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_D1;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_D2;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_D3;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_D4;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_D5;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_D6;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_DO5;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_DO6;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_D_CY;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X50Y128_D_XOR;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_A;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_A1;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_A2;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_A3;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_A4;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_A5;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_A6;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_AO5;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_AO6;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_A_CY;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_A_XOR;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_B;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_B1;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_B2;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_B3;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_B4;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_B5;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_B6;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_BO5;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_BO6;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_B_CY;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_B_XOR;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_C;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_C1;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_C2;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_C3;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_C4;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_C5;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_C6;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_CO5;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_CO6;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_C_CY;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_C_XOR;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_D;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_D1;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_D2;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_D3;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_D4;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_D5;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_D6;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_DO5;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_DO6;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_D_CY;
  wire [0:0] CLBLL_L_X34Y128_SLICE_X51Y128_D_XOR;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_A;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_A1;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_A2;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_A3;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_A4;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_A5;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_A6;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_AO5;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_A_CY;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_A_XOR;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_B;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_B1;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_B2;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_B3;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_B4;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_B5;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_B6;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_BO5;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_BO6;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_B_CY;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_B_XOR;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_C;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_C1;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_C2;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_C3;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_C4;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_C5;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_C6;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_CO5;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_CO6;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_C_CY;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_C_XOR;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_D;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_D1;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_D2;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_D3;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_D4;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_D5;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_D6;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_DO5;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_DO6;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_D_CY;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X50Y129_D_XOR;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_A;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_A1;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_A2;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_A3;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_A4;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_A5;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_A6;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_AO5;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_AO6;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_A_CY;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_A_XOR;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_B;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_B1;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_B2;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_B3;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_B4;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_B5;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_B6;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_BO5;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_BO6;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_B_CY;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_B_XOR;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_C;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_C1;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_C2;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_C3;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_C4;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_C5;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_C6;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_CO5;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_CO6;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_C_CY;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_C_XOR;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_D;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_D1;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_D2;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_D3;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_D4;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_D5;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_D6;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_DO5;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_DO6;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_D_CY;
  wire [0:0] CLBLL_L_X34Y129_SLICE_X51Y129_D_XOR;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_A;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_A1;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_A2;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_A3;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_A4;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_A5;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_A6;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_AMUX;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_AO5;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_AO6;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_A_CY;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_A_XOR;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_B;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_B1;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_B2;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_B3;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_B4;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_B5;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_B6;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_BO5;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_BO6;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_B_CY;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_B_XOR;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_C;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_C1;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_C2;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_C3;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_C4;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_C5;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_C6;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_CO5;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_CO6;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_C_CY;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_C_XOR;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_D;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_D1;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_D2;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_D3;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_D4;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_D5;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_D6;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_DO5;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_DO6;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_D_CY;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X54Y115_D_XOR;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_A;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_A1;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_A2;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_A3;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_A4;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_A5;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_A6;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_AO5;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_AO6;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_A_CY;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_A_XOR;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_B;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_B1;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_B2;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_B3;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_B4;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_B5;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_B6;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_BO5;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_BO6;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_B_CY;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_B_XOR;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_C;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_C1;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_C2;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_C3;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_C4;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_C5;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_C6;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_CO5;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_CO6;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_C_CY;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_C_XOR;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_D;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_D1;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_D2;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_D3;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_D4;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_D5;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_D6;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_DO5;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_DO6;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_D_CY;
  wire [0:0] CLBLL_L_X36Y115_SLICE_X55Y115_D_XOR;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_A;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_A1;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_A2;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_A3;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_A4;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_A5;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_A6;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_AMUX;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_AO5;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_AO6;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_A_CY;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_A_XOR;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_B;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_B1;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_B2;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_B3;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_B4;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_B5;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_B6;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_BMUX;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_BO5;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_BO6;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_B_CY;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_B_XOR;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_C;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_C1;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_C2;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_C3;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_C4;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_C5;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_C6;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_CMUX;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_CO5;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_CO6;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_C_CY;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_C_XOR;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_D;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_D1;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_D2;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_D3;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_D4;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_D5;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_D6;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_DO5;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_DO6;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_D_CY;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X54Y116_D_XOR;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_A;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_A1;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_A2;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_A3;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_A4;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_A5;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_A6;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_AMUX;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_AO5;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_AO6;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_A_CY;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_A_XOR;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_B;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_B1;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_B2;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_B3;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_B4;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_B5;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_B6;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_BO5;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_BO6;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_B_CY;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_B_XOR;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_C;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_C1;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_C2;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_C3;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_C4;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_C5;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_C6;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_CO5;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_CO6;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_C_CY;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_C_XOR;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_D;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_D1;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_D2;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_D3;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_D4;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_D5;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_D6;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_DO5;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_DO6;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_D_CY;
  wire [0:0] CLBLL_L_X36Y116_SLICE_X55Y116_D_XOR;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_A;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_A1;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_A2;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_A3;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_A4;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_A5;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_A6;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_AO5;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_AO6;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_A_CY;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_A_XOR;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_B;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_B1;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_B2;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_B3;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_B4;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_B5;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_B6;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_BO5;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_BO6;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_B_CY;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_B_XOR;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_C;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_C1;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_C2;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_C3;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_C4;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_C5;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_C6;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_CO5;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_CO6;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_C_CY;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_C_XOR;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_D;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_D1;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_D2;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_D3;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_D4;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_D5;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_D6;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_DO5;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_DO6;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_D_CY;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X54Y117_D_XOR;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_A;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_A1;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_A2;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_A3;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_A4;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_A5;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_A6;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_AMUX;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_AO5;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_AO6;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_A_CY;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_A_XOR;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_B;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_B1;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_B2;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_B3;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_B4;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_B5;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_B6;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_BMUX;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_BO5;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_BO6;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_B_CY;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_B_XOR;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_C;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_C1;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_C2;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_C3;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_C4;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_C5;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_C6;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_CO5;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_CO6;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_C_CY;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_C_XOR;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_D;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_D1;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_D2;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_D3;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_D4;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_D5;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_D6;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_DO5;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_DO6;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_D_CY;
  wire [0:0] CLBLL_L_X36Y117_SLICE_X55Y117_D_XOR;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_A;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_A1;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_A2;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_A3;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_A4;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_A5;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_A6;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_AO5;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_AO6;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_A_CY;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_A_XOR;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_B;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_B1;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_B2;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_B3;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_B4;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_B5;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_B6;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_BO5;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_BO6;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_B_CY;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_B_XOR;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_C;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_C1;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_C2;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_C3;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_C4;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_C5;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_C6;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_CO5;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_CO6;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_C_CY;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_C_XOR;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_D;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_D1;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_D2;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_D3;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_D4;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_D5;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_D6;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_DO5;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_DO6;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_D_CY;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X54Y118_D_XOR;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_A;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_A1;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_A2;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_A3;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_A4;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_A5;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_A6;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_AMUX;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_AO5;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_AO6;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_A_CY;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_A_XOR;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_B;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_B1;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_B2;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_B3;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_B4;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_B5;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_B6;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_BO5;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_BO6;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_B_CY;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_B_XOR;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_C;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_C1;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_C2;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_C3;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_C4;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_C5;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_C6;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_CMUX;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_CO5;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_CO6;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_C_CY;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_C_XOR;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_D;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_D1;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_D2;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_D3;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_D4;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_D5;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_D6;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_DO5;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_DO6;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_D_CY;
  wire [0:0] CLBLL_L_X36Y118_SLICE_X55Y118_D_XOR;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_A;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_A1;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_A2;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_A3;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_A4;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_A5;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_A6;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_AO5;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_AO6;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_A_CY;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_A_XOR;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_B;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_B1;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_B2;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_B3;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_B4;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_B5;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_B6;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_BO5;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_BO6;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_B_CY;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_B_XOR;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_C;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_C1;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_C2;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_C3;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_C4;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_C5;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_C6;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_CO5;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_CO6;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_C_CY;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_C_XOR;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_D;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_D1;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_D2;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_D3;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_D4;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_D5;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_D6;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_DO5;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_DO6;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_D_CY;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X54Y119_D_XOR;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_A;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_A1;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_A2;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_A3;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_A4;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_A5;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_A6;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_AO5;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_AO6;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_A_CY;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_A_XOR;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_B;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_B1;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_B2;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_B3;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_B4;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_B5;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_B6;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_BO5;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_BO6;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_B_CY;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_B_XOR;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_C;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_C1;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_C2;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_C3;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_C4;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_C5;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_C6;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_CO5;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_CO6;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_C_CY;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_C_XOR;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_D;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_D1;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_D2;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_D3;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_D4;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_D5;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_D6;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_DO5;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_DO6;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_D_CY;
  wire [0:0] CLBLL_L_X36Y119_SLICE_X55Y119_D_XOR;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_A;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_A1;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_A2;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_A3;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_A4;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_A5;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_A6;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_AO5;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_AO6;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_A_CY;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_A_XOR;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_B;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_B1;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_B2;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_B3;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_B4;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_B5;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_B6;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_BO5;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_BO6;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_B_CY;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_B_XOR;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_C;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_C1;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_C2;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_C3;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_C4;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_C5;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_C6;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_CO5;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_CO6;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_C_CY;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_C_XOR;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_D;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_D1;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_D2;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_D3;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_D4;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_D5;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_D6;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_DO5;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_DO6;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_D_CY;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X54Y120_D_XOR;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_A;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_A1;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_A2;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_A3;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_A4;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_A5;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_A6;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_AO5;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_AO6;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_A_CY;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_A_XOR;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_B;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_B1;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_B2;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_B3;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_B4;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_B5;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_B6;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_BO5;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_BO6;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_B_CY;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_B_XOR;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_C;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_C1;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_C2;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_C3;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_C4;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_C5;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_C6;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_CO5;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_CO6;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_C_CY;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_C_XOR;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_D;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_D1;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_D2;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_D3;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_D4;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_D5;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_D6;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_DO5;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_DO6;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_D_CY;
  wire [0:0] CLBLL_L_X36Y120_SLICE_X55Y120_D_XOR;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_A;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_A1;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_A2;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_A3;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_A4;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_A5;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_A6;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_AMUX;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_AO5;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_AO6;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_A_CY;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_A_XOR;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_B;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_B1;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_B2;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_B3;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_B4;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_B5;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_B6;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_BO5;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_BO6;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_B_CY;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_B_XOR;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_C;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_C1;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_C2;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_C3;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_C4;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_C5;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_C6;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_CO5;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_CO6;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_C_CY;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_C_XOR;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_D;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_D1;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_D2;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_D3;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_D4;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_D5;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_D6;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_DO5;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_DO6;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_D_CY;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X54Y121_D_XOR;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_A;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_A1;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_A2;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_A3;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_A4;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_A5;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_A6;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_AMUX;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_AO5;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_AO6;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_A_CY;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_A_XOR;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_B;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_B1;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_B2;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_B3;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_B4;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_B5;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_B6;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_BO5;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_BO6;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_B_CY;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_B_XOR;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_C;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_C1;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_C2;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_C3;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_C4;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_C5;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_C6;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_CO5;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_CO6;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_C_CY;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_C_XOR;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_D;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_D1;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_D2;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_D3;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_D4;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_D5;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_D6;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_DO5;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_DO6;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_D_CY;
  wire [0:0] CLBLL_L_X36Y121_SLICE_X55Y121_D_XOR;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_A;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_A1;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_A2;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_A3;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_A4;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_A5;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_A6;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_AMUX;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_AO5;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_AO6;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_A_CY;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_A_XOR;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_B;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_B1;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_B2;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_B3;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_B4;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_B5;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_B6;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_BO5;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_BO6;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_B_CY;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_B_XOR;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_C;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_C1;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_C2;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_C3;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_C4;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_C5;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_C6;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_CO5;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_CO6;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_C_CY;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_C_XOR;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_D;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_D1;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_D2;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_D3;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_D4;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_D5;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_D6;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_DO5;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_DO6;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_D_CY;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X54Y122_D_XOR;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_A;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_A1;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_A2;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_A3;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_A4;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_A5;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_A6;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_AMUX;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_AO5;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_AO6;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_A_CY;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_A_XOR;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_B;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_B1;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_B2;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_B3;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_B4;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_B5;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_B6;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_BO5;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_BO6;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_B_CY;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_B_XOR;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_C;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_C1;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_C2;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_C3;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_C4;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_C5;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_C6;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_CO5;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_CO6;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_C_CY;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_C_XOR;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_D;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_D1;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_D2;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_D3;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_D4;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_D5;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_D6;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_DO5;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_DO6;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_D_CY;
  wire [0:0] CLBLL_L_X36Y122_SLICE_X55Y122_D_XOR;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_A;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_A1;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_A2;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_A3;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_A4;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_A5;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_A6;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_AMUX;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_AO5;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_AO6;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_A_CY;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_A_XOR;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_B;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_B1;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_B2;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_B3;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_B4;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_B5;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_B6;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_BO5;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_BO6;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_B_CY;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_B_XOR;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_C;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_C1;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_C2;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_C3;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_C4;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_C5;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_C6;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_CO5;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_CO6;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_C_CY;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_C_XOR;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_D;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_D1;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_D2;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_D3;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_D4;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_D5;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_D6;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_DO5;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_DO6;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_D_CY;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X54Y123_D_XOR;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_A;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_A1;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_A2;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_A3;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_A4;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_A5;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_A6;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_AO5;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_AO6;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_A_CY;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_A_XOR;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_B;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_B1;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_B2;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_B3;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_B4;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_B5;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_B6;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_BO5;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_BO6;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_B_CY;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_B_XOR;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_C;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_C1;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_C2;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_C3;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_C4;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_C5;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_C6;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_CO5;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_CO6;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_C_CY;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_C_XOR;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_D;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_D1;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_D2;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_D3;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_D4;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_D5;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_D6;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_DO5;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_DO6;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_D_CY;
  wire [0:0] CLBLL_L_X36Y123_SLICE_X55Y123_D_XOR;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_A;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_A1;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_A2;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_A3;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_A4;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_A5;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_A6;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_AO5;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_AO6;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_A_CY;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_A_XOR;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_B;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_B1;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_B2;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_B3;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_B4;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_B5;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_B6;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_BO5;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_BO6;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_B_CY;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_B_XOR;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_C;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_C1;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_C2;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_C3;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_C4;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_C5;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_C6;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_CO5;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_CO6;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_C_CY;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_C_XOR;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_D;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_D1;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_D2;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_D3;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_D4;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_D5;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_D6;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_DO5;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_DO6;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_D_CY;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_D_XOR;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_A;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_A1;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_A2;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_A3;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_A4;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_A5;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_A6;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_AO5;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_AO6;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_A_CY;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_A_XOR;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_B;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_B1;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_B2;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_B3;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_B4;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_B5;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_B6;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_BMUX;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_BO5;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_BO6;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_B_CY;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_B_XOR;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_C;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_C1;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_C2;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_C3;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_C4;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_C5;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_C6;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_CMUX;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_CO5;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_CO6;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_C_CY;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_C_XOR;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_D;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_D1;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_D2;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_D3;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_D4;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_D5;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_D6;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_DO5;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_DO6;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_D_CY;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_D_XOR;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_A;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_A1;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_A2;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_A3;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_A4;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_A5;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_A6;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_AO5;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_AO6;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_A_CY;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_A_XOR;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_B;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_B1;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_B2;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_B3;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_B4;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_B5;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_B6;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_BO5;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_BO6;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_B_CY;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_B_XOR;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_C;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_C1;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_C2;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_C3;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_C4;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_C5;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_C6;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_CO5;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_CO6;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_C_CY;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_C_XOR;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_D;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_D1;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_D2;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_D3;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_D4;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_D5;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_D6;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_DO5;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_DO6;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_D_CY;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X54Y125_D_XOR;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_A;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_A1;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_A2;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_A3;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_A4;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_A5;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_A6;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_AMUX;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_AO5;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_AO6;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_A_CY;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_A_XOR;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_B;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_B1;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_B2;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_B3;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_B4;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_B5;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_B6;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_BMUX;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_BO5;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_BO6;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_B_CY;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_B_XOR;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_C;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_C1;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_C2;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_C3;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_C4;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_C5;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_C6;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_CMUX;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_CO5;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_CO6;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_C_CY;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_C_XOR;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_D;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_D1;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_D2;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_D3;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_D4;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_D5;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_D6;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_DO5;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_DO6;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_D_CY;
  wire [0:0] CLBLL_L_X36Y125_SLICE_X55Y125_D_XOR;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_A;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_A1;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_A2;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_A3;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_A4;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_A5;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_A6;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_AO5;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_AO6;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_A_CY;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_A_XOR;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_B;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_B1;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_B2;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_B3;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_B4;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_B5;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_B6;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_BO5;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_BO6;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_B_CY;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_B_XOR;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_C;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_C1;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_C2;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_C3;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_C4;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_C5;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_C6;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_CMUX;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_CO5;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_CO6;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_C_CY;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_C_XOR;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_D;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_D1;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_D2;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_D3;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_D4;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_D5;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_D6;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_DO5;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_DO6;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_D_CY;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X54Y126_D_XOR;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_A;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_A1;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_A2;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_A3;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_A4;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_A5;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_A6;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_AO5;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_AO6;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_A_CY;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_A_XOR;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_B;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_B1;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_B2;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_B3;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_B4;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_B5;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_B6;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_BO5;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_BO6;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_B_CY;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_B_XOR;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_C;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_C1;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_C2;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_C3;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_C4;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_C5;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_C6;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_CO5;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_CO6;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_C_CY;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_C_XOR;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_D;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_D1;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_D2;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_D3;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_D4;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_D5;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_D6;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_DO5;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_DO6;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_D_CY;
  wire [0:0] CLBLL_L_X36Y126_SLICE_X55Y126_D_XOR;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_A;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_A1;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_A2;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_A3;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_A4;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_A5;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_A6;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_AO5;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_AO6;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_A_CY;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_A_XOR;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_B;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_B1;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_B2;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_B3;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_B4;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_B5;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_B6;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_BO5;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_BO6;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_B_CY;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_B_XOR;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_C;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_C1;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_C2;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_C3;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_C4;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_C5;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_C6;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_CO5;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_CO6;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_C_CY;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_C_XOR;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_D;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_D1;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_D2;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_D3;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_D4;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_D5;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_D6;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_DO5;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_DO6;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_D_CY;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_D_XOR;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_A;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_A1;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_A2;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_A3;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_A4;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_A5;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_A6;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_AO5;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_AO6;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_A_CY;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_A_XOR;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_B;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_B1;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_B2;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_B3;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_B4;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_B5;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_B6;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_BO5;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_BO6;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_B_CY;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_B_XOR;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_C;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_C1;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_C2;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_C3;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_C4;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_C5;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_C6;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_CO5;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_CO6;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_C_CY;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_C_XOR;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_D;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_D1;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_D2;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_D3;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_D4;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_D5;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_D6;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_DO5;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_DO6;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_D_CY;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_D_XOR;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_A;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_A1;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_A2;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_A3;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_A4;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_A5;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_A6;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_AO5;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_AO6;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_A_CY;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_A_XOR;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_B;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_B1;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_B2;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_B3;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_B4;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_B5;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_B6;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_BO5;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_BO6;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_B_CY;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_B_XOR;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_C;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_C1;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_C2;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_C3;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_C4;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_C5;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_C6;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_CO5;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_CO6;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_C_CY;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_C_XOR;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_D;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_D1;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_D2;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_D3;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_D4;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_D5;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_D6;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_DO5;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_DO6;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_D_CY;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X54Y128_D_XOR;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_A;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_A1;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_A2;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_A3;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_A4;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_A5;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_A6;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_AO5;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_AO6;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_A_CY;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_A_XOR;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_B;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_B1;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_B2;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_B3;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_B4;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_B5;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_B6;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_BO5;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_BO6;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_B_CY;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_B_XOR;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_C;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_C1;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_C2;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_C3;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_C4;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_C5;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_C6;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_CO5;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_CO6;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_C_CY;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_C_XOR;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_D;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_D1;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_D2;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_D3;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_D4;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_D5;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_D6;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_DO5;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_DO6;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_D_CY;
  wire [0:0] CLBLL_L_X36Y128_SLICE_X55Y128_D_XOR;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_A;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_A1;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_A2;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_A3;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_A4;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_A5;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_A6;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_AO5;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_AO6;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_A_CY;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_A_XOR;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_B;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_B1;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_B2;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_B3;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_B4;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_B5;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_B6;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_BO5;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_BO6;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_B_CY;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_B_XOR;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_C;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_C1;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_C2;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_C3;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_C4;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_C5;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_C6;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_CO5;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_CO6;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_C_CY;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_C_XOR;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_D;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_D1;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_D2;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_D3;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_D4;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_D5;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_D6;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_DO5;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_DO6;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_D_CY;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X54Y129_D_XOR;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_A;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_A1;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_A2;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_A3;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_A4;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_A5;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_A6;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_AO5;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_AO6;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_A_CY;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_A_XOR;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_B;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_B1;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_B2;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_B3;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_B4;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_B5;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_B6;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_BO5;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_BO6;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_B_CY;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_B_XOR;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_C;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_C1;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_C2;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_C3;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_C4;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_C5;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_C6;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_CO5;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_CO6;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_C_CY;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_C_XOR;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_D;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_D1;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_D2;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_D3;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_D4;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_D5;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_D6;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_DO5;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_DO6;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_D_CY;
  wire [0:0] CLBLL_L_X36Y129_SLICE_X55Y129_D_XOR;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_A;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_A1;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_A2;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_A3;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_A4;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_A5;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_A6;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_AMUX;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_AO5;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_AO6;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_A_CY;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_A_XOR;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_B;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_B1;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_B2;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_B3;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_B4;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_B5;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_B6;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_BO5;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_BO6;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_B_CY;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_B_XOR;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_C;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_C1;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_C2;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_C3;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_C4;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_C5;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_C6;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_CO5;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_CO6;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_C_CY;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_C_XOR;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_D;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_D1;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_D2;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_D3;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_D4;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_D5;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_D6;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_DO5;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_DO6;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_D_CY;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X58Y118_D_XOR;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_A;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_A1;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_A2;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_A3;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_A4;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_A5;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_A6;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_AO5;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_AO6;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_A_CY;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_A_XOR;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_B;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_B1;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_B2;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_B3;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_B4;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_B5;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_B6;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_BO5;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_BO6;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_B_CY;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_B_XOR;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_C;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_C1;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_C2;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_C3;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_C4;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_C5;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_C6;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_CO5;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_CO6;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_C_CY;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_C_XOR;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_D;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_D1;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_D2;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_D3;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_D4;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_D5;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_D6;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_DO5;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_DO6;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_D_CY;
  wire [0:0] CLBLL_L_X38Y118_SLICE_X59Y118_D_XOR;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_A;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_A1;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_A2;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_A3;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_A4;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_A5;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_A6;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_AO5;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_AO6;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_A_CY;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_A_XOR;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_B;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_B1;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_B2;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_B3;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_B4;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_B5;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_B6;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_BO5;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_BO6;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_B_CY;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_B_XOR;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_C;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_C1;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_C2;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_C3;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_C4;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_C5;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_C6;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_CO5;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_CO6;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_C_CY;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_C_XOR;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_D;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_D1;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_D2;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_D3;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_D4;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_D5;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_D6;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_DO5;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_DO6;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_D_CY;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X58Y119_D_XOR;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_A;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_A1;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_A2;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_A3;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_A4;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_A5;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_A6;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_AO5;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_AO6;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_A_CY;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_A_XOR;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_B;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_B1;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_B2;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_B3;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_B4;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_B5;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_B6;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_BO5;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_BO6;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_B_CY;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_B_XOR;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_C;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_C1;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_C2;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_C3;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_C4;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_C5;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_C6;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_CO5;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_CO6;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_C_CY;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_C_XOR;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_D;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_D1;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_D2;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_D3;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_D4;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_D5;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_D6;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_DO5;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_DO6;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_D_CY;
  wire [0:0] CLBLL_L_X38Y119_SLICE_X59Y119_D_XOR;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_A;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_A1;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_A2;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_A3;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_A4;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_A5;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_A6;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_AO5;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_AO6;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_A_CY;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_A_XOR;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_B;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_B1;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_B2;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_B3;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_B4;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_B5;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_B6;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_BO5;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_BO6;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_B_CY;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_B_XOR;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_C;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_C1;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_C2;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_C3;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_C4;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_C5;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_C6;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_CO5;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_CO6;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_C_CY;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_C_XOR;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_D;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_D1;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_D2;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_D3;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_D4;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_D5;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_D6;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_DO5;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_DO6;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_D_CY;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X58Y121_D_XOR;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_A;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_A1;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_A2;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_A3;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_A4;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_A5;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_A6;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_AO5;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_AO6;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_A_CY;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_A_XOR;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_B;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_B1;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_B2;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_B3;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_B4;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_B5;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_B6;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_BO5;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_BO6;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_B_CY;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_B_XOR;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_C;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_C1;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_C2;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_C3;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_C4;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_C5;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_C6;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_CO5;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_CO6;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_C_CY;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_C_XOR;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_D;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_D1;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_D2;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_D3;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_D4;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_D5;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_D6;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_DO5;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_DO6;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_D_CY;
  wire [0:0] CLBLL_L_X38Y121_SLICE_X59Y121_D_XOR;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_A;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_A1;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_A2;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_A3;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_A4;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_A5;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_A6;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_AO5;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_AO6;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_A_CY;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_A_XOR;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_B;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_B1;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_B2;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_B3;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_B4;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_B5;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_B6;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_BO5;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_BO6;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_B_CY;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_B_XOR;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_C;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_C1;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_C2;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_C3;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_C4;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_C5;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_C6;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_CO5;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_CO6;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_C_CY;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_C_XOR;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_D;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_D1;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_D2;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_D3;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_D4;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_D5;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_D6;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_DO5;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_DO6;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_D_CY;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X58Y123_D_XOR;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_A;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_A1;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_A2;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_A3;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_A4;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_A5;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_A6;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_AO5;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_AO6;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_A_CY;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_A_XOR;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_B;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_B1;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_B2;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_B3;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_B4;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_B5;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_B6;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_BO5;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_BO6;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_B_CY;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_B_XOR;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_C;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_C1;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_C2;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_C3;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_C4;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_C5;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_C6;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_CO5;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_CO6;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_C_CY;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_C_XOR;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_D;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_D1;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_D2;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_D3;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_D4;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_D5;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_D6;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_DO5;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_DO6;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_D_CY;
  wire [0:0] CLBLL_L_X38Y123_SLICE_X59Y123_D_XOR;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_A;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_A1;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_A2;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_A3;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_A4;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_A5;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_A6;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_AMUX;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_AO5;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_AO6;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_A_CY;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_A_XOR;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_B;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_B1;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_B2;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_B3;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_B4;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_B5;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_B6;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_BO5;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_BO6;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_B_CY;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_B_XOR;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_C;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_C1;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_C2;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_C3;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_C4;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_C5;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_C6;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_CO5;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_CO6;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_C_CY;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_C_XOR;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_D;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_D1;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_D2;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_D3;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_D4;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_D5;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_D6;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_DO5;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_DO6;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_D_CY;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X58Y124_D_XOR;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_A;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_A1;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_A2;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_A3;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_A4;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_A5;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_A6;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_AO5;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_AO6;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_A_CY;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_A_XOR;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_B;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_B1;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_B2;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_B3;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_B4;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_B5;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_B6;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_BO5;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_BO6;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_B_CY;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_B_XOR;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_C;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_C1;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_C2;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_C3;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_C4;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_C5;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_C6;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_CO5;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_CO6;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_C_CY;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_C_XOR;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_D;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_D1;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_D2;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_D3;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_D4;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_D5;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_D6;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_DO5;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_DO6;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_D_CY;
  wire [0:0] CLBLL_L_X38Y124_SLICE_X59Y124_D_XOR;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_A;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_A1;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_A2;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_A3;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_A4;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_A5;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_A6;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_AO5;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_AO6;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_A_CY;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_A_XOR;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_B;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_B1;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_B2;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_B3;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_B4;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_B5;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_B6;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_BO5;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_BO6;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_B_CY;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_B_XOR;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_C;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_C1;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_C2;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_C3;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_C4;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_C5;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_C6;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_CO5;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_CO6;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_C_CY;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_C_XOR;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_D;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_D1;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_D2;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_D3;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_D4;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_D5;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_D6;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_DO5;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_DO6;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_D_CY;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X58Y126_D_XOR;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_A;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_A1;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_A2;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_A3;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_A4;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_A5;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_A6;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_AO5;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_AO6;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_A_CY;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_A_XOR;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_B;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_B1;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_B2;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_B3;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_B4;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_B5;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_B6;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_BO5;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_BO6;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_B_CY;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_B_XOR;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_C;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_C1;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_C2;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_C3;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_C4;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_C5;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_C6;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_CO5;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_CO6;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_C_CY;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_C_XOR;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_D;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_D1;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_D2;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_D3;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_D4;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_D5;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_D6;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_DO5;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_DO6;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_D_CY;
  wire [0:0] CLBLL_L_X38Y126_SLICE_X59Y126_D_XOR;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_A;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_A1;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_A2;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_A3;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_A4;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_A5;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_A6;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_AO5;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_AO6;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_A_CY;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_A_XOR;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_B;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_B1;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_B2;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_B3;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_B4;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_B5;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_B6;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_BO5;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_BO6;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_B_CY;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_B_XOR;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_C;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_C1;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_C2;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_C3;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_C4;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_C5;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_C6;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_CO5;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_CO6;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_C_CY;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_C_XOR;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_D;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_D1;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_D2;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_D3;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_D4;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_D5;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_D6;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_DO5;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_DO6;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_D_CY;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X46Y116_D_XOR;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_A;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_A1;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_A2;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_A3;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_A4;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_A5;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_A6;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_AO5;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_AO6;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_A_CY;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_A_XOR;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_B;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_B1;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_B2;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_B3;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_B4;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_B5;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_B6;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_BO5;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_BO6;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_B_CY;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_B_XOR;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_C;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_C1;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_C2;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_C3;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_C4;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_C5;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_C6;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_CO5;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_CO6;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_C_CY;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_C_XOR;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_D;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_D1;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_D2;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_D3;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_D4;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_D5;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_D6;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_DO5;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_DO6;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_D_CY;
  wire [0:0] CLBLM_L_X32Y116_SLICE_X47Y116_D_XOR;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_A;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_A1;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_A2;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_A3;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_A4;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_A5;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_A6;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_AO5;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_AO6;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_A_CY;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_A_XOR;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_B;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_B1;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_B2;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_B3;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_B4;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_B5;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_B6;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_BO5;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_BO6;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_B_CY;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_B_XOR;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_C;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_C1;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_C2;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_C3;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_C4;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_C5;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_C6;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_CO5;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_CO6;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_C_CY;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_C_XOR;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_D;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_D1;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_D2;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_D3;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_D4;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_D5;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_D6;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_DO5;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_DO6;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_D_CY;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X46Y117_D_XOR;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_A;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_A1;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_A2;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_A3;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_A4;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_A5;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_A6;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_AO5;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_AO6;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_A_CY;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_A_XOR;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_B;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_B1;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_B2;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_B3;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_B4;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_B5;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_B6;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_BO5;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_BO6;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_B_CY;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_B_XOR;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_C;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_C1;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_C2;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_C3;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_C4;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_C5;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_C6;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_CO5;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_CO6;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_C_CY;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_C_XOR;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_D;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_D1;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_D2;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_D3;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_D4;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_D5;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_D6;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_DO5;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_DO6;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_D_CY;
  wire [0:0] CLBLM_L_X32Y117_SLICE_X47Y117_D_XOR;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_A;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_A1;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_A2;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_A3;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_A4;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_A5;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_A6;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_AO5;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_AO6;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_A_CY;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_A_XOR;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_B;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_B1;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_B2;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_B3;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_B4;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_B5;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_B6;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_BO5;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_BO6;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_B_CY;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_B_XOR;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_C;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_C1;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_C2;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_C3;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_C4;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_C5;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_C6;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_CO5;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_CO6;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_C_CY;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_C_XOR;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_D;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_D1;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_D2;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_D3;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_D4;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_D5;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_D6;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_DO5;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_DO6;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_D_CY;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X46Y123_D_XOR;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_A;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_A1;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_A2;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_A3;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_A4;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_A5;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_A6;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_AMUX;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_AO5;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_AO6;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_A_CY;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_A_XOR;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_B;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_B1;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_B2;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_B3;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_B4;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_B5;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_B6;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_BO5;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_BO6;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_B_CY;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_B_XOR;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_C;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_C1;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_C2;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_C3;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_C4;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_C5;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_C6;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_CO5;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_CO6;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_C_CY;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_C_XOR;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_D;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_D1;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_D2;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_D3;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_D4;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_D5;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_D6;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_DO5;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_DO6;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_D_CY;
  wire [0:0] CLBLM_L_X32Y123_SLICE_X47Y123_D_XOR;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_A;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_A1;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_A2;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_A3;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_A4;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_A5;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_A6;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_AO5;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_AO6;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_A_CY;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_A_XOR;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_B;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_B1;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_B2;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_B3;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_B4;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_B5;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_B6;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_BO5;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_BO6;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_B_CY;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_B_XOR;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_C;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_C1;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_C2;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_C3;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_C4;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_C5;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_C6;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_CO5;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_CO6;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_C_CY;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_C_XOR;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_D;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_D1;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_D2;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_D3;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_D4;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_D5;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_D6;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_DO5;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_DO6;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_D_CY;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X48Y115_D_XOR;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_A;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_A1;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_A2;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_A3;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_A4;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_A5;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_A6;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_AMUX;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_AO5;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_AO6;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_A_CY;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_A_XOR;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_B;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_B1;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_B2;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_B3;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_B4;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_B5;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_B6;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_BO5;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_BO6;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_B_CY;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_B_XOR;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_C;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_C1;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_C2;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_C3;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_C4;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_C5;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_C6;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_CO5;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_CO6;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_C_CY;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_C_XOR;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_D;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_D1;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_D2;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_D3;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_D4;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_D5;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_D6;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_DO5;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_DO6;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_D_CY;
  wire [0:0] CLBLM_R_X33Y115_SLICE_X49Y115_D_XOR;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_A;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_A1;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_A2;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_A3;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_A4;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_A5;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_A6;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_AO5;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_AO6;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_A_CY;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_A_XOR;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_B;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_B1;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_B2;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_B3;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_B4;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_B5;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_B6;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_BO5;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_BO6;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_B_CY;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_B_XOR;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_C;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_C1;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_C2;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_C3;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_C4;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_C5;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_C6;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_CO5;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_CO6;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_C_CY;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_C_XOR;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_D;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_D1;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_D2;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_D3;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_D4;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_D5;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_D6;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_DO5;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_DO6;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_D_CY;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X48Y116_D_XOR;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_A;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_A1;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_A2;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_A3;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_A4;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_A5;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_A6;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_AO5;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_AO6;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_A_CY;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_A_XOR;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_B;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_B1;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_B2;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_B3;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_B4;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_B5;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_B6;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_BO5;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_BO6;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_B_CY;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_B_XOR;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_C;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_C1;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_C2;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_C3;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_C4;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_C5;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_C6;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_CO5;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_CO6;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_C_CY;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_C_XOR;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_D;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_D1;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_D2;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_D3;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_D4;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_D5;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_D6;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_DMUX;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_DO5;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_DO6;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_D_CY;
  wire [0:0] CLBLM_R_X33Y116_SLICE_X49Y116_D_XOR;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_A;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_A1;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_A2;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_A3;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_A4;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_A5;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_A6;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_AO5;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_AO6;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_A_CY;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_A_XOR;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_B;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_B1;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_B2;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_B3;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_B4;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_B5;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_B6;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_BO5;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_BO6;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_B_CY;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_B_XOR;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_C;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_C1;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_C2;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_C3;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_C4;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_C5;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_C6;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_CO5;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_CO6;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_C_CY;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_C_XOR;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_D;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_D1;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_D2;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_D3;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_D4;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_D5;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_D6;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_DO5;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_DO6;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_D_CY;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X48Y117_D_XOR;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_A;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_A1;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_A2;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_A3;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_A4;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_A5;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_A6;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_AO5;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_AO6;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_A_CY;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_A_XOR;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_B;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_B1;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_B2;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_B3;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_B4;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_B5;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_B6;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_BO5;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_BO6;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_B_CY;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_B_XOR;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_C;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_C1;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_C2;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_C3;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_C4;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_C5;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_C6;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_CO5;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_CO6;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_C_CY;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_C_XOR;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_D;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_D1;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_D2;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_D3;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_D4;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_D5;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_D6;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_DO5;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_DO6;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_D_CY;
  wire [0:0] CLBLM_R_X33Y117_SLICE_X49Y117_D_XOR;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_A;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_A1;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_A2;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_A3;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_A4;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_A5;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_A6;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_AMUX;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_AO5;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_AO6;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_A_CY;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_A_XOR;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_B;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_B1;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_B2;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_B3;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_B4;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_B5;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_B6;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_BO5;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_BO6;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_B_CY;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_B_XOR;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_C;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_C1;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_C2;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_C3;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_C4;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_C5;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_C6;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_CO5;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_CO6;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_C_CY;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_C_XOR;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_D;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_D1;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_D2;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_D3;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_D4;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_D5;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_D6;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_DO5;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_DO6;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_D_CY;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X48Y118_D_XOR;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_A;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_A1;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_A2;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_A3;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_A4;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_A5;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_A6;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_AO5;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_AO6;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_A_CY;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_A_XOR;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_B;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_B1;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_B2;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_B3;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_B4;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_B5;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_B6;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_BO5;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_BO6;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_B_CY;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_B_XOR;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_C;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_C1;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_C2;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_C3;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_C4;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_C5;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_C6;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_CO5;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_CO6;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_C_CY;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_C_XOR;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_D;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_D1;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_D2;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_D3;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_D4;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_D5;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_D6;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_DO5;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_DO6;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_D_CY;
  wire [0:0] CLBLM_R_X33Y118_SLICE_X49Y118_D_XOR;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_A;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_A1;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_A2;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_A3;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_A4;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_A5;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_A6;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_AO5;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_AO6;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_A_CY;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_A_XOR;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_B;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_B1;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_B2;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_B3;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_B4;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_B5;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_B6;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_BO5;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_BO6;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_B_CY;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_B_XOR;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_C;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_C1;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_C2;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_C3;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_C4;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_C5;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_C6;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_CO5;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_CO6;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_C_CY;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_C_XOR;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_D;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_D1;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_D2;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_D3;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_D4;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_D5;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_D6;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_DO5;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_DO6;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_D_CY;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X48Y119_D_XOR;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_A;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_A1;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_A2;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_A3;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_A4;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_A5;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_A6;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_AMUX;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_AO5;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_AO6;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_A_CY;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_A_XOR;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_B;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_B1;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_B2;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_B3;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_B4;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_B5;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_B6;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_BMUX;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_BO5;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_BO6;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_B_CY;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_B_XOR;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_C;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_C1;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_C2;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_C3;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_C4;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_C5;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_C6;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_CO5;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_CO6;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_C_CY;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_C_XOR;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_D;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_D1;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_D2;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_D3;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_D4;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_D5;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_D6;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_DO5;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_DO6;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_D_CY;
  wire [0:0] CLBLM_R_X33Y119_SLICE_X49Y119_D_XOR;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_A;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_A1;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_A2;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_A3;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_A4;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_A5;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_A6;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_AO5;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_AO6;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_A_CY;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_A_XOR;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_B;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_B1;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_B2;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_B3;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_B4;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_B5;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_B6;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_BO5;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_BO6;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_B_CY;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_B_XOR;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_C;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_C1;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_C2;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_C3;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_C4;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_C5;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_C6;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_CO5;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_CO6;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_C_CY;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_C_XOR;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_D;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_D1;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_D2;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_D3;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_D4;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_D5;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_D6;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_DMUX;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_DO5;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_DO6;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_D_CY;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X48Y121_D_XOR;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_A;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_A1;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_A2;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_A3;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_A4;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_A5;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_A6;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_AO5;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_AO6;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_A_CY;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_A_XOR;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_B;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_B1;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_B2;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_B3;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_B4;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_B5;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_B6;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_BO5;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_BO6;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_B_CY;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_B_XOR;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_C;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_C1;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_C2;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_C3;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_C4;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_C5;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_C6;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_CO5;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_CO6;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_C_CY;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_C_XOR;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_D;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_D1;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_D2;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_D3;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_D4;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_D5;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_D6;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_DO5;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_DO6;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_D_CY;
  wire [0:0] CLBLM_R_X33Y121_SLICE_X49Y121_D_XOR;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_A;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_A1;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_A2;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_A3;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_A4;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_A5;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_A6;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_AMUX;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_AO5;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_AO6;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_A_CY;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_A_XOR;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_B;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_B1;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_B2;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_B3;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_B4;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_B5;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_B6;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_BO5;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_BO6;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_B_CY;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_B_XOR;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_C;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_C1;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_C2;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_C3;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_C4;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_C5;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_C6;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_CO5;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_CO6;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_C_CY;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_C_XOR;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_D;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_D1;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_D2;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_D3;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_D4;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_D5;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_D6;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_DO5;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_DO6;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_D_CY;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X48Y122_D_XOR;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_A;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_A1;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_A2;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_A3;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_A4;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_A5;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_A6;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_AO5;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_AO6;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_A_CY;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_A_XOR;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_B;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_B1;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_B2;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_B3;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_B4;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_B5;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_B6;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_BO5;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_BO6;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_B_CY;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_B_XOR;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_C;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_C1;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_C2;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_C3;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_C4;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_C5;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_C6;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_CO5;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_CO6;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_C_CY;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_C_XOR;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_D;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_D1;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_D2;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_D3;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_D4;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_D5;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_D6;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_DO5;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_DO6;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_D_CY;
  wire [0:0] CLBLM_R_X33Y122_SLICE_X49Y122_D_XOR;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_A;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_A1;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_A2;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_A3;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_A4;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_A5;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_A6;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_AO5;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_AO6;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_A_CY;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_A_XOR;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_B;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_B1;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_B2;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_B3;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_B4;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_B5;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_B6;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_BO5;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_BO6;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_B_CY;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_B_XOR;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_C;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_C1;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_C2;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_C3;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_C4;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_C5;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_C6;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_CO5;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_CO6;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_C_CY;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_C_XOR;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_D;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_D1;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_D2;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_D3;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_D4;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_D5;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_D6;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_DMUX;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_DO5;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_DO6;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_D_CY;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X48Y123_D_XOR;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_A;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_A1;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_A2;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_A3;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_A4;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_A5;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_A6;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_AO5;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_AO6;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_A_CY;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_A_XOR;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_B;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_B1;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_B2;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_B3;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_B4;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_B5;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_B6;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_BO5;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_BO6;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_B_CY;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_B_XOR;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_C;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_C1;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_C2;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_C3;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_C4;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_C5;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_C6;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_CO5;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_CO6;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_C_CY;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_C_XOR;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_D;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_D1;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_D2;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_D3;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_D4;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_D5;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_D6;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_DO5;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_DO6;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_D_CY;
  wire [0:0] CLBLM_R_X33Y123_SLICE_X49Y123_D_XOR;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_A;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_A1;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_A2;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_A3;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_A4;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_A5;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_A6;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_AMUX;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_AO5;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_AO6;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_A_CY;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_A_XOR;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_B;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_B1;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_B2;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_B3;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_B4;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_B5;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_B6;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_BO5;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_BO6;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_B_CY;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_B_XOR;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_C;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_C1;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_C2;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_C3;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_C4;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_C5;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_C6;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_CO5;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_CO6;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_C_CY;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_C_XOR;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_D;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_D1;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_D2;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_D3;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_D4;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_D5;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_D6;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_DO5;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_DO6;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_D_CY;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X48Y124_D_XOR;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_A;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_A1;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_A2;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_A3;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_A4;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_A5;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_A6;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_AMUX;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_AO5;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_AO6;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_A_CY;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_A_XOR;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_B;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_B1;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_B2;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_B3;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_B4;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_B5;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_B6;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_BO5;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_BO6;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_B_CY;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_B_XOR;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_C;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_C1;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_C2;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_C3;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_C4;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_C5;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_C6;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_CO5;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_CO6;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_C_CY;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_C_XOR;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_D;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_D1;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_D2;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_D3;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_D4;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_D5;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_D6;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_DO5;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_DO6;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_D_CY;
  wire [0:0] CLBLM_R_X33Y124_SLICE_X49Y124_D_XOR;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_A;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_A1;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_A2;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_A3;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_A4;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_A5;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_A6;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_AO5;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_AO6;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_A_CY;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_A_XOR;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_B;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_B1;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_B2;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_B3;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_B4;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_B5;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_B6;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_BO5;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_BO6;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_B_CY;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_B_XOR;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_C;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_C1;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_C2;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_C3;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_C4;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_C5;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_C6;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_CO5;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_CO6;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_C_CY;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_C_XOR;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_D;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_D1;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_D2;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_D3;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_D4;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_D5;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_D6;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_DO5;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_DO6;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_D_CY;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X48Y125_D_XOR;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_A;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_A1;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_A2;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_A3;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_A4;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_A5;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_A6;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_AMUX;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_AO5;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_AO6;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_A_CY;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_A_XOR;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_B;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_B1;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_B2;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_B3;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_B4;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_B5;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_B6;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_BMUX;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_BO5;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_BO6;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_B_CY;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_B_XOR;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_C;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_C1;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_C2;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_C3;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_C4;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_C5;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_C6;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_CO5;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_CO6;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_C_CY;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_C_XOR;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_D;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_D1;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_D2;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_D3;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_D4;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_D5;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_D6;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_DO5;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_DO6;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_D_CY;
  wire [0:0] CLBLM_R_X33Y125_SLICE_X49Y125_D_XOR;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_A;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_A1;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_A2;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_A3;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_A4;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_A5;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_A6;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_AO5;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_AO6;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_A_CY;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_A_XOR;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_B;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_B1;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_B2;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_B3;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_B4;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_B5;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_B6;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_BO5;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_BO6;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_B_CY;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_B_XOR;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_C;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_C1;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_C2;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_C3;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_C4;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_C5;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_C6;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_CO5;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_CO6;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_C_CY;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_C_XOR;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_D;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_D1;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_D2;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_D3;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_D4;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_D5;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_D6;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_DO5;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_DO6;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_D_CY;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X52Y114_D_XOR;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_A;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_A1;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_A2;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_A3;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_A4;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_A5;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_A6;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_AO5;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_AO6;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_A_CY;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_A_XOR;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_B;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_B1;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_B2;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_B3;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_B4;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_B5;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_B6;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_BO5;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_BO6;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_B_CY;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_B_XOR;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_C;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_C1;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_C2;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_C3;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_C4;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_C5;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_C6;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_CO5;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_CO6;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_C_CY;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_C_XOR;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_D;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_D1;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_D2;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_D3;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_D4;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_D5;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_D6;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_DO5;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_DO6;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_D_CY;
  wire [0:0] CLBLM_R_X35Y114_SLICE_X53Y114_D_XOR;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_A;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_A1;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_A2;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_A3;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_A4;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_A5;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_A6;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_AMUX;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_AO5;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_AO6;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_A_CY;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_A_XOR;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_B;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_B1;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_B2;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_B3;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_B4;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_B5;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_B6;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_BO5;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_BO6;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_B_CY;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_B_XOR;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_C;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_C1;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_C2;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_C3;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_C4;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_C5;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_C6;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_CO5;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_CO6;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_C_CY;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_C_XOR;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_D;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_D1;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_D2;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_D3;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_D4;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_D5;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_D6;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_DO5;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_DO6;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_D_CY;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X52Y115_D_XOR;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_A;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_A1;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_A2;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_A3;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_A4;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_A5;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_A6;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_AO5;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_AO6;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_A_CY;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_A_XOR;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_B;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_B1;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_B2;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_B3;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_B4;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_B5;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_B6;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_BO5;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_BO6;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_B_CY;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_B_XOR;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_C;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_C1;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_C2;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_C3;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_C4;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_C5;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_C6;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_CMUX;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_CO5;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_CO6;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_C_CY;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_C_XOR;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_D;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_D1;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_D2;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_D3;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_D4;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_D5;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_D6;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_DO5;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_DO6;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_D_CY;
  wire [0:0] CLBLM_R_X35Y115_SLICE_X53Y115_D_XOR;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_A;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_A1;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_A2;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_A3;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_A4;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_A5;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_A6;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_AMUX;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_AO5;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_AO6;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_A_CY;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_A_XOR;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_B;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_B1;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_B2;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_B3;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_B4;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_B5;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_B6;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_BO5;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_BO6;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_B_CY;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_B_XOR;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_C;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_C1;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_C2;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_C3;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_C4;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_C5;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_C6;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_CO5;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_CO6;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_C_CY;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_C_XOR;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_D;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_D1;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_D2;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_D3;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_D4;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_D5;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_D6;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_DO5;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_DO6;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_D_CY;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X52Y116_D_XOR;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_A;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_A1;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_A2;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_A3;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_A4;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_A5;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_A6;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_AO5;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_AO6;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_A_CY;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_A_XOR;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_B;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_B1;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_B2;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_B3;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_B4;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_B5;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_B6;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_BO5;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_BO6;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_B_CY;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_B_XOR;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_C;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_C1;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_C2;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_C3;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_C4;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_C5;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_C6;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_CO5;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_CO6;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_C_CY;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_C_XOR;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_D;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_D1;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_D2;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_D3;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_D4;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_D5;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_D6;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_DO5;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_DO6;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_D_CY;
  wire [0:0] CLBLM_R_X35Y116_SLICE_X53Y116_D_XOR;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_A;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_A1;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_A2;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_A3;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_A4;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_A5;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_A6;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_AMUX;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_AO5;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_AO6;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_A_CY;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_A_XOR;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_B;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_B1;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_B2;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_B3;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_B4;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_B5;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_B6;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_BO5;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_BO6;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_B_CY;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_B_XOR;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_C;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_C1;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_C2;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_C3;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_C4;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_C5;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_C6;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_CO5;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_CO6;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_C_CY;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_C_XOR;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_D;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_D1;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_D2;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_D3;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_D4;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_D5;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_D6;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_DO5;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_DO6;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_D_CY;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X52Y117_D_XOR;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_A;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_A1;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_A2;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_A3;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_A4;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_A5;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_A6;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_AO5;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_AO6;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_A_CY;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_A_XOR;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_B;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_B1;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_B2;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_B3;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_B4;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_B5;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_B6;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_BMUX;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_BO5;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_BO6;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_B_CY;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_B_XOR;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_C;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_C1;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_C2;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_C3;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_C4;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_C5;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_C6;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_CO5;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_CO6;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_C_CY;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_C_XOR;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_D;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_D1;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_D2;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_D3;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_D4;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_D5;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_D6;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_DO5;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_DO6;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_D_CY;
  wire [0:0] CLBLM_R_X35Y117_SLICE_X53Y117_D_XOR;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_A;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_A1;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_A2;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_A3;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_A4;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_A5;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_A6;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_AMUX;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_AO5;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_AO6;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_AX;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_A_CY;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_A_XOR;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_B;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_B1;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_B2;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_B3;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_B4;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_B5;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_B6;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_BMUX;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_BO5;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_BO6;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_BX;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_B_CY;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_B_XOR;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_C;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_C1;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_C2;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_C3;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_C4;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_C5;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_C6;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_CMUX;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_CO5;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_CO6;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_COUT;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_CX;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_C_CY;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_C_XOR;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_D;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_D1;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_D2;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_D3;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_D4;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_D5;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_D6;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_DMUX;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_DO5;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_DO6;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_DX;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_D_CY;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X52Y118_D_XOR;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_A;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_A1;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_A2;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_A3;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_A4;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_A5;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_A6;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_AMUX;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_AO5;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_AO6;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_A_CY;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_A_XOR;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_B;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_B1;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_B2;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_B3;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_B4;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_B5;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_B6;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_BMUX;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_BO5;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_BO6;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_B_CY;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_B_XOR;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_C;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_C1;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_C2;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_C3;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_C4;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_C5;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_C6;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_CO5;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_CO6;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_C_CY;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_C_XOR;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_D;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_D1;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_D2;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_D3;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_D4;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_D5;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_D6;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_DO5;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_DO6;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_D_CY;
  wire [0:0] CLBLM_R_X35Y118_SLICE_X53Y118_D_XOR;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_A;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_A1;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_A2;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_A3;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_A4;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_A5;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_A6;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_AMUX;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_AO5;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_AO6;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_AX;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_A_CY;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_A_XOR;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_B;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_B1;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_B2;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_B3;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_B4;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_B5;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_B6;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_BMUX;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_BO5;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_BO6;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_BX;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_B_CY;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_B_XOR;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_C;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_C1;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_C2;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_C3;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_C4;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_C5;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_C6;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_CIN;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_CMUX;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_CO5;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_CO6;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_COUT;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_CX;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_C_CY;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_C_XOR;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_D;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_D1;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_D2;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_D3;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_D4;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_D5;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_D6;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_DMUX;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_DO5;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_DO6;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_DX;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_D_CY;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X52Y119_D_XOR;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_A;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_A1;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_A2;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_A3;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_A4;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_A5;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_A6;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_AO5;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_AO6;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_A_CY;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_A_XOR;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_B;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_B1;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_B2;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_B3;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_B4;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_B5;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_B6;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_BO5;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_BO6;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_B_CY;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_B_XOR;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_C;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_C1;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_C2;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_C3;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_C4;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_C5;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_C6;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_CO5;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_CO6;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_C_CY;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_C_XOR;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_D;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_D1;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_D2;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_D3;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_D4;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_D5;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_D6;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_DO5;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_DO6;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_D_CY;
  wire [0:0] CLBLM_R_X35Y119_SLICE_X53Y119_D_XOR;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_A;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_A1;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_A2;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_A3;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_A4;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_A5;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_A6;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_AMUX;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_AO5;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_AO6;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_AX;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_A_CY;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_A_XOR;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_B;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_B1;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_B2;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_B3;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_B4;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_B5;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_B6;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_BMUX;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_BO5;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_BO6;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_BX;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_B_CY;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_B_XOR;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_C;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_C1;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_C2;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_C3;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_C4;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_C5;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_C6;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_CIN;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_CMUX;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_CO5;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_CO6;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_COUT;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_CX;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_C_CY;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_C_XOR;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_D;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_D1;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_D2;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_D3;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_D4;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_D5;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_D6;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_DMUX;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_DO5;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_DO6;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_DX;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_D_CY;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X52Y120_D_XOR;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_A;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_A1;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_A2;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_A3;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_A4;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_A5;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_A6;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_AMUX;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_AO5;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_AO6;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_AX;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_A_CY;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_A_XOR;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_B;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_B1;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_B2;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_B3;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_B4;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_B5;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_B6;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_BMUX;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_BO5;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_BO6;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_BX;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_B_CY;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_B_XOR;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_C;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_C1;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_C2;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_C3;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_C4;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_C5;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_C6;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_CMUX;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_CO5;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_CO6;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_COUT;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_CX;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_C_CY;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_C_XOR;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_D;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_D1;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_D2;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_D3;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_D4;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_D5;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_D6;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_DMUX;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_DO5;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_DO6;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_DX;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_D_CY;
  wire [0:0] CLBLM_R_X35Y120_SLICE_X53Y120_D_XOR;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_A;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_A1;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_A2;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_A3;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_A4;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_A5;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_A6;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_AMUX;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_AO5;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_AO6;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_AX;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_A_CY;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_A_XOR;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_B;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_B1;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_B2;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_B3;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_B4;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_B5;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_B6;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_BMUX;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_BO5;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_BO6;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_BX;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_B_CY;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_B_XOR;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_C;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_C1;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_C2;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_C3;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_C4;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_C5;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_C6;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_CIN;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_CMUX;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_CO5;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_CO6;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_COUT;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_CX;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_C_CY;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_C_XOR;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_D;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_D1;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_D2;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_D3;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_D4;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_D5;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_D6;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_DMUX;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_DO5;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_DO6;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_DX;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_D_CY;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X52Y121_D_XOR;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_A;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_A1;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_A2;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_A3;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_A4;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_A5;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_A6;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_AMUX;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_AO5;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_AO6;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_AX;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_A_CY;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_A_XOR;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_B;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_B1;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_B2;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_B3;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_B4;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_B5;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_B6;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_BMUX;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_BO5;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_BO6;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_BX;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_B_CY;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_B_XOR;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_C;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_C1;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_C2;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_C3;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_C4;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_C5;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_C6;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_CIN;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_CMUX;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_CO5;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_CO6;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_COUT;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_CX;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_C_CY;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_C_XOR;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_D;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_D1;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_D2;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_D3;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_D4;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_D5;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_D6;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_DMUX;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_DO5;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_DO6;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_DX;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_D_CY;
  wire [0:0] CLBLM_R_X35Y121_SLICE_X53Y121_D_XOR;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_A;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_A1;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_A2;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_A3;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_A4;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_A5;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_A6;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_AMUX;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_AO5;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_AO6;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_AX;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_A_CY;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_A_XOR;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_B;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_B1;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_B2;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_B3;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_B4;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_B5;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_B6;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_BMUX;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_BO5;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_BO6;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_BX;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_B_CY;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_B_XOR;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_C;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_C1;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_C2;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_C3;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_C4;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_C5;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_C6;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_CIN;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_CMUX;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_CO5;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_CO6;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_COUT;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_CX;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_C_CY;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_C_XOR;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_D;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_D1;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_D2;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_D3;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_D4;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_D5;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_D6;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_DMUX;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_DO5;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_DO6;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_DX;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_D_CY;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X52Y122_D_XOR;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_A;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_A1;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_A2;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_A3;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_A4;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_A5;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_A6;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_AMUX;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_AO5;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_AO6;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_AX;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_A_CY;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_A_XOR;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_B;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_B1;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_B2;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_B3;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_B4;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_B5;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_B6;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_BMUX;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_BO5;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_BO6;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_BX;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_B_CY;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_B_XOR;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_C;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_C1;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_C2;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_C3;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_C4;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_C5;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_C6;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_CIN;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_CMUX;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_CO5;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_CO6;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_COUT;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_CX;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_C_CY;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_C_XOR;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_D;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_D1;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_D2;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_D3;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_D4;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_D5;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_D6;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_DMUX;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_DO5;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_DO6;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_DX;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_D_CY;
  wire [0:0] CLBLM_R_X35Y122_SLICE_X53Y122_D_XOR;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_A;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_A1;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_A2;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_A3;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_A4;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_A5;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_A6;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_AMUX;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_AO5;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_AO6;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_AX;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_A_CY;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_A_XOR;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_B;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_B1;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_B2;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_B3;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_B4;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_B5;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_B6;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_BMUX;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_BO5;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_BO6;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_BX;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_B_CY;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_B_XOR;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_C;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_C1;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_C2;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_C3;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_C4;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_C5;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_C6;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_CIN;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_CMUX;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_CO5;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_CO6;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_COUT;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_CX;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_C_CY;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_C_XOR;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_D;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_D1;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_D2;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_D3;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_D4;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_D5;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_D6;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_DMUX;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_DO5;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_DO6;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_DX;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_D_CY;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X52Y123_D_XOR;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_A;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_A1;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_A2;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_A3;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_A4;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_A5;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_A6;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_AMUX;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_AO5;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_AO6;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_AX;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_A_CY;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_A_XOR;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_B;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_B1;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_B2;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_B3;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_B4;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_B5;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_B6;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_BMUX;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_BO5;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_BO6;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_BX;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_B_CY;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_B_XOR;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_C;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_C1;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_C2;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_C3;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_C4;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_C5;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_C6;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_CIN;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_CMUX;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_CO5;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_CO6;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_COUT;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_CX;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_C_CY;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_C_XOR;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_D;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_D1;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_D2;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_D3;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_D4;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_D5;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_D6;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_DMUX;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_DO5;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_DO6;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_DX;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_D_CY;
  wire [0:0] CLBLM_R_X35Y123_SLICE_X53Y123_D_XOR;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_A;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_A1;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_A2;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_A3;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_A4;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_A5;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_A6;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_AMUX;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_AO5;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_AO6;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_AX;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_A_CY;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_A_XOR;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_B;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_B1;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_B2;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_B3;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_B4;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_B5;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_B6;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_BMUX;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_BO5;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_BO6;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_BX;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_B_CY;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_B_XOR;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_C;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_C1;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_C2;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_C3;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_C4;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_C5;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_C6;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_CIN;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_CMUX;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_CO5;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_CO6;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_COUT;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_CX;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_C_CY;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_C_XOR;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_D;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_D1;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_D2;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_D3;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_D4;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_D5;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_D6;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_DMUX;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_DO5;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_DO6;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_DX;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_D_CY;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X52Y124_D_XOR;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_A;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_A1;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_A2;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_A3;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_A4;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_A5;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_A6;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_AMUX;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_AO5;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_AO6;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_AX;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_A_CY;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_A_XOR;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_B;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_B1;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_B2;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_B3;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_B4;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_B5;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_B6;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_BMUX;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_BO5;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_BO6;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_BX;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_B_CY;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_B_XOR;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_C;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_C1;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_C2;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_C3;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_C4;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_C5;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_C6;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_CIN;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_CMUX;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_CO5;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_CO6;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_COUT;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_CX;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_C_CY;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_C_XOR;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_D;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_D1;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_D2;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_D3;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_D4;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_D5;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_D6;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_DMUX;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_DO5;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_DO6;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_DX;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_D_CY;
  wire [0:0] CLBLM_R_X35Y124_SLICE_X53Y124_D_XOR;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_A;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_A1;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_A2;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_A3;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_A4;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_A5;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_A6;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_AMUX;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_AO5;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_AO6;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_AX;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_A_CY;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_A_XOR;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_B;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_B1;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_B2;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_B3;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_B4;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_B5;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_B6;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_BMUX;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_BO5;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_BO6;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_BX;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_B_CY;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_B_XOR;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_C;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_C1;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_C2;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_C3;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_C4;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_C5;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_C6;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_CIN;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_CMUX;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_CO5;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_CO6;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_COUT;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_CX;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_C_CY;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_C_XOR;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_D;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_D1;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_D2;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_D3;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_D4;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_D5;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_D6;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_DMUX;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_DO5;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_DO6;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_DX;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_D_CY;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X52Y125_D_XOR;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_A;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_A1;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_A2;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_A3;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_A4;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_A5;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_A6;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_AMUX;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_AO5;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_AO6;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_AX;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_A_CY;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_A_XOR;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_B;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_B1;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_B2;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_B3;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_B4;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_B5;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_B6;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_BMUX;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_BO5;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_BO6;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_BX;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_B_CY;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_B_XOR;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_C;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_C1;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_C2;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_C3;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_C4;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_C5;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_C6;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_CIN;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_CMUX;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_CO5;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_CO6;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_COUT;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_CX;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_C_CY;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_C_XOR;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_D;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_D1;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_D2;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_D3;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_D4;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_D5;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_D6;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_DMUX;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_DO5;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_DO6;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_DX;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_D_CY;
  wire [0:0] CLBLM_R_X35Y125_SLICE_X53Y125_D_XOR;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_A;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_A1;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_A2;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_A3;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_A4;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_A5;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_A6;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_AO5;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_AO6;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_A_CY;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_A_XOR;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_B;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_B1;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_B2;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_B3;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_B4;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_B5;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_B6;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_BO5;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_BO6;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_B_CY;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_B_XOR;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_C;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_C1;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_C2;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_C3;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_C4;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_C5;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_C6;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_CO5;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_CO6;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_C_CY;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_C_XOR;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_D;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_D1;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_D2;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_D3;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_D4;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_D5;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_D6;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_DO5;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_DO6;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_D_CY;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X52Y126_D_XOR;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_A;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_A1;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_A2;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_A3;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_A4;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_A5;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_A6;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_AMUX;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_AO5;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_AO6;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_AX;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_A_CY;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_A_XOR;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_B;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_B1;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_B2;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_B3;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_B4;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_B5;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_B6;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_BMUX;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_BO5;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_BO6;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_BX;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_B_CY;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_B_XOR;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_C;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_C1;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_C2;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_C3;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_C4;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_C5;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_C6;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_CIN;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_CMUX;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_CO5;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_CO6;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_COUT;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_CX;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_C_CY;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_C_XOR;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_D;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_D1;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_D2;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_D3;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_D4;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_D5;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_D6;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_DMUX;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_DO5;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_DO6;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_DX;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_D_CY;
  wire [0:0] CLBLM_R_X35Y126_SLICE_X53Y126_D_XOR;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_A;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_A1;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_A2;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_A3;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_A4;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_A5;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_A6;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_AO5;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_AO6;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_A_CY;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_A_XOR;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_B;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_B1;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_B2;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_B3;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_B4;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_B5;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_B6;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_BO5;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_BO6;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_B_CY;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_B_XOR;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_C;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_C1;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_C2;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_C3;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_C4;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_C5;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_C6;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_CO5;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_CO6;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_C_CY;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_C_XOR;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_D;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_D1;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_D2;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_D3;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_D4;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_D5;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_D6;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_DMUX;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_DO5;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_DO6;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_D_CY;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X52Y127_D_XOR;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_A;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_A1;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_A2;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_A3;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_A4;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_A5;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_A6;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_AMUX;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_AO5;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_AO6;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_AX;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_A_CY;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_A_XOR;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_B;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_B1;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_B2;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_B3;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_B4;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_B5;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_B6;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_BMUX;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_BO5;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_BO6;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_BX;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_B_CY;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_B_XOR;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_C;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_C1;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_C2;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_C3;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_C4;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_C5;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_C6;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_CIN;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_CMUX;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_CO5;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_CO6;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_COUT;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_CX;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_C_CY;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_C_XOR;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_D;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_D1;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_D2;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_D3;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_D4;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_D5;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_D6;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_DMUX;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_DO5;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_DO6;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_DX;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_D_CY;
  wire [0:0] CLBLM_R_X35Y127_SLICE_X53Y127_D_XOR;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_A;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_A1;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_A2;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_A3;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_A4;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_A5;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_A6;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_AO5;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_AO6;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_A_CY;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_A_XOR;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_B;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_B1;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_B2;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_B3;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_B4;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_B5;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_B6;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_BMUX;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_BO5;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_BO6;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_B_CY;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_B_XOR;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_C;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_C1;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_C2;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_C3;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_C4;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_C5;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_C6;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_CO5;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_CO6;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_C_CY;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_C_XOR;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_D;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_D1;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_D2;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_D3;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_D4;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_D5;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_D6;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_DO5;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_DO6;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_D_CY;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X52Y128_D_XOR;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_A;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_A1;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_A2;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_A3;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_A4;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_A5;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_A6;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_AO5;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_AO6;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_A_CY;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_A_XOR;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_B;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_B1;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_B2;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_B3;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_B4;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_B5;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_B6;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_BMUX;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_BO5;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_BO6;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_B_CY;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_B_XOR;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_C;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_C1;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_C2;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_C3;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_C4;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_C5;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_C6;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_CO5;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_CO6;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_C_CY;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_C_XOR;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_D;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_D1;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_D2;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_D3;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_D4;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_D5;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_D6;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_DO5;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_DO6;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_D_CY;
  wire [0:0] CLBLM_R_X35Y128_SLICE_X53Y128_D_XOR;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_A;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_A1;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_A2;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_A3;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_A4;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_A5;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_A6;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_AO5;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_AO6;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_A_CY;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_A_XOR;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_B;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_B1;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_B2;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_B3;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_B4;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_B5;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_B6;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_BO5;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_BO6;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_B_CY;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_B_XOR;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_C;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_C1;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_C2;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_C3;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_C4;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_C5;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_C6;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_CO5;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_CO6;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_C_CY;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_C_XOR;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_D;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_D1;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_D2;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_D3;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_D4;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_D5;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_D6;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_DO5;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_DO6;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_D_CY;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X52Y129_D_XOR;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_A;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_A1;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_A2;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_A3;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_A4;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_A5;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_A6;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_AO5;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_AO6;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_A_CY;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_A_XOR;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_B;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_B1;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_B2;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_B3;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_B4;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_B5;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_B6;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_BO5;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_BO6;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_B_CY;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_B_XOR;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_C;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_C1;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_C2;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_C3;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_C4;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_C5;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_C6;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_CO5;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_CO6;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_C_CY;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_C_XOR;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_D;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_D1;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_D2;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_D3;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_D4;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_D5;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_D6;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_DO5;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_DO6;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_D_CY;
  wire [0:0] CLBLM_R_X35Y129_SLICE_X53Y129_D_XOR;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_A;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_A1;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_A2;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_A3;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_A4;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_A5;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_A6;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_AMUX;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_AO5;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_AO6;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_A_CY;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_A_XOR;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_B;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_B1;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_B2;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_B3;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_B4;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_B5;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_B6;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_BO5;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_BO6;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_B_CY;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_B_XOR;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_C;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_C1;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_C2;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_C3;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_C4;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_C5;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_C6;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_CO5;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_CO6;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_C_CY;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_C_XOR;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_D;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_D1;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_D2;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_D3;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_D4;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_D5;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_D6;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_DO5;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_DO6;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_D_CY;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_D_XOR;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_A;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_A1;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_A2;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_A3;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_A4;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_A5;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_A6;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_AO5;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_AO6;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_A_CY;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_A_XOR;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_B;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_B1;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_B2;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_B3;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_B4;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_B5;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_B6;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_BO5;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_BO6;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_B_CY;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_B_XOR;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_C;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_C1;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_C2;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_C3;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_C4;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_C5;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_C6;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_CO5;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_CO6;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_C_CY;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_C_XOR;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_D;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_D1;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_D2;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_D3;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_D4;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_D5;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_D6;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_DO5;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_DO6;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_D_CY;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_D_XOR;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_A;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_A1;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_A2;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_A3;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_A4;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_A5;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_A6;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_AO5;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_AO6;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_A_CY;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_A_XOR;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_B;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_B1;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_B2;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_B3;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_B4;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_B5;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_B6;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_BO5;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_BO6;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_B_CY;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_B_XOR;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_C;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_C1;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_C2;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_C3;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_C4;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_C5;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_C6;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_CO5;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_CO6;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_C_CY;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_C_XOR;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_D;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_D1;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_D2;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_D3;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_D4;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_D5;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_D6;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_DO5;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_DO6;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_D_CY;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X56Y118_D_XOR;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_A;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_A1;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_A2;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_A3;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_A4;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_A5;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_A6;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_AMUX;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_AO5;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_AO6;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_A_CY;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_A_XOR;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_B;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_B1;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_B2;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_B3;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_B4;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_B5;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_B6;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_BMUX;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_BO5;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_BO6;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_B_CY;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_B_XOR;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_C;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_C1;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_C2;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_C3;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_C4;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_C5;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_C6;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_CO5;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_CO6;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_C_CY;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_C_XOR;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_D;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_D1;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_D2;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_D3;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_D4;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_D5;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_D6;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_DO5;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_DO6;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_D_CY;
  wire [0:0] CLBLM_R_X37Y118_SLICE_X57Y118_D_XOR;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_A;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_A1;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_A2;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_A3;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_A4;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_A5;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_A6;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_AO5;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_AO6;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_A_CY;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_A_XOR;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_B;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_B1;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_B2;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_B3;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_B4;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_B5;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_B6;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_BO5;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_BO6;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_B_CY;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_B_XOR;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_C;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_C1;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_C2;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_C3;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_C4;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_C5;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_C6;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_CO5;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_CO6;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_C_CY;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_C_XOR;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_D;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_D1;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_D2;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_D3;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_D4;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_D5;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_D6;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_DO5;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_DO6;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_D_CY;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_D_XOR;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_A;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_A1;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_A2;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_A3;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_A4;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_A5;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_A6;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_AO5;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_AO6;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_A_CY;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_A_XOR;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_B;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_B1;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_B2;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_B3;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_B4;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_B5;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_B6;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_BMUX;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_BO5;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_BO6;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_B_CY;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_B_XOR;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_C;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_C1;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_C2;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_C3;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_C4;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_C5;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_C6;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_CO5;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_CO6;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_C_CY;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_C_XOR;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_D;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_D1;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_D2;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_D3;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_D4;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_D5;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_D6;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_DO5;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_DO6;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_D_CY;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_D_XOR;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_A;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_A1;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_A2;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_A3;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_A4;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_A5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_A6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_AO5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_AO6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_A_CY;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_A_XOR;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_B;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_B1;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_B2;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_B3;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_B4;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_B5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_B6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_BO5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_BO6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_B_CY;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_B_XOR;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_C;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_C1;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_C2;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_C3;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_C4;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_C5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_C6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_CO5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_CO6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_C_CY;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_C_XOR;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_D;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_D1;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_D2;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_D3;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_D4;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_D5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_D6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_DO5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_DO6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_D_CY;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_D_XOR;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_A;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_A1;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_A2;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_A3;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_A4;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_A5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_A6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_AO5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_AO6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_A_CY;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_A_XOR;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_B;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_B1;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_B2;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_B3;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_B4;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_B5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_B6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_BO5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_BO6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_B_CY;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_B_XOR;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_C;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_C1;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_C2;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_C3;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_C4;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_C5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_C6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_CO5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_CO6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_C_CY;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_C_XOR;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_D;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_D1;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_D2;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_D3;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_D4;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_D5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_D6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_DO5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_DO6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_D_CY;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_D_XOR;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_A;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_A1;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_A2;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_A3;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_A4;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_A5;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_A6;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_AO5;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_AO6;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_A_CY;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_A_XOR;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_B;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_B1;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_B2;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_B3;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_B4;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_B5;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_B6;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_BO5;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_BO6;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_B_CY;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_B_XOR;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_C;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_C1;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_C2;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_C3;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_C4;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_C5;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_C6;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_CO5;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_CO6;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_C_CY;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_C_XOR;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_D;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_D1;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_D2;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_D3;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_D4;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_D5;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_D6;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_DO5;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_DO6;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_D_CY;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X56Y121_D_XOR;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_A;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_A1;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_A2;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_A3;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_A4;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_A5;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_A6;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_AO5;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_AO6;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_A_CY;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_A_XOR;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_B;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_B1;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_B2;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_B3;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_B4;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_B5;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_B6;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_BMUX;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_BO5;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_BO6;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_B_CY;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_B_XOR;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_C;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_C1;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_C2;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_C3;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_C4;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_C5;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_C6;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_CO5;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_CO6;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_C_CY;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_C_XOR;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_D;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_D1;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_D2;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_D3;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_D4;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_D5;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_D6;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_DMUX;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_DO5;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_DO6;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_D_CY;
  wire [0:0] CLBLM_R_X37Y121_SLICE_X57Y121_D_XOR;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_A;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_A1;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_A2;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_A3;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_A4;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_A5;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_A6;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_AO5;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_AO6;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_A_CY;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_A_XOR;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_B;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_B1;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_B2;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_B3;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_B4;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_B5;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_B6;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_BO5;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_BO6;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_B_CY;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_B_XOR;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_C;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_C1;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_C2;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_C3;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_C4;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_C5;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_C6;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_CO5;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_CO6;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_C_CY;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_C_XOR;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_D;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_D1;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_D2;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_D3;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_D4;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_D5;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_D6;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_DO5;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_DO6;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_D_CY;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X56Y122_D_XOR;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_A;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_A1;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_A2;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_A3;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_A4;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_A5;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_A6;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_AO5;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_AO6;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_A_CY;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_A_XOR;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_B;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_B1;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_B2;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_B3;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_B4;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_B5;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_B6;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_BO5;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_BO6;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_B_CY;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_B_XOR;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_C;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_C1;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_C2;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_C3;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_C4;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_C5;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_C6;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_CMUX;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_CO5;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_CO6;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_C_CY;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_C_XOR;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_D;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_D1;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_D2;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_D3;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_D4;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_D5;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_D6;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_DO5;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_DO6;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_D_CY;
  wire [0:0] CLBLM_R_X37Y122_SLICE_X57Y122_D_XOR;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_A;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_A1;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_A2;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_A3;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_A4;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_A5;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_A6;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_AO5;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_AO6;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_A_CY;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_A_XOR;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_B;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_B1;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_B2;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_B3;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_B4;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_B5;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_B6;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_BO5;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_BO6;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_B_CY;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_B_XOR;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_C;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_C1;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_C2;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_C3;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_C4;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_C5;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_C6;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_CMUX;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_CO5;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_CO6;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_C_CY;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_C_XOR;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_D;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_D1;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_D2;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_D3;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_D4;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_D5;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_D6;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_DMUX;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_DO5;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_DO6;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_D_CY;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X56Y123_D_XOR;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_A;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_A1;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_A2;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_A3;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_A4;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_A5;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_A6;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_AO5;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_AO6;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_A_CY;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_A_XOR;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_B;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_B1;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_B2;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_B3;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_B4;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_B5;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_B6;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_BMUX;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_BO5;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_BO6;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_B_CY;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_B_XOR;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_C;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_C1;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_C2;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_C3;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_C4;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_C5;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_C6;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_CO5;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_CO6;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_C_CY;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_C_XOR;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_D;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_D1;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_D2;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_D3;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_D4;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_D5;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_D6;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_DMUX;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_DO5;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_DO6;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_D_CY;
  wire [0:0] CLBLM_R_X37Y123_SLICE_X57Y123_D_XOR;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_A;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_A1;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_A2;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_A3;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_A4;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_A5;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_A6;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_AO5;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_AO6;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_A_CY;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_A_XOR;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_B;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_B1;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_B2;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_B3;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_B4;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_B5;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_B6;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_BMUX;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_BO5;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_BO6;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_B_CY;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_B_XOR;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_C;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_C1;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_C2;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_C3;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_C4;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_C5;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_C6;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_CO5;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_CO6;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_C_CY;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_C_XOR;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_D;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_D1;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_D2;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_D3;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_D4;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_D5;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_D6;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_DO5;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_DO6;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_D_CY;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X56Y124_D_XOR;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_A;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_A1;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_A2;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_A3;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_A4;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_A5;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_A6;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_AO5;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_AO6;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_A_CY;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_A_XOR;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_B;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_B1;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_B2;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_B3;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_B4;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_B5;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_B6;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_BO5;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_BO6;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_B_CY;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_B_XOR;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_C;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_C1;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_C2;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_C3;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_C4;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_C5;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_C6;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_CO5;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_CO6;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_C_CY;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_C_XOR;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_D;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_D1;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_D2;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_D3;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_D4;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_D5;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_D6;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_DO5;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_DO6;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_D_CY;
  wire [0:0] CLBLM_R_X37Y124_SLICE_X57Y124_D_XOR;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_A;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_A1;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_A2;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_A3;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_A4;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_A5;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_A6;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_AO5;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_AO6;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_A_CY;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_A_XOR;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_B;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_B1;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_B2;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_B3;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_B4;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_B5;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_B6;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_BO5;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_BO6;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_B_CY;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_B_XOR;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_C;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_C1;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_C2;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_C3;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_C4;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_C5;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_C6;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_CO5;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_CO6;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_C_CY;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_C_XOR;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_D;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_D1;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_D2;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_D3;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_D4;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_D5;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_D6;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_DO5;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_DO6;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_D_CY;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X56Y125_D_XOR;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_A;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_A1;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_A2;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_A3;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_A4;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_A5;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_A6;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_AO5;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_AO6;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_A_CY;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_A_XOR;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_B;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_B1;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_B2;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_B3;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_B4;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_B5;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_B6;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_BO5;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_BO6;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_B_CY;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_B_XOR;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_C;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_C1;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_C2;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_C3;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_C4;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_C5;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_C6;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_CO5;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_CO6;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_C_CY;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_C_XOR;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_D;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_D1;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_D2;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_D3;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_D4;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_D5;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_D6;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_DO5;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_DO6;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_D_CY;
  wire [0:0] CLBLM_R_X37Y125_SLICE_X57Y125_D_XOR;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_A;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_A1;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_A2;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_A3;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_A4;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_A5;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_A6;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_AMUX;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_AO5;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_AO6;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_A_CY;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_A_XOR;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_B;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_B1;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_B2;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_B3;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_B4;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_B5;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_B6;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_BO5;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_BO6;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_B_CY;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_B_XOR;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_C;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_C1;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_C2;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_C3;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_C4;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_C5;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_C6;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_CO5;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_CO6;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_C_CY;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_C_XOR;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_D;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_D1;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_D2;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_D3;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_D4;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_D5;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_D6;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_DO5;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_DO6;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_D_CY;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X56Y126_D_XOR;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_A;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_A1;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_A2;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_A3;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_A4;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_A5;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_A6;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_AO5;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_AO6;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_A_CY;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_A_XOR;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_B;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_B1;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_B2;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_B3;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_B4;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_B5;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_B6;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_BO5;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_BO6;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_B_CY;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_B_XOR;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_C;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_C1;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_C2;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_C3;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_C4;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_C5;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_C6;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_CMUX;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_CO5;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_CO6;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_C_CY;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_C_XOR;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_D;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_D1;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_D2;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_D3;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_D4;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_D5;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_D6;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_DO5;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_DO6;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_D_CY;
  wire [0:0] CLBLM_R_X37Y126_SLICE_X57Y126_D_XOR;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_A;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_A1;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_A2;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_A3;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_A4;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_A5;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_A6;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_AO5;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_AO6;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_A_CY;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_A_XOR;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_B;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_B1;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_B2;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_B3;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_B4;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_B5;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_B6;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_BO5;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_BO6;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_B_CY;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_B_XOR;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_C;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_C1;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_C2;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_C3;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_C4;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_C5;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_C6;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_CO5;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_CO6;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_C_CY;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_C_XOR;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_D;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_D1;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_D2;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_D3;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_D4;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_D5;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_D6;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_DO5;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_DO6;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_D_CY;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X56Y127_D_XOR;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_A;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_A1;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_A2;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_A3;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_A4;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_A5;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_A6;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_AO5;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_AO6;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_A_CY;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_A_XOR;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_B;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_B1;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_B2;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_B3;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_B4;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_B5;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_B6;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_BO5;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_BO6;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_B_CY;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_B_XOR;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_C;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_C1;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_C2;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_C3;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_C4;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_C5;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_C6;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_CO5;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_CO6;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_C_CY;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_C_XOR;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_D;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_D1;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_D2;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_D3;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_D4;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_D5;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_D6;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_DO5;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_DO6;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_D_CY;
  wire [0:0] CLBLM_R_X37Y127_SLICE_X57Y127_D_XOR;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_A;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_A1;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_A2;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_A3;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_A4;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_A5;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_A6;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_AO5;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_AO6;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_A_CY;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_A_XOR;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_B;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_B1;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_B2;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_B3;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_B4;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_B5;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_B6;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_BO5;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_BO6;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_B_CY;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_B_XOR;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_C;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_C1;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_C2;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_C3;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_C4;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_C5;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_C6;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_CO5;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_CO6;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_C_CY;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_C_XOR;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_D;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_D1;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_D2;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_D3;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_D4;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_D5;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_D6;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_DO5;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_DO6;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_D_CY;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X56Y128_D_XOR;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_A;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_A1;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_A2;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_A3;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_A4;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_A5;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_A6;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_AO5;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_AO6;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_A_CY;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_A_XOR;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_B;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_B1;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_B2;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_B3;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_B4;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_B5;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_B6;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_BO5;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_BO6;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_B_CY;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_B_XOR;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_C;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_C1;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_C2;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_C3;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_C4;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_C5;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_C6;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_CO5;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_CO6;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_C_CY;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_C_XOR;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_D;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_D1;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_D2;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_D3;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_D4;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_D5;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_D6;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_DO5;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_DO6;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_D_CY;
  wire [0:0] CLBLM_R_X37Y128_SLICE_X57Y128_D_XOR;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_I;
  wire [0:0] LIOB33_SING_X0Y149_IOB_X0Y149_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_I;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_I;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_I;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_I;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_I;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_I;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_I;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_I;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_I;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_I;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_I;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_I;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_I;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_I;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_I;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_I;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_I;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_I;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_I;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y129_I;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y130_I;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y131_I;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y132_I;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y133_I;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y134_I;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y135_I;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y136_I;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_I;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y138_I;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y139_I;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y140_I;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y141_I;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y142_I;
  wire [0:0] LIOB33_X0Y143_IOB_X0Y143_I;
  wire [0:0] LIOB33_X0Y143_IOB_X0Y144_I;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y145_I;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y146_I;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y147_I;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y148_I;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y65_O;
  wire [0:0] LIOI3_SING_X0Y100_ILOGIC_X0Y100_D;
  wire [0:0] LIOI3_SING_X0Y100_ILOGIC_X0Y100_O;
  wire [0:0] LIOI3_SING_X0Y149_ILOGIC_X0Y149_D;
  wire [0:0] LIOI3_SING_X0Y149_ILOGIC_X0Y149_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y119_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y119_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y120_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y120_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y131_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y131_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y132_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y132_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_ILOGIC_X0Y143_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_ILOGIC_X0Y143_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_ILOGIC_X0Y144_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_ILOGIC_X0Y144_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y138_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y138_O;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_O;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_O;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_D;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_O;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y110_D;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y110_O;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y111_D;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y111_O;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_D;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_O;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y115_D;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y115_O;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y116_D;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y116_O;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y117_D;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y117_O;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y118_D;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y118_O;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y121_D;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y121_O;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y122_D;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y122_O;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y123_D;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y123_O;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y124_D;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y124_O;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y125_D;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y125_O;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y126_D;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y126_O;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y127_D;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y127_O;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y128_D;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y128_O;
  wire [0:0] LIOI3_X0Y129_ILOGIC_X0Y129_D;
  wire [0:0] LIOI3_X0Y129_ILOGIC_X0Y129_O;
  wire [0:0] LIOI3_X0Y129_ILOGIC_X0Y130_D;
  wire [0:0] LIOI3_X0Y129_ILOGIC_X0Y130_O;
  wire [0:0] LIOI3_X0Y133_ILOGIC_X0Y133_D;
  wire [0:0] LIOI3_X0Y133_ILOGIC_X0Y133_O;
  wire [0:0] LIOI3_X0Y133_ILOGIC_X0Y134_D;
  wire [0:0] LIOI3_X0Y133_ILOGIC_X0Y134_O;
  wire [0:0] LIOI3_X0Y135_ILOGIC_X0Y135_D;
  wire [0:0] LIOI3_X0Y135_ILOGIC_X0Y135_O;
  wire [0:0] LIOI3_X0Y135_ILOGIC_X0Y136_D;
  wire [0:0] LIOI3_X0Y135_ILOGIC_X0Y136_O;
  wire [0:0] LIOI3_X0Y139_ILOGIC_X0Y139_D;
  wire [0:0] LIOI3_X0Y139_ILOGIC_X0Y139_O;
  wire [0:0] LIOI3_X0Y139_ILOGIC_X0Y140_D;
  wire [0:0] LIOI3_X0Y139_ILOGIC_X0Y140_O;
  wire [0:0] LIOI3_X0Y141_ILOGIC_X0Y141_D;
  wire [0:0] LIOI3_X0Y141_ILOGIC_X0Y141_O;
  wire [0:0] LIOI3_X0Y141_ILOGIC_X0Y142_D;
  wire [0:0] LIOI3_X0Y141_ILOGIC_X0Y142_O;
  wire [0:0] LIOI3_X0Y145_ILOGIC_X0Y145_D;
  wire [0:0] LIOI3_X0Y145_ILOGIC_X0Y145_O;
  wire [0:0] LIOI3_X0Y145_ILOGIC_X0Y146_D;
  wire [0:0] LIOI3_X0Y145_ILOGIC_X0Y146_O;
  wire [0:0] LIOI3_X0Y147_ILOGIC_X0Y147_D;
  wire [0:0] LIOI3_X0Y147_ILOGIC_X0Y147_O;
  wire [0:0] LIOI3_X0Y147_ILOGIC_X0Y148_D;
  wire [0:0] LIOI3_X0Y147_ILOGIC_X0Y148_O;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y65_D1;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y65_OQ;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y65_T1;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y65_TQ;
  wire [0:0] RIOB33_SING_X105Y100_IOB_X1Y100_I;
  wire [0:0] RIOB33_SING_X105Y149_IOB_X1Y149_O;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y101_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y102_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y103_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y104_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y105_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y106_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y107_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y108_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y109_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y110_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y111_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y112_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y113_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y114_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y115_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y116_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y117_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y118_O;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y119_O;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y120_O;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y121_O;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y122_O;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y123_O;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y124_O;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y125_O;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y126_O;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y127_O;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y128_O;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y129_O;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y130_O;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y131_O;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y132_O;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y133_O;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y134_O;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y135_O;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y136_O;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y137_O;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y138_O;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y139_O;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y140_O;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y141_O;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y142_O;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y143_O;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y144_O;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y145_O;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y146_O;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y147_O;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y148_O;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_D;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_O;
  wire [0:0] RIOI3_SING_X105Y149_OLOGIC_X1Y149_D1;
  wire [0:0] RIOI3_SING_X105Y149_OLOGIC_X1Y149_OQ;
  wire [0:0] RIOI3_SING_X105Y149_OLOGIC_X1Y149_T1;
  wire [0:0] RIOI3_SING_X105Y149_OLOGIC_X1Y149_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_TQ;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_O;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_O;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y118_D1;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y118_OQ;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y118_T1;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y118_TQ;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y121_D1;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y121_OQ;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y121_T1;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y121_TQ;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y122_D1;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y122_OQ;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y122_T1;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y122_TQ;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y123_D1;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y123_OQ;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y123_T1;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y123_TQ;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y124_D1;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y124_OQ;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y124_T1;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y124_TQ;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y125_D1;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y125_OQ;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y125_T1;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y125_TQ;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y126_D1;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y126_OQ;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y126_T1;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y126_TQ;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_D1;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_OQ;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_T1;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_TQ;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y128_D1;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y128_OQ;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y128_T1;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y128_TQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_D1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_OQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_T1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_TQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_D1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_OQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_T1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_TQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_D1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_OQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_T1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_TQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_D1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_OQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_T1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_TQ;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_D1;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_OQ;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_T1;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_TQ;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y136_D1;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y136_OQ;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y136_T1;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y136_TQ;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y139_D1;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y139_OQ;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y139_T1;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y139_TQ;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y140_D1;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y140_OQ;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y140_T1;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y140_TQ;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y141_D1;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y141_OQ;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y141_T1;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y141_TQ;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y142_D1;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y142_OQ;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y142_T1;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y142_TQ;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y145_D1;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y145_OQ;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y145_T1;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y145_TQ;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y146_D1;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y146_OQ;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y146_T1;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y146_TQ;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y147_D1;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y147_OQ;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y147_T1;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y147_TQ;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y148_D1;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y148_OQ;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y148_T1;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y148_TQ;


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y114_SLICE_X50Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y114_SLICE_X50Y114_DO5),
.O6(CLBLL_L_X34Y114_SLICE_X50Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y114_SLICE_X50Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y114_SLICE_X50Y114_CO5),
.O6(CLBLL_L_X34Y114_SLICE_X50Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y114_SLICE_X50Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y114_SLICE_X50Y114_BO5),
.O6(CLBLL_L_X34Y114_SLICE_X50Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y114_SLICE_X50Y114_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y114_SLICE_X50Y114_AO5),
.O6(CLBLL_L_X34Y114_SLICE_X50Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0000ffff0000ff)
  ) CLBLL_L_X34Y114_SLICE_X51Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(LIOB33_X0Y117_IOB_X0Y118_I),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(1'b1),
.O5(CLBLL_L_X34Y114_SLICE_X51Y114_DO5),
.O6(CLBLL_L_X34Y114_SLICE_X51Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaccaaf0fff000)
  ) CLBLL_L_X34Y114_SLICE_X51Y114_CLUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(RIOB33_X105Y113_IOB_X1Y114_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(LIOB33_X0Y117_IOB_X0Y118_I),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLL_L_X34Y114_SLICE_X51Y114_CO5),
.O6(CLBLL_L_X34Y114_SLICE_X51Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00bb00b800b80088)
  ) CLBLL_L_X34Y114_SLICE_X51Y114_BLUT (
.I0(CLBLM_R_X35Y120_SLICE_X53Y120_A_XOR),
.I1(LIOB33_X0Y147_IOB_X0Y147_I),
.I2(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I3(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I4(LIOB33_X0Y145_IOB_X0Y146_I),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLL_L_X34Y114_SLICE_X51Y114_BO5),
.O6(CLBLL_L_X34Y114_SLICE_X51Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaaccfff000f0)
  ) CLBLL_L_X34Y114_SLICE_X51Y114_ALUT (
.I0(RIOB33_X105Y115_IOB_X1Y115_I),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(LIOB33_X0Y117_IOB_X0Y118_I),
.O5(CLBLL_L_X34Y114_SLICE_X51Y114_AO5),
.O6(CLBLL_L_X34Y114_SLICE_X51Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaeefa4450ee5044)
  ) CLBLL_L_X34Y115_SLICE_X50Y115_DLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(RIOB33_X105Y111_IOB_X1Y111_I),
.I3(LIOB33_X0Y117_IOB_X0Y118_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(RIOB33_X105Y117_IOB_X1Y117_I),
.O5(CLBLL_L_X34Y115_SLICE_X50Y115_DO5),
.O6(CLBLL_L_X34Y115_SLICE_X50Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbfef104000000000)
  ) CLBLL_L_X34Y115_SLICE_X50Y115_CLUT (
.I0(LIOB33_X0Y147_IOB_X0Y147_I),
.I1(LIOB33_X0Y117_IOB_X0Y118_I),
.I2(LIOB33_X0Y145_IOB_X0Y146_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(CLBLM_R_X35Y121_SLICE_X53Y121_A_XOR),
.I5(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.O5(CLBLL_L_X34Y115_SLICE_X50Y115_CO5),
.O6(CLBLL_L_X34Y115_SLICE_X50Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccc088c000c088c0)
  ) CLBLL_L_X34Y115_SLICE_X50Y115_BLUT (
.I0(CLBLM_R_X33Y117_SLICE_X48Y117_CO6),
.I1(CLBLL_L_X34Y128_SLICE_X50Y128_AO6),
.I2(CLBLM_R_X35Y121_SLICE_X53Y121_A_XOR),
.I3(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I4(LIOB33_X0Y147_IOB_X0Y147_I),
.I5(CLBLL_L_X34Y116_SLICE_X50Y116_AO5),
.O5(CLBLL_L_X34Y115_SLICE_X50Y115_BO5),
.O6(CLBLL_L_X34Y115_SLICE_X50Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacacacaff0ff000)
  ) CLBLL_L_X34Y115_SLICE_X50Y115_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(LIOB33_X0Y117_IOB_X0Y118_I),
.O5(CLBLL_L_X34Y115_SLICE_X50Y115_AO5),
.O6(CLBLL_L_X34Y115_SLICE_X50Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb0b0f4f472507250)
  ) CLBLL_L_X34Y115_SLICE_X51Y115_DLUT (
.I0(LIOB33_X0Y147_IOB_X0Y147_I),
.I1(LIOB33_X0Y145_IOB_X0Y146_I),
.I2(CLBLM_R_X35Y121_SLICE_X53Y121_A_XOR),
.I3(CLBLM_R_X35Y119_SLICE_X52Y119_A_XOR),
.I4(CLBLL_L_X34Y114_SLICE_X51Y114_DO6),
.I5(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.O5(CLBLL_L_X34Y115_SLICE_X51Y115_DO5),
.O6(CLBLL_L_X34Y115_SLICE_X51Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00000e080e08)
  ) CLBLL_L_X34Y115_SLICE_X51Y115_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I2(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.I3(LIOB33_X0Y117_IOB_X0Y118_I),
.I4(CLBLL_L_X34Y115_SLICE_X51Y115_DO6),
.I5(LIOB33_X0Y147_IOB_X0Y148_I),
.O5(CLBLL_L_X34Y115_SLICE_X51Y115_CO5),
.O6(CLBLL_L_X34Y115_SLICE_X51Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc8c8ccc88888cc88)
  ) CLBLL_L_X34Y115_SLICE_X51Y115_BLUT (
.I0(CLBLL_L_X34Y115_SLICE_X50Y115_CO6),
.I1(LIOB33_X0Y147_IOB_X0Y148_I),
.I2(CLBLL_L_X36Y122_SLICE_X55Y122_AO6),
.I3(CLBLM_R_X35Y121_SLICE_X53Y121_A_XOR),
.I4(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.I5(CLBLM_R_X35Y119_SLICE_X52Y119_A_XOR),
.O5(CLBLL_L_X34Y115_SLICE_X51Y115_BO5),
.O6(CLBLL_L_X34Y115_SLICE_X51Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbffbb33b8fcb830)
  ) CLBLL_L_X34Y115_SLICE_X51Y115_ALUT (
.I0(CLBLM_R_X35Y115_SLICE_X52Y115_AO5),
.I1(LIOB33_X0Y147_IOB_X0Y148_I),
.I2(CLBLL_L_X34Y114_SLICE_X51Y114_BO6),
.I3(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I4(CLBLL_L_X34Y118_SLICE_X51Y118_DO6),
.I5(CLBLL_L_X34Y116_SLICE_X50Y116_BO6),
.O5(CLBLL_L_X34Y115_SLICE_X51Y115_AO5),
.O6(CLBLL_L_X34Y115_SLICE_X51Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0033003300000000)
  ) CLBLL_L_X34Y116_SLICE_X50Y116_DLUT (
.I0(1'b1),
.I1(LIOB33_X0Y145_IOB_X0Y146_I),
.I2(1'b1),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(1'b1),
.I5(CLBLL_L_X34Y117_SLICE_X50Y117_AO6),
.O5(CLBLL_L_X34Y116_SLICE_X50Y116_DO5),
.O6(CLBLL_L_X34Y116_SLICE_X50Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc4c4c4808080c480)
  ) CLBLL_L_X34Y116_SLICE_X50Y116_CLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(CLBLL_L_X34Y116_SLICE_X51Y116_AO5),
.I2(CLBLL_L_X34Y117_SLICE_X50Y117_DO6),
.I3(CLBLL_L_X34Y115_SLICE_X50Y115_AO6),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(CLBLL_L_X34Y114_SLICE_X51Y114_CO6),
.O5(CLBLL_L_X34Y116_SLICE_X50Y116_CO5),
.O6(CLBLL_L_X34Y116_SLICE_X50Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0c080c000)
  ) CLBLL_L_X34Y116_SLICE_X50Y116_BLUT (
.I0(CLBLL_L_X34Y117_SLICE_X50Y117_AO6),
.I1(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I2(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.I3(CLBLL_L_X34Y117_SLICE_X51Y117_AO6),
.I4(CLBLL_L_X34Y116_SLICE_X50Y116_AO6),
.I5(CLBLL_L_X34Y116_SLICE_X50Y116_CO6),
.O5(CLBLL_L_X34Y116_SLICE_X50Y116_BO5),
.O6(CLBLL_L_X34Y116_SLICE_X50Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0c0c0cfef20e02)
  ) CLBLL_L_X34Y116_SLICE_X50Y116_ALUT (
.I0(CLBLL_L_X34Y117_SLICE_X51Y117_CO6),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(LIOB33_X0Y145_IOB_X0Y146_I),
.I3(CLBLL_L_X34Y116_SLICE_X51Y116_DO6),
.I4(CLBLM_R_X35Y121_SLICE_X53Y121_A_XOR),
.I5(1'b1),
.O5(CLBLL_L_X34Y116_SLICE_X50Y116_AO5),
.O6(CLBLL_L_X34Y116_SLICE_X50Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafa0a0cfc0cfc0)
  ) CLBLL_L_X34Y116_SLICE_X51Y116_DLUT (
.I0(CLBLM_R_X35Y116_SLICE_X53Y116_AO6),
.I1(CLBLL_L_X34Y115_SLICE_X50Y115_DO6),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(CLBLL_L_X34Y114_SLICE_X51Y114_AO6),
.I4(CLBLM_R_X35Y117_SLICE_X52Y117_AO6),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLL_L_X34Y116_SLICE_X51Y116_DO5),
.O6(CLBLL_L_X34Y116_SLICE_X51Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h88c0cccc88c00000)
  ) CLBLL_L_X34Y116_SLICE_X51Y116_CLUT (
.I0(CLBLL_L_X34Y116_SLICE_X51Y116_AO6),
.I1(CLBLL_L_X34Y128_SLICE_X50Y128_AO6),
.I2(CLBLM_R_X33Y117_SLICE_X49Y117_CO6),
.I3(LIOB33_X0Y147_IOB_X0Y147_I),
.I4(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I5(CLBLM_R_X35Y121_SLICE_X53Y121_B_XOR),
.O5(CLBLL_L_X34Y116_SLICE_X51Y116_CO5),
.O6(CLBLL_L_X34Y116_SLICE_X51Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd555800000000000)
  ) CLBLL_L_X34Y116_SLICE_X51Y116_BLUT (
.I0(LIOB33_X0Y145_IOB_X0Y146_I),
.I1(CLBLL_L_X36Y116_SLICE_X54Y116_BO5),
.I2(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I3(CLBLL_L_X36Y121_SLICE_X54Y121_AO5),
.I4(CLBLM_R_X33Y117_SLICE_X49Y117_AO6),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLL_L_X34Y116_SLICE_X51Y116_BO5),
.O6(CLBLL_L_X34Y116_SLICE_X51Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hef45ea4005050505)
  ) CLBLL_L_X34Y116_SLICE_X51Y116_ALUT (
.I0(LIOB33_X0Y145_IOB_X0Y146_I),
.I1(CLBLL_L_X34Y118_SLICE_X51Y118_CO6),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(CLBLM_R_X35Y121_SLICE_X53Y121_B_XOR),
.I4(CLBLL_L_X34Y116_SLICE_X51Y116_DO6),
.I5(1'b1),
.O5(CLBLL_L_X34Y116_SLICE_X51Y116_AO5),
.O6(CLBLL_L_X34Y116_SLICE_X51Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f5f5a0a0a0a0)
  ) CLBLL_L_X34Y117_SLICE_X50Y117_DLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(1'b1),
.I2(CLBLL_L_X34Y117_SLICE_X51Y117_BO6),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X33Y117_SLICE_X48Y117_AO6),
.O5(CLBLL_L_X34Y117_SLICE_X50Y117_DO5),
.O6(CLBLL_L_X34Y117_SLICE_X50Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0ddddf5a08888)
  ) CLBLL_L_X34Y117_SLICE_X50Y117_CLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(CLBLM_R_X35Y117_SLICE_X52Y117_AO6),
.I2(CLBLL_L_X34Y115_SLICE_X50Y115_DO6),
.I3(CLBLL_L_X34Y114_SLICE_X51Y114_AO6),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(CLBLL_L_X34Y119_SLICE_X50Y119_BO6),
.O5(CLBLL_L_X34Y117_SLICE_X50Y117_CO5),
.O6(CLBLL_L_X34Y117_SLICE_X50Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4ffaae4e45500)
  ) CLBLL_L_X34Y117_SLICE_X50Y117_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(CLBLL_L_X34Y117_SLICE_X51Y117_BO6),
.I2(CLBLL_L_X34Y119_SLICE_X51Y119_CO6),
.I3(CLBLM_R_X33Y117_SLICE_X48Y117_AO6),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(CLBLL_L_X34Y114_SLICE_X51Y114_CO6),
.O5(CLBLL_L_X34Y117_SLICE_X50Y117_BO5),
.O6(CLBLL_L_X34Y117_SLICE_X50Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddddfa508888fa50)
  ) CLBLL_L_X34Y117_SLICE_X50Y117_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(CLBLM_R_X35Y117_SLICE_X52Y117_AO6),
.I2(CLBLL_L_X34Y119_SLICE_X50Y119_AO6),
.I3(CLBLL_L_X34Y119_SLICE_X50Y119_BO6),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(CLBLL_L_X34Y114_SLICE_X51Y114_AO6),
.O5(CLBLL_L_X34Y117_SLICE_X50Y117_AO5),
.O6(CLBLL_L_X34Y117_SLICE_X50Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3e323e320e020e02)
  ) CLBLL_L_X34Y117_SLICE_X51Y117_DLUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_X0Y117_IOB_X0Y118_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(1'b1),
.I5(RIOB33_X105Y113_IOB_X1Y114_I),
.O5(CLBLL_L_X34Y117_SLICE_X51Y117_DO5),
.O6(CLBLL_L_X34Y117_SLICE_X51Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3bb88c0c0bb88)
  ) CLBLL_L_X34Y117_SLICE_X51Y117_CLUT (
.I0(CLBLL_L_X34Y119_SLICE_X51Y119_CO6),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(CLBLM_R_X33Y118_SLICE_X49Y118_AO6),
.I3(CLBLL_L_X34Y114_SLICE_X51Y114_CO6),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(CLBLL_L_X34Y117_SLICE_X51Y117_BO6),
.O5(CLBLL_L_X34Y117_SLICE_X51Y117_CO5),
.O6(CLBLL_L_X34Y117_SLICE_X51Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf0f0ff00cccc)
  ) CLBLL_L_X34Y117_SLICE_X51Y117_BLUT (
.I0(RIOB33_X105Y115_IOB_X1Y116_I),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(LIOB33_X0Y117_IOB_X0Y118_I),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLL_L_X34Y117_SLICE_X51Y117_BO5),
.O6(CLBLL_L_X34Y117_SLICE_X51Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h888800c088880000)
  ) CLBLL_L_X34Y117_SLICE_X51Y117_ALUT (
.I0(CLBLM_R_X35Y120_SLICE_X53Y120_A_XOR),
.I1(LIOB33_X0Y145_IOB_X0Y146_I),
.I2(CLBLL_L_X36Y116_SLICE_X54Y116_BO5),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y147_IOB_X0Y147_I),
.I5(CLBLL_L_X34Y119_SLICE_X51Y119_AO5),
.O5(CLBLL_L_X34Y117_SLICE_X51Y117_AO5),
.O6(CLBLL_L_X34Y117_SLICE_X51Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaf0ffccaaf000)
  ) CLBLL_L_X34Y118_SLICE_X50Y118_DLUT (
.I0(CLBLM_R_X33Y118_SLICE_X49Y118_AO6),
.I1(CLBLM_R_X35Y118_SLICE_X53Y118_CO6),
.I2(CLBLL_L_X34Y118_SLICE_X51Y118_AO6),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(CLBLL_L_X34Y119_SLICE_X51Y119_CO6),
.O5(CLBLL_L_X34Y118_SLICE_X50Y118_DO5),
.O6(CLBLL_L_X34Y118_SLICE_X50Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaee50eefa445044)
  ) CLBLL_L_X34Y118_SLICE_X50Y118_CLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(CLBLL_L_X34Y114_SLICE_X51Y114_AO6),
.I2(CLBLL_L_X34Y119_SLICE_X50Y119_DO6),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(CLBLM_R_X33Y121_SLICE_X49Y121_CO6),
.I5(CLBLM_R_X35Y117_SLICE_X52Y117_AO6),
.O5(CLBLL_L_X34Y118_SLICE_X50Y118_CO5),
.O6(CLBLL_L_X34Y118_SLICE_X50Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff00aaaacccc)
  ) CLBLL_L_X34Y118_SLICE_X50Y118_BLUT (
.I0(CLBLL_L_X34Y114_SLICE_X51Y114_AO6),
.I1(CLBLL_L_X34Y119_SLICE_X50Y119_BO6),
.I2(CLBLL_L_X34Y119_SLICE_X50Y119_DO6),
.I3(CLBLM_R_X35Y117_SLICE_X52Y117_AO6),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLL_L_X34Y118_SLICE_X50Y118_BO5),
.O6(CLBLL_L_X34Y118_SLICE_X50Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00aaaaf0f0cccc)
  ) CLBLL_L_X34Y118_SLICE_X50Y118_ALUT (
.I0(CLBLM_R_X35Y118_SLICE_X53Y118_CO6),
.I1(CLBLM_R_X33Y118_SLICE_X49Y118_AO6),
.I2(CLBLL_L_X34Y118_SLICE_X51Y118_AO6),
.I3(CLBLM_R_X37Y118_SLICE_X57Y118_AO5),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLL_L_X34Y118_SLICE_X50Y118_AO5),
.O6(CLBLL_L_X34Y118_SLICE_X50Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbfbc8c83b3b0808)
  ) CLBLL_L_X34Y118_SLICE_X51Y118_DLUT (
.I0(CLBLM_R_X35Y118_SLICE_X52Y118_A_XOR),
.I1(LIOB33_X0Y147_IOB_X0Y147_I),
.I2(LIOB33_X0Y145_IOB_X0Y146_I),
.I3(1'b1),
.I4(CLBLM_R_X35Y120_SLICE_X53Y120_A_XOR),
.I5(CLBLL_L_X34Y126_SLICE_X51Y126_D_CY),
.O5(CLBLL_L_X34Y118_SLICE_X51Y118_DO5),
.O6(CLBLL_L_X34Y118_SLICE_X51Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafcfa0cfafc0a0c0)
  ) CLBLL_L_X34Y118_SLICE_X51Y118_CLUT (
.I0(CLBLL_L_X34Y118_SLICE_X51Y118_AO6),
.I1(CLBLL_L_X34Y119_SLICE_X51Y119_CO6),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(CLBLM_R_X33Y118_SLICE_X49Y118_AO6),
.I5(CLBLL_L_X34Y117_SLICE_X51Y117_BO6),
.O5(CLBLL_L_X34Y118_SLICE_X51Y118_CO5),
.O6(CLBLL_L_X34Y118_SLICE_X51Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0cfc0afafa0a0)
  ) CLBLL_L_X34Y118_SLICE_X51Y118_BLUT (
.I0(CLBLM_R_X35Y118_SLICE_X53Y118_CO6),
.I1(CLBLL_L_X36Y115_SLICE_X54Y115_AO6),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(CLBLM_R_X37Y118_SLICE_X57Y118_AO5),
.I4(CLBLL_L_X34Y118_SLICE_X51Y118_AO6),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLL_L_X34Y118_SLICE_X51Y118_BO5),
.O6(CLBLL_L_X34Y118_SLICE_X51Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfd5df858ad0da808)
  ) CLBLL_L_X34Y118_SLICE_X51Y118_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(LIOB33_X0Y117_IOB_X0Y118_I),
.I3(RIOB33_X105Y117_IOB_X1Y117_I),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(RIOB33_X105Y113_IOB_X1Y114_I),
.O5(CLBLL_L_X34Y118_SLICE_X51Y118_AO5),
.O6(CLBLL_L_X34Y118_SLICE_X51Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33003300fcfc3030)
  ) CLBLL_L_X34Y119_SLICE_X50Y119_DLUT (
.I0(1'b1),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(LIOB33_X0Y117_IOB_X0Y118_I),
.O5(CLBLL_L_X34Y119_SLICE_X50Y119_DO5),
.O6(CLBLL_L_X34Y119_SLICE_X50Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000ccaaccaa)
  ) CLBLL_L_X34Y119_SLICE_X50Y119_CLUT (
.I0(CLBLM_R_X35Y117_SLICE_X52Y117_AO6),
.I1(CLBLM_R_X33Y121_SLICE_X49Y121_CO6),
.I2(CLBLL_L_X34Y121_SLICE_X51Y121_DO6),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(CLBLL_L_X34Y119_SLICE_X50Y119_DO6),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLL_L_X34Y119_SLICE_X50Y119_CO5),
.O6(CLBLL_L_X34Y119_SLICE_X50Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50fa50dddd8888)
  ) CLBLL_L_X34Y119_SLICE_X50Y119_BLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(LIOB33_X0Y111_IOB_X0Y111_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(LIOB33_X0Y117_IOB_X0Y118_I),
.O5(CLBLL_L_X34Y119_SLICE_X50Y119_BO5),
.O6(CLBLL_L_X34Y119_SLICE_X50Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa5500d8d8d8d8)
  ) CLBLL_L_X34Y119_SLICE_X50Y119_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(LIOB33_X0Y117_IOB_X0Y118_I),
.O5(CLBLL_L_X34Y119_SLICE_X50Y119_AO5),
.O6(CLBLL_L_X34Y119_SLICE_X50Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he222e222ee222222)
  ) CLBLL_L_X34Y119_SLICE_X51Y119_DLUT (
.I0(CLBLM_R_X35Y118_SLICE_X53Y118_BO6),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(CLBLL_L_X36Y121_SLICE_X54Y121_AO5),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLL_L_X34Y119_SLICE_X51Y119_DO5),
.O6(CLBLL_L_X34Y119_SLICE_X51Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbcb3b0bf8c83808)
  ) CLBLL_L_X34Y119_SLICE_X51Y119_CLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(LIOB33_X0Y117_IOB_X0Y118_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(RIOB33_X105Y117_IOB_X1Y117_I),
.I5(LIOB33_X0Y107_IOB_X0Y108_I),
.O5(CLBLL_L_X34Y119_SLICE_X51Y119_CO5),
.O6(CLBLL_L_X34Y119_SLICE_X51Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cfafafc0c0a0a)
  ) CLBLL_L_X34Y119_SLICE_X51Y119_BLUT (
.I0(CLBLL_L_X34Y121_SLICE_X51Y121_DO6),
.I1(CLBLM_R_X35Y118_SLICE_X53Y118_AO5),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(CLBLM_R_X37Y117_SLICE_X56Y117_AO5),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(CLBLL_L_X36Y121_SLICE_X55Y121_AO6),
.O5(CLBLL_L_X34Y119_SLICE_X51Y119_BO5),
.O6(CLBLL_L_X34Y119_SLICE_X51Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1e0f1e011110000)
  ) CLBLL_L_X34Y119_SLICE_X51Y119_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(LIOB33_X0Y117_IOB_X0Y118_I),
.I2(RIOB33_X105Y117_IOB_X1Y117_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(1'b1),
.O5(CLBLL_L_X34Y119_SLICE_X51Y119_AO5),
.O6(CLBLL_L_X34Y119_SLICE_X51Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffd8d80000d8d8)
  ) CLBLL_L_X34Y120_SLICE_X50Y120_DLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(CLBLL_L_X34Y118_SLICE_X50Y118_DO6),
.I2(CLBLM_R_X35Y117_SLICE_X52Y117_CO6),
.I3(1'b1),
.I4(LIOB33_X0Y145_IOB_X0Y146_I),
.I5(CLBLM_R_X35Y121_SLICE_X53Y121_D_XOR),
.O5(CLBLL_L_X34Y120_SLICE_X50Y120_DO5),
.O6(CLBLL_L_X34Y120_SLICE_X50Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5dda0ddf588a088)
  ) CLBLL_L_X34Y120_SLICE_X50Y120_CLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(CLBLM_R_X33Y121_SLICE_X49Y121_CO6),
.I2(CLBLL_L_X36Y121_SLICE_X55Y121_AO6),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(CLBLL_L_X34Y121_SLICE_X51Y121_DO6),
.I5(CLBLL_L_X34Y119_SLICE_X50Y119_DO6),
.O5(CLBLL_L_X34Y120_SLICE_X50Y120_CO5),
.O6(CLBLL_L_X34Y120_SLICE_X50Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbf8c0000b3800000)
  ) CLBLL_L_X34Y120_SLICE_X50Y120_BLUT (
.I0(CLBLL_L_X34Y120_SLICE_X50Y120_DO6),
.I1(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I2(LIOB33_X0Y147_IOB_X0Y147_I),
.I3(CLBLM_R_X35Y121_SLICE_X53Y121_D_XOR),
.I4(CLBLL_L_X34Y128_SLICE_X50Y128_AO6),
.I5(CLBLM_R_X33Y119_SLICE_X49Y119_CO6),
.O5(CLBLL_L_X34Y120_SLICE_X50Y120_BO5),
.O6(CLBLL_L_X34Y120_SLICE_X50Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff00aaaacccc)
  ) CLBLL_L_X34Y120_SLICE_X50Y120_ALUT (
.I0(CLBLL_L_X34Y121_SLICE_X51Y121_DO6),
.I1(CLBLM_R_X33Y121_SLICE_X49Y121_CO6),
.I2(CLBLM_R_X35Y118_SLICE_X53Y118_AO5),
.I3(CLBLL_L_X36Y121_SLICE_X55Y121_AO6),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLL_L_X34Y120_SLICE_X50Y120_AO5),
.O6(CLBLL_L_X34Y120_SLICE_X50Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5e4e4a0a0e4e4)
  ) CLBLL_L_X34Y120_SLICE_X51Y120_DLUT (
.I0(LIOB33_X0Y145_IOB_X0Y146_I),
.I1(CLBLL_L_X34Y118_SLICE_X51Y118_CO6),
.I2(CLBLM_R_X35Y121_SLICE_X53Y121_C_XOR),
.I3(1'b1),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(CLBLM_R_X35Y117_SLICE_X52Y117_CO6),
.O5(CLBLL_L_X34Y120_SLICE_X51Y120_DO5),
.O6(CLBLL_L_X34Y120_SLICE_X51Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfef000010200000)
  ) CLBLL_L_X34Y120_SLICE_X51Y120_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(LIOB33_X0Y147_IOB_X0Y147_I),
.I2(LIOB33_X0Y145_IOB_X0Y146_I),
.I3(LIOB33_X0Y121_IOB_X0Y121_I),
.I4(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I5(CLBLM_R_X35Y121_SLICE_X53Y121_D_XOR),
.O5(CLBLL_L_X34Y120_SLICE_X51Y120_CO5),
.O6(CLBLL_L_X34Y120_SLICE_X51Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaaa080808)
  ) CLBLL_L_X34Y120_SLICE_X51Y120_BLUT (
.I0(LIOB33_X0Y147_IOB_X0Y148_I),
.I1(CLBLM_R_X35Y121_SLICE_X53Y121_D_XOR),
.I2(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.I3(CLBLM_R_X35Y119_SLICE_X52Y119_D_XOR),
.I4(CLBLL_L_X36Y122_SLICE_X55Y122_AO6),
.I5(CLBLL_L_X34Y120_SLICE_X51Y120_CO6),
.O5(CLBLL_L_X34Y120_SLICE_X51Y120_BO5),
.O6(CLBLL_L_X34Y120_SLICE_X51Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffeffecffccffcc)
  ) CLBLL_L_X34Y120_SLICE_X51Y120_ALUT (
.I0(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I1(CLBLL_L_X34Y120_SLICE_X50Y120_BO6),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(CLBLL_L_X34Y120_SLICE_X51Y120_BO6),
.I4(LIOB33_X0Y121_IOB_X0Y121_I),
.I5(CLBLL_L_X36Y116_SLICE_X55Y116_AO5),
.O5(CLBLL_L_X34Y120_SLICE_X51Y120_AO5),
.O6(CLBLL_L_X34Y120_SLICE_X51Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hefec2320efec2320)
  ) CLBLL_L_X34Y121_SLICE_X50Y121_DLUT (
.I0(CLBLL_L_X34Y118_SLICE_X50Y118_AO6),
.I1(LIOB33_X0Y145_IOB_X0Y146_I),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(CLBLM_R_X35Y117_SLICE_X52Y117_DO6),
.I4(CLBLM_R_X35Y122_SLICE_X53Y122_B_XOR),
.I5(1'b1),
.O5(CLBLL_L_X34Y121_SLICE_X50Y121_DO5),
.O6(CLBLL_L_X34Y121_SLICE_X50Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd8ddd8dd888d888)
  ) CLBLL_L_X34Y121_SLICE_X50Y121_CLUT (
.I0(LIOB33_X0Y145_IOB_X0Y146_I),
.I1(CLBLM_R_X35Y122_SLICE_X53Y122_A_XOR),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(CLBLM_R_X35Y117_SLICE_X52Y117_DO6),
.I4(1'b1),
.I5(CLBLL_L_X34Y118_SLICE_X50Y118_DO6),
.O5(CLBLL_L_X34Y121_SLICE_X50Y121_CO5),
.O6(CLBLL_L_X34Y121_SLICE_X50Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0ddddf5a08888)
  ) CLBLL_L_X34Y121_SLICE_X50Y121_BLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(CLBLM_R_X33Y118_SLICE_X49Y118_BO6),
.I2(CLBLM_R_X33Y121_SLICE_X49Y121_BO6),
.I3(CLBLM_R_X33Y122_SLICE_X49Y122_BO6),
.I4(LIOB33_X0Y145_IOB_X0Y146_I),
.I5(CLBLL_L_X34Y120_SLICE_X50Y120_CO6),
.O5(CLBLL_L_X34Y121_SLICE_X50Y121_BO5),
.O6(CLBLL_L_X34Y121_SLICE_X50Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb080b080f0f00000)
  ) CLBLL_L_X34Y121_SLICE_X50Y121_ALUT (
.I0(CLBLL_L_X34Y121_SLICE_X50Y121_DO6),
.I1(LIOB33_X0Y147_IOB_X0Y147_I),
.I2(CLBLL_L_X34Y128_SLICE_X50Y128_AO6),
.I3(CLBLL_L_X34Y121_SLICE_X50Y121_BO6),
.I4(CLBLM_R_X35Y122_SLICE_X53Y122_B_XOR),
.I5(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.O5(CLBLL_L_X34Y121_SLICE_X50Y121_AO5),
.O6(CLBLL_L_X34Y121_SLICE_X50Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333e2e20000e2e2)
  ) CLBLL_L_X34Y121_SLICE_X51Y121_DLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(LIOB33_X0Y117_IOB_X0Y118_I),
.I2(RIOB33_X105Y115_IOB_X1Y115_I),
.I3(1'b1),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(RIOB33_X105Y107_IOB_X1Y107_I),
.O5(CLBLL_L_X34Y121_SLICE_X51Y121_DO5),
.O6(CLBLL_L_X34Y121_SLICE_X51Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf066f0f000000000)
  ) CLBLL_L_X34Y121_SLICE_X51Y121_CLUT (
.I0(LIOB33_X0Y123_IOB_X0Y123_I),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(CLBLM_R_X35Y122_SLICE_X53Y122_B_XOR),
.I3(LIOB33_X0Y147_IOB_X0Y147_I),
.I4(LIOB33_X0Y145_IOB_X0Y146_I),
.I5(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.O5(CLBLL_L_X34Y121_SLICE_X51Y121_CO5),
.O6(CLBLL_L_X34Y121_SLICE_X51Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000a0ec0000)
  ) CLBLL_L_X34Y121_SLICE_X51Y121_BLUT (
.I0(CLBLL_L_X36Y122_SLICE_X55Y122_AO6),
.I1(CLBLM_R_X35Y122_SLICE_X53Y122_B_XOR),
.I2(CLBLM_R_X35Y120_SLICE_X52Y120_B_XOR),
.I3(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.I4(LIOB33_X0Y147_IOB_X0Y148_I),
.I5(CLBLL_L_X34Y121_SLICE_X51Y121_CO6),
.O5(CLBLL_L_X34Y121_SLICE_X51Y121_BO5),
.O6(CLBLL_L_X34Y121_SLICE_X51Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffefff8fff0fff0)
  ) CLBLL_L_X34Y121_SLICE_X51Y121_ALUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I2(CLBLL_L_X34Y121_SLICE_X50Y121_AO6),
.I3(CLBLL_L_X34Y121_SLICE_X51Y121_BO6),
.I4(LIOB33_X0Y123_IOB_X0Y123_I),
.I5(CLBLL_L_X36Y116_SLICE_X55Y116_AO5),
.O5(CLBLL_L_X34Y121_SLICE_X51Y121_AO5),
.O6(CLBLL_L_X34Y121_SLICE_X51Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00e2e2e2e2)
  ) CLBLL_L_X34Y122_SLICE_X50Y122_DLUT (
.I0(CLBLM_R_X35Y117_SLICE_X52Y117_BO6),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(CLBLL_L_X34Y118_SLICE_X51Y118_BO6),
.I3(CLBLM_R_X35Y122_SLICE_X53Y122_D_XOR),
.I4(1'b1),
.I5(LIOB33_X0Y145_IOB_X0Y146_I),
.O5(CLBLL_L_X34Y122_SLICE_X50Y122_DO5),
.O6(CLBLL_L_X34Y122_SLICE_X50Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccff00aaaaf0f0)
  ) CLBLL_L_X34Y122_SLICE_X50Y122_CLUT (
.I0(CLBLM_R_X35Y117_SLICE_X53Y117_AO6),
.I1(CLBLL_L_X36Y122_SLICE_X54Y122_AO5),
.I2(CLBLL_L_X34Y120_SLICE_X50Y120_AO6),
.I3(CLBLL_L_X36Y123_SLICE_X54Y123_AO6),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(LIOB33_X0Y145_IOB_X0Y146_I),
.O5(CLBLL_L_X34Y122_SLICE_X50Y122_CO5),
.O6(CLBLL_L_X34Y122_SLICE_X50Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8c80ccc08c800c00)
  ) CLBLL_L_X34Y122_SLICE_X50Y122_BLUT (
.I0(CLBLL_L_X34Y122_SLICE_X50Y122_DO6),
.I1(CLBLL_L_X34Y128_SLICE_X50Y128_AO6),
.I2(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I3(CLBLM_R_X35Y122_SLICE_X53Y122_D_XOR),
.I4(LIOB33_X0Y147_IOB_X0Y147_I),
.I5(CLBLL_L_X34Y122_SLICE_X50Y122_CO6),
.O5(CLBLL_L_X34Y122_SLICE_X50Y122_BO5),
.O6(CLBLL_L_X34Y122_SLICE_X50Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee2222f3c0f3c0)
  ) CLBLL_L_X34Y122_SLICE_X50Y122_ALUT (
.I0(CLBLL_L_X36Y122_SLICE_X54Y122_AO5),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(CLBLL_L_X34Y120_SLICE_X50Y120_AO6),
.I3(CLBLM_R_X33Y118_SLICE_X49Y118_BO6),
.I4(CLBLM_R_X33Y122_SLICE_X49Y122_BO6),
.I5(LIOB33_X0Y145_IOB_X0Y146_I),
.O5(CLBLL_L_X34Y122_SLICE_X50Y122_AO5),
.O6(CLBLL_L_X34Y122_SLICE_X50Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33dd11ee22cc00)
  ) CLBLL_L_X34Y122_SLICE_X51Y122_DLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(LIOB33_X0Y145_IOB_X0Y146_I),
.I2(1'b1),
.I3(CLBLM_R_X35Y123_SLICE_X53Y123_A_XOR),
.I4(CLBLL_L_X36Y117_SLICE_X55Y117_CO6),
.I5(CLBLL_L_X34Y118_SLICE_X51Y118_BO6),
.O5(CLBLL_L_X34Y122_SLICE_X51Y122_DO5),
.O6(CLBLL_L_X34Y122_SLICE_X51Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacacacafff00f00)
  ) CLBLL_L_X34Y122_SLICE_X51Y122_CLUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(RIOB33_X105Y115_IOB_X1Y116_I),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(LIOB33_X0Y117_IOB_X0Y118_I),
.O5(CLBLL_L_X34Y122_SLICE_X51Y122_CO5),
.O6(CLBLL_L_X34Y122_SLICE_X51Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffb8ccb833b800b8)
  ) CLBLL_L_X34Y122_SLICE_X51Y122_BLUT (
.I0(CLBLM_R_X33Y123_SLICE_X49Y123_DO6),
.I1(LIOB33_X0Y145_IOB_X0Y146_I),
.I2(CLBLM_R_X35Y117_SLICE_X53Y117_AO6),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(CLBLL_L_X34Y119_SLICE_X51Y119_BO6),
.I5(CLBLL_L_X36Y123_SLICE_X54Y123_AO6),
.O5(CLBLL_L_X34Y122_SLICE_X51Y122_BO5),
.O6(CLBLL_L_X34Y122_SLICE_X51Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb800ff00b8000000)
  ) CLBLL_L_X34Y122_SLICE_X51Y122_ALUT (
.I0(CLBLL_L_X34Y122_SLICE_X51Y122_DO6),
.I1(LIOB33_X0Y147_IOB_X0Y147_I),
.I2(CLBLL_L_X34Y122_SLICE_X51Y122_BO6),
.I3(CLBLL_L_X34Y128_SLICE_X50Y128_AO6),
.I4(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I5(CLBLM_R_X35Y123_SLICE_X53Y123_A_XOR),
.O5(CLBLL_L_X34Y122_SLICE_X51Y122_AO5),
.O6(CLBLL_L_X34Y122_SLICE_X51Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50fa50ee44ee44)
  ) CLBLL_L_X34Y123_SLICE_X50Y123_DLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(CLBLM_R_X33Y125_SLICE_X49Y125_BO6),
.I2(CLBLM_L_X32Y123_SLICE_X47Y123_AO6),
.I3(CLBLL_L_X34Y123_SLICE_X50Y123_CO6),
.I4(1'b1),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLL_L_X34Y123_SLICE_X50Y123_DO5),
.O6(CLBLL_L_X34Y123_SLICE_X50Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000022220000fc30)
  ) CLBLL_L_X34Y123_SLICE_X50Y123_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(LIOB33_X0Y117_IOB_X0Y118_I),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLL_L_X34Y123_SLICE_X50Y123_CO5),
.O6(CLBLL_L_X34Y123_SLICE_X50Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3120312073516240)
  ) CLBLL_L_X34Y123_SLICE_X50Y123_BLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(LIOB33_X0Y117_IOB_X0Y118_I),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(1'b1),
.O5(CLBLL_L_X34Y123_SLICE_X50Y123_BO5),
.O6(CLBLL_L_X34Y123_SLICE_X50Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f500a050ee5044)
  ) CLBLL_L_X34Y123_SLICE_X50Y123_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(RIOB33_X105Y107_IOB_X1Y108_I),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(LIOB33_X0Y117_IOB_X0Y118_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(1'b1),
.O5(CLBLL_L_X34Y123_SLICE_X50Y123_AO5),
.O6(CLBLL_L_X34Y123_SLICE_X50Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_L_X34Y123_SLICE_X51Y123_CARRY4 (
.CI(1'b0),
.CO({CLBLL_L_X34Y123_SLICE_X51Y123_D_CY, CLBLL_L_X34Y123_SLICE_X51Y123_C_CY, CLBLL_L_X34Y123_SLICE_X51Y123_B_CY, CLBLL_L_X34Y123_SLICE_X51Y123_A_CY}),
.CYINIT(1'b0),
.DI({CLBLL_L_X34Y123_SLICE_X51Y123_DO5, CLBLL_L_X34Y123_SLICE_X51Y123_CO5, CLBLL_L_X34Y123_SLICE_X51Y123_BO5, CLBLL_L_X34Y123_SLICE_X51Y123_AO5}),
.O({CLBLL_L_X34Y123_SLICE_X51Y123_D_XOR, CLBLL_L_X34Y123_SLICE_X51Y123_C_XOR, CLBLL_L_X34Y123_SLICE_X51Y123_B_XOR, CLBLL_L_X34Y123_SLICE_X51Y123_A_XOR}),
.S({CLBLL_L_X34Y123_SLICE_X51Y123_DO6, CLBLL_L_X34Y123_SLICE_X51Y123_CO6, CLBLL_L_X34Y123_SLICE_X51Y123_BO6, CLBLL_L_X34Y123_SLICE_X51Y123_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8484212173731010)
  ) CLBLL_L_X34Y123_SLICE_X51Y123_DLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(LIOB33_X0Y119_IOB_X0Y120_I),
.I3(1'b1),
.I4(LIOB33_X0Y121_IOB_X0Y121_I),
.I5(1'b1),
.O5(CLBLL_L_X34Y123_SLICE_X51Y123_DO5),
.O6(CLBLL_L_X34Y123_SLICE_X51Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8822441177551100)
  ) CLBLL_L_X34Y123_SLICE_X51Y123_CLUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(1'b1),
.I3(LIOB33_X0Y117_IOB_X0Y118_I),
.I4(LIOB33_X0Y119_IOB_X0Y119_I),
.I5(1'b1),
.O5(CLBLL_L_X34Y123_SLICE_X51Y123_CO5),
.O6(CLBLL_L_X34Y123_SLICE_X51Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h990000992222bb22)
  ) CLBLL_L_X34Y123_SLICE_X51Y123_BLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(1'b1),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(1'b1),
.O5(CLBLL_L_X34Y123_SLICE_X51Y123_BO5),
.O6(CLBLL_L_X34Y123_SLICE_X51Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha00a500500f0a0fa)
  ) CLBLL_L_X34Y123_SLICE_X51Y123_ALUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(1'b1),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(1'b1),
.O5(CLBLL_L_X34Y123_SLICE_X51Y123_AO5),
.O6(CLBLL_L_X34Y123_SLICE_X51Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff00ccccaaaa)
  ) CLBLL_L_X34Y124_SLICE_X50Y124_DLUT (
.I0(CLBLM_R_X33Y124_SLICE_X49Y124_DO6),
.I1(CLBLL_L_X34Y123_SLICE_X50Y123_AO5),
.I2(CLBLM_R_X33Y124_SLICE_X48Y124_AO5),
.I3(CLBLM_R_X33Y125_SLICE_X49Y125_AO5),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLL_L_X34Y124_SLICE_X50Y124_DO5),
.O6(CLBLL_L_X34Y124_SLICE_X50Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf060f0f000600000)
  ) CLBLL_L_X34Y124_SLICE_X50Y124_CLUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(LIOB33_X0Y125_IOB_X0Y126_I),
.I2(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I3(LIOB33_X0Y147_IOB_X0Y147_I),
.I4(LIOB33_X0Y145_IOB_X0Y146_I),
.I5(CLBLM_R_X35Y123_SLICE_X53Y123_A_XOR),
.O5(CLBLL_L_X34Y124_SLICE_X50Y124_CO5),
.O6(CLBLL_L_X34Y124_SLICE_X50Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa8a0aaaaa8800)
  ) CLBLL_L_X34Y124_SLICE_X50Y124_BLUT (
.I0(LIOB33_X0Y147_IOB_X0Y148_I),
.I1(CLBLL_L_X36Y122_SLICE_X55Y122_AO6),
.I2(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.I3(CLBLM_R_X35Y121_SLICE_X52Y121_A_XOR),
.I4(CLBLL_L_X34Y124_SLICE_X50Y124_CO6),
.I5(CLBLM_R_X35Y123_SLICE_X53Y123_A_XOR),
.O5(CLBLL_L_X34Y124_SLICE_X50Y124_BO5),
.O6(CLBLL_L_X34Y124_SLICE_X50Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffafff8fff8fff0)
  ) CLBLL_L_X34Y124_SLICE_X50Y124_ALUT (
.I0(CLBLL_L_X36Y116_SLICE_X55Y116_AO5),
.I1(LIOB33_X0Y125_IOB_X0Y126_I),
.I2(CLBLL_L_X34Y122_SLICE_X51Y122_AO6),
.I3(CLBLL_L_X34Y124_SLICE_X50Y124_BO6),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.O5(CLBLL_L_X34Y124_SLICE_X50Y124_AO5),
.O6(CLBLL_L_X34Y124_SLICE_X50Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_L_X34Y124_SLICE_X51Y124_CARRY4 (
.CI(CLBLL_L_X34Y123_SLICE_X51Y123_D_CY),
.CO({CLBLL_L_X34Y124_SLICE_X51Y124_D_CY, CLBLL_L_X34Y124_SLICE_X51Y124_C_CY, CLBLL_L_X34Y124_SLICE_X51Y124_B_CY, CLBLL_L_X34Y124_SLICE_X51Y124_A_CY}),
.CYINIT(1'b0),
.DI({CLBLL_L_X34Y124_SLICE_X51Y124_DO5, CLBLL_L_X34Y124_SLICE_X51Y124_CO5, CLBLL_L_X34Y124_SLICE_X51Y124_BO5, CLBLL_L_X34Y124_SLICE_X51Y124_AO5}),
.O({CLBLL_L_X34Y124_SLICE_X51Y124_D_XOR, CLBLL_L_X34Y124_SLICE_X51Y124_C_XOR, CLBLL_L_X34Y124_SLICE_X51Y124_B_XOR, CLBLL_L_X34Y124_SLICE_X51Y124_A_XOR}),
.S({CLBLL_L_X34Y124_SLICE_X51Y124_DO6, CLBLL_L_X34Y124_SLICE_X51Y124_CO6, CLBLL_L_X34Y124_SLICE_X51Y124_BO6, CLBLL_L_X34Y124_SLICE_X51Y124_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8822441100cc88ee)
  ) CLBLL_L_X34Y124_SLICE_X51Y124_DLUT (
.I0(LIOB33_X0Y127_IOB_X0Y128_I),
.I1(LIOB33_X0Y129_IOB_X0Y129_I),
.I2(1'b1),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(1'b1),
.O5(CLBLL_L_X34Y124_SLICE_X51Y124_DO5),
.O6(CLBLL_L_X34Y124_SLICE_X51Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha50000a55050f550)
  ) CLBLL_L_X34Y124_SLICE_X51Y124_CLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(1'b1),
.I2(LIOB33_X0Y127_IOB_X0Y127_I),
.I3(LIOB33_X0Y125_IOB_X0Y126_I),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(1'b1),
.O5(CLBLL_L_X34Y124_SLICE_X51Y124_CO5),
.O6(CLBLL_L_X34Y124_SLICE_X51Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h882244113300bb22)
  ) CLBLL_L_X34Y124_SLICE_X51Y124_BLUT (
.I0(LIOB33_X0Y123_IOB_X0Y124_I),
.I1(LIOB33_X0Y111_IOB_X0Y111_I),
.I2(1'b1),
.I3(LIOB33_X0Y125_IOB_X0Y125_I),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(1'b1),
.O5(CLBLL_L_X34Y124_SLICE_X51Y124_BO5),
.O6(CLBLL_L_X34Y124_SLICE_X51Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha50000a50aff000a)
  ) CLBLL_L_X34Y124_SLICE_X51Y124_ALUT (
.I0(LIOB33_X0Y121_IOB_X0Y122_I),
.I1(1'b1),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(LIOB33_X0Y123_IOB_X0Y123_I),
.I5(1'b1),
.O5(CLBLL_L_X34Y124_SLICE_X51Y124_AO5),
.O6(CLBLL_L_X34Y124_SLICE_X51Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc30fc30bbbb8888)
  ) CLBLL_L_X34Y125_SLICE_X50Y125_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(RIOB33_X105Y113_IOB_X1Y114_I),
.I5(LIOB33_X0Y117_IOB_X0Y118_I),
.O5(CLBLL_L_X34Y125_SLICE_X50Y125_DO5),
.O6(CLBLL_L_X34Y125_SLICE_X50Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafacfc00a0acfc0)
  ) CLBLL_L_X34Y125_SLICE_X50Y125_CLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(RIOB33_X105Y115_IOB_X1Y115_I),
.I4(LIOB33_X0Y117_IOB_X0Y118_I),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLL_L_X34Y125_SLICE_X50Y125_CO5),
.O6(CLBLL_L_X34Y125_SLICE_X50Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfedc7654ba983210)
  ) CLBLL_L_X34Y125_SLICE_X50Y125_BLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(LIOB33_X0Y117_IOB_X0Y118_I),
.I2(RIOB33_X105Y111_IOB_X1Y111_I),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLL_L_X34Y125_SLICE_X50Y125_BO5),
.O6(CLBLL_L_X34Y125_SLICE_X50Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacff0facacf000)
  ) CLBLL_L_X34Y125_SLICE_X50Y125_ALUT (
.I0(CLBLM_R_X33Y125_SLICE_X49Y125_AO5),
.I1(CLBLM_R_X33Y124_SLICE_X49Y124_DO6),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(CLBLL_L_X34Y123_SLICE_X50Y123_AO5),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(CLBLM_R_X33Y125_SLICE_X49Y125_DO6),
.O5(CLBLL_L_X34Y125_SLICE_X50Y125_AO5),
.O6(CLBLL_L_X34Y125_SLICE_X50Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_L_X34Y125_SLICE_X51Y125_CARRY4 (
.CI(CLBLL_L_X34Y124_SLICE_X51Y124_D_CY),
.CO({CLBLL_L_X34Y125_SLICE_X51Y125_D_CY, CLBLL_L_X34Y125_SLICE_X51Y125_C_CY, CLBLL_L_X34Y125_SLICE_X51Y125_B_CY, CLBLL_L_X34Y125_SLICE_X51Y125_A_CY}),
.CYINIT(1'b0),
.DI({CLBLL_L_X34Y125_SLICE_X51Y125_DO5, CLBLL_L_X34Y125_SLICE_X51Y125_CO5, CLBLL_L_X34Y125_SLICE_X51Y125_BO5, CLBLL_L_X34Y125_SLICE_X51Y125_AO5}),
.O({CLBLL_L_X34Y125_SLICE_X51Y125_D_XOR, CLBLL_L_X34Y125_SLICE_X51Y125_C_XOR, CLBLL_L_X34Y125_SLICE_X51Y125_B_XOR, CLBLL_L_X34Y125_SLICE_X51Y125_A_XOR}),
.S({CLBLL_L_X34Y125_SLICE_X51Y125_DO6, CLBLL_L_X34Y125_SLICE_X51Y125_CO6, CLBLL_L_X34Y125_SLICE_X51Y125_BO6, CLBLL_L_X34Y125_SLICE_X51Y125_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h828241412020baba)
  ) CLBLL_L_X34Y125_SLICE_X51Y125_DLUT (
.I0(LIOB33_X0Y137_IOB_X0Y137_I),
.I1(RIOB33_X105Y107_IOB_X1Y108_I),
.I2(LIOB33_X0Y135_IOB_X0Y136_I),
.I3(1'b1),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(1'b1),
.O5(CLBLL_L_X34Y125_SLICE_X51Y125_DO5),
.O6(CLBLL_L_X34Y125_SLICE_X51Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0500a055000f5f0)
  ) CLBLL_L_X34Y125_SLICE_X51Y125_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(1'b1),
.I2(LIOB33_X0Y135_IOB_X0Y135_I),
.I3(LIOB33_X0Y133_IOB_X0Y134_I),
.I4(RIOB33_X105Y107_IOB_X1Y107_I),
.I5(1'b1),
.O5(CLBLL_L_X34Y125_SLICE_X51Y125_CO5),
.O6(CLBLL_L_X34Y125_SLICE_X51Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8844221100aa88ee)
  ) CLBLL_L_X34Y125_SLICE_X51Y125_BLUT (
.I0(LIOB33_X0Y133_IOB_X0Y133_I),
.I1(LIOB33_X0Y131_IOB_X0Y132_I),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(1'b1),
.O5(CLBLL_L_X34Y125_SLICE_X51Y125_BO5),
.O6(CLBLL_L_X34Y125_SLICE_X51Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc00c300333f30030)
  ) CLBLL_L_X34Y125_SLICE_X51Y125_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(LIOB33_X0Y129_IOB_X0Y130_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(LIOB33_X0Y131_IOB_X0Y131_I),
.I5(1'b1),
.O5(CLBLL_L_X34Y125_SLICE_X51Y125_AO5),
.O6(CLBLL_L_X34Y125_SLICE_X51Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haafff0ccaa00f0cc)
  ) CLBLL_L_X34Y126_SLICE_X50Y126_DLUT (
.I0(CLBLM_R_X33Y124_SLICE_X49Y124_DO6),
.I1(CLBLL_L_X34Y122_SLICE_X51Y122_CO6),
.I2(CLBLM_R_X33Y125_SLICE_X49Y125_DO6),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(CLBLL_L_X34Y125_SLICE_X50Y125_DO6),
.O5(CLBLL_L_X34Y126_SLICE_X50Y126_DO5),
.O6(CLBLL_L_X34Y126_SLICE_X50Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccaaaaf0f0ff00)
  ) CLBLL_L_X34Y126_SLICE_X50Y126_CLUT (
.I0(CLBLM_R_X33Y124_SLICE_X49Y124_DO6),
.I1(CLBLL_L_X34Y123_SLICE_X50Y123_AO5),
.I2(CLBLM_R_X33Y125_SLICE_X49Y125_DO6),
.I3(CLBLL_L_X34Y125_SLICE_X50Y125_DO6),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLL_L_X34Y126_SLICE_X50Y126_CO5),
.O6(CLBLL_L_X34Y126_SLICE_X50Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he2ffe233e2cce200)
  ) CLBLL_L_X34Y126_SLICE_X50Y126_BLUT (
.I0(CLBLL_L_X34Y123_SLICE_X50Y123_BO5),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(CLBLM_R_X33Y125_SLICE_X49Y125_BO5),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(CLBLL_L_X34Y125_SLICE_X50Y125_BO6),
.I5(CLBLM_R_X33Y125_SLICE_X49Y125_CO6),
.O5(CLBLL_L_X34Y126_SLICE_X50Y126_BO5),
.O6(CLBLL_L_X34Y126_SLICE_X50Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc30fc30bbbb8888)
  ) CLBLL_L_X34Y126_SLICE_X50Y126_ALUT (
.I0(CLBLL_L_X34Y123_SLICE_X50Y123_BO5),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(CLBLM_R_X33Y125_SLICE_X49Y125_BO5),
.I3(CLBLM_R_X33Y122_SLICE_X48Y122_AO5),
.I4(CLBLL_L_X34Y125_SLICE_X50Y125_BO6),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLL_L_X34Y126_SLICE_X50Y126_AO5),
.O6(CLBLL_L_X34Y126_SLICE_X50Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_L_X34Y126_SLICE_X51Y126_CARRY4 (
.CI(CLBLL_L_X34Y125_SLICE_X51Y125_D_CY),
.CO({CLBLL_L_X34Y126_SLICE_X51Y126_D_CY, CLBLL_L_X34Y126_SLICE_X51Y126_C_CY, CLBLL_L_X34Y126_SLICE_X51Y126_B_CY, CLBLL_L_X34Y126_SLICE_X51Y126_A_CY}),
.CYINIT(1'b0),
.DI({CLBLL_L_X34Y126_SLICE_X51Y126_DO5, CLBLL_L_X34Y126_SLICE_X51Y126_CO5, CLBLL_L_X34Y126_SLICE_X51Y126_BO5, CLBLL_L_X34Y126_SLICE_X51Y126_AO5}),
.O({CLBLL_L_X34Y126_SLICE_X51Y126_D_XOR, CLBLL_L_X34Y126_SLICE_X51Y126_C_XOR, CLBLL_L_X34Y126_SLICE_X51Y126_B_XOR, CLBLL_L_X34Y126_SLICE_X51Y126_A_XOR}),
.S({CLBLL_L_X34Y126_SLICE_X51Y126_DO6, CLBLL_L_X34Y126_SLICE_X51Y126_CO6, CLBLL_L_X34Y126_SLICE_X51Y126_BO6, CLBLL_L_X34Y126_SLICE_X51Y126_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8421842108ce08ce)
  ) CLBLL_L_X34Y126_SLICE_X51Y126_DLUT (
.I0(LIOB33_X0Y143_IOB_X0Y144_I),
.I1(RIOB33_X105Y117_IOB_X1Y117_I),
.I2(RIOB33_X105Y115_IOB_X1Y116_I),
.I3(LIOB33_X0Y145_IOB_X0Y145_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y126_SLICE_X51Y126_DO5),
.O6(CLBLL_L_X34Y126_SLICE_X51Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h990000994444dd44)
  ) CLBLL_L_X34Y126_SLICE_X51Y126_CLUT (
.I0(RIOB33_X105Y115_IOB_X1Y115_I),
.I1(LIOB33_X0Y143_IOB_X0Y143_I),
.I2(1'b1),
.I3(LIOB33_X0Y141_IOB_X0Y142_I),
.I4(RIOB33_X105Y113_IOB_X1Y114_I),
.I5(1'b1),
.O5(CLBLL_L_X34Y126_SLICE_X51Y126_CO5),
.O6(CLBLL_L_X34Y126_SLICE_X51Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h909009094f4f0404)
  ) CLBLL_L_X34Y126_SLICE_X51Y126_BLUT (
.I0(RIOB33_X105Y111_IOB_X1Y112_I),
.I1(LIOB33_X0Y139_IOB_X0Y140_I),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(1'b1),
.I4(LIOB33_X0Y141_IOB_X0Y141_I),
.I5(1'b1),
.O5(CLBLL_L_X34Y126_SLICE_X51Y126_BO5),
.O6(CLBLL_L_X34Y126_SLICE_X51Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h824182410c8e0c8e)
  ) CLBLL_L_X34Y126_SLICE_X51Y126_ALUT (
.I0(LIOB33_X0Y137_IOB_X0Y138_I),
.I1(LIOB33_X0Y139_IOB_X0Y139_I),
.I2(RIOB33_X105Y111_IOB_X1Y111_I),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y126_SLICE_X51Y126_AO5),
.O6(CLBLL_L_X34Y126_SLICE_X51Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00ffaaffaa)
  ) CLBLL_L_X34Y127_SLICE_X50Y127_DLUT (
.I0(LIOB33_X0Y145_IOB_X0Y146_I),
.I1(1'b1),
.I2(1'b1),
.I3(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I4(1'b1),
.I5(LIOB33_X0Y147_IOB_X0Y147_I),
.O5(CLBLL_L_X34Y127_SLICE_X50Y127_DO5),
.O6(CLBLL_L_X34Y127_SLICE_X50Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafcfa0cfafc0a0c0)
  ) CLBLL_L_X34Y127_SLICE_X50Y127_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(LIOB33_X0Y117_IOB_X0Y118_I),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(RIOB33_X105Y117_IOB_X1Y117_I),
.O5(CLBLL_L_X34Y127_SLICE_X50Y127_CO5),
.O6(CLBLL_L_X34Y127_SLICE_X50Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e2ff33e2e2cc00)
  ) CLBLL_L_X34Y127_SLICE_X50Y127_BLUT (
.I0(CLBLL_L_X34Y125_SLICE_X50Y125_CO6),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(CLBLL_L_X34Y125_SLICE_X50Y125_BO6),
.I3(CLBLM_R_X33Y125_SLICE_X49Y125_CO6),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(CLBLL_L_X34Y127_SLICE_X50Y127_CO6),
.O5(CLBLL_L_X34Y127_SLICE_X50Y127_BO5),
.O6(CLBLL_L_X34Y127_SLICE_X50Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb88f3f3bb88c0c0)
  ) CLBLL_L_X34Y127_SLICE_X50Y127_ALUT (
.I0(CLBLL_L_X34Y123_SLICE_X50Y123_BO5),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(CLBLL_L_X34Y125_SLICE_X50Y125_BO6),
.I3(CLBLM_R_X33Y125_SLICE_X49Y125_CO6),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(CLBLL_L_X34Y125_SLICE_X50Y125_CO6),
.O5(CLBLL_L_X34Y127_SLICE_X50Y127_AO5),
.O6(CLBLL_L_X34Y127_SLICE_X50Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y127_SLICE_X51Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y127_SLICE_X51Y127_DO5),
.O6(CLBLL_L_X34Y127_SLICE_X51Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y127_SLICE_X51Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y127_SLICE_X51Y127_CO5),
.O6(CLBLL_L_X34Y127_SLICE_X51Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y127_SLICE_X51Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y127_SLICE_X51Y127_BO5),
.O6(CLBLL_L_X34Y127_SLICE_X51Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y127_SLICE_X51Y127_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y127_SLICE_X51Y127_AO5),
.O6(CLBLL_L_X34Y127_SLICE_X51Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y128_SLICE_X50Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y128_SLICE_X50Y128_DO5),
.O6(CLBLL_L_X34Y128_SLICE_X50Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y128_SLICE_X50Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y128_SLICE_X50Y128_CO5),
.O6(CLBLL_L_X34Y128_SLICE_X50Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y128_SLICE_X50Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y128_SLICE_X50Y128_BO5),
.O6(CLBLL_L_X34Y128_SLICE_X50Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffff0000f0f0)
  ) CLBLL_L_X34Y128_SLICE_X50Y128_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y147_IOB_X0Y147_I),
.I3(1'b1),
.I4(LIOB33_X0Y147_IOB_X0Y148_I),
.I5(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.O5(CLBLL_L_X34Y128_SLICE_X50Y128_AO5),
.O6(CLBLL_L_X34Y128_SLICE_X50Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y128_SLICE_X51Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y128_SLICE_X51Y128_DO5),
.O6(CLBLL_L_X34Y128_SLICE_X51Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y128_SLICE_X51Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y128_SLICE_X51Y128_CO5),
.O6(CLBLL_L_X34Y128_SLICE_X51Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y128_SLICE_X51Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y128_SLICE_X51Y128_BO5),
.O6(CLBLL_L_X34Y128_SLICE_X51Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y128_SLICE_X51Y128_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y128_SLICE_X51Y128_AO5),
.O6(CLBLL_L_X34Y128_SLICE_X51Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y129_SLICE_X50Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y129_SLICE_X50Y129_DO5),
.O6(CLBLL_L_X34Y129_SLICE_X50Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y129_SLICE_X50Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y129_SLICE_X50Y129_CO5),
.O6(CLBLL_L_X34Y129_SLICE_X50Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y129_SLICE_X50Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y129_SLICE_X50Y129_BO5),
.O6(CLBLL_L_X34Y129_SLICE_X50Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff0f0fffff0f0)
  ) CLBLL_L_X34Y129_SLICE_X50Y129_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y147_IOB_X0Y147_I),
.I3(1'b1),
.I4(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I5(1'b1),
.O5(CLBLL_L_X34Y129_SLICE_X50Y129_AO5),
.O6(CLBLL_L_X34Y129_SLICE_X50Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y129_SLICE_X51Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y129_SLICE_X51Y129_DO5),
.O6(CLBLL_L_X34Y129_SLICE_X51Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y129_SLICE_X51Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y129_SLICE_X51Y129_CO5),
.O6(CLBLL_L_X34Y129_SLICE_X51Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y129_SLICE_X51Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y129_SLICE_X51Y129_BO5),
.O6(CLBLL_L_X34Y129_SLICE_X51Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X34Y129_SLICE_X51Y129_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X34Y129_SLICE_X51Y129_AO5),
.O6(CLBLL_L_X34Y129_SLICE_X51Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X36Y115_SLICE_X54Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y115_SLICE_X54Y115_DO5),
.O6(CLBLL_L_X36Y115_SLICE_X54Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000073516240)
  ) CLBLL_L_X36Y115_SLICE_X54Y115_CLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(RIOB33_X105Y115_IOB_X1Y116_I),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(LIOB33_X0Y117_IOB_X0Y118_I),
.O5(CLBLL_L_X36Y115_SLICE_X54Y115_CO5),
.O6(CLBLL_L_X36Y115_SLICE_X54Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000075316420)
  ) CLBLL_L_X36Y115_SLICE_X54Y115_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(RIOB33_X105Y113_IOB_X1Y114_I),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(LIOB33_X0Y117_IOB_X0Y118_I),
.O5(CLBLL_L_X36Y115_SLICE_X54Y115_BO5),
.O6(CLBLL_L_X36Y115_SLICE_X54Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccaa00f000aa)
  ) CLBLL_L_X36Y115_SLICE_X54Y115_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(RIOB33_X105Y117_IOB_X1Y117_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(LIOB33_X0Y117_IOB_X0Y118_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(1'b1),
.O5(CLBLL_L_X36Y115_SLICE_X54Y115_AO5),
.O6(CLBLL_L_X36Y115_SLICE_X54Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X36Y115_SLICE_X55Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y115_SLICE_X55Y115_DO5),
.O6(CLBLL_L_X36Y115_SLICE_X55Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X36Y115_SLICE_X55Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y115_SLICE_X55Y115_CO5),
.O6(CLBLL_L_X36Y115_SLICE_X55Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X36Y115_SLICE_X55Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y115_SLICE_X55Y115_BO5),
.O6(CLBLL_L_X36Y115_SLICE_X55Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X36Y115_SLICE_X55Y115_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y115_SLICE_X55Y115_AO5),
.O6(CLBLL_L_X36Y115_SLICE_X55Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he0e0ff002020ff00)
  ) CLBLL_L_X36Y116_SLICE_X54Y116_DLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(CLBLL_L_X36Y121_SLICE_X54Y121_AO5),
.I3(CLBLL_L_X36Y115_SLICE_X54Y115_CO6),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(RIOB33_X105Y113_IOB_X1Y114_I),
.O5(CLBLL_L_X36Y116_SLICE_X54Y116_DO5),
.O6(CLBLL_L_X36Y116_SLICE_X54Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8d8d8aa55aa55)
  ) CLBLL_L_X36Y116_SLICE_X54Y116_CLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(CLBLL_L_X36Y115_SLICE_X54Y115_CO6),
.I2(CLBLL_L_X36Y115_SLICE_X54Y115_BO6),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y116_SLICE_X54Y116_CO5),
.O6(CLBLL_L_X36Y116_SLICE_X54Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe0ef40405050505)
  ) CLBLL_L_X36Y116_SLICE_X54Y116_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(CLBLL_L_X36Y115_SLICE_X54Y115_AO5),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(CLBLL_L_X36Y115_SLICE_X54Y115_BO6),
.I4(CLBLL_L_X36Y116_SLICE_X54Y116_AO6),
.I5(1'b1),
.O5(CLBLL_L_X36Y116_SLICE_X54Y116_BO5),
.O6(CLBLL_L_X36Y116_SLICE_X54Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h30303300b8b8bb88)
  ) CLBLL_L_X36Y116_SLICE_X54Y116_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y117_I),
.I1(LIOB33_X0Y117_IOB_X0Y118_I),
.I2(RIOB33_X105Y115_IOB_X1Y116_I),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(1'b1),
.O5(CLBLL_L_X36Y116_SLICE_X54Y116_AO5),
.O6(CLBLL_L_X36Y116_SLICE_X54Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X36Y116_SLICE_X55Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y116_SLICE_X55Y116_DO5),
.O6(CLBLL_L_X36Y116_SLICE_X55Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X36Y116_SLICE_X55Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y116_SLICE_X55Y116_CO5),
.O6(CLBLL_L_X36Y116_SLICE_X55Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0cafa00c0cafa0)
  ) CLBLL_L_X36Y116_SLICE_X55Y116_BLUT (
.I0(RIOB33_X105Y107_IOB_X1Y108_I),
.I1(RIOB33_X105Y115_IOB_X1Y116_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(LIOB33_X0Y117_IOB_X0Y118_I),
.I5(1'b1),
.O5(CLBLL_L_X36Y116_SLICE_X55Y116_BO5),
.O6(CLBLL_L_X36Y116_SLICE_X55Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f00000050005)
  ) CLBLL_L_X36Y116_SLICE_X55Y116_ALUT (
.I0(LIOB33_X0Y147_IOB_X0Y148_I),
.I1(1'b1),
.I2(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I3(LIOB33_X0Y147_IOB_X0Y147_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y116_SLICE_X55Y116_AO5),
.O6(CLBLL_L_X36Y116_SLICE_X55Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888b8b822eeaaaa)
  ) CLBLL_L_X36Y117_SLICE_X54Y117_DLUT (
.I0(CLBLM_R_X35Y120_SLICE_X53Y120_B_XOR),
.I1(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I2(CLBLM_R_X35Y118_SLICE_X52Y118_B_XOR),
.I3(CLBLL_L_X36Y116_SLICE_X54Y116_CO5),
.I4(LIOB33_X0Y145_IOB_X0Y146_I),
.I5(LIOB33_X0Y147_IOB_X0Y147_I),
.O5(CLBLL_L_X36Y117_SLICE_X54Y117_DO5),
.O6(CLBLL_L_X36Y117_SLICE_X54Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff540054ff400040)
  ) CLBLL_L_X36Y117_SLICE_X54Y117_CLUT (
.I0(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(CLBLL_L_X36Y117_SLICE_X54Y117_DO6),
.I5(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.O5(CLBLL_L_X36Y117_SLICE_X54Y117_CO5),
.O6(CLBLL_L_X36Y117_SLICE_X54Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa5050ee44ee44)
  ) CLBLL_L_X36Y117_SLICE_X54Y117_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(CLBLM_R_X37Y118_SLICE_X57Y118_AO6),
.I2(CLBLL_L_X36Y117_SLICE_X55Y117_AO6),
.I3(CLBLL_L_X36Y115_SLICE_X54Y115_AO5),
.I4(CLBLL_L_X36Y116_SLICE_X54Y116_AO6),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLL_L_X36Y117_SLICE_X54Y117_BO5),
.O6(CLBLL_L_X36Y117_SLICE_X54Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a0dddd8888)
  ) CLBLL_L_X36Y117_SLICE_X54Y117_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(CLBLM_R_X37Y118_SLICE_X57Y118_AO6),
.I2(CLBLL_L_X36Y117_SLICE_X55Y117_AO6),
.I3(CLBLL_L_X36Y115_SLICE_X54Y115_AO5),
.I4(CLBLL_L_X36Y116_SLICE_X55Y116_BO6),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLL_L_X36Y117_SLICE_X54Y117_AO5),
.O6(CLBLL_L_X36Y117_SLICE_X54Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffe0302fcfe0002)
  ) CLBLL_L_X36Y117_SLICE_X55Y117_DLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_X0Y117_IOB_X0Y118_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(RIOB33_X105Y117_IOB_X1Y117_I),
.I5(RIOB33_X105Y113_IOB_X1Y114_I),
.O5(CLBLL_L_X36Y117_SLICE_X55Y117_DO5),
.O6(CLBLL_L_X36Y117_SLICE_X55Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b8ffccb8b83300)
  ) CLBLL_L_X36Y117_SLICE_X55Y117_CLUT (
.I0(CLBLM_R_X37Y117_SLICE_X56Y117_AO6),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(CLBLL_L_X36Y121_SLICE_X55Y121_AO5),
.I3(CLBLM_R_X35Y117_SLICE_X53Y117_BO6),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(CLBLM_R_X35Y118_SLICE_X53Y118_AO6),
.O5(CLBLL_L_X36Y117_SLICE_X55Y117_CO5),
.O6(CLBLL_L_X36Y117_SLICE_X55Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000acacaaaaacac)
  ) CLBLL_L_X36Y117_SLICE_X55Y117_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y117_I),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(1'b1),
.I4(LIOB33_X0Y117_IOB_X0Y118_I),
.I5(1'b1),
.O5(CLBLL_L_X36Y117_SLICE_X55Y117_BO5),
.O6(CLBLL_L_X36Y117_SLICE_X55Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00fc000caafcaa0c)
  ) CLBLL_L_X36Y117_SLICE_X55Y117_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y117_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(LIOB33_X0Y117_IOB_X0Y118_I),
.I4(RIOB33_X105Y113_IOB_X1Y114_I),
.I5(1'b1),
.O5(CLBLL_L_X36Y117_SLICE_X55Y117_AO5),
.O6(CLBLL_L_X36Y117_SLICE_X55Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaccccff00f0f0)
  ) CLBLL_L_X36Y118_SLICE_X54Y118_DLUT (
.I0(CLBLL_L_X36Y117_SLICE_X55Y117_BO6),
.I1(CLBLL_L_X36Y118_SLICE_X55Y118_AO6),
.I2(CLBLM_R_X35Y118_SLICE_X53Y118_AO5),
.I3(CLBLM_R_X37Y117_SLICE_X56Y117_AO5),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLL_L_X36Y118_SLICE_X54Y118_DO5),
.O6(CLBLL_L_X36Y118_SLICE_X54Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hddf588f5dda088a0)
  ) CLBLL_L_X36Y118_SLICE_X54Y118_CLUT (
.I0(LIOB33_X0Y145_IOB_X0Y146_I),
.I1(CLBLM_L_X32Y123_SLICE_X47Y123_BO6),
.I2(CLBLM_R_X33Y124_SLICE_X49Y124_CO6),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(CLBLL_L_X36Y118_SLICE_X54Y118_DO6),
.I5(CLBLL_L_X36Y117_SLICE_X54Y117_BO6),
.O5(CLBLL_L_X36Y118_SLICE_X54Y118_CO5),
.O6(CLBLL_L_X36Y118_SLICE_X54Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44f5f5a0a0)
  ) CLBLL_L_X36Y118_SLICE_X54Y118_BLUT (
.I0(LIOB33_X0Y145_IOB_X0Y146_I),
.I1(CLBLL_L_X36Y117_SLICE_X54Y117_BO6),
.I2(CLBLM_L_X32Y123_SLICE_X47Y123_BO6),
.I3(CLBLM_R_X33Y124_SLICE_X49Y124_BO6),
.I4(CLBLL_L_X36Y118_SLICE_X54Y118_AO6),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLL_L_X36Y118_SLICE_X54Y118_BO5),
.O6(CLBLL_L_X36Y118_SLICE_X54Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5a0a0dd88dd88)
  ) CLBLL_L_X36Y118_SLICE_X54Y118_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(CLBLM_R_X35Y118_SLICE_X53Y118_AO5),
.I2(CLBLL_L_X36Y118_SLICE_X55Y118_AO6),
.I3(CLBLL_L_X36Y121_SLICE_X55Y121_AO6),
.I4(CLBLM_R_X37Y117_SLICE_X56Y117_AO5),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLL_L_X36Y118_SLICE_X54Y118_AO5),
.O6(CLBLL_L_X36Y118_SLICE_X54Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaff0a0ffaf00a00)
  ) CLBLL_L_X36Y118_SLICE_X55Y118_DLUT (
.I0(CLBLL_L_X34Y119_SLICE_X51Y119_AO6),
.I1(1'b1),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(CLBLL_L_X36Y117_SLICE_X55Y117_DO6),
.I5(CLBLL_L_X36Y116_SLICE_X54Y116_AO5),
.O5(CLBLL_L_X36Y118_SLICE_X55Y118_DO5),
.O6(CLBLL_L_X36Y118_SLICE_X55Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafacafaca0aca0ac)
  ) CLBLL_L_X36Y118_SLICE_X55Y118_CLUT (
.I0(CLBLL_L_X38Y119_SLICE_X58Y119_AO6),
.I1(CLBLM_R_X37Y117_SLICE_X56Y117_AO5),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(1'b1),
.I5(CLBLL_L_X36Y117_SLICE_X55Y117_BO6),
.O5(CLBLL_L_X36Y118_SLICE_X55Y118_CO5),
.O6(CLBLL_L_X36Y118_SLICE_X55Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hef4fe545ea4ae040)
  ) CLBLL_L_X36Y118_SLICE_X55Y118_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(CLBLM_R_X35Y118_SLICE_X53Y118_AO6),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(CLBLL_L_X36Y118_SLICE_X55Y118_AO5),
.I4(CLBLM_R_X37Y117_SLICE_X56Y117_AO6),
.I5(CLBLL_L_X36Y121_SLICE_X55Y121_AO5),
.O5(CLBLL_L_X36Y118_SLICE_X55Y118_BO5),
.O6(CLBLL_L_X36Y118_SLICE_X55Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f000c0cafa0acac)
  ) CLBLL_L_X36Y118_SLICE_X55Y118_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y117_I),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(LIOB33_X0Y117_IOB_X0Y118_I),
.I3(RIOB33_X105Y115_IOB_X1Y115_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(1'b1),
.O5(CLBLL_L_X36Y118_SLICE_X55Y118_AO5),
.O6(CLBLL_L_X36Y118_SLICE_X55Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaffccaaaa00cc)
  ) CLBLL_L_X36Y119_SLICE_X54Y119_DLUT (
.I0(CLBLM_R_X35Y123_SLICE_X53Y123_C_XOR),
.I1(CLBLM_R_X35Y118_SLICE_X53Y118_DO6),
.I2(1'b1),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y145_IOB_X0Y146_I),
.I5(CLBLL_L_X36Y118_SLICE_X55Y118_BO6),
.O5(CLBLL_L_X36Y119_SLICE_X54Y119_DO5),
.O6(CLBLL_L_X36Y119_SLICE_X54Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbcb3b0bf8c83808)
  ) CLBLL_L_X36Y119_SLICE_X54Y119_CLUT (
.I0(CLBLL_L_X36Y116_SLICE_X54Y116_BO6),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(LIOB33_X0Y145_IOB_X0Y146_I),
.I3(CLBLM_L_X32Y123_SLICE_X47Y123_CO6),
.I4(CLBLM_R_X33Y124_SLICE_X49Y124_CO6),
.I5(CLBLL_L_X36Y118_SLICE_X54Y118_DO6),
.O5(CLBLL_L_X36Y119_SLICE_X54Y119_CO5),
.O6(CLBLL_L_X36Y119_SLICE_X54Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccc088c044c000c0)
  ) CLBLL_L_X36Y119_SLICE_X54Y119_BLUT (
.I0(LIOB33_X0Y147_IOB_X0Y147_I),
.I1(CLBLL_L_X34Y128_SLICE_X50Y128_AO6),
.I2(CLBLM_R_X35Y123_SLICE_X53Y123_D_XOR),
.I3(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I4(CLBLL_L_X36Y118_SLICE_X54Y118_BO6),
.I5(CLBLM_R_X37Y119_SLICE_X56Y119_BO6),
.O5(CLBLL_L_X36Y119_SLICE_X54Y119_BO5),
.O6(CLBLL_L_X36Y119_SLICE_X54Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaddfa8850dd5088)
  ) CLBLL_L_X36Y119_SLICE_X54Y119_ALUT (
.I0(LIOB33_X0Y145_IOB_X0Y146_I),
.I1(CLBLM_R_X33Y124_SLICE_X49Y124_BO6),
.I2(CLBLL_L_X36Y118_SLICE_X54Y118_AO6),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(CLBLL_L_X36Y117_SLICE_X54Y117_AO6),
.I5(CLBLL_L_X34Y123_SLICE_X50Y123_DO6),
.O5(CLBLL_L_X36Y119_SLICE_X54Y119_AO5),
.O6(CLBLL_L_X36Y119_SLICE_X54Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfef000010200000)
  ) CLBLL_L_X36Y119_SLICE_X55Y119_DLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(LIOB33_X0Y147_IOB_X0Y147_I),
.I2(LIOB33_X0Y145_IOB_X0Y146_I),
.I3(LIOB33_X0Y119_IOB_X0Y120_I),
.I4(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I5(CLBLM_R_X35Y121_SLICE_X53Y121_C_XOR),
.O5(CLBLL_L_X36Y119_SLICE_X55Y119_DO5),
.O6(CLBLL_L_X36Y119_SLICE_X55Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff008f00ff008800)
  ) CLBLL_L_X36Y119_SLICE_X55Y119_CLUT (
.I0(CLBLL_L_X36Y122_SLICE_X55Y122_AO6),
.I1(CLBLM_R_X35Y119_SLICE_X52Y119_C_XOR),
.I2(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(CLBLL_L_X36Y119_SLICE_X55Y119_DO6),
.I5(CLBLM_R_X35Y121_SLICE_X53Y121_C_XOR),
.O5(CLBLL_L_X36Y119_SLICE_X55Y119_CO5),
.O6(CLBLL_L_X36Y119_SLICE_X55Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffaf8f8f0)
  ) CLBLL_L_X36Y119_SLICE_X55Y119_BLUT (
.I0(CLBLL_L_X36Y116_SLICE_X55Y116_AO5),
.I1(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I2(CLBLM_R_X35Y119_SLICE_X53Y119_DO6),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(LIOB33_X0Y119_IOB_X0Y120_I),
.I5(CLBLL_L_X36Y119_SLICE_X55Y119_CO6),
.O5(CLBLL_L_X36Y119_SLICE_X55Y119_BO5),
.O6(CLBLL_L_X36Y119_SLICE_X55Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc884400c480c480)
  ) CLBLL_L_X36Y119_SLICE_X55Y119_ALUT (
.I0(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I1(CLBLL_L_X34Y128_SLICE_X50Y128_AO6),
.I2(CLBLL_L_X36Y119_SLICE_X54Y119_AO6),
.I3(CLBLM_R_X35Y123_SLICE_X53Y123_C_XOR),
.I4(CLBLL_L_X36Y119_SLICE_X54Y119_DO6),
.I5(LIOB33_X0Y147_IOB_X0Y147_I),
.O5(CLBLL_L_X36Y119_SLICE_X55Y119_AO5),
.O6(CLBLL_L_X36Y119_SLICE_X55Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaff0faaaaf000)
  ) CLBLL_L_X36Y120_SLICE_X54Y120_DLUT (
.I0(CLBLM_R_X35Y123_SLICE_X53Y123_B_XOR),
.I1(1'b1),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(CLBLM_R_X35Y118_SLICE_X53Y118_DO6),
.I4(LIOB33_X0Y145_IOB_X0Y146_I),
.I5(CLBLL_L_X36Y117_SLICE_X55Y117_CO6),
.O5(CLBLL_L_X36Y120_SLICE_X54Y120_DO5),
.O6(CLBLL_L_X36Y120_SLICE_X54Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00aaaaf0f0cccc)
  ) CLBLL_L_X36Y120_SLICE_X54Y120_CLUT (
.I0(CLBLL_L_X36Y118_SLICE_X55Y118_CO6),
.I1(CLBLL_L_X36Y116_SLICE_X54Y116_BO6),
.I2(CLBLM_R_X33Y123_SLICE_X48Y123_BO6),
.I3(CLBLM_L_X32Y123_SLICE_X47Y123_CO6),
.I4(LIOB33_X0Y145_IOB_X0Y146_I),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLL_L_X36Y120_SLICE_X54Y120_CO5),
.O6(CLBLL_L_X36Y120_SLICE_X54Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdec7564b9a83120)
  ) CLBLL_L_X36Y120_SLICE_X54Y120_BLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(LIOB33_X0Y145_IOB_X0Y146_I),
.I2(CLBLL_L_X36Y117_SLICE_X54Y117_AO6),
.I3(CLBLL_L_X34Y119_SLICE_X51Y119_BO6),
.I4(CLBLM_R_X33Y123_SLICE_X49Y123_DO6),
.I5(CLBLL_L_X34Y123_SLICE_X50Y123_DO6),
.O5(CLBLL_L_X36Y120_SLICE_X54Y120_BO5),
.O6(CLBLL_L_X36Y120_SLICE_X54Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b80000fc300000)
  ) CLBLL_L_X36Y120_SLICE_X54Y120_ALUT (
.I0(CLBLL_L_X36Y120_SLICE_X54Y120_DO6),
.I1(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I2(CLBLM_R_X35Y123_SLICE_X53Y123_B_XOR),
.I3(CLBLL_L_X36Y120_SLICE_X54Y120_BO6),
.I4(CLBLL_L_X34Y128_SLICE_X50Y128_AO6),
.I5(LIOB33_X0Y147_IOB_X0Y147_I),
.O5(CLBLL_L_X36Y120_SLICE_X54Y120_AO5),
.O6(CLBLL_L_X36Y120_SLICE_X54Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccfa50fa50)
  ) CLBLL_L_X36Y120_SLICE_X55Y120_DLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(CLBLM_R_X35Y125_SLICE_X53Y125_A_XOR),
.I2(CLBLM_R_X37Y118_SLICE_X57Y118_DO6),
.I3(CLBLM_R_X37Y119_SLICE_X56Y119_DO6),
.I4(1'b1),
.I5(LIOB33_X0Y145_IOB_X0Y146_I),
.O5(CLBLL_L_X36Y120_SLICE_X55Y120_DO5),
.O6(CLBLL_L_X36Y120_SLICE_X55Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeaef4a45e0e5404)
  ) CLBLL_L_X36Y120_SLICE_X55Y120_CLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(CLBLL_L_X36Y116_SLICE_X54Y116_CO6),
.I2(LIOB33_X0Y145_IOB_X0Y146_I),
.I3(CLBLM_R_X33Y123_SLICE_X48Y123_CO6),
.I4(CLBLM_R_X37Y119_SLICE_X57Y119_DO6),
.I5(CLBLM_L_X32Y123_SLICE_X47Y123_DO6),
.O5(CLBLL_L_X36Y120_SLICE_X55Y120_CO5),
.O6(CLBLL_L_X36Y120_SLICE_X55Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0f0c0c0a000c0c0)
  ) CLBLL_L_X36Y120_SLICE_X55Y120_BLUT (
.I0(CLBLL_L_X36Y120_SLICE_X55Y120_DO6),
.I1(CLBLM_R_X35Y125_SLICE_X53Y125_A_XOR),
.I2(CLBLL_L_X34Y128_SLICE_X50Y128_AO6),
.I3(LIOB33_X0Y147_IOB_X0Y147_I),
.I4(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I5(CLBLL_L_X36Y120_SLICE_X55Y120_CO6),
.O5(CLBLL_L_X36Y120_SLICE_X55Y120_BO5),
.O6(CLBLL_L_X36Y120_SLICE_X55Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccf0ffaaccf000)
  ) CLBLL_L_X36Y120_SLICE_X55Y120_ALUT (
.I0(CLBLM_R_X33Y123_SLICE_X48Y123_BO6),
.I1(CLBLM_L_X32Y123_SLICE_X47Y123_DO6),
.I2(CLBLL_L_X36Y116_SLICE_X54Y116_CO6),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y145_IOB_X0Y146_I),
.I5(CLBLL_L_X36Y118_SLICE_X55Y118_CO6),
.O5(CLBLL_L_X36Y120_SLICE_X55Y120_AO5),
.O6(CLBLL_L_X36Y120_SLICE_X55Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he222e222ee222222)
  ) CLBLL_L_X36Y121_SLICE_X54Y121_DLUT (
.I0(CLBLL_L_X36Y121_SLICE_X54Y121_AO6),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(RIOB33_X105Y115_IOB_X1Y116_I),
.I3(CLBLL_L_X36Y121_SLICE_X54Y121_AO5),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLL_L_X36Y121_SLICE_X54Y121_DO5),
.O6(CLBLL_L_X36Y121_SLICE_X54Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa2a8a00002080)
  ) CLBLL_L_X36Y121_SLICE_X54Y121_CLUT (
.I0(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I1(LIOB33_X0Y125_IOB_X0Y125_I),
.I2(LIOB33_X0Y145_IOB_X0Y146_I),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(LIOB33_X0Y147_IOB_X0Y147_I),
.I5(CLBLM_R_X35Y122_SLICE_X53Y122_D_XOR),
.O5(CLBLL_L_X36Y121_SLICE_X54Y121_CO5),
.O6(CLBLL_L_X36Y121_SLICE_X54Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0d0c05000)
  ) CLBLL_L_X36Y121_SLICE_X54Y121_BLUT (
.I0(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.I1(CLBLM_R_X35Y120_SLICE_X52Y120_D_XOR),
.I2(LIOB33_X0Y147_IOB_X0Y148_I),
.I3(CLBLM_R_X35Y122_SLICE_X53Y122_D_XOR),
.I4(CLBLL_L_X36Y122_SLICE_X55Y122_AO6),
.I5(CLBLL_L_X36Y121_SLICE_X54Y121_CO6),
.O5(CLBLL_L_X36Y121_SLICE_X54Y121_BO5),
.O6(CLBLL_L_X36Y121_SLICE_X54Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000541000005555)
  ) CLBLL_L_X36Y121_SLICE_X54Y121_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(RIOB33_X105Y113_IOB_X1Y114_I),
.I4(LIOB33_X0Y117_IOB_X0Y118_I),
.I5(1'b1),
.O5(CLBLL_L_X36Y121_SLICE_X54Y121_AO5),
.O6(CLBLL_L_X36Y121_SLICE_X54Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a030a0c0a0)
  ) CLBLL_L_X36Y121_SLICE_X55Y121_DLUT (
.I0(CLBLM_R_X35Y123_SLICE_X53Y123_C_XOR),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I3(LIOB33_X0Y145_IOB_X0Y146_I),
.I4(LIOB33_X0Y127_IOB_X0Y128_I),
.I5(LIOB33_X0Y147_IOB_X0Y147_I),
.O5(CLBLL_L_X36Y121_SLICE_X55Y121_DO5),
.O6(CLBLL_L_X36Y121_SLICE_X55Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ce00ff000a00)
  ) CLBLL_L_X36Y121_SLICE_X55Y121_CLUT (
.I0(CLBLM_R_X35Y123_SLICE_X53Y123_C_XOR),
.I1(CLBLL_L_X36Y122_SLICE_X55Y122_AO6),
.I2(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(CLBLL_L_X36Y121_SLICE_X55Y121_DO6),
.I5(CLBLM_R_X35Y121_SLICE_X52Y121_C_XOR),
.O5(CLBLL_L_X36Y121_SLICE_X55Y121_CO5),
.O6(CLBLL_L_X36Y121_SLICE_X55Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffef0f8f0)
  ) CLBLL_L_X36Y121_SLICE_X55Y121_BLUT (
.I0(LIOB33_X0Y127_IOB_X0Y128_I),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(CLBLL_L_X36Y119_SLICE_X55Y119_AO6),
.I3(CLBLL_L_X36Y116_SLICE_X55Y116_AO5),
.I4(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I5(CLBLL_L_X36Y121_SLICE_X55Y121_CO6),
.O5(CLBLL_L_X36Y121_SLICE_X55Y121_BO5),
.O6(CLBLL_L_X36Y121_SLICE_X55Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4444f5a0ccccf5a0)
  ) CLBLL_L_X36Y121_SLICE_X55Y121_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(RIOB33_X105Y117_IOB_X1Y117_I),
.I2(RIOB33_X105Y109_IOB_X1Y109_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(LIOB33_X0Y117_IOB_X0Y118_I),
.I5(1'b1),
.O5(CLBLL_L_X36Y121_SLICE_X55Y121_AO5),
.O6(CLBLL_L_X36Y121_SLICE_X55Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00003aca0000)
  ) CLBLL_L_X36Y122_SLICE_X54Y122_DLUT (
.I0(CLBLM_R_X35Y123_SLICE_X53Y123_D_XOR),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(LIOB33_X0Y145_IOB_X0Y146_I),
.I3(LIOB33_X0Y129_IOB_X0Y129_I),
.I4(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I5(LIOB33_X0Y147_IOB_X0Y147_I),
.O5(CLBLL_L_X36Y122_SLICE_X54Y122_DO5),
.O6(CLBLL_L_X36Y122_SLICE_X54Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffc0ea00000000)
  ) CLBLL_L_X36Y122_SLICE_X54Y122_CLUT (
.I0(CLBLM_R_X35Y123_SLICE_X53Y123_D_XOR),
.I1(CLBLM_R_X35Y121_SLICE_X52Y121_D_XOR),
.I2(CLBLL_L_X36Y122_SLICE_X55Y122_AO6),
.I3(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.I4(CLBLL_L_X36Y122_SLICE_X54Y122_DO6),
.I5(LIOB33_X0Y147_IOB_X0Y148_I),
.O5(CLBLL_L_X36Y122_SLICE_X54Y122_CO5),
.O6(CLBLL_L_X36Y122_SLICE_X54Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffeeecffffeccc)
  ) CLBLL_L_X36Y122_SLICE_X54Y122_BLUT (
.I0(CLBLL_L_X36Y116_SLICE_X55Y116_AO5),
.I1(CLBLL_L_X34Y122_SLICE_X50Y122_BO6),
.I2(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I3(LIOB33_X0Y125_IOB_X0Y125_I),
.I4(CLBLL_L_X36Y121_SLICE_X54Y121_BO6),
.I5(LIOB33_X0Y111_IOB_X0Y111_I),
.O5(CLBLL_L_X36Y122_SLICE_X54Y122_BO5),
.O6(CLBLL_L_X36Y122_SLICE_X54Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c0afa0afa0)
  ) CLBLL_L_X36Y122_SLICE_X54Y122_ALUT (
.I0(CLBLM_R_X33Y122_SLICE_X49Y122_CO6),
.I1(CLBLM_R_X37Y123_SLICE_X56Y123_CO6),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(CLBLM_L_X32Y123_SLICE_X46Y123_AO6),
.I4(CLBLM_R_X37Y119_SLICE_X57Y119_BO6),
.I5(1'b1),
.O5(CLBLL_L_X36Y122_SLICE_X54Y122_AO5),
.O6(CLBLL_L_X36Y122_SLICE_X54Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00002a8a2080)
  ) CLBLL_L_X36Y122_SLICE_X55Y122_DLUT (
.I0(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I1(LIOB33_X0Y131_IOB_X0Y132_I),
.I2(LIOB33_X0Y145_IOB_X0Y146_I),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(CLBLM_R_X35Y124_SLICE_X53Y124_C_XOR),
.I5(LIOB33_X0Y147_IOB_X0Y147_I),
.O5(CLBLL_L_X36Y122_SLICE_X55Y122_DO5),
.O6(CLBLL_L_X36Y122_SLICE_X55Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff88f800000000)
  ) CLBLL_L_X36Y122_SLICE_X55Y122_CLUT (
.I0(CLBLL_L_X36Y122_SLICE_X55Y122_AO6),
.I1(CLBLM_R_X35Y122_SLICE_X52Y122_C_XOR),
.I2(CLBLM_R_X35Y124_SLICE_X53Y124_C_XOR),
.I3(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.I4(CLBLL_L_X36Y122_SLICE_X55Y122_DO6),
.I5(LIOB33_X0Y147_IOB_X0Y148_I),
.O5(CLBLL_L_X36Y122_SLICE_X55Y122_CO5),
.O6(CLBLL_L_X36Y122_SLICE_X55Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeeffecffecffcc)
  ) CLBLL_L_X36Y122_SLICE_X55Y122_BLUT (
.I0(CLBLL_L_X36Y116_SLICE_X55Y116_AO5),
.I1(CLBLL_L_X36Y119_SLICE_X54Y119_BO6),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(CLBLL_L_X36Y122_SLICE_X54Y122_CO6),
.I4(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I5(LIOB33_X0Y129_IOB_X0Y129_I),
.O5(CLBLL_L_X36Y122_SLICE_X55Y122_BO5),
.O6(CLBLL_L_X36Y122_SLICE_X55Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000550000ff00aa)
  ) CLBLL_L_X36Y122_SLICE_X55Y122_ALUT (
.I0(LIOB33_X0Y145_IOB_X0Y146_I),
.I1(1'b1),
.I2(1'b1),
.I3(LIOB33_X0Y147_IOB_X0Y147_I),
.I4(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I5(1'b1),
.O5(CLBLL_L_X36Y122_SLICE_X55Y122_AO5),
.O6(CLBLL_L_X36Y122_SLICE_X55Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfd5df858ad0da808)
  ) CLBLL_L_X36Y123_SLICE_X54Y123_DLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(CLBLL_L_X36Y121_SLICE_X54Y121_DO6),
.I2(LIOB33_X0Y145_IOB_X0Y146_I),
.I3(CLBLM_R_X33Y123_SLICE_X48Y123_DO6),
.I4(CLBLM_R_X37Y119_SLICE_X57Y119_AO6),
.I5(CLBLM_R_X33Y124_SLICE_X48Y124_BO6),
.O5(CLBLL_L_X36Y123_SLICE_X54Y123_DO5),
.O6(CLBLL_L_X36Y123_SLICE_X54Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a02288a0a0)
  ) CLBLL_L_X36Y123_SLICE_X54Y123_CLUT (
.I0(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(CLBLM_R_X35Y125_SLICE_X53Y125_B_XOR),
.I3(LIOB33_X0Y135_IOB_X0Y135_I),
.I4(LIOB33_X0Y145_IOB_X0Y146_I),
.I5(LIOB33_X0Y147_IOB_X0Y147_I),
.O5(CLBLL_L_X36Y123_SLICE_X54Y123_CO5),
.O6(CLBLL_L_X36Y123_SLICE_X54Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0f0202020)
  ) CLBLL_L_X36Y123_SLICE_X54Y123_BLUT (
.I0(CLBLM_R_X35Y125_SLICE_X53Y125_B_XOR),
.I1(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.I2(LIOB33_X0Y147_IOB_X0Y148_I),
.I3(CLBLM_R_X35Y123_SLICE_X52Y123_B_XOR),
.I4(CLBLL_L_X36Y122_SLICE_X55Y122_AO6),
.I5(CLBLL_L_X36Y123_SLICE_X54Y123_CO6),
.O5(CLBLL_L_X36Y123_SLICE_X54Y123_BO5),
.O6(CLBLL_L_X36Y123_SLICE_X54Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ccccf0f0aaaa)
  ) CLBLL_L_X36Y123_SLICE_X54Y123_ALUT (
.I0(CLBLL_L_X36Y117_SLICE_X55Y117_DO6),
.I1(CLBLL_L_X34Y123_SLICE_X50Y123_CO6),
.I2(CLBLM_R_X37Y123_SLICE_X56Y123_DO6),
.I3(CLBLM_R_X33Y123_SLICE_X48Y123_AO6),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(1'b1),
.O5(CLBLL_L_X36Y123_SLICE_X54Y123_AO5),
.O6(CLBLL_L_X36Y123_SLICE_X54Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff000f0ffcc00cc)
  ) CLBLL_L_X36Y123_SLICE_X55Y123_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X37Y119_SLICE_X56Y119_DO6),
.I2(CLBLL_L_X36Y118_SLICE_X55Y118_DO6),
.I3(LIOB33_X0Y145_IOB_X0Y146_I),
.I4(CLBLM_R_X35Y125_SLICE_X53Y125_B_XOR),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLL_L_X36Y123_SLICE_X55Y123_DO5),
.O6(CLBLL_L_X36Y123_SLICE_X55Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaccffcc00)
  ) CLBLL_L_X36Y123_SLICE_X55Y123_CLUT (
.I0(CLBLM_R_X37Y119_SLICE_X57Y119_AO6),
.I1(CLBLM_R_X33Y123_SLICE_X48Y123_DO6),
.I2(CLBLM_R_X33Y122_SLICE_X48Y122_BO6),
.I3(LIOB33_X0Y145_IOB_X0Y146_I),
.I4(CLBLL_L_X36Y116_SLICE_X54Y116_DO6),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLL_L_X36Y123_SLICE_X55Y123_CO5),
.O6(CLBLL_L_X36Y123_SLICE_X55Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ff000acacacac)
  ) CLBLL_L_X36Y123_SLICE_X55Y123_BLUT (
.I0(CLBLL_L_X36Y116_SLICE_X54Y116_DO6),
.I1(CLBLM_R_X37Y119_SLICE_X57Y119_DO6),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(CLBLM_R_X33Y123_SLICE_X48Y123_CO6),
.I4(CLBLM_R_X33Y122_SLICE_X48Y122_BO6),
.I5(LIOB33_X0Y145_IOB_X0Y146_I),
.O5(CLBLL_L_X36Y123_SLICE_X55Y123_BO5),
.O6(CLBLL_L_X36Y123_SLICE_X55Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888cc00c0c0c0c0)
  ) CLBLL_L_X36Y123_SLICE_X55Y123_ALUT (
.I0(CLBLL_L_X36Y123_SLICE_X55Y123_DO6),
.I1(CLBLL_L_X34Y128_SLICE_X50Y128_AO6),
.I2(CLBLM_R_X35Y125_SLICE_X53Y125_B_XOR),
.I3(CLBLL_L_X36Y123_SLICE_X55Y123_BO6),
.I4(LIOB33_X0Y147_IOB_X0Y147_I),
.I5(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.O5(CLBLL_L_X36Y123_SLICE_X55Y123_AO5),
.O6(CLBLL_L_X36Y123_SLICE_X55Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffa0a0000fa0a)
  ) CLBLL_L_X36Y124_SLICE_X54Y124_DLUT (
.I0(CLBLL_L_X36Y122_SLICE_X54Y122_AO6),
.I1(1'b1),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(CLBLL_L_X36Y123_SLICE_X54Y123_AO5),
.I4(LIOB33_X0Y145_IOB_X0Y146_I),
.I5(CLBLM_R_X35Y125_SLICE_X53Y125_D_XOR),
.O5(CLBLL_L_X36Y124_SLICE_X54Y124_DO5),
.O6(CLBLL_L_X36Y124_SLICE_X54Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4c0c480844044000)
  ) CLBLL_L_X36Y124_SLICE_X54Y124_CLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(CLBLL_L_X36Y121_SLICE_X54Y121_AO5),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(RIOB33_X105Y115_IOB_X1Y116_I),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(RIOB33_X105Y113_IOB_X1Y114_I),
.O5(CLBLL_L_X36Y124_SLICE_X54Y124_CO5),
.O6(CLBLL_L_X36Y124_SLICE_X54Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffe455e4aae400e4)
  ) CLBLL_L_X36Y124_SLICE_X54Y124_BLUT (
.I0(LIOB33_X0Y145_IOB_X0Y146_I),
.I1(CLBLL_L_X38Y121_SLICE_X58Y121_AO6),
.I2(CLBLL_L_X34Y126_SLICE_X50Y126_AO6),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(CLBLL_L_X34Y124_SLICE_X50Y124_DO6),
.I5(CLBLL_L_X36Y124_SLICE_X54Y124_CO6),
.O5(CLBLL_L_X36Y124_SLICE_X54Y124_BO5),
.O6(CLBLL_L_X36Y124_SLICE_X54Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeef5a04444f5a0)
  ) CLBLL_L_X36Y124_SLICE_X54Y124_ALUT (
.I0(LIOB33_X0Y145_IOB_X0Y146_I),
.I1(CLBLL_L_X38Y121_SLICE_X58Y121_AO6),
.I2(CLBLL_L_X34Y124_SLICE_X50Y124_DO6),
.I3(CLBLL_L_X36Y121_SLICE_X54Y121_DO6),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(CLBLM_R_X33Y124_SLICE_X48Y124_BO6),
.O5(CLBLL_L_X36Y124_SLICE_X54Y124_AO5),
.O6(CLBLL_L_X36Y124_SLICE_X54Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccdcdccccc8c8)
  ) CLBLL_L_X36Y124_SLICE_X55Y124_DLUT (
.I0(LIOB33_X0Y117_IOB_X0Y118_I),
.I1(RIOB33_X105Y117_IOB_X1Y117_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(1'b1),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(RIOB33_X105Y115_IOB_X1Y115_I),
.O5(CLBLL_L_X36Y124_SLICE_X55Y124_DO5),
.O6(CLBLL_L_X36Y124_SLICE_X55Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff00f00fcfc0c0c)
  ) CLBLL_L_X36Y124_SLICE_X55Y124_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X36Y118_SLICE_X55Y118_DO6),
.I2(LIOB33_X0Y145_IOB_X0Y146_I),
.I3(CLBLL_L_X36Y122_SLICE_X54Y122_AO6),
.I4(CLBLM_R_X35Y125_SLICE_X53Y125_C_XOR),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLL_L_X36Y124_SLICE_X55Y124_CO5),
.O6(CLBLL_L_X36Y124_SLICE_X55Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0acf0ac000000000)
  ) CLBLL_L_X36Y124_SLICE_X55Y124_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y117_I),
.I1(RIOB33_X105Y115_IOB_X1Y115_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(CLBLL_L_X36Y121_SLICE_X54Y121_AO5),
.O5(CLBLL_L_X36Y124_SLICE_X55Y124_BO5),
.O6(CLBLL_L_X36Y124_SLICE_X55Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0c03000a0a0a0a0)
  ) CLBLL_L_X36Y124_SLICE_X55Y124_ALUT (
.I0(CLBLM_R_X35Y125_SLICE_X53Y125_C_XOR),
.I1(LIOB33_X0Y147_IOB_X0Y147_I),
.I2(CLBLL_L_X34Y128_SLICE_X50Y128_AO6),
.I3(CLBLL_L_X36Y123_SLICE_X55Y123_CO6),
.I4(CLBLL_L_X36Y124_SLICE_X55Y124_CO6),
.I5(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.O5(CLBLL_L_X36Y124_SLICE_X55Y124_AO5),
.O6(CLBLL_L_X36Y124_SLICE_X55Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf5ccf5cca0cca0)
  ) CLBLL_L_X36Y125_SLICE_X54Y125_DLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(CLBLM_R_X35Y126_SLICE_X53Y126_A_XOR),
.I2(CLBLL_L_X36Y125_SLICE_X55Y125_AO6),
.I3(LIOB33_X0Y145_IOB_X0Y146_I),
.I4(1'b1),
.I5(CLBLL_L_X36Y123_SLICE_X54Y123_AO5),
.O5(CLBLL_L_X36Y125_SLICE_X54Y125_DO5),
.O6(CLBLL_L_X36Y125_SLICE_X54Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0aacc00f0aacc)
  ) CLBLL_L_X36Y125_SLICE_X54Y125_CLUT (
.I0(CLBLL_L_X34Y125_SLICE_X50Y125_AO6),
.I1(CLBLL_L_X36Y124_SLICE_X54Y124_CO6),
.I2(CLBLL_L_X36Y124_SLICE_X55Y124_BO6),
.I3(LIOB33_X0Y145_IOB_X0Y146_I),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(CLBLL_L_X34Y126_SLICE_X50Y126_AO6),
.O5(CLBLL_L_X36Y125_SLICE_X54Y125_CO5),
.O6(CLBLL_L_X36Y125_SLICE_X54Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb00f3008800c000)
  ) CLBLL_L_X36Y125_SLICE_X54Y125_BLUT (
.I0(CLBLL_L_X36Y125_SLICE_X54Y125_DO6),
.I1(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I2(CLBLL_L_X36Y124_SLICE_X54Y124_AO6),
.I3(CLBLL_L_X34Y128_SLICE_X50Y128_AO6),
.I4(LIOB33_X0Y147_IOB_X0Y147_I),
.I5(CLBLM_R_X35Y126_SLICE_X53Y126_A_XOR),
.O5(CLBLL_L_X36Y125_SLICE_X54Y125_BO5),
.O6(CLBLL_L_X36Y125_SLICE_X54Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ae00ae00ae00)
  ) CLBLL_L_X36Y125_SLICE_X54Y125_ALUT (
.I0(CLBLM_R_X35Y126_SLICE_X52Y126_AO6),
.I1(CLBLM_R_X35Y126_SLICE_X53Y126_A_XOR),
.I2(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(CLBLL_L_X36Y122_SLICE_X55Y122_AO6),
.I5(CLBLM_R_X35Y124_SLICE_X52Y124_A_XOR),
.O5(CLBLL_L_X36Y125_SLICE_X54Y125_AO5),
.O6(CLBLL_L_X36Y125_SLICE_X54Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he2c0c0c000000000)
  ) CLBLL_L_X36Y125_SLICE_X55Y125_DLUT (
.I0(RIOB33_X105Y115_IOB_X1Y116_I),
.I1(LIOB33_X0Y145_IOB_X0Y146_I),
.I2(CLBLL_L_X34Y126_SLICE_X50Y126_CO6),
.I3(CLBLL_L_X36Y121_SLICE_X54Y121_AO5),
.I4(CLBLL_L_X36Y116_SLICE_X54Y116_BO5),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLL_L_X36Y125_SLICE_X55Y125_DO5),
.O6(CLBLL_L_X36Y125_SLICE_X55Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbf8fbc8cb383b080)
  ) CLBLL_L_X36Y125_SLICE_X55Y125_CLUT (
.I0(CLBLL_L_X34Y125_SLICE_X50Y125_AO6),
.I1(LIOB33_X0Y145_IOB_X0Y146_I),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(CLBLM_R_X37Y125_SLICE_X56Y125_BO6),
.I4(CLBLL_L_X36Y124_SLICE_X55Y124_BO6),
.I5(CLBLL_L_X34Y126_SLICE_X50Y126_BO6),
.O5(CLBLL_L_X36Y125_SLICE_X55Y125_CO5),
.O6(CLBLL_L_X36Y125_SLICE_X55Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00500050f0f1f0e0)
  ) CLBLL_L_X36Y125_SLICE_X55Y125_BLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(RIOB33_X105Y117_IOB_X1Y117_I),
.I3(LIOB33_X0Y117_IOB_X0Y118_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(1'b1),
.O5(CLBLL_L_X36Y125_SLICE_X55Y125_BO5),
.O6(CLBLL_L_X36Y125_SLICE_X55Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0afa0cacacaca)
  ) CLBLL_L_X36Y125_SLICE_X55Y125_ALUT (
.I0(CLBLL_L_X36Y125_SLICE_X55Y125_BO5),
.I1(CLBLL_L_X36Y124_SLICE_X55Y124_DO6),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(CLBLM_R_X37Y123_SLICE_X56Y123_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y125_SLICE_X55Y125_AO5),
.O6(CLBLL_L_X36Y125_SLICE_X55Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffb8ffb800b800b8)
  ) CLBLL_L_X36Y126_SLICE_X54Y126_DLUT (
.I0(CLBLL_L_X36Y125_SLICE_X55Y125_AO5),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(CLBLM_R_X37Y126_SLICE_X56Y126_AO6),
.I3(LIOB33_X0Y145_IOB_X0Y146_I),
.I4(1'b1),
.I5(CLBLM_R_X35Y126_SLICE_X53Y126_C_XOR),
.O5(CLBLL_L_X36Y126_SLICE_X54Y126_DO5),
.O6(CLBLL_L_X36Y126_SLICE_X54Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcfffc000cf00c0)
  ) CLBLL_L_X36Y126_SLICE_X54Y126_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X37Y126_SLICE_X56Y126_AO6),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(LIOB33_X0Y145_IOB_X0Y146_I),
.I4(CLBLL_L_X36Y125_SLICE_X55Y125_AO6),
.I5(CLBLM_R_X35Y126_SLICE_X53Y126_B_XOR),
.O5(CLBLL_L_X36Y126_SLICE_X54Y126_CO5),
.O6(CLBLL_L_X36Y126_SLICE_X54Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb0b08080f000f000)
  ) CLBLL_L_X36Y126_SLICE_X54Y126_BLUT (
.I0(CLBLL_L_X36Y126_SLICE_X54Y126_DO6),
.I1(LIOB33_X0Y147_IOB_X0Y147_I),
.I2(CLBLL_L_X34Y128_SLICE_X50Y128_AO6),
.I3(CLBLM_R_X35Y126_SLICE_X53Y126_C_XOR),
.I4(CLBLL_L_X36Y125_SLICE_X54Y125_CO6),
.I5(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.O5(CLBLL_L_X36Y126_SLICE_X54Y126_BO5),
.O6(CLBLL_L_X36Y126_SLICE_X54Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0d07050a0802000)
  ) CLBLL_L_X36Y126_SLICE_X54Y126_ALUT (
.I0(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I1(LIOB33_X0Y147_IOB_X0Y147_I),
.I2(CLBLL_L_X34Y128_SLICE_X50Y128_AO6),
.I3(CLBLL_L_X36Y124_SLICE_X54Y124_BO6),
.I4(CLBLL_L_X36Y126_SLICE_X54Y126_CO6),
.I5(CLBLM_R_X35Y126_SLICE_X53Y126_B_XOR),
.O5(CLBLL_L_X36Y126_SLICE_X54Y126_AO5),
.O6(CLBLL_L_X36Y126_SLICE_X54Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeeccee33220022)
  ) CLBLL_L_X36Y126_SLICE_X55Y126_DLUT (
.I0(CLBLL_L_X36Y125_SLICE_X55Y125_AO5),
.I1(LIOB33_X0Y145_IOB_X0Y146_I),
.I2(1'b1),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(CLBLM_R_X37Y126_SLICE_X56Y126_AO5),
.I5(CLBLM_R_X35Y126_SLICE_X53Y126_D_XOR),
.O5(CLBLL_L_X36Y126_SLICE_X55Y126_DO5),
.O6(CLBLL_L_X36Y126_SLICE_X55Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0e0f0c0c0e0c0)
  ) CLBLL_L_X36Y126_SLICE_X55Y126_CLUT (
.I0(CLBLL_L_X34Y127_SLICE_X50Y127_AO6),
.I1(CLBLL_L_X36Y125_SLICE_X55Y125_DO6),
.I2(CLBLL_L_X36Y122_SLICE_X55Y122_AO5),
.I3(LIOB33_X0Y145_IOB_X0Y146_I),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(CLBLM_R_X37Y127_SLICE_X56Y127_AO6),
.O5(CLBLL_L_X36Y126_SLICE_X55Y126_CO5),
.O6(CLBLL_L_X36Y126_SLICE_X55Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8d8d8ff55aa00)
  ) CLBLL_L_X36Y126_SLICE_X55Y126_BLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(CLBLL_L_X34Y126_SLICE_X50Y126_BO6),
.I2(CLBLL_L_X34Y126_SLICE_X50Y126_CO6),
.I3(CLBLM_R_X37Y127_SLICE_X56Y127_AO6),
.I4(CLBLM_R_X37Y125_SLICE_X56Y125_BO6),
.I5(LIOB33_X0Y145_IOB_X0Y146_I),
.O5(CLBLL_L_X36Y126_SLICE_X55Y126_BO5),
.O6(CLBLL_L_X36Y126_SLICE_X55Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb008800f000f000)
  ) CLBLL_L_X36Y126_SLICE_X55Y126_ALUT (
.I0(CLBLL_L_X36Y126_SLICE_X55Y126_DO6),
.I1(LIOB33_X0Y147_IOB_X0Y147_I),
.I2(CLBLM_R_X35Y126_SLICE_X53Y126_D_XOR),
.I3(CLBLL_L_X34Y128_SLICE_X50Y128_AO6),
.I4(CLBLL_L_X36Y125_SLICE_X55Y125_CO6),
.I5(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.O5(CLBLL_L_X36Y126_SLICE_X55Y126_AO5),
.O6(CLBLL_L_X36Y126_SLICE_X55Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a030c0a0a0)
  ) CLBLL_L_X36Y127_SLICE_X54Y127_DLUT (
.I0(CLBLM_R_X35Y126_SLICE_X53Y126_B_XOR),
.I1(LIOB33_X0Y139_IOB_X0Y139_I),
.I2(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(LIOB33_X0Y145_IOB_X0Y146_I),
.I5(LIOB33_X0Y147_IOB_X0Y147_I),
.O5(CLBLL_L_X36Y127_SLICE_X54Y127_DO5),
.O6(CLBLL_L_X36Y127_SLICE_X54Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00b300ff00a000)
  ) CLBLL_L_X36Y127_SLICE_X54Y127_CLUT (
.I0(CLBLL_L_X36Y122_SLICE_X55Y122_AO6),
.I1(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.I2(CLBLM_R_X35Y124_SLICE_X52Y124_B_XOR),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(CLBLL_L_X36Y127_SLICE_X54Y127_DO6),
.I5(CLBLM_R_X35Y126_SLICE_X53Y126_B_XOR),
.O5(CLBLL_L_X36Y127_SLICE_X54Y127_CO5),
.O6(CLBLL_L_X36Y127_SLICE_X54Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffe800)
  ) CLBLL_L_X36Y127_SLICE_X54Y127_BLUT (
.I0(LIOB33_X0Y139_IOB_X0Y139_I),
.I1(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I2(RIOB33_X105Y111_IOB_X1Y111_I),
.I3(CLBLL_L_X36Y116_SLICE_X55Y116_AO5),
.I4(CLBLL_L_X36Y126_SLICE_X54Y126_AO6),
.I5(CLBLL_L_X36Y127_SLICE_X54Y127_CO6),
.O5(CLBLL_L_X36Y127_SLICE_X54Y127_BO5),
.O6(CLBLL_L_X36Y127_SLICE_X54Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffaf8fffff8f0)
  ) CLBLL_L_X36Y127_SLICE_X54Y127_ALUT (
.I0(CLBLL_L_X36Y116_SLICE_X55Y116_AO5),
.I1(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I2(CLBLL_L_X36Y125_SLICE_X54Y125_BO6),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(CLBLL_L_X36Y125_SLICE_X54Y125_AO6),
.I5(LIOB33_X0Y137_IOB_X0Y138_I),
.O5(CLBLL_L_X36Y127_SLICE_X54Y127_AO5),
.O6(CLBLL_L_X36Y127_SLICE_X54Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000300)
  ) CLBLL_L_X36Y127_SLICE_X55Y127_DLUT (
.I0(1'b1),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(RIOB33_X105Y115_IOB_X1Y116_I),
.I4(LIOB33_X0Y117_IOB_X0Y118_I),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLL_L_X36Y127_SLICE_X55Y127_DO5),
.O6(CLBLL_L_X36Y127_SLICE_X55Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcaffca0fcaf0ca00)
  ) CLBLL_L_X36Y127_SLICE_X55Y127_CLUT (
.I0(CLBLL_L_X34Y127_SLICE_X50Y127_AO6),
.I1(CLBLL_L_X34Y126_SLICE_X50Y126_CO6),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(LIOB33_X0Y145_IOB_X0Y146_I),
.I4(CLBLL_L_X36Y127_SLICE_X55Y127_DO6),
.I5(CLBLM_R_X37Y127_SLICE_X56Y127_AO6),
.O5(CLBLL_L_X36Y127_SLICE_X55Y127_CO5),
.O6(CLBLL_L_X36Y127_SLICE_X55Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heef044f0eee444e4)
  ) CLBLL_L_X36Y127_SLICE_X55Y127_BLUT (
.I0(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I1(CLBLM_R_X35Y127_SLICE_X53Y127_A_XOR),
.I2(CLBLL_L_X36Y126_SLICE_X55Y126_BO6),
.I3(LIOB33_X0Y147_IOB_X0Y147_I),
.I4(CLBLL_L_X36Y128_SLICE_X55Y128_DO6),
.I5(LIOB33_X0Y145_IOB_X0Y146_I),
.O5(CLBLL_L_X36Y127_SLICE_X55Y127_BO5),
.O6(CLBLL_L_X36Y127_SLICE_X55Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccccccdccc8)
  ) CLBLL_L_X36Y127_SLICE_X55Y127_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(RIOB33_X105Y117_IOB_X1Y117_I),
.I2(LIOB33_X0Y117_IOB_X0Y118_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(RIOB33_X105Y115_IOB_X1Y115_I),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLL_L_X36Y127_SLICE_X55Y127_AO5),
.O6(CLBLL_L_X36Y127_SLICE_X55Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc30fc30ee22ee22)
  ) CLBLL_L_X36Y128_SLICE_X54Y128_DLUT (
.I0(CLBLL_L_X36Y127_SLICE_X55Y127_AO6),
.I1(LIOB33_X0Y145_IOB_X0Y146_I),
.I2(CLBLM_R_X37Y127_SLICE_X56Y127_BO6),
.I3(CLBLM_R_X35Y127_SLICE_X53Y127_B_XOR),
.I4(1'b1),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLL_L_X36Y128_SLICE_X54Y128_DO5),
.O6(CLBLL_L_X36Y128_SLICE_X54Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0c03000a0a0a0a0)
  ) CLBLL_L_X36Y128_SLICE_X54Y128_CLUT (
.I0(CLBLM_R_X35Y127_SLICE_X53Y127_B_XOR),
.I1(LIOB33_X0Y147_IOB_X0Y147_I),
.I2(CLBLL_L_X34Y128_SLICE_X50Y128_AO6),
.I3(CLBLL_L_X36Y127_SLICE_X55Y127_CO6),
.I4(CLBLL_L_X36Y128_SLICE_X54Y128_DO6),
.I5(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.O5(CLBLL_L_X36Y128_SLICE_X54Y128_CO5),
.O6(CLBLL_L_X36Y128_SLICE_X54Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8a8a8a80808a8080)
  ) CLBLL_L_X36Y128_SLICE_X54Y128_BLUT (
.I0(CLBLL_L_X36Y116_SLICE_X55Y116_AO6),
.I1(CLBLM_R_X35Y127_SLICE_X53Y127_B_XOR),
.I2(LIOB33_X0Y145_IOB_X0Y146_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(CLBLL_L_X36Y127_SLICE_X55Y127_AO6),
.I5(CLBLM_R_X37Y127_SLICE_X56Y127_BO6),
.O5(CLBLL_L_X36Y128_SLICE_X54Y128_BO5),
.O6(CLBLL_L_X36Y128_SLICE_X54Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff0f0fff4f0f0)
  ) CLBLL_L_X36Y128_SLICE_X54Y128_ALUT (
.I0(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I1(CLBLM_R_X35Y127_SLICE_X53Y127_B_XOR),
.I2(CLBLM_R_X35Y127_SLICE_X52Y127_AO6),
.I3(CLBLL_L_X36Y128_SLICE_X54Y128_BO6),
.I4(CLBLL_L_X34Y128_SLICE_X50Y128_AO6),
.I5(CLBLL_L_X36Y126_SLICE_X55Y126_CO6),
.O5(CLBLL_L_X36Y128_SLICE_X54Y128_AO5),
.O6(CLBLL_L_X36Y128_SLICE_X54Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbbff8800bb0088)
  ) CLBLL_L_X36Y128_SLICE_X55Y128_DLUT (
.I0(CLBLL_L_X36Y127_SLICE_X55Y127_AO6),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(1'b1),
.I3(LIOB33_X0Y145_IOB_X0Y146_I),
.I4(CLBLM_R_X37Y126_SLICE_X56Y126_AO5),
.I5(CLBLM_R_X35Y127_SLICE_X53Y127_A_XOR),
.O5(CLBLL_L_X36Y128_SLICE_X55Y128_DO5),
.O6(CLBLL_L_X36Y128_SLICE_X55Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000101000001013)
  ) CLBLL_L_X36Y128_SLICE_X55Y128_CLUT (
.I0(CLBLM_R_X35Y129_SLICE_X53Y129_AO6),
.I1(CLBLL_L_X36Y128_SLICE_X54Y128_CO6),
.I2(LIOB33_X0Y147_IOB_X0Y148_I),
.I3(CLBLM_R_X35Y128_SLICE_X52Y128_BO6),
.I4(CLBLM_R_X35Y127_SLICE_X52Y127_AO6),
.I5(CLBLM_R_X35Y129_SLICE_X53Y129_BO6),
.O5(CLBLL_L_X36Y128_SLICE_X55Y128_CO5),
.O6(CLBLL_L_X36Y128_SLICE_X55Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000ff00cd)
  ) CLBLL_L_X36Y128_SLICE_X55Y128_BLUT (
.I0(CLBLM_R_X35Y129_SLICE_X52Y129_AO6),
.I1(CLBLM_R_X35Y128_SLICE_X52Y128_CO6),
.I2(CLBLL_L_X36Y126_SLICE_X55Y126_AO6),
.I3(CLBLL_L_X36Y128_SLICE_X54Y128_CO6),
.I4(CLBLL_L_X36Y128_SLICE_X55Y128_AO6),
.I5(CLBLM_R_X35Y127_SLICE_X52Y127_AO6),
.O5(CLBLL_L_X36Y128_SLICE_X55Y128_BO5),
.O6(CLBLL_L_X36Y128_SLICE_X55Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hacff0000ac000000)
  ) CLBLL_L_X36Y128_SLICE_X55Y128_ALUT (
.I0(CLBLL_L_X36Y128_SLICE_X55Y128_DO6),
.I1(CLBLL_L_X36Y126_SLICE_X55Y126_BO6),
.I2(LIOB33_X0Y147_IOB_X0Y147_I),
.I3(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I4(CLBLL_L_X34Y128_SLICE_X50Y128_AO6),
.I5(CLBLM_R_X35Y127_SLICE_X53Y127_A_XOR),
.O5(CLBLL_L_X36Y128_SLICE_X55Y128_AO5),
.O6(CLBLL_L_X36Y128_SLICE_X55Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X36Y129_SLICE_X54Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y129_SLICE_X54Y129_DO5),
.O6(CLBLL_L_X36Y129_SLICE_X54Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbf00fb0004004000)
  ) CLBLL_L_X36Y129_SLICE_X54Y129_CLUT (
.I0(LIOB33_X0Y147_IOB_X0Y147_I),
.I1(LIOB33_X0Y145_IOB_X0Y146_I),
.I2(RIOB33_X105Y113_IOB_X1Y114_I),
.I3(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I4(LIOB33_X0Y141_IOB_X0Y142_I),
.I5(CLBLM_R_X35Y127_SLICE_X53Y127_A_XOR),
.O5(CLBLL_L_X36Y129_SLICE_X54Y129_CO5),
.O6(CLBLL_L_X36Y129_SLICE_X54Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa8080aa80)
  ) CLBLL_L_X36Y129_SLICE_X54Y129_BLUT (
.I0(LIOB33_X0Y147_IOB_X0Y148_I),
.I1(CLBLM_R_X35Y125_SLICE_X52Y125_A_XOR),
.I2(CLBLL_L_X36Y122_SLICE_X55Y122_AO6),
.I3(CLBLM_R_X35Y127_SLICE_X53Y127_A_XOR),
.I4(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.I5(CLBLL_L_X36Y129_SLICE_X54Y129_CO6),
.O5(CLBLL_L_X36Y129_SLICE_X54Y129_BO5),
.O6(CLBLL_L_X36Y129_SLICE_X54Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeeffecffecffcc)
  ) CLBLL_L_X36Y129_SLICE_X54Y129_ALUT (
.I0(CLBLL_L_X36Y116_SLICE_X55Y116_AO5),
.I1(CLBLL_L_X36Y128_SLICE_X55Y128_AO6),
.I2(RIOB33_X105Y113_IOB_X1Y114_I),
.I3(CLBLL_L_X36Y129_SLICE_X54Y129_BO6),
.I4(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I5(LIOB33_X0Y141_IOB_X0Y142_I),
.O5(CLBLL_L_X36Y129_SLICE_X54Y129_AO5),
.O6(CLBLL_L_X36Y129_SLICE_X54Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffafffa0f0a0f0a)
  ) CLBLL_L_X36Y129_SLICE_X55Y129_DLUT (
.I0(CLBLM_R_X35Y128_SLICE_X52Y128_BO6),
.I1(1'b1),
.I2(LIOB33_X0Y147_IOB_X0Y148_I),
.I3(CLBLM_R_X35Y129_SLICE_X53Y129_BO6),
.I4(1'b1),
.I5(CLBLM_R_X35Y129_SLICE_X53Y129_AO6),
.O5(CLBLL_L_X36Y129_SLICE_X55Y129_DO5),
.O6(CLBLL_L_X36Y129_SLICE_X55Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbf00fb0004004000)
  ) CLBLL_L_X36Y129_SLICE_X55Y129_CLUT (
.I0(LIOB33_X0Y147_IOB_X0Y147_I),
.I1(LIOB33_X0Y145_IOB_X0Y146_I),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I4(LIOB33_X0Y141_IOB_X0Y141_I),
.I5(CLBLM_R_X35Y126_SLICE_X53Y126_D_XOR),
.O5(CLBLL_L_X36Y129_SLICE_X55Y129_CO5),
.O6(CLBLL_L_X36Y129_SLICE_X55Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaaa080808)
  ) CLBLL_L_X36Y129_SLICE_X55Y129_BLUT (
.I0(LIOB33_X0Y147_IOB_X0Y148_I),
.I1(CLBLM_R_X35Y126_SLICE_X53Y126_D_XOR),
.I2(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.I3(CLBLL_L_X36Y122_SLICE_X55Y122_AO6),
.I4(CLBLM_R_X35Y124_SLICE_X52Y124_D_XOR),
.I5(CLBLL_L_X36Y129_SLICE_X55Y129_CO6),
.O5(CLBLL_L_X36Y129_SLICE_X55Y129_BO5),
.O6(CLBLL_L_X36Y129_SLICE_X55Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffa8ffffff80)
  ) CLBLL_L_X36Y129_SLICE_X55Y129_ALUT (
.I0(CLBLL_L_X36Y116_SLICE_X55Y116_AO5),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I3(CLBLL_L_X36Y129_SLICE_X55Y129_BO6),
.I4(CLBLL_L_X36Y126_SLICE_X55Y126_AO6),
.I5(LIOB33_X0Y141_IOB_X0Y141_I),
.O5(CLBLL_L_X36Y129_SLICE_X55Y129_AO5),
.O6(CLBLL_L_X36Y129_SLICE_X55Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X38Y118_SLICE_X58Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X38Y118_SLICE_X58Y118_DO5),
.O6(CLBLL_L_X38Y118_SLICE_X58Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X38Y118_SLICE_X58Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X38Y118_SLICE_X58Y118_CO5),
.O6(CLBLL_L_X38Y118_SLICE_X58Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X38Y118_SLICE_X58Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X38Y118_SLICE_X58Y118_BO5),
.O6(CLBLL_L_X38Y118_SLICE_X58Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaafa0aaaaacac)
  ) CLBLL_L_X38Y118_SLICE_X58Y118_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y117_I),
.I1(RIOB33_X105Y111_IOB_X1Y111_I),
.I2(LIOB33_X0Y117_IOB_X0Y118_I),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(1'b1),
.O5(CLBLL_L_X38Y118_SLICE_X58Y118_AO5),
.O6(CLBLL_L_X38Y118_SLICE_X58Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X38Y118_SLICE_X59Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X38Y118_SLICE_X59Y118_DO5),
.O6(CLBLL_L_X38Y118_SLICE_X59Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X38Y118_SLICE_X59Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X38Y118_SLICE_X59Y118_CO5),
.O6(CLBLL_L_X38Y118_SLICE_X59Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X38Y118_SLICE_X59Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X38Y118_SLICE_X59Y118_BO5),
.O6(CLBLL_L_X38Y118_SLICE_X59Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X38Y118_SLICE_X59Y118_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X38Y118_SLICE_X59Y118_AO5),
.O6(CLBLL_L_X38Y118_SLICE_X59Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X38Y119_SLICE_X58Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X38Y119_SLICE_X58Y119_DO5),
.O6(CLBLL_L_X38Y119_SLICE_X58Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X38Y119_SLICE_X58Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X38Y119_SLICE_X58Y119_CO5),
.O6(CLBLL_L_X38Y119_SLICE_X58Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X38Y119_SLICE_X58Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X38Y119_SLICE_X58Y119_BO5),
.O6(CLBLL_L_X38Y119_SLICE_X58Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00005e0e00005404)
  ) CLBLL_L_X38Y119_SLICE_X58Y119_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(RIOB33_X105Y115_IOB_X1Y115_I),
.I4(LIOB33_X0Y117_IOB_X0Y118_I),
.I5(RIOB33_X105Y111_IOB_X1Y111_I),
.O5(CLBLL_L_X38Y119_SLICE_X58Y119_AO5),
.O6(CLBLL_L_X38Y119_SLICE_X58Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X38Y119_SLICE_X59Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X38Y119_SLICE_X59Y119_DO5),
.O6(CLBLL_L_X38Y119_SLICE_X59Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X38Y119_SLICE_X59Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X38Y119_SLICE_X59Y119_CO5),
.O6(CLBLL_L_X38Y119_SLICE_X59Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X38Y119_SLICE_X59Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X38Y119_SLICE_X59Y119_BO5),
.O6(CLBLL_L_X38Y119_SLICE_X59Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X38Y119_SLICE_X59Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X38Y119_SLICE_X59Y119_AO5),
.O6(CLBLL_L_X38Y119_SLICE_X59Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0405040504000400)
  ) CLBLL_L_X38Y121_SLICE_X58Y121_DLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(RIOB33_X105Y115_IOB_X1Y115_I),
.I2(LIOB33_X0Y117_IOB_X0Y118_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(1'b1),
.I5(RIOB33_X105Y111_IOB_X1Y111_I),
.O5(CLBLL_L_X38Y121_SLICE_X58Y121_DO5),
.O6(CLBLL_L_X38Y121_SLICE_X58Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h882ebbaa882e88aa)
  ) CLBLL_L_X38Y121_SLICE_X58Y121_CLUT (
.I0(CLBLM_R_X35Y123_SLICE_X53Y123_C_XOR),
.I1(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I2(CLBLM_R_X37Y121_SLICE_X57Y121_DO5),
.I3(LIOB33_X0Y147_IOB_X0Y147_I),
.I4(LIOB33_X0Y145_IOB_X0Y146_I),
.I5(CLBLM_R_X35Y121_SLICE_X52Y121_C_XOR),
.O5(CLBLL_L_X38Y121_SLICE_X58Y121_CO5),
.O6(CLBLL_L_X38Y121_SLICE_X58Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f2f2f003020200)
  ) CLBLL_L_X38Y121_SLICE_X58Y121_BLUT (
.I0(LIOB33_X0Y127_IOB_X0Y128_I),
.I1(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.I2(LIOB33_X0Y147_IOB_X0Y148_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I5(CLBLL_L_X38Y121_SLICE_X58Y121_CO6),
.O5(CLBLL_L_X38Y121_SLICE_X58Y121_BO5),
.O6(CLBLL_L_X38Y121_SLICE_X58Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcaca0a0afa0a0a0a)
  ) CLBLL_L_X38Y121_SLICE_X58Y121_ALUT (
.I0(CLBLL_L_X38Y121_SLICE_X58Y121_DO6),
.I1(RIOB33_X105Y117_IOB_X1Y117_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(CLBLL_L_X36Y121_SLICE_X54Y121_AO5),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLL_L_X38Y121_SLICE_X58Y121_AO5),
.O6(CLBLL_L_X38Y121_SLICE_X58Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X38Y121_SLICE_X59Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X38Y121_SLICE_X59Y121_DO5),
.O6(CLBLL_L_X38Y121_SLICE_X59Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X38Y121_SLICE_X59Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X38Y121_SLICE_X59Y121_CO5),
.O6(CLBLL_L_X38Y121_SLICE_X59Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X38Y121_SLICE_X59Y121_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X38Y121_SLICE_X59Y121_BO5),
.O6(CLBLL_L_X38Y121_SLICE_X59Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X38Y121_SLICE_X59Y121_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X38Y121_SLICE_X59Y121_AO5),
.O6(CLBLL_L_X38Y121_SLICE_X59Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X38Y123_SLICE_X58Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X38Y123_SLICE_X58Y123_DO5),
.O6(CLBLL_L_X38Y123_SLICE_X58Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X38Y123_SLICE_X58Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X38Y123_SLICE_X58Y123_CO5),
.O6(CLBLL_L_X38Y123_SLICE_X58Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X38Y123_SLICE_X58Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X38Y123_SLICE_X58Y123_BO5),
.O6(CLBLL_L_X38Y123_SLICE_X58Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X38Y123_SLICE_X58Y123_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X38Y123_SLICE_X58Y123_AO5),
.O6(CLBLL_L_X38Y123_SLICE_X58Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X38Y123_SLICE_X59Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X38Y123_SLICE_X59Y123_DO5),
.O6(CLBLL_L_X38Y123_SLICE_X59Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X38Y123_SLICE_X59Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X38Y123_SLICE_X59Y123_CO5),
.O6(CLBLL_L_X38Y123_SLICE_X59Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X38Y123_SLICE_X59Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X38Y123_SLICE_X59Y123_BO5),
.O6(CLBLL_L_X38Y123_SLICE_X59Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000310000003131)
  ) CLBLL_L_X38Y123_SLICE_X59Y123_ALUT (
.I0(CLBLL_L_X34Y121_SLICE_X51Y121_AO6),
.I1(CLBLM_R_X33Y121_SLICE_X48Y121_AO6),
.I2(CLBLM_R_X33Y123_SLICE_X49Y123_AO6),
.I3(CLBLL_L_X34Y120_SLICE_X51Y120_AO6),
.I4(CLBLL_L_X36Y122_SLICE_X54Y122_BO6),
.I5(CLBLL_L_X36Y119_SLICE_X55Y119_BO6),
.O5(CLBLL_L_X38Y123_SLICE_X59Y123_AO5),
.O6(CLBLL_L_X38Y123_SLICE_X59Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X38Y124_SLICE_X58Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X38Y124_SLICE_X58Y124_DO5),
.O6(CLBLL_L_X38Y124_SLICE_X58Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf00ff00ff00ff00f)
  ) CLBLL_L_X38Y124_SLICE_X58Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y133_IOB_X0Y134_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X38Y124_SLICE_X58Y124_CO5),
.O6(CLBLL_L_X38Y124_SLICE_X58Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc00ccaccc0fccacc)
  ) CLBLL_L_X38Y124_SLICE_X58Y124_BLUT (
.I0(CLBLM_R_X35Y123_SLICE_X52Y123_A_XOR),
.I1(CLBLM_R_X35Y125_SLICE_X53Y125_A_XOR),
.I2(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I3(LIOB33_X0Y147_IOB_X0Y147_I),
.I4(LIOB33_X0Y145_IOB_X0Y146_I),
.I5(CLBLL_L_X38Y124_SLICE_X58Y124_CO6),
.O5(CLBLL_L_X38Y124_SLICE_X58Y124_BO5),
.O6(CLBLL_L_X38Y124_SLICE_X58Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000fe0ef808)
  ) CLBLL_L_X38Y124_SLICE_X58Y124_ALUT (
.I0(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I1(LIOB33_X0Y133_IOB_X0Y134_I),
.I2(LIOB33_X0Y147_IOB_X0Y148_I),
.I3(CLBLL_L_X38Y124_SLICE_X58Y124_BO6),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.O5(CLBLL_L_X38Y124_SLICE_X58Y124_AO5),
.O6(CLBLL_L_X38Y124_SLICE_X58Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X38Y124_SLICE_X59Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X38Y124_SLICE_X59Y124_DO5),
.O6(CLBLL_L_X38Y124_SLICE_X59Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X38Y124_SLICE_X59Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X38Y124_SLICE_X59Y124_CO5),
.O6(CLBLL_L_X38Y124_SLICE_X59Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X38Y124_SLICE_X59Y124_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X38Y124_SLICE_X59Y124_BO5),
.O6(CLBLL_L_X38Y124_SLICE_X59Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X38Y124_SLICE_X59Y124_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X38Y124_SLICE_X59Y124_AO5),
.O6(CLBLL_L_X38Y124_SLICE_X59Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X38Y126_SLICE_X58Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X38Y126_SLICE_X58Y126_DO5),
.O6(CLBLL_L_X38Y126_SLICE_X58Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a030a0a0a0c0a0)
  ) CLBLL_L_X38Y126_SLICE_X58Y126_CLUT (
.I0(CLBLM_R_X35Y125_SLICE_X53Y125_D_XOR),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I3(LIOB33_X0Y145_IOB_X0Y146_I),
.I4(LIOB33_X0Y147_IOB_X0Y147_I),
.I5(LIOB33_X0Y137_IOB_X0Y137_I),
.O5(CLBLL_L_X38Y126_SLICE_X58Y126_CO5),
.O6(CLBLL_L_X38Y126_SLICE_X58Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaaa202020)
  ) CLBLL_L_X38Y126_SLICE_X58Y126_BLUT (
.I0(LIOB33_X0Y147_IOB_X0Y148_I),
.I1(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.I2(CLBLM_R_X35Y125_SLICE_X53Y125_D_XOR),
.I3(CLBLM_R_X35Y123_SLICE_X52Y123_D_XOR),
.I4(CLBLL_L_X36Y122_SLICE_X55Y122_AO6),
.I5(CLBLL_L_X38Y126_SLICE_X58Y126_CO6),
.O5(CLBLL_L_X38Y126_SLICE_X58Y126_BO5),
.O6(CLBLL_L_X38Y126_SLICE_X58Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffafff8fff8fff0)
  ) CLBLL_L_X38Y126_SLICE_X58Y126_ALUT (
.I0(CLBLL_L_X36Y116_SLICE_X55Y116_AO5),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(CLBLM_R_X37Y125_SLICE_X57Y125_DO6),
.I3(CLBLL_L_X38Y126_SLICE_X58Y126_BO6),
.I4(LIOB33_X0Y137_IOB_X0Y137_I),
.I5(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.O5(CLBLL_L_X38Y126_SLICE_X58Y126_AO5),
.O6(CLBLL_L_X38Y126_SLICE_X58Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X38Y126_SLICE_X59Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X38Y126_SLICE_X59Y126_DO5),
.O6(CLBLL_L_X38Y126_SLICE_X59Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000051005151)
  ) CLBLL_L_X38Y126_SLICE_X59Y126_CLUT (
.I0(CLBLM_R_X37Y122_SLICE_X57Y122_AO6),
.I1(CLBLL_L_X36Y122_SLICE_X55Y122_BO6),
.I2(CLBLM_R_X37Y121_SLICE_X57Y121_AO6),
.I3(CLBLM_R_X35Y119_SLICE_X53Y119_AO6),
.I4(CLBLL_L_X34Y124_SLICE_X50Y124_AO6),
.I5(CLBLL_L_X36Y121_SLICE_X55Y121_BO6),
.O5(CLBLL_L_X38Y126_SLICE_X59Y126_CO5),
.O6(CLBLL_L_X38Y126_SLICE_X59Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLL_L_X38Y126_SLICE_X59Y126_BLUT (
.I0(CLBLM_R_X37Y123_SLICE_X57Y123_AO6),
.I1(CLBLM_R_X37Y125_SLICE_X56Y125_AO6),
.I2(CLBLM_R_X37Y125_SLICE_X57Y125_AO6),
.I3(CLBLL_L_X38Y126_SLICE_X58Y126_AO6),
.I4(CLBLM_R_X37Y123_SLICE_X56Y123_BO6),
.I5(CLBLM_R_X37Y126_SLICE_X56Y126_BO6),
.O5(CLBLL_L_X38Y126_SLICE_X59Y126_BO5),
.O6(CLBLL_L_X38Y126_SLICE_X59Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLL_L_X38Y126_SLICE_X59Y126_ALUT (
.I0(CLBLM_R_X35Y116_SLICE_X53Y116_DO6),
.I1(CLBLM_R_X37Y124_SLICE_X56Y124_DO6),
.I2(CLBLM_R_X37Y128_SLICE_X56Y128_AO6),
.I3(CLBLL_L_X38Y126_SLICE_X59Y126_BO6),
.I4(CLBLL_L_X38Y123_SLICE_X59Y123_AO6),
.I5(CLBLL_L_X38Y126_SLICE_X59Y126_CO6),
.O5(CLBLL_L_X38Y126_SLICE_X59Y126_AO5),
.O6(CLBLL_L_X38Y126_SLICE_X59Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X32Y116_SLICE_X46Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X32Y116_SLICE_X46Y116_DO5),
.O6(CLBLM_L_X32Y116_SLICE_X46Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X32Y116_SLICE_X46Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X32Y116_SLICE_X46Y116_CO5),
.O6(CLBLM_L_X32Y116_SLICE_X46Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X32Y116_SLICE_X46Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X32Y116_SLICE_X46Y116_BO5),
.O6(CLBLM_L_X32Y116_SLICE_X46Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X32Y116_SLICE_X46Y116_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X32Y116_SLICE_X46Y116_AO5),
.O6(CLBLM_L_X32Y116_SLICE_X46Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X32Y116_SLICE_X47Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X32Y116_SLICE_X47Y116_DO5),
.O6(CLBLM_L_X32Y116_SLICE_X47Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X32Y116_SLICE_X47Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X32Y116_SLICE_X47Y116_CO5),
.O6(CLBLM_L_X32Y116_SLICE_X47Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X32Y116_SLICE_X47Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X32Y116_SLICE_X47Y116_BO5),
.O6(CLBLM_L_X32Y116_SLICE_X47Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000011100100)
  ) CLBLM_L_X32Y116_SLICE_X47Y116_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(LIOB33_X0Y117_IOB_X0Y118_I),
.O5(CLBLM_L_X32Y116_SLICE_X47Y116_AO5),
.O6(CLBLM_L_X32Y116_SLICE_X47Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X32Y117_SLICE_X46Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X32Y117_SLICE_X46Y117_DO5),
.O6(CLBLM_L_X32Y117_SLICE_X46Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X32Y117_SLICE_X46Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X32Y117_SLICE_X46Y117_CO5),
.O6(CLBLM_L_X32Y117_SLICE_X46Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X32Y117_SLICE_X46Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X32Y117_SLICE_X46Y117_BO5),
.O6(CLBLM_L_X32Y117_SLICE_X46Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X32Y117_SLICE_X46Y117_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X32Y117_SLICE_X46Y117_AO5),
.O6(CLBLM_L_X32Y117_SLICE_X46Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X32Y117_SLICE_X47Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X32Y117_SLICE_X47Y117_DO5),
.O6(CLBLM_L_X32Y117_SLICE_X47Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X32Y117_SLICE_X47Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X32Y117_SLICE_X47Y117_CO5),
.O6(CLBLM_L_X32Y117_SLICE_X47Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X32Y117_SLICE_X47Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X32Y117_SLICE_X47Y117_BO5),
.O6(CLBLM_L_X32Y117_SLICE_X47Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000510040)
  ) CLBLM_L_X32Y117_SLICE_X47Y117_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(LIOB33_X0Y117_IOB_X0Y118_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_L_X32Y117_SLICE_X47Y117_AO5),
.O6(CLBLM_L_X32Y117_SLICE_X47Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X32Y123_SLICE_X46Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X32Y123_SLICE_X46Y123_DO5),
.O6(CLBLM_L_X32Y123_SLICE_X46Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X32Y123_SLICE_X46Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X32Y123_SLICE_X46Y123_CO5),
.O6(CLBLM_L_X32Y123_SLICE_X46Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X32Y123_SLICE_X46Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X32Y123_SLICE_X46Y123_BO5),
.O6(CLBLM_L_X32Y123_SLICE_X46Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0705030106040200)
  ) CLBLM_L_X32Y123_SLICE_X46Y123_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_X0Y117_IOB_X0Y118_I),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_L_X32Y123_SLICE_X46Y123_AO5),
.O6(CLBLM_L_X32Y123_SLICE_X46Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacff0facacf000)
  ) CLBLM_L_X32Y123_SLICE_X47Y123_DLUT (
.I0(CLBLM_R_X33Y125_SLICE_X49Y125_BO6),
.I1(CLBLL_L_X34Y123_SLICE_X50Y123_BO6),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(CLBLM_L_X32Y123_SLICE_X47Y123_AO5),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(CLBLM_R_X33Y122_SLICE_X48Y122_AO5),
.O5(CLBLM_L_X32Y123_SLICE_X47Y123_DO5),
.O6(CLBLM_L_X32Y123_SLICE_X47Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafcfc0a0a0cfc0)
  ) CLBLM_L_X32Y123_SLICE_X47Y123_CLUT (
.I0(CLBLM_R_X33Y122_SLICE_X48Y122_AO6),
.I1(CLBLL_L_X34Y123_SLICE_X50Y123_BO6),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(CLBLM_L_X32Y123_SLICE_X47Y123_AO5),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(CLBLM_R_X33Y125_SLICE_X49Y125_BO6),
.O5(CLBLM_L_X32Y123_SLICE_X47Y123_CO5),
.O6(CLBLM_L_X32Y123_SLICE_X47Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa5500e4e4e4e4)
  ) CLBLM_L_X32Y123_SLICE_X47Y123_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(CLBLL_L_X34Y123_SLICE_X50Y123_BO6),
.I2(CLBLM_R_X33Y122_SLICE_X48Y122_AO6),
.I3(CLBLM_R_X33Y125_SLICE_X49Y125_BO6),
.I4(CLBLM_L_X32Y123_SLICE_X47Y123_AO6),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLM_L_X32Y123_SLICE_X47Y123_BO5),
.O6(CLBLM_L_X32Y123_SLICE_X47Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000e4e45050dd88)
  ) CLBLM_L_X32Y123_SLICE_X47Y123_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(LIOB33_X0Y117_IOB_X0Y118_I),
.I5(1'b1),
.O5(CLBLM_L_X32Y123_SLICE_X47Y123_AO5),
.O6(CLBLM_L_X32Y123_SLICE_X47Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X33Y115_SLICE_X48Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X33Y115_SLICE_X48Y115_DO5),
.O6(CLBLM_R_X33Y115_SLICE_X48Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X33Y115_SLICE_X48Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X33Y115_SLICE_X48Y115_CO5),
.O6(CLBLM_R_X33Y115_SLICE_X48Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X33Y115_SLICE_X48Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X33Y115_SLICE_X48Y115_BO5),
.O6(CLBLM_R_X33Y115_SLICE_X48Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa0000fcc0)
  ) CLBLM_R_X33Y115_SLICE_X48Y115_ALUT (
.I0(CLBLM_R_X33Y118_SLICE_X48Y118_CO6),
.I1(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.I5(LIOB33_X0Y147_IOB_X0Y148_I),
.O5(CLBLM_R_X33Y115_SLICE_X48Y115_AO5),
.O6(CLBLM_R_X33Y115_SLICE_X48Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4e4e4ff00ee44)
  ) CLBLM_R_X33Y115_SLICE_X49Y115_DLUT (
.I0(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I1(CLBLM_R_X35Y121_SLICE_X53Y121_A_XOR),
.I2(CLBLL_L_X34Y116_SLICE_X50Y116_AO5),
.I3(CLBLM_R_X33Y117_SLICE_X48Y117_CO6),
.I4(LIOB33_X0Y145_IOB_X0Y146_I),
.I5(LIOB33_X0Y147_IOB_X0Y147_I),
.O5(CLBLM_R_X33Y115_SLICE_X49Y115_DO5),
.O6(CLBLM_R_X33Y115_SLICE_X49Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50fa50ccccd8d8)
  ) CLBLM_R_X33Y115_SLICE_X49Y115_CLUT (
.I0(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I1(CLBLM_R_X33Y116_SLICE_X49Y116_CO6),
.I2(CLBLM_R_X35Y120_SLICE_X53Y120_C_XOR),
.I3(CLBLM_R_X33Y116_SLICE_X49Y116_DO6),
.I4(LIOB33_X0Y145_IOB_X0Y146_I),
.I5(LIOB33_X0Y147_IOB_X0Y147_I),
.O5(CLBLM_R_X33Y115_SLICE_X49Y115_CO5),
.O6(CLBLM_R_X33Y115_SLICE_X49Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0300030303010303)
  ) CLBLM_R_X33Y115_SLICE_X49Y115_BLUT (
.I0(CLBLM_R_X33Y115_SLICE_X49Y115_DO6),
.I1(CLBLL_L_X34Y115_SLICE_X51Y115_CO6),
.I2(CLBLM_R_X33Y115_SLICE_X48Y115_AO6),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.I5(CLBLM_R_X33Y115_SLICE_X49Y115_CO6),
.O5(CLBLM_R_X33Y115_SLICE_X49Y115_BO5),
.O6(CLBLM_R_X33Y115_SLICE_X49Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0001000011110000)
  ) CLBLM_R_X33Y115_SLICE_X49Y115_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y118_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(1'b1),
.O5(CLBLM_R_X33Y115_SLICE_X49Y115_AO5),
.O6(CLBLM_R_X33Y115_SLICE_X49Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hefeaefea45404540)
  ) CLBLM_R_X33Y116_SLICE_X48Y116_DLUT (
.I0(LIOB33_X0Y145_IOB_X0Y146_I),
.I1(CLBLL_L_X34Y117_SLICE_X51Y117_CO6),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(CLBLL_L_X34Y117_SLICE_X50Y117_CO6),
.I4(1'b1),
.I5(CLBLM_R_X35Y120_SLICE_X53Y120_D_XOR),
.O5(CLBLM_R_X33Y116_SLICE_X48Y116_DO5),
.O6(CLBLM_R_X33Y116_SLICE_X48Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha8aa08aaa8000800)
  ) CLBLM_R_X33Y116_SLICE_X48Y116_CLUT (
.I0(CLBLL_L_X34Y128_SLICE_X50Y128_AO6),
.I1(CLBLM_R_X33Y117_SLICE_X48Y117_BO6),
.I2(LIOB33_X0Y147_IOB_X0Y147_I),
.I3(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I4(CLBLM_R_X33Y116_SLICE_X48Y116_DO6),
.I5(CLBLM_R_X35Y120_SLICE_X53Y120_D_XOR),
.O5(CLBLM_R_X33Y116_SLICE_X48Y116_CO5),
.O6(CLBLM_R_X33Y116_SLICE_X48Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb0f4f4b000000000)
  ) CLBLM_R_X33Y116_SLICE_X48Y116_BLUT (
.I0(LIOB33_X0Y147_IOB_X0Y147_I),
.I1(LIOB33_X0Y145_IOB_X0Y146_I),
.I2(CLBLM_R_X35Y120_SLICE_X53Y120_C_XOR),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.O5(CLBLM_R_X33Y116_SLICE_X48Y116_BO5),
.O6(CLBLM_R_X33Y116_SLICE_X48Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff4ff4400000000)
  ) CLBLM_R_X33Y116_SLICE_X48Y116_ALUT (
.I0(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.I1(CLBLM_R_X35Y120_SLICE_X53Y120_C_XOR),
.I2(CLBLM_R_X35Y118_SLICE_X52Y118_C_XOR),
.I3(CLBLM_R_X33Y116_SLICE_X48Y116_BO6),
.I4(CLBLL_L_X36Y122_SLICE_X55Y122_AO6),
.I5(LIOB33_X0Y147_IOB_X0Y148_I),
.O5(CLBLM_R_X33Y116_SLICE_X48Y116_AO5),
.O6(CLBLM_R_X33Y116_SLICE_X48Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4f5f5e4e4a0a0)
  ) CLBLM_R_X33Y116_SLICE_X49Y116_DLUT (
.I0(LIOB33_X0Y145_IOB_X0Y146_I),
.I1(CLBLL_L_X34Y117_SLICE_X50Y117_CO6),
.I2(CLBLM_R_X35Y120_SLICE_X53Y120_C_XOR),
.I3(1'b1),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(CLBLL_L_X34Y117_SLICE_X50Y117_BO6),
.O5(CLBLM_R_X33Y116_SLICE_X49Y116_DO5),
.O6(CLBLM_R_X33Y116_SLICE_X49Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaff00f0f0cccc)
  ) CLBLM_R_X33Y116_SLICE_X49Y116_CLUT (
.I0(CLBLM_R_X33Y115_SLICE_X49Y115_AO6),
.I1(CLBLM_R_X33Y117_SLICE_X49Y117_AO6),
.I2(CLBLL_L_X34Y118_SLICE_X50Y118_BO6),
.I3(CLBLM_L_X32Y116_SLICE_X47Y116_AO6),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(LIOB33_X0Y145_IOB_X0Y146_I),
.O5(CLBLM_R_X33Y116_SLICE_X49Y116_CO5),
.O6(CLBLM_R_X33Y116_SLICE_X49Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hef4fe04000000000)
  ) CLBLM_R_X33Y116_SLICE_X49Y116_BLUT (
.I0(LIOB33_X0Y147_IOB_X0Y147_I),
.I1(CLBLM_R_X33Y116_SLICE_X49Y116_CO6),
.I2(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I3(CLBLM_R_X33Y116_SLICE_X49Y116_DO6),
.I4(CLBLM_R_X35Y120_SLICE_X53Y120_C_XOR),
.I5(CLBLL_L_X34Y128_SLICE_X50Y128_AO6),
.O5(CLBLM_R_X33Y116_SLICE_X49Y116_BO5),
.O6(CLBLM_R_X33Y116_SLICE_X49Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffafff8fff8fff0)
  ) CLBLM_R_X33Y116_SLICE_X49Y116_ALUT (
.I0(CLBLL_L_X36Y116_SLICE_X55Y116_AO5),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(CLBLM_R_X33Y116_SLICE_X48Y116_AO6),
.I3(CLBLM_R_X33Y116_SLICE_X49Y116_BO6),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.O5(CLBLM_R_X33Y116_SLICE_X49Y116_AO5),
.O6(CLBLM_R_X33Y116_SLICE_X49Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3300b8b800000000)
  ) CLBLM_R_X33Y117_SLICE_X48Y117_DLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(CLBLL_L_X36Y121_SLICE_X54Y121_AO5),
.O5(CLBLM_R_X33Y117_SLICE_X48Y117_DO5),
.O6(CLBLM_R_X33Y117_SLICE_X48Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hefeae5e04f4a4540)
  ) CLBLM_R_X33Y117_SLICE_X48Y117_CLUT (
.I0(LIOB33_X0Y145_IOB_X0Y146_I),
.I1(CLBLL_L_X34Y118_SLICE_X50Y118_CO6),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(CLBLM_R_X33Y117_SLICE_X49Y117_BO6),
.I4(CLBLM_R_X33Y117_SLICE_X48Y117_DO6),
.I5(CLBLM_L_X32Y117_SLICE_X47Y117_AO6),
.O5(CLBLM_R_X33Y117_SLICE_X48Y117_CO5),
.O6(CLBLM_R_X33Y117_SLICE_X48Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdf85d58ada80d08)
  ) CLBLM_R_X33Y117_SLICE_X48Y117_BLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(CLBLM_R_X33Y117_SLICE_X49Y117_BO6),
.I2(LIOB33_X0Y145_IOB_X0Y146_I),
.I3(CLBLL_L_X34Y118_SLICE_X50Y118_BO6),
.I4(CLBLM_L_X32Y116_SLICE_X47Y116_AO6),
.I5(CLBLM_L_X32Y117_SLICE_X47Y117_AO6),
.O5(CLBLM_R_X33Y117_SLICE_X48Y117_BO5),
.O6(CLBLM_R_X33Y117_SLICE_X48Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffd855d8aad800d8)
  ) CLBLM_R_X33Y117_SLICE_X48Y117_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(LIOB33_X0Y117_IOB_X0Y118_I),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(RIOB33_X105Y103_IOB_X1Y104_I),
.O5(CLBLM_R_X33Y117_SLICE_X48Y117_AO5),
.O6(CLBLM_R_X33Y117_SLICE_X48Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0c0c0cfafa0a0a)
  ) CLBLM_R_X33Y117_SLICE_X49Y117_DLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(1'b1),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(LIOB33_X0Y117_IOB_X0Y118_I),
.O5(CLBLM_R_X33Y117_SLICE_X49Y117_DO5),
.O6(CLBLM_R_X33Y117_SLICE_X49Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4ffaae4e45500)
  ) CLBLM_R_X33Y117_SLICE_X49Y117_CLUT (
.I0(LIOB33_X0Y145_IOB_X0Y146_I),
.I1(CLBLM_R_X33Y118_SLICE_X49Y118_CO6),
.I2(CLBLM_R_X33Y117_SLICE_X48Y117_DO6),
.I3(CLBLL_L_X34Y118_SLICE_X50Y118_CO6),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(CLBLM_R_X33Y119_SLICE_X49Y119_BO6),
.O5(CLBLM_R_X33Y117_SLICE_X49Y117_CO5),
.O6(CLBLM_R_X33Y117_SLICE_X49Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafcfa0c0afc0a0c)
  ) CLBLM_R_X33Y117_SLICE_X49Y117_BLUT (
.I0(CLBLM_R_X33Y117_SLICE_X49Y117_DO6),
.I1(CLBLL_L_X34Y114_SLICE_X51Y114_CO6),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(CLBLL_L_X34Y117_SLICE_X51Y117_BO6),
.I5(CLBLM_R_X33Y118_SLICE_X48Y118_DO6),
.O5(CLBLM_R_X33Y117_SLICE_X49Y117_BO5),
.O6(CLBLM_R_X33Y117_SLICE_X49Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaaccfff000f0)
  ) CLBLM_R_X33Y117_SLICE_X49Y117_ALUT (
.I0(CLBLM_R_X33Y117_SLICE_X49Y117_DO6),
.I1(CLBLL_L_X34Y114_SLICE_X51Y114_CO6),
.I2(CLBLM_R_X33Y117_SLICE_X48Y117_AO6),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(CLBLL_L_X34Y117_SLICE_X51Y117_BO6),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLM_R_X33Y117_SLICE_X49Y117_AO5),
.O6(CLBLM_R_X33Y117_SLICE_X49Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0000afa0afa0)
  ) CLBLM_R_X33Y118_SLICE_X48Y118_DLUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(1'b1),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(LIOB33_X0Y117_IOB_X0Y118_I),
.O5(CLBLM_R_X33Y118_SLICE_X48Y118_DO5),
.O6(CLBLM_R_X33Y118_SLICE_X48Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5ff000a4f4f4040)
  ) CLBLM_R_X33Y118_SLICE_X48Y118_CLUT (
.I0(LIOB33_X0Y145_IOB_X0Y146_I),
.I1(CLBLM_R_X35Y118_SLICE_X52Y118_C_XOR),
.I2(LIOB33_X0Y147_IOB_X0Y147_I),
.I3(CLBLM_R_X33Y118_SLICE_X48Y118_AO5),
.I4(CLBLM_R_X35Y120_SLICE_X53Y120_C_XOR),
.I5(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.O5(CLBLM_R_X33Y118_SLICE_X48Y118_CO5),
.O6(CLBLM_R_X33Y118_SLICE_X48Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8fcf80c08f0f8000)
  ) CLBLM_R_X33Y118_SLICE_X48Y118_BLUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(CLBLL_L_X36Y121_SLICE_X54Y121_AO5),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(CLBLM_R_X33Y118_SLICE_X48Y118_AO6),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_R_X33Y118_SLICE_X48Y118_BO5),
.O6(CLBLM_R_X33Y118_SLICE_X48Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h10101100f0f00f0f)
  ) CLBLM_R_X33Y118_SLICE_X48Y118_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(LIOB33_X0Y117_IOB_X0Y118_I),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(1'b1),
.O5(CLBLM_R_X33Y118_SLICE_X48Y118_AO5),
.O6(CLBLM_R_X33Y118_SLICE_X48Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88f5f5dd88a0a0)
  ) CLBLM_R_X33Y118_SLICE_X49Y118_DLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(CLBLL_L_X36Y116_SLICE_X55Y116_BO6),
.I2(CLBLM_R_X33Y118_SLICE_X48Y118_DO6),
.I3(CLBLL_L_X34Y117_SLICE_X51Y117_DO6),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(CLBLM_R_X33Y117_SLICE_X49Y117_DO6),
.O5(CLBLM_R_X33Y118_SLICE_X49Y118_DO5),
.O6(CLBLM_R_X33Y118_SLICE_X49Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50eeeefa504444)
  ) CLBLM_R_X33Y118_SLICE_X49Y118_CLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(CLBLL_L_X34Y117_SLICE_X51Y117_BO6),
.I2(CLBLM_R_X33Y118_SLICE_X48Y118_DO6),
.I3(CLBLL_L_X34Y117_SLICE_X51Y117_DO6),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(CLBLM_R_X33Y117_SLICE_X49Y117_DO6),
.O5(CLBLM_R_X33Y118_SLICE_X49Y118_CO5),
.O6(CLBLM_R_X33Y118_SLICE_X49Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0acfcffa0ac0c0)
  ) CLBLM_R_X33Y118_SLICE_X49Y118_BLUT (
.I0(CLBLL_L_X34Y117_SLICE_X51Y117_DO6),
.I1(CLBLL_L_X36Y116_SLICE_X55Y116_BO6),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(CLBLM_R_X37Y118_SLICE_X57Y118_AO6),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(CLBLM_R_X33Y118_SLICE_X48Y118_DO6),
.O5(CLBLM_R_X33Y118_SLICE_X49Y118_BO5),
.O6(CLBLM_R_X33Y118_SLICE_X49Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5dda0ddf588a088)
  ) CLBLM_R_X33Y118_SLICE_X49Y118_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(RIOB33_X105Y117_IOB_X1Y117_I),
.I3(LIOB33_X0Y117_IOB_X0Y118_I),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_R_X33Y118_SLICE_X49Y118_AO5),
.O6(CLBLM_R_X33Y118_SLICE_X49Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X33Y119_SLICE_X48Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X33Y119_SLICE_X48Y119_DO5),
.O6(CLBLM_R_X33Y119_SLICE_X48Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X33Y119_SLICE_X48Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X33Y119_SLICE_X48Y119_CO5),
.O6(CLBLM_R_X33Y119_SLICE_X48Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X33Y119_SLICE_X48Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X33Y119_SLICE_X48Y119_BO5),
.O6(CLBLM_R_X33Y119_SLICE_X48Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X33Y119_SLICE_X48Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X33Y119_SLICE_X48Y119_AO5),
.O6(CLBLM_R_X33Y119_SLICE_X48Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X33Y119_SLICE_X49Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X33Y119_SLICE_X49Y119_DO5),
.O6(CLBLM_R_X33Y119_SLICE_X49Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafaee445050ee44)
  ) CLBLM_R_X33Y119_SLICE_X49Y119_CLUT (
.I0(LIOB33_X0Y145_IOB_X0Y146_I),
.I1(CLBLL_L_X34Y119_SLICE_X50Y119_CO6),
.I2(CLBLM_R_X33Y118_SLICE_X49Y118_DO6),
.I3(CLBLL_L_X34Y119_SLICE_X51Y119_DO6),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(CLBLM_R_X33Y118_SLICE_X48Y118_BO6),
.O5(CLBLM_R_X33Y119_SLICE_X49Y119_CO5),
.O6(CLBLM_R_X33Y119_SLICE_X49Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7300510062004000)
  ) CLBLM_R_X33Y119_SLICE_X49Y119_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(CLBLL_L_X36Y121_SLICE_X54Y121_AO5),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLM_R_X33Y119_SLICE_X49Y119_BO5),
.O6(CLBLM_R_X33Y119_SLICE_X49Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0cfcfafa0c0c0)
  ) CLBLM_R_X33Y119_SLICE_X49Y119_ALUT (
.I0(CLBLM_R_X33Y119_SLICE_X49Y119_BO6),
.I1(CLBLL_L_X34Y119_SLICE_X50Y119_CO6),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(CLBLM_R_X33Y118_SLICE_X48Y118_BO6),
.I4(LIOB33_X0Y145_IOB_X0Y146_I),
.I5(CLBLM_R_X33Y118_SLICE_X49Y118_CO6),
.O5(CLBLM_R_X33Y119_SLICE_X49Y119_AO5),
.O6(CLBLM_R_X33Y119_SLICE_X49Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc48cccc00480000)
  ) CLBLM_R_X33Y121_SLICE_X48Y121_DLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I2(LIOB33_X0Y121_IOB_X0Y122_I),
.I3(LIOB33_X0Y147_IOB_X0Y147_I),
.I4(LIOB33_X0Y145_IOB_X0Y146_I),
.I5(CLBLM_R_X35Y122_SLICE_X53Y122_A_XOR),
.O5(CLBLM_R_X33Y121_SLICE_X48Y121_DO5),
.O6(CLBLM_R_X33Y121_SLICE_X48Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he0e0e04040e04040)
  ) CLBLM_R_X33Y121_SLICE_X48Y121_CLUT (
.I0(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I1(CLBLM_R_X35Y122_SLICE_X53Y122_A_XOR),
.I2(CLBLL_L_X34Y128_SLICE_X50Y128_AO6),
.I3(LIOB33_X0Y147_IOB_X0Y147_I),
.I4(CLBLM_R_X33Y121_SLICE_X49Y121_AO6),
.I5(CLBLL_L_X34Y121_SLICE_X50Y121_CO6),
.O5(CLBLM_R_X33Y121_SLICE_X48Y121_CO5),
.O6(CLBLM_R_X33Y121_SLICE_X48Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc80cccccc80cc80)
  ) CLBLM_R_X33Y121_SLICE_X48Y121_BLUT (
.I0(CLBLL_L_X36Y122_SLICE_X55Y122_AO6),
.I1(LIOB33_X0Y147_IOB_X0Y148_I),
.I2(CLBLM_R_X35Y120_SLICE_X52Y120_A_XOR),
.I3(CLBLM_R_X33Y121_SLICE_X48Y121_DO6),
.I4(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.I5(CLBLM_R_X35Y122_SLICE_X53Y122_A_XOR),
.O5(CLBLM_R_X33Y121_SLICE_X48Y121_BO5),
.O6(CLBLM_R_X33Y121_SLICE_X48Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffc8ff80)
  ) CLBLM_R_X33Y121_SLICE_X48Y121_ALUT (
.I0(LIOB33_X0Y121_IOB_X0Y122_I),
.I1(CLBLL_L_X36Y116_SLICE_X55Y116_AO5),
.I2(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I3(CLBLM_R_X33Y121_SLICE_X48Y121_BO6),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(CLBLM_R_X33Y121_SLICE_X48Y121_CO6),
.O5(CLBLM_R_X33Y121_SLICE_X48Y121_AO5),
.O6(CLBLM_R_X33Y121_SLICE_X48Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X33Y121_SLICE_X49Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X33Y121_SLICE_X49Y121_DO5),
.O6(CLBLM_R_X33Y121_SLICE_X49Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0000fa0afa0a)
  ) CLBLM_R_X33Y121_SLICE_X49Y121_CLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(1'b1),
.I2(LIOB33_X0Y117_IOB_X0Y118_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X33Y121_SLICE_X49Y121_CO5),
.O6(CLBLM_R_X33Y121_SLICE_X49Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0ff008888ff00)
  ) CLBLM_R_X33Y121_SLICE_X49Y121_BLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLL_L_X36Y121_SLICE_X54Y121_AO5),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(CLBLM_R_X33Y122_SLICE_X49Y122_CO6),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLM_R_X33Y121_SLICE_X49Y121_BO5),
.O6(CLBLM_R_X33Y121_SLICE_X49Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff00f00cacacaca)
  ) CLBLM_R_X33Y121_SLICE_X49Y121_ALUT (
.I0(CLBLM_R_X33Y118_SLICE_X49Y118_DO6),
.I1(CLBLL_L_X34Y120_SLICE_X50Y120_CO6),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(CLBLM_R_X33Y121_SLICE_X49Y121_BO6),
.I4(CLBLL_L_X34Y119_SLICE_X51Y119_DO6),
.I5(LIOB33_X0Y145_IOB_X0Y146_I),
.O5(CLBLM_R_X33Y121_SLICE_X49Y121_AO5),
.O6(CLBLM_R_X33Y121_SLICE_X49Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X33Y122_SLICE_X48Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X33Y122_SLICE_X48Y122_DO5),
.O6(CLBLM_R_X33Y122_SLICE_X48Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X33Y122_SLICE_X48Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X33Y122_SLICE_X48Y122_CO5),
.O6(CLBLM_R_X33Y122_SLICE_X48Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00f0f0ccccaaaa)
  ) CLBLM_R_X33Y122_SLICE_X48Y122_BLUT (
.I0(CLBLM_R_X33Y125_SLICE_X49Y125_BO5),
.I1(CLBLM_R_X33Y122_SLICE_X48Y122_AO5),
.I2(CLBLM_L_X32Y123_SLICE_X47Y123_AO5),
.I3(CLBLL_L_X34Y123_SLICE_X50Y123_BO6),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLM_R_X33Y122_SLICE_X48Y122_BO5),
.O6(CLBLM_R_X33Y122_SLICE_X48Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cf00c00cfa0c0a)
  ) CLBLM_R_X33Y122_SLICE_X48Y122_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(LIOB33_X0Y117_IOB_X0Y118_I),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(1'b1),
.O5(CLBLM_R_X33Y122_SLICE_X48Y122_AO5),
.O6(CLBLM_R_X33Y122_SLICE_X48Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffdd880000dd88)
  ) CLBLM_R_X33Y122_SLICE_X49Y122_DLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(CLBLM_R_X35Y117_SLICE_X52Y117_BO6),
.I2(1'b1),
.I3(CLBLL_L_X34Y118_SLICE_X50Y118_AO6),
.I4(LIOB33_X0Y145_IOB_X0Y146_I),
.I5(CLBLM_R_X35Y122_SLICE_X53Y122_C_XOR),
.O5(CLBLM_R_X33Y122_SLICE_X49Y122_DO5),
.O6(CLBLM_R_X33Y122_SLICE_X49Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000022f3000022c0)
  ) CLBLM_R_X33Y122_SLICE_X49Y122_CLUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y117_IOB_X0Y118_I),
.I5(LIOB33_X0Y107_IOB_X0Y108_I),
.O5(CLBLM_R_X33Y122_SLICE_X49Y122_CO5),
.O6(CLBLM_R_X33Y122_SLICE_X49Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd558800f555a000)
  ) CLBLM_R_X33Y122_SLICE_X49Y122_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(CLBLL_L_X36Y121_SLICE_X54Y121_AO5),
.I4(CLBLM_R_X33Y123_SLICE_X48Y123_AO6),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLM_R_X33Y122_SLICE_X49Y122_BO5),
.O6(CLBLM_R_X33Y122_SLICE_X49Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc840c840cccc0000)
  ) CLBLM_R_X33Y122_SLICE_X49Y122_ALUT (
.I0(LIOB33_X0Y147_IOB_X0Y147_I),
.I1(CLBLL_L_X34Y128_SLICE_X50Y128_AO6),
.I2(CLBLL_L_X34Y122_SLICE_X50Y122_AO6),
.I3(CLBLM_R_X33Y122_SLICE_X49Y122_DO6),
.I4(CLBLM_R_X35Y122_SLICE_X53Y122_C_XOR),
.I5(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.O5(CLBLM_R_X33Y122_SLICE_X49Y122_AO5),
.O6(CLBLM_R_X33Y122_SLICE_X49Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfd75b931ec64a820)
  ) CLBLM_R_X33Y123_SLICE_X48Y123_DLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(CLBLM_R_X33Y125_SLICE_X49Y125_AO5),
.I3(CLBLM_R_X33Y124_SLICE_X49Y124_AO6),
.I4(CLBLM_R_X33Y124_SLICE_X48Y124_AO5),
.I5(CLBLL_L_X34Y123_SLICE_X50Y123_AO5),
.O5(CLBLM_R_X33Y123_SLICE_X48Y123_DO5),
.O6(CLBLM_R_X33Y123_SLICE_X48Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffd855d8aad800d8)
  ) CLBLM_R_X33Y123_SLICE_X48Y123_CLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(CLBLM_R_X33Y124_SLICE_X48Y124_AO5),
.I2(CLBLM_R_X33Y125_SLICE_X49Y125_AO5),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(CLBLL_L_X34Y123_SLICE_X50Y123_AO6),
.I5(CLBLM_R_X33Y124_SLICE_X49Y124_AO6),
.O5(CLBLM_R_X33Y123_SLICE_X48Y123_CO5),
.O6(CLBLM_R_X33Y123_SLICE_X48Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hefe32f23ece02c20)
  ) CLBLM_R_X33Y123_SLICE_X48Y123_BLUT (
.I0(CLBLL_L_X34Y123_SLICE_X50Y123_AO6),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(CLBLM_R_X33Y124_SLICE_X49Y124_AO6),
.I4(CLBLM_R_X33Y125_SLICE_X49Y125_AO6),
.I5(CLBLM_R_X33Y124_SLICE_X48Y124_AO5),
.O5(CLBLM_R_X33Y123_SLICE_X48Y123_BO5),
.O6(CLBLM_R_X33Y123_SLICE_X48Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h030e000e03020002)
  ) CLBLM_R_X33Y123_SLICE_X48Y123_ALUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(LIOB33_X0Y117_IOB_X0Y118_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLM_R_X33Y123_SLICE_X48Y123_AO5),
.O6(CLBLM_R_X33Y123_SLICE_X48Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffe2e20000e2e2)
  ) CLBLM_R_X33Y123_SLICE_X49Y123_DLUT (
.I0(CLBLM_R_X33Y125_SLICE_X49Y125_AO6),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(CLBLM_R_X33Y124_SLICE_X49Y124_AO5),
.I3(1'b1),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(CLBLM_L_X32Y123_SLICE_X46Y123_AO6),
.O5(CLBLM_R_X33Y123_SLICE_X49Y123_DO5),
.O6(CLBLM_R_X33Y123_SLICE_X49Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdf00ef0010002000)
  ) CLBLM_R_X33Y123_SLICE_X49Y123_CLUT (
.I0(LIOB33_X0Y123_IOB_X0Y124_I),
.I1(LIOB33_X0Y147_IOB_X0Y147_I),
.I2(LIOB33_X0Y145_IOB_X0Y146_I),
.I3(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(CLBLM_R_X35Y122_SLICE_X53Y122_C_XOR),
.O5(CLBLM_R_X33Y123_SLICE_X49Y123_CO5),
.O6(CLBLM_R_X33Y123_SLICE_X49Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000dc500000)
  ) CLBLM_R_X33Y123_SLICE_X49Y123_BLUT (
.I0(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.I1(CLBLL_L_X36Y122_SLICE_X55Y122_AO6),
.I2(CLBLM_R_X35Y122_SLICE_X53Y122_C_XOR),
.I3(CLBLM_R_X35Y120_SLICE_X52Y120_C_XOR),
.I4(LIOB33_X0Y147_IOB_X0Y148_I),
.I5(CLBLM_R_X33Y123_SLICE_X49Y123_CO6),
.O5(CLBLM_R_X33Y123_SLICE_X49Y123_BO5),
.O6(CLBLM_R_X33Y123_SLICE_X49Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffa8ffffff80)
  ) CLBLM_R_X33Y123_SLICE_X49Y123_ALUT (
.I0(CLBLL_L_X36Y116_SLICE_X55Y116_AO5),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(LIOB33_X0Y123_IOB_X0Y124_I),
.I3(CLBLM_R_X33Y123_SLICE_X49Y123_BO6),
.I4(CLBLM_R_X33Y122_SLICE_X49Y122_AO6),
.I5(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.O5(CLBLM_R_X33Y123_SLICE_X49Y123_AO5),
.O6(CLBLM_R_X33Y123_SLICE_X49Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X33Y124_SLICE_X48Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X33Y124_SLICE_X48Y124_DO5),
.O6(CLBLM_R_X33Y124_SLICE_X48Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X33Y124_SLICE_X48Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X33Y124_SLICE_X48Y124_CO5),
.O6(CLBLM_R_X33Y124_SLICE_X48Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0afcfcfa0a0c0c)
  ) CLBLM_R_X33Y124_SLICE_X48Y124_BLUT (
.I0(CLBLM_R_X33Y125_SLICE_X49Y125_BO5),
.I1(CLBLL_L_X34Y123_SLICE_X50Y123_BO5),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(CLBLM_L_X32Y123_SLICE_X47Y123_AO5),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(CLBLM_R_X33Y122_SLICE_X48Y122_AO5),
.O5(CLBLM_R_X33Y124_SLICE_X48Y124_BO5),
.O6(CLBLM_R_X33Y124_SLICE_X48Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0c03003e320e02)
  ) CLBLM_R_X33Y124_SLICE_X48Y124_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_X0Y117_IOB_X0Y118_I),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(1'b1),
.O5(CLBLM_R_X33Y124_SLICE_X48Y124_AO5),
.O6(CLBLM_R_X33Y124_SLICE_X48Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaccf000aaccf0)
  ) CLBLM_R_X33Y124_SLICE_X49Y124_DLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y117_IOB_X0Y118_I),
.I5(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.O5(CLBLM_R_X33Y124_SLICE_X49Y124_DO5),
.O6(CLBLM_R_X33Y124_SLICE_X49Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc00ccf0aaf0aa)
  ) CLBLM_R_X33Y124_SLICE_X49Y124_CLUT (
.I0(CLBLM_R_X33Y124_SLICE_X49Y124_AO6),
.I1(CLBLM_R_X33Y125_SLICE_X49Y125_AO6),
.I2(CLBLL_L_X34Y123_SLICE_X50Y123_AO6),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(CLBLM_R_X33Y124_SLICE_X48Y124_AO6),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLM_R_X33Y124_SLICE_X49Y124_CO5),
.O6(CLBLM_R_X33Y124_SLICE_X49Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfafc0a0cfa0c0a)
  ) CLBLM_R_X33Y124_SLICE_X49Y124_BLUT (
.I0(CLBLL_L_X34Y123_SLICE_X50Y123_AO6),
.I1(CLBLM_R_X33Y124_SLICE_X48Y124_AO6),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(CLBLM_R_X33Y125_SLICE_X49Y125_AO6),
.I5(CLBLM_R_X33Y124_SLICE_X49Y124_AO5),
.O5(CLBLM_R_X33Y124_SLICE_X49Y124_BO5),
.O6(CLBLM_R_X33Y124_SLICE_X49Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5050ee440000f5a0)
  ) CLBLM_R_X33Y124_SLICE_X49Y124_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(LIOB33_X0Y117_IOB_X0Y118_I),
.I5(1'b1),
.O5(CLBLM_R_X33Y124_SLICE_X49Y124_AO5),
.O6(CLBLM_R_X33Y124_SLICE_X49Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X33Y125_SLICE_X48Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X33Y125_SLICE_X48Y125_DO5),
.O6(CLBLM_R_X33Y125_SLICE_X48Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X33Y125_SLICE_X48Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X33Y125_SLICE_X48Y125_CO5),
.O6(CLBLM_R_X33Y125_SLICE_X48Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X33Y125_SLICE_X48Y125_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X33Y125_SLICE_X48Y125_BO5),
.O6(CLBLM_R_X33Y125_SLICE_X48Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X33Y125_SLICE_X48Y125_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X33Y125_SLICE_X48Y125_AO5),
.O6(CLBLM_R_X33Y125_SLICE_X48Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7e6b3a2d5c49180)
  ) CLBLM_R_X33Y125_SLICE_X49Y125_DLUT (
.I0(LIOB33_X0Y117_IOB_X0Y118_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_R_X33Y125_SLICE_X49Y125_DO5),
.O6(CLBLM_R_X33Y125_SLICE_X49Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b8b8b8ff33cc00)
  ) CLBLM_R_X33Y125_SLICE_X49Y125_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(LIOB33_X0Y117_IOB_X0Y118_I),
.O5(CLBLM_R_X33Y125_SLICE_X49Y125_CO5),
.O6(CLBLM_R_X33Y125_SLICE_X49Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000f3c03030ee22)
  ) CLBLM_R_X33Y125_SLICE_X49Y125_BLUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(LIOB33_X0Y113_IOB_X0Y113_I),
.I4(LIOB33_X0Y117_IOB_X0Y118_I),
.I5(1'b1),
.O5(CLBLM_R_X33Y125_SLICE_X49Y125_BO5),
.O6(CLBLM_R_X33Y125_SLICE_X49Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00bb008822fc2230)
  ) CLBLM_R_X33Y125_SLICE_X49Y125_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(LIOB33_X0Y117_IOB_X0Y118_I),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(1'b1),
.O5(CLBLM_R_X33Y125_SLICE_X49Y125_AO5),
.O6(CLBLM_R_X33Y125_SLICE_X49Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X35Y114_SLICE_X52Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y114_SLICE_X52Y114_DO5),
.O6(CLBLM_R_X35Y114_SLICE_X52Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X35Y114_SLICE_X52Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y114_SLICE_X52Y114_CO5),
.O6(CLBLM_R_X35Y114_SLICE_X52Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X35Y114_SLICE_X52Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y114_SLICE_X52Y114_BO5),
.O6(CLBLM_R_X35Y114_SLICE_X52Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a5a5a5a5a5a5a5)
  ) CLBLM_R_X35Y114_SLICE_X52Y114_ALUT (
.I0(LIOB33_X0Y119_IOB_X0Y119_I),
.I1(1'b1),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y114_SLICE_X52Y114_AO5),
.O6(CLBLM_R_X35Y114_SLICE_X52Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X35Y114_SLICE_X53Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y114_SLICE_X53Y114_DO5),
.O6(CLBLM_R_X35Y114_SLICE_X53Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X35Y114_SLICE_X53Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y114_SLICE_X53Y114_CO5),
.O6(CLBLM_R_X35Y114_SLICE_X53Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X35Y114_SLICE_X53Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y114_SLICE_X53Y114_BO5),
.O6(CLBLM_R_X35Y114_SLICE_X53Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X35Y114_SLICE_X53Y114_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y114_SLICE_X53Y114_AO5),
.O6(CLBLM_R_X35Y114_SLICE_X53Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0f3e2c0c0e2c0)
  ) CLBLM_R_X35Y115_SLICE_X52Y115_DLUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(LIOB33_X0Y147_IOB_X0Y148_I),
.I2(CLBLM_R_X35Y116_SLICE_X52Y116_DO6),
.I3(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I4(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.I5(LIOB33_X0Y119_IOB_X0Y119_I),
.O5(CLBLM_R_X35Y115_SLICE_X52Y115_DO5),
.O6(CLBLM_R_X35Y115_SLICE_X52Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000ee000000ef)
  ) CLBLM_R_X35Y115_SLICE_X52Y115_CLUT (
.I0(CLBLL_L_X34Y115_SLICE_X51Y115_CO6),
.I1(CLBLL_L_X34Y115_SLICE_X50Y115_BO6),
.I2(CLBLM_R_X35Y115_SLICE_X53Y115_DO6),
.I3(CLBLL_L_X34Y116_SLICE_X51Y116_CO6),
.I4(CLBLM_R_X35Y115_SLICE_X52Y115_DO6),
.I5(CLBLM_R_X33Y116_SLICE_X48Y116_CO6),
.O5(CLBLM_R_X35Y115_SLICE_X52Y115_CO5),
.O6(CLBLM_R_X35Y115_SLICE_X52Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffafff8fff8fff0)
  ) CLBLM_R_X35Y115_SLICE_X52Y115_BLUT (
.I0(CLBLL_L_X36Y116_SLICE_X55Y116_AO5),
.I1(LIOB33_X0Y117_IOB_X0Y118_I),
.I2(CLBLL_L_X34Y115_SLICE_X51Y115_BO6),
.I3(CLBLL_L_X34Y115_SLICE_X50Y115_BO6),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.O5(CLBLM_R_X35Y115_SLICE_X52Y115_BO5),
.O6(CLBLM_R_X35Y115_SLICE_X52Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000aaaaf072f0d8)
  ) CLBLM_R_X35Y115_SLICE_X52Y115_ALUT (
.I0(LIOB33_X0Y145_IOB_X0Y146_I),
.I1(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I2(CLBLM_R_X35Y120_SLICE_X53Y120_A_XOR),
.I3(LIOB33_X0Y147_IOB_X0Y147_I),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(1'b1),
.O5(CLBLM_R_X35Y115_SLICE_X52Y115_AO5),
.O6(CLBLM_R_X35Y115_SLICE_X52Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0f0acccc0a00)
  ) CLBLM_R_X35Y115_SLICE_X53Y115_DLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(CLBLM_R_X35Y116_SLICE_X53Y116_CO6),
.I2(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.I3(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I4(LIOB33_X0Y147_IOB_X0Y148_I),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X35Y115_SLICE_X53Y115_DO5),
.O6(CLBLM_R_X35Y115_SLICE_X53Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdf001000ef002000)
  ) CLBLM_R_X35Y115_SLICE_X53Y115_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(LIOB33_X0Y147_IOB_X0Y147_I),
.I2(LIOB33_X0Y145_IOB_X0Y146_I),
.I3(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I4(CLBLM_R_X35Y120_SLICE_X53Y120_D_XOR),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X35Y115_SLICE_X53Y115_CO5),
.O6(CLBLM_R_X35Y115_SLICE_X53Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffce0a00000000)
  ) CLBLM_R_X35Y115_SLICE_X53Y115_BLUT (
.I0(CLBLM_R_X35Y120_SLICE_X53Y120_D_XOR),
.I1(CLBLM_R_X35Y118_SLICE_X52Y118_D_XOR),
.I2(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.I3(CLBLL_L_X36Y122_SLICE_X55Y122_AO6),
.I4(CLBLM_R_X35Y115_SLICE_X53Y115_CO6),
.I5(LIOB33_X0Y147_IOB_X0Y148_I),
.O5(CLBLM_R_X35Y115_SLICE_X53Y115_BO5),
.O6(CLBLM_R_X35Y115_SLICE_X53Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffeffccffecffcc)
  ) CLBLM_R_X35Y115_SLICE_X53Y115_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_R_X33Y116_SLICE_X48Y116_CO6),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(CLBLM_R_X35Y115_SLICE_X53Y115_BO6),
.I4(CLBLL_L_X36Y116_SLICE_X55Y116_AO5),
.I5(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.O5(CLBLM_R_X35Y115_SLICE_X53Y115_AO5),
.O6(CLBLM_R_X35Y115_SLICE_X53Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd11ff003300f3c0)
  ) CLBLM_R_X35Y116_SLICE_X52Y116_DLUT (
.I0(CLBLM_R_X35Y114_SLICE_X52Y114_AO6),
.I1(LIOB33_X0Y147_IOB_X0Y147_I),
.I2(CLBLM_R_X35Y119_SLICE_X52Y119_B_XOR),
.I3(CLBLM_R_X35Y121_SLICE_X53Y121_B_XOR),
.I4(LIOB33_X0Y145_IOB_X0Y146_I),
.I5(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.O5(CLBLM_R_X35Y116_SLICE_X52Y116_DO5),
.O6(CLBLM_R_X35Y116_SLICE_X52Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hde12ff0000000000)
  ) CLBLM_R_X35Y116_SLICE_X52Y116_CLUT (
.I0(LIOB33_X0Y119_IOB_X0Y119_I),
.I1(LIOB33_X0Y147_IOB_X0Y147_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(CLBLM_R_X35Y121_SLICE_X53Y121_B_XOR),
.I4(LIOB33_X0Y145_IOB_X0Y146_I),
.I5(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.O5(CLBLM_R_X35Y116_SLICE_X52Y116_CO5),
.O6(CLBLM_R_X35Y116_SLICE_X52Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00ae000c00)
  ) CLBLM_R_X35Y116_SLICE_X52Y116_BLUT (
.I0(CLBLM_R_X35Y119_SLICE_X52Y119_B_XOR),
.I1(CLBLM_R_X35Y121_SLICE_X53Y121_B_XOR),
.I2(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(CLBLL_L_X36Y122_SLICE_X55Y122_AO6),
.I5(CLBLM_R_X35Y116_SLICE_X52Y116_CO6),
.O5(CLBLM_R_X35Y116_SLICE_X52Y116_BO5),
.O6(CLBLM_R_X35Y116_SLICE_X52Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccccccc8000)
  ) CLBLM_R_X35Y116_SLICE_X52Y116_ALUT (
.I0(CLBLL_L_X36Y116_SLICE_X54Y116_BO5),
.I1(CLBLL_L_X36Y122_SLICE_X55Y122_AO5),
.I2(CLBLM_R_X35Y115_SLICE_X52Y115_AO6),
.I3(CLBLM_R_X33Y115_SLICE_X49Y115_AO5),
.I4(CLBLL_L_X34Y116_SLICE_X51Y116_BO6),
.I5(CLBLL_L_X34Y116_SLICE_X50Y116_DO6),
.O5(CLBLM_R_X35Y116_SLICE_X52Y116_AO5),
.O6(CLBLM_R_X35Y116_SLICE_X52Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000008)
  ) CLBLM_R_X35Y116_SLICE_X53Y116_DLUT (
.I0(CLBLM_R_X35Y115_SLICE_X52Y115_CO6),
.I1(CLBLM_R_X33Y115_SLICE_X49Y115_BO6),
.I2(CLBLL_L_X34Y120_SLICE_X51Y120_AO6),
.I3(CLBLM_R_X35Y117_SLICE_X53Y117_CO6),
.I4(CLBLL_L_X34Y115_SLICE_X51Y115_AO6),
.I5(CLBLM_R_X35Y116_SLICE_X53Y116_BO6),
.O5(CLBLM_R_X35Y116_SLICE_X53Y116_DO5),
.O6(CLBLM_R_X35Y116_SLICE_X53Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haf5dff5d00085008)
  ) CLBLM_R_X35Y116_SLICE_X53Y116_CLUT (
.I0(LIOB33_X0Y147_IOB_X0Y147_I),
.I1(CLBLM_R_X35Y118_SLICE_X52Y118_D_XOR),
.I2(LIOB33_X0Y145_IOB_X0Y146_I),
.I3(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I4(CLBLM_R_X35Y118_SLICE_X53Y118_BO5),
.I5(CLBLM_R_X35Y120_SLICE_X53Y120_D_XOR),
.O5(CLBLM_R_X35Y116_SLICE_X53Y116_CO5),
.O6(CLBLM_R_X35Y116_SLICE_X53Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffeeecffffeccc)
  ) CLBLM_R_X35Y116_SLICE_X53Y116_BLUT (
.I0(CLBLL_L_X36Y116_SLICE_X55Y116_AO5),
.I1(CLBLM_R_X35Y116_SLICE_X52Y116_BO6),
.I2(LIOB33_X0Y119_IOB_X0Y119_I),
.I3(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I4(CLBLL_L_X34Y116_SLICE_X51Y116_CO6),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLM_R_X35Y116_SLICE_X53Y116_BO5),
.O6(CLBLM_R_X35Y116_SLICE_X53Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd8888fa50fa50)
  ) CLBLM_R_X35Y116_SLICE_X53Y116_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y118_I),
.I1(RIOB33_X105Y117_IOB_X1Y117_I),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X35Y116_SLICE_X53Y116_AO5),
.O6(CLBLM_R_X35Y116_SLICE_X53Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc3030bb88bb88)
  ) CLBLM_R_X35Y117_SLICE_X52Y117_DLUT (
.I0(CLBLM_R_X35Y116_SLICE_X53Y116_AO6),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(CLBLM_R_X35Y117_SLICE_X53Y117_BO6),
.I3(CLBLL_L_X34Y115_SLICE_X50Y115_DO6),
.I4(CLBLL_L_X36Y121_SLICE_X55Y121_AO5),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLM_R_X35Y117_SLICE_X52Y117_DO5),
.O6(CLBLM_R_X35Y117_SLICE_X52Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaffcc00cc)
  ) CLBLM_R_X35Y117_SLICE_X52Y117_CLUT (
.I0(CLBLM_R_X35Y116_SLICE_X53Y116_AO6),
.I1(CLBLM_R_X35Y117_SLICE_X52Y117_AO6),
.I2(CLBLM_R_X35Y117_SLICE_X53Y117_BO6),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(CLBLL_L_X34Y115_SLICE_X50Y115_DO6),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLM_R_X35Y117_SLICE_X52Y117_CO5),
.O6(CLBLM_R_X35Y117_SLICE_X52Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc00ccaaf0aaf0)
  ) CLBLM_R_X35Y117_SLICE_X52Y117_BLUT (
.I0(CLBLL_L_X36Y121_SLICE_X55Y121_AO5),
.I1(CLBLM_R_X35Y117_SLICE_X53Y117_BO6),
.I2(CLBLM_R_X35Y116_SLICE_X53Y116_AO6),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(CLBLM_R_X35Y118_SLICE_X53Y118_AO6),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLM_R_X35Y117_SLICE_X52Y117_BO5),
.O6(CLBLM_R_X35Y117_SLICE_X52Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaffcc00cc)
  ) CLBLM_R_X35Y117_SLICE_X52Y117_ALUT (
.I0(RIOB33_X105Y109_IOB_X1Y109_I),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(RIOB33_X105Y117_IOB_X1Y117_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(LIOB33_X0Y117_IOB_X0Y118_I),
.O5(CLBLM_R_X35Y117_SLICE_X52Y117_AO5),
.O6(CLBLM_R_X35Y117_SLICE_X52Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbeaeaea00000000)
  ) CLBLM_R_X35Y117_SLICE_X53Y117_DLUT (
.I0(CLBLL_L_X34Y116_SLICE_X50Y116_DO6),
.I1(LIOB33_X0Y145_IOB_X0Y146_I),
.I2(CLBLM_R_X35Y120_SLICE_X53Y120_B_XOR),
.I3(CLBLL_L_X34Y117_SLICE_X50Y117_BO6),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(CLBLL_L_X36Y116_SLICE_X55Y116_AO6),
.O5(CLBLM_R_X35Y117_SLICE_X53Y117_DO5),
.O6(CLBLM_R_X35Y117_SLICE_X53Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffcccccc40)
  ) CLBLM_R_X35Y117_SLICE_X53Y117_CLUT (
.I0(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I1(CLBLL_L_X34Y128_SLICE_X50Y128_AO6),
.I2(CLBLM_R_X35Y120_SLICE_X53Y120_B_XOR),
.I3(CLBLM_R_X35Y116_SLICE_X52Y116_AO6),
.I4(CLBLM_R_X35Y117_SLICE_X53Y117_DO6),
.I5(CLBLL_L_X36Y117_SLICE_X54Y117_CO6),
.O5(CLBLM_R_X35Y117_SLICE_X53Y117_CO5),
.O6(CLBLM_R_X35Y117_SLICE_X53Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa00aaccf0ccf0)
  ) CLBLM_R_X35Y117_SLICE_X53Y117_BLUT (
.I0(RIOB33_X105Y115_IOB_X1Y115_I),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(RIOB33_X105Y117_IOB_X1Y117_I),
.I5(LIOB33_X0Y117_IOB_X0Y118_I),
.O5(CLBLM_R_X35Y117_SLICE_X53Y117_BO5),
.O6(CLBLM_R_X35Y117_SLICE_X53Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfadd50ddfa885088)
  ) CLBLM_R_X35Y117_SLICE_X53Y117_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(CLBLL_L_X36Y116_SLICE_X55Y116_BO6),
.I2(CLBLM_R_X37Y118_SLICE_X57Y118_AO6),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(CLBLL_L_X36Y115_SLICE_X54Y115_AO5),
.I5(CLBLL_L_X34Y117_SLICE_X51Y117_DO6),
.O5(CLBLM_R_X35Y117_SLICE_X53Y117_AO5),
.O6(CLBLM_R_X35Y117_SLICE_X53Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X35Y118_SLICE_X52Y118_CARRY4 (
.CI(1'b0),
.CO({CLBLM_R_X35Y118_SLICE_X52Y118_D_CY, CLBLM_R_X35Y118_SLICE_X52Y118_C_CY, CLBLM_R_X35Y118_SLICE_X52Y118_B_CY, CLBLM_R_X35Y118_SLICE_X52Y118_A_CY}),
.CYINIT(1'b1),
.DI({LIOB33_X0Y103_IOB_X0Y103_I, LIOB33_X0Y101_IOB_X0Y102_I, LIOB33_X0Y101_IOB_X0Y101_I, LIOB33_SING_X0Y100_IOB_X0Y100_I}),
.O({CLBLM_R_X35Y118_SLICE_X52Y118_D_XOR, CLBLM_R_X35Y118_SLICE_X52Y118_C_XOR, CLBLM_R_X35Y118_SLICE_X52Y118_B_XOR, CLBLM_R_X35Y118_SLICE_X52Y118_A_XOR}),
.S({CLBLM_R_X35Y118_SLICE_X52Y118_DO6, CLBLM_R_X35Y118_SLICE_X52Y118_CO6, CLBLM_R_X35Y118_SLICE_X52Y118_BO6, CLBLM_R_X35Y118_SLICE_X52Y118_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a5a5a5a5a5a5a5)
  ) CLBLM_R_X35Y118_SLICE_X52Y118_DLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(1'b1),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y118_SLICE_X52Y118_DO5),
.O6(CLBLM_R_X35Y118_SLICE_X52Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00f0ff0f00f0f)
  ) CLBLM_R_X35Y118_SLICE_X52Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(1'b1),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(1'b1),
.O5(CLBLM_R_X35Y118_SLICE_X52Y118_CO5),
.O6(CLBLM_R_X35Y118_SLICE_X52Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc33333333)
  ) CLBLM_R_X35Y118_SLICE_X52Y118_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLM_R_X35Y118_SLICE_X52Y118_BO5),
.O6(CLBLM_R_X35Y118_SLICE_X52Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa5555aaaa5555)
  ) CLBLM_R_X35Y118_SLICE_X52Y118_ALUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(1'b1),
.O5(CLBLM_R_X35Y118_SLICE_X52Y118_AO5),
.O6(CLBLM_R_X35Y118_SLICE_X52Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfda8f8ad5d08580)
  ) CLBLM_R_X35Y118_SLICE_X53Y118_DLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(CLBLL_L_X36Y117_SLICE_X55Y117_AO5),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(CLBLM_R_X35Y118_SLICE_X53Y118_CO6),
.I4(CLBLM_R_X37Y118_SLICE_X57Y118_AO5),
.I5(CLBLL_L_X36Y115_SLICE_X54Y115_AO6),
.O5(CLBLM_R_X35Y118_SLICE_X53Y118_DO5),
.O6(CLBLM_R_X35Y118_SLICE_X53Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff00f00cacacaca)
  ) CLBLM_R_X35Y118_SLICE_X53Y118_CLUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(RIOB33_X105Y107_IOB_X1Y108_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(RIOB33_X105Y115_IOB_X1Y116_I),
.I4(RIOB33_X105Y117_IOB_X1Y117_I),
.I5(LIOB33_X0Y117_IOB_X0Y118_I),
.O5(CLBLM_R_X35Y118_SLICE_X53Y118_CO5),
.O6(CLBLM_R_X35Y118_SLICE_X53Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h10101100a5a5a5a5)
  ) CLBLM_R_X35Y118_SLICE_X53Y118_BLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(LIOB33_X0Y117_IOB_X0Y118_I),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(1'b1),
.O5(CLBLM_R_X35Y118_SLICE_X53Y118_BO5),
.O6(CLBLM_R_X35Y118_SLICE_X53Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ddf08800dd0088)
  ) CLBLM_R_X35Y118_SLICE_X53Y118_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(RIOB33_X105Y111_IOB_X1Y111_I),
.I2(RIOB33_X105Y117_IOB_X1Y117_I),
.I3(LIOB33_X0Y117_IOB_X0Y118_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(1'b1),
.O5(CLBLM_R_X35Y118_SLICE_X53Y118_AO5),
.O6(CLBLM_R_X35Y118_SLICE_X53Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X35Y119_SLICE_X52Y119_CARRY4 (
.CI(CLBLM_R_X35Y118_SLICE_X52Y118_D_CY),
.CO({CLBLM_R_X35Y119_SLICE_X52Y119_D_CY, CLBLM_R_X35Y119_SLICE_X52Y119_C_CY, CLBLM_R_X35Y119_SLICE_X52Y119_B_CY, CLBLM_R_X35Y119_SLICE_X52Y119_A_CY}),
.CYINIT(1'b0),
.DI({LIOB33_X0Y107_IOB_X0Y107_I, LIOB33_X0Y105_IOB_X0Y106_I, LIOB33_X0Y105_IOB_X0Y105_I, LIOB33_X0Y103_IOB_X0Y104_I}),
.O({CLBLM_R_X35Y119_SLICE_X52Y119_D_XOR, CLBLM_R_X35Y119_SLICE_X52Y119_C_XOR, CLBLM_R_X35Y119_SLICE_X52Y119_B_XOR, CLBLM_R_X35Y119_SLICE_X52Y119_A_XOR}),
.S({CLBLM_R_X35Y119_SLICE_X52Y119_DO6, CLBLM_R_X35Y119_SLICE_X52Y119_CO6, CLBLM_R_X35Y119_SLICE_X52Y119_BO6, CLBLM_R_X35Y119_SLICE_X52Y119_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0000ff00ff)
  ) CLBLM_R_X35Y119_SLICE_X52Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(LIOB33_X0Y121_IOB_X0Y121_I),
.I4(1'b1),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLM_R_X35Y119_SLICE_X52Y119_DO5),
.O6(CLBLM_R_X35Y119_SLICE_X52Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa55aa55aa55aa55)
  ) CLBLM_R_X35Y119_SLICE_X52Y119_CLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(1'b1),
.I2(1'b1),
.I3(LIOB33_X0Y119_IOB_X0Y120_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y119_SLICE_X52Y119_CO5),
.O6(CLBLM_R_X35Y119_SLICE_X52Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc33333333)
  ) CLBLM_R_X35Y119_SLICE_X52Y119_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y119_IOB_X0Y119_I),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLM_R_X35Y119_SLICE_X52Y119_BO5),
.O6(CLBLM_R_X35Y119_SLICE_X52Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc33333333)
  ) CLBLM_R_X35Y119_SLICE_X52Y119_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y117_IOB_X0Y118_I),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_R_X35Y119_SLICE_X52Y119_AO5),
.O6(CLBLM_R_X35Y119_SLICE_X52Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e20000ee220000)
  ) CLBLM_R_X35Y119_SLICE_X53Y119_DLUT (
.I0(CLBLM_R_X35Y121_SLICE_X53Y121_C_XOR),
.I1(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I2(CLBLL_L_X34Y120_SLICE_X51Y120_DO6),
.I3(CLBLM_R_X33Y119_SLICE_X49Y119_AO6),
.I4(CLBLL_L_X34Y128_SLICE_X50Y128_AO6),
.I5(LIOB33_X0Y147_IOB_X0Y147_I),
.O5(CLBLM_R_X35Y119_SLICE_X53Y119_DO5),
.O6(CLBLM_R_X35Y119_SLICE_X53Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8a00ba00ba008a00)
  ) CLBLM_R_X35Y119_SLICE_X53Y119_CLUT (
.I0(CLBLM_R_X35Y123_SLICE_X53Y123_B_XOR),
.I1(LIOB33_X0Y147_IOB_X0Y147_I),
.I2(LIOB33_X0Y145_IOB_X0Y146_I),
.I3(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I4(LIOB33_X0Y127_IOB_X0Y127_I),
.I5(LIOB33_X0Y113_IOB_X0Y113_I),
.O5(CLBLM_R_X35Y119_SLICE_X53Y119_CO5),
.O6(CLBLM_R_X35Y119_SLICE_X53Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccccc404040)
  ) CLBLM_R_X35Y119_SLICE_X53Y119_BLUT (
.I0(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.I1(LIOB33_X0Y147_IOB_X0Y148_I),
.I2(CLBLM_R_X35Y123_SLICE_X53Y123_B_XOR),
.I3(CLBLM_R_X35Y121_SLICE_X52Y121_B_XOR),
.I4(CLBLL_L_X36Y122_SLICE_X55Y122_AO6),
.I5(CLBLM_R_X35Y119_SLICE_X53Y119_CO6),
.O5(CLBLM_R_X35Y119_SLICE_X53Y119_BO5),
.O6(CLBLM_R_X35Y119_SLICE_X53Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffa8ffffff80)
  ) CLBLM_R_X35Y119_SLICE_X53Y119_ALUT (
.I0(CLBLL_L_X36Y116_SLICE_X55Y116_AO5),
.I1(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(CLBLM_R_X35Y119_SLICE_X53Y119_BO6),
.I4(CLBLL_L_X36Y120_SLICE_X54Y120_AO6),
.I5(LIOB33_X0Y127_IOB_X0Y127_I),
.O5(CLBLM_R_X35Y119_SLICE_X53Y119_AO5),
.O6(CLBLM_R_X35Y119_SLICE_X53Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X35Y120_SLICE_X52Y120_CARRY4 (
.CI(CLBLM_R_X35Y119_SLICE_X52Y119_D_CY),
.CO({CLBLM_R_X35Y120_SLICE_X52Y120_D_CY, CLBLM_R_X35Y120_SLICE_X52Y120_C_CY, CLBLM_R_X35Y120_SLICE_X52Y120_B_CY, CLBLM_R_X35Y120_SLICE_X52Y120_A_CY}),
.CYINIT(1'b0),
.DI({LIOB33_X0Y111_IOB_X0Y111_I, LIOB33_X0Y109_IOB_X0Y110_I, LIOB33_X0Y109_IOB_X0Y109_I, LIOB33_X0Y107_IOB_X0Y108_I}),
.O({CLBLM_R_X35Y120_SLICE_X52Y120_D_XOR, CLBLM_R_X35Y120_SLICE_X52Y120_C_XOR, CLBLM_R_X35Y120_SLICE_X52Y120_B_XOR, CLBLM_R_X35Y120_SLICE_X52Y120_A_XOR}),
.S({CLBLM_R_X35Y120_SLICE_X52Y120_DO6, CLBLM_R_X35Y120_SLICE_X52Y120_CO6, CLBLM_R_X35Y120_SLICE_X52Y120_BO6, CLBLM_R_X35Y120_SLICE_X52Y120_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa55555555)
  ) CLBLM_R_X35Y120_SLICE_X52Y120_DLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y125_IOB_X0Y125_I),
.O5(CLBLM_R_X35Y120_SLICE_X52Y120_DO5),
.O6(CLBLM_R_X35Y120_SLICE_X52Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf00ff00ff00ff00f)
  ) CLBLM_R_X35Y120_SLICE_X52Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(LIOB33_X0Y123_IOB_X0Y124_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y120_SLICE_X52Y120_CO5),
.O6(CLBLM_R_X35Y120_SLICE_X52Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f00f0f0f0f)
  ) CLBLM_R_X35Y120_SLICE_X52Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y123_IOB_X0Y123_I),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLM_R_X35Y120_SLICE_X52Y120_BO5),
.O6(CLBLM_R_X35Y120_SLICE_X52Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc33cc33cc33cc33)
  ) CLBLM_R_X35Y120_SLICE_X52Y120_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(1'b1),
.I3(LIOB33_X0Y121_IOB_X0Y122_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y120_SLICE_X52Y120_AO5),
.O6(CLBLM_R_X35Y120_SLICE_X52Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X35Y120_SLICE_X53Y120_CARRY4 (
.CI(1'b0),
.CO({CLBLM_R_X35Y120_SLICE_X53Y120_D_CY, CLBLM_R_X35Y120_SLICE_X53Y120_C_CY, CLBLM_R_X35Y120_SLICE_X53Y120_B_CY, CLBLM_R_X35Y120_SLICE_X53Y120_A_CY}),
.CYINIT(1'b0),
.DI({LIOB33_X0Y103_IOB_X0Y103_I, LIOB33_X0Y101_IOB_X0Y102_I, LIOB33_X0Y101_IOB_X0Y101_I, LIOB33_SING_X0Y100_IOB_X0Y100_I}),
.O({CLBLM_R_X35Y120_SLICE_X53Y120_D_XOR, CLBLM_R_X35Y120_SLICE_X53Y120_C_XOR, CLBLM_R_X35Y120_SLICE_X53Y120_B_XOR, CLBLM_R_X35Y120_SLICE_X53Y120_A_XOR}),
.S({CLBLM_R_X35Y120_SLICE_X53Y120_DO6, CLBLM_R_X35Y120_SLICE_X53Y120_CO6, CLBLM_R_X35Y120_SLICE_X53Y120_BO6, CLBLM_R_X35Y120_SLICE_X53Y120_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0ff0f0f0f0)
  ) CLBLM_R_X35Y120_SLICE_X53Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X35Y120_SLICE_X53Y120_DO5),
.O6(CLBLM_R_X35Y120_SLICE_X53Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33cc33cc33cc33cc)
  ) CLBLM_R_X35Y120_SLICE_X53Y120_CLUT (
.I0(1'b1),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(1'b1),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y120_SLICE_X53Y120_CO5),
.O6(CLBLM_R_X35Y120_SLICE_X53Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c3c3c3c3c3c)
  ) CLBLM_R_X35Y120_SLICE_X53Y120_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y120_SLICE_X53Y120_BO5),
.O6(CLBLM_R_X35Y120_SLICE_X53Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555555aaaaaaaa)
  ) CLBLM_R_X35Y120_SLICE_X53Y120_ALUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLM_R_X35Y120_SLICE_X53Y120_AO5),
.O6(CLBLM_R_X35Y120_SLICE_X53Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X35Y121_SLICE_X52Y121_CARRY4 (
.CI(CLBLM_R_X35Y120_SLICE_X52Y120_D_CY),
.CO({CLBLM_R_X35Y121_SLICE_X52Y121_D_CY, CLBLM_R_X35Y121_SLICE_X52Y121_C_CY, CLBLM_R_X35Y121_SLICE_X52Y121_B_CY, CLBLM_R_X35Y121_SLICE_X52Y121_A_CY}),
.CYINIT(1'b0),
.DI({RIOB33_X105Y101_IOB_X1Y101_I, RIOB33_SING_X105Y100_IOB_X1Y100_I, LIOB33_X0Y113_IOB_X0Y113_I, LIOB33_X0Y111_IOB_X0Y112_I}),
.O({CLBLM_R_X35Y121_SLICE_X52Y121_D_XOR, CLBLM_R_X35Y121_SLICE_X52Y121_C_XOR, CLBLM_R_X35Y121_SLICE_X52Y121_B_XOR, CLBLM_R_X35Y121_SLICE_X52Y121_A_XOR}),
.S({CLBLM_R_X35Y121_SLICE_X52Y121_DO6, CLBLM_R_X35Y121_SLICE_X52Y121_CO6, CLBLM_R_X35Y121_SLICE_X52Y121_BO6, CLBLM_R_X35Y121_SLICE_X52Y121_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf00ff00ff00ff00f)
  ) CLBLM_R_X35Y121_SLICE_X52Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(LIOB33_X0Y129_IOB_X0Y129_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y121_SLICE_X52Y121_DO5),
.O6(CLBLM_R_X35Y121_SLICE_X52Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa5555aaaa5555)
  ) CLBLM_R_X35Y121_SLICE_X52Y121_CLUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(LIOB33_X0Y127_IOB_X0Y128_I),
.I5(1'b1),
.O5(CLBLM_R_X35Y121_SLICE_X52Y121_CO5),
.O6(CLBLM_R_X35Y121_SLICE_X52Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a5a5a5a5a5a5a5)
  ) CLBLM_R_X35Y121_SLICE_X52Y121_BLUT (
.I0(LIOB33_X0Y127_IOB_X0Y127_I),
.I1(1'b1),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y121_SLICE_X52Y121_BO5),
.O6(CLBLM_R_X35Y121_SLICE_X52Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0000ffff0000ff)
  ) CLBLM_R_X35Y121_SLICE_X52Y121_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(LIOB33_X0Y125_IOB_X0Y126_I),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(1'b1),
.O5(CLBLM_R_X35Y121_SLICE_X52Y121_AO5),
.O6(CLBLM_R_X35Y121_SLICE_X52Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X35Y121_SLICE_X53Y121_CARRY4 (
.CI(CLBLM_R_X35Y120_SLICE_X53Y120_D_CY),
.CO({CLBLM_R_X35Y121_SLICE_X53Y121_D_CY, CLBLM_R_X35Y121_SLICE_X53Y121_C_CY, CLBLM_R_X35Y121_SLICE_X53Y121_B_CY, CLBLM_R_X35Y121_SLICE_X53Y121_A_CY}),
.CYINIT(1'b0),
.DI({LIOB33_X0Y107_IOB_X0Y107_I, LIOB33_X0Y105_IOB_X0Y106_I, LIOB33_X0Y105_IOB_X0Y105_I, LIOB33_X0Y103_IOB_X0Y104_I}),
.O({CLBLM_R_X35Y121_SLICE_X53Y121_D_XOR, CLBLM_R_X35Y121_SLICE_X53Y121_C_XOR, CLBLM_R_X35Y121_SLICE_X53Y121_B_XOR, CLBLM_R_X35Y121_SLICE_X53Y121_A_XOR}),
.S({CLBLM_R_X35Y121_SLICE_X53Y121_DO6, CLBLM_R_X35Y121_SLICE_X53Y121_CO6, CLBLM_R_X35Y121_SLICE_X53Y121_BO6, CLBLM_R_X35Y121_SLICE_X53Y121_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c3c3c3c3c3c)
  ) CLBLM_R_X35Y121_SLICE_X53Y121_DLUT (
.I0(1'b1),
.I1(LIOB33_X0Y121_IOB_X0Y121_I),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y121_SLICE_X53Y121_DO5),
.O6(CLBLM_R_X35Y121_SLICE_X53Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a5a5a5a5a5a)
  ) CLBLM_R_X35Y121_SLICE_X53Y121_CLUT (
.I0(LIOB33_X0Y119_IOB_X0Y120_I),
.I1(1'b1),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y121_SLICE_X53Y121_CO5),
.O6(CLBLM_R_X35Y121_SLICE_X53Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c3c3c3c3c3c)
  ) CLBLM_R_X35Y121_SLICE_X53Y121_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y119_IOB_X0Y119_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y121_SLICE_X53Y121_BO5),
.O6(CLBLM_R_X35Y121_SLICE_X53Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333333cccccccc)
  ) CLBLM_R_X35Y121_SLICE_X53Y121_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y117_IOB_X0Y118_I),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_R_X35Y121_SLICE_X53Y121_AO5),
.O6(CLBLM_R_X35Y121_SLICE_X53Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X35Y122_SLICE_X52Y122_CARRY4 (
.CI(CLBLM_R_X35Y121_SLICE_X52Y121_D_CY),
.CO({CLBLM_R_X35Y122_SLICE_X52Y122_D_CY, CLBLM_R_X35Y122_SLICE_X52Y122_C_CY, CLBLM_R_X35Y122_SLICE_X52Y122_B_CY, CLBLM_R_X35Y122_SLICE_X52Y122_A_CY}),
.CYINIT(1'b0),
.DI({RIOB33_X105Y105_IOB_X1Y105_I, RIOB33_X105Y103_IOB_X1Y104_I, RIOB33_X105Y103_IOB_X1Y103_I, RIOB33_X105Y101_IOB_X1Y102_I}),
.O({CLBLM_R_X35Y122_SLICE_X52Y122_D_XOR, CLBLM_R_X35Y122_SLICE_X52Y122_C_XOR, CLBLM_R_X35Y122_SLICE_X52Y122_B_XOR, CLBLM_R_X35Y122_SLICE_X52Y122_A_XOR}),
.S({CLBLM_R_X35Y122_SLICE_X52Y122_DO6, CLBLM_R_X35Y122_SLICE_X52Y122_CO6, CLBLM_R_X35Y122_SLICE_X52Y122_BO6, CLBLM_R_X35Y122_SLICE_X52Y122_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a5a5a5a5a5a5a5)
  ) CLBLM_R_X35Y122_SLICE_X52Y122_DLUT (
.I0(LIOB33_X0Y133_IOB_X0Y133_I),
.I1(1'b1),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y122_SLICE_X52Y122_DO5),
.O6(CLBLM_R_X35Y122_SLICE_X52Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f00f0f0f0f)
  ) CLBLM_R_X35Y122_SLICE_X52Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y131_IOB_X0Y132_I),
.O5(CLBLM_R_X35Y122_SLICE_X52Y122_CO5),
.O6(CLBLM_R_X35Y122_SLICE_X52Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9999999999999999)
  ) CLBLM_R_X35Y122_SLICE_X52Y122_BLUT (
.I0(LIOB33_X0Y131_IOB_X0Y131_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y122_SLICE_X52Y122_BO5),
.O6(CLBLM_R_X35Y122_SLICE_X52Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf00ff00ff00ff00f)
  ) CLBLM_R_X35Y122_SLICE_X52Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y129_IOB_X0Y130_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y122_SLICE_X52Y122_AO5),
.O6(CLBLM_R_X35Y122_SLICE_X52Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X35Y122_SLICE_X53Y122_CARRY4 (
.CI(CLBLM_R_X35Y121_SLICE_X53Y121_D_CY),
.CO({CLBLM_R_X35Y122_SLICE_X53Y122_D_CY, CLBLM_R_X35Y122_SLICE_X53Y122_C_CY, CLBLM_R_X35Y122_SLICE_X53Y122_B_CY, CLBLM_R_X35Y122_SLICE_X53Y122_A_CY}),
.CYINIT(1'b0),
.DI({LIOB33_X0Y111_IOB_X0Y111_I, LIOB33_X0Y109_IOB_X0Y110_I, LIOB33_X0Y109_IOB_X0Y109_I, LIOB33_X0Y107_IOB_X0Y108_I}),
.O({CLBLM_R_X35Y122_SLICE_X53Y122_D_XOR, CLBLM_R_X35Y122_SLICE_X53Y122_C_XOR, CLBLM_R_X35Y122_SLICE_X53Y122_B_XOR, CLBLM_R_X35Y122_SLICE_X53Y122_A_XOR}),
.S({CLBLM_R_X35Y122_SLICE_X53Y122_DO6, CLBLM_R_X35Y122_SLICE_X53Y122_CO6, CLBLM_R_X35Y122_SLICE_X53Y122_BO6, CLBLM_R_X35Y122_SLICE_X53Y122_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ffff00ff00)
  ) CLBLM_R_X35Y122_SLICE_X53Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(1'b1),
.I5(LIOB33_X0Y125_IOB_X0Y125_I),
.O5(CLBLM_R_X35Y122_SLICE_X53Y122_DO5),
.O6(CLBLM_R_X35Y122_SLICE_X53Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333333cccccccc)
  ) CLBLM_R_X35Y122_SLICE_X53Y122_CLUT (
.I0(1'b1),
.I1(LIOB33_X0Y123_IOB_X0Y124_I),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_R_X35Y122_SLICE_X53Y122_CO5),
.O6(CLBLM_R_X35Y122_SLICE_X53Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333333cccccccc)
  ) CLBLM_R_X35Y122_SLICE_X53Y122_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y123_IOB_X0Y123_I),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLM_R_X35Y122_SLICE_X53Y122_BO5),
.O6(CLBLM_R_X35Y122_SLICE_X53Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33cc33cc33cc33cc)
  ) CLBLM_R_X35Y122_SLICE_X53Y122_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y121_IOB_X0Y122_I),
.I2(1'b1),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y122_SLICE_X53Y122_AO5),
.O6(CLBLM_R_X35Y122_SLICE_X53Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X35Y123_SLICE_X52Y123_CARRY4 (
.CI(CLBLM_R_X35Y122_SLICE_X52Y122_D_CY),
.CO({CLBLM_R_X35Y123_SLICE_X52Y123_D_CY, CLBLM_R_X35Y123_SLICE_X52Y123_C_CY, CLBLM_R_X35Y123_SLICE_X52Y123_B_CY, CLBLM_R_X35Y123_SLICE_X52Y123_A_CY}),
.CYINIT(1'b0),
.DI({RIOB33_X105Y109_IOB_X1Y109_I, RIOB33_X105Y107_IOB_X1Y108_I, RIOB33_X105Y107_IOB_X1Y107_I, RIOB33_X105Y105_IOB_X1Y106_I}),
.O({CLBLM_R_X35Y123_SLICE_X52Y123_D_XOR, CLBLM_R_X35Y123_SLICE_X52Y123_C_XOR, CLBLM_R_X35Y123_SLICE_X52Y123_B_XOR, CLBLM_R_X35Y123_SLICE_X52Y123_A_XOR}),
.S({CLBLM_R_X35Y123_SLICE_X52Y123_DO6, CLBLM_R_X35Y123_SLICE_X52Y123_CO6, CLBLM_R_X35Y123_SLICE_X52Y123_BO6, CLBLM_R_X35Y123_SLICE_X52Y123_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc3c3c3c3c3c3c3c3)
  ) CLBLM_R_X35Y123_SLICE_X52Y123_DLUT (
.I0(1'b1),
.I1(LIOB33_X0Y137_IOB_X0Y137_I),
.I2(RIOB33_X105Y109_IOB_X1Y109_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y123_SLICE_X52Y123_DO5),
.O6(CLBLM_R_X35Y123_SLICE_X52Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f00f0f0f0f)
  ) CLBLM_R_X35Y123_SLICE_X52Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y135_IOB_X0Y136_I),
.O5(CLBLM_R_X35Y123_SLICE_X52Y123_CO5),
.O6(CLBLM_R_X35Y123_SLICE_X52Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0000ff00ff)
  ) CLBLM_R_X35Y123_SLICE_X52Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(1'b1),
.I5(LIOB33_X0Y135_IOB_X0Y135_I),
.O5(CLBLM_R_X35Y123_SLICE_X52Y123_BO5),
.O6(CLBLM_R_X35Y123_SLICE_X52Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa55aa55aa55aa55)
  ) CLBLM_R_X35Y123_SLICE_X52Y123_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(1'b1),
.I2(1'b1),
.I3(LIOB33_X0Y133_IOB_X0Y134_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y123_SLICE_X52Y123_AO5),
.O6(CLBLM_R_X35Y123_SLICE_X52Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X35Y123_SLICE_X53Y123_CARRY4 (
.CI(CLBLM_R_X35Y122_SLICE_X53Y122_D_CY),
.CO({CLBLM_R_X35Y123_SLICE_X53Y123_D_CY, CLBLM_R_X35Y123_SLICE_X53Y123_C_CY, CLBLM_R_X35Y123_SLICE_X53Y123_B_CY, CLBLM_R_X35Y123_SLICE_X53Y123_A_CY}),
.CYINIT(1'b0),
.DI({RIOB33_X105Y101_IOB_X1Y101_I, RIOB33_SING_X105Y100_IOB_X1Y100_I, LIOB33_X0Y113_IOB_X0Y113_I, LIOB33_X0Y111_IOB_X0Y112_I}),
.O({CLBLM_R_X35Y123_SLICE_X53Y123_D_XOR, CLBLM_R_X35Y123_SLICE_X53Y123_C_XOR, CLBLM_R_X35Y123_SLICE_X53Y123_B_XOR, CLBLM_R_X35Y123_SLICE_X53Y123_A_XOR}),
.S({CLBLM_R_X35Y123_SLICE_X53Y123_DO6, CLBLM_R_X35Y123_SLICE_X53Y123_CO6, CLBLM_R_X35Y123_SLICE_X53Y123_BO6, CLBLM_R_X35Y123_SLICE_X53Y123_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333cccc3333cccc)
  ) CLBLM_R_X35Y123_SLICE_X53Y123_DLUT (
.I0(1'b1),
.I1(LIOB33_X0Y129_IOB_X0Y129_I),
.I2(1'b1),
.I3(1'b1),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(1'b1),
.O5(CLBLM_R_X35Y123_SLICE_X53Y123_DO5),
.O6(CLBLM_R_X35Y123_SLICE_X53Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0ff0f00f0ff0f0)
  ) CLBLM_R_X35Y123_SLICE_X53Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y127_IOB_X0Y128_I),
.I3(1'b1),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(1'b1),
.O5(CLBLM_R_X35Y123_SLICE_X53Y123_CO5),
.O6(CLBLM_R_X35Y123_SLICE_X53Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333cccc3333cccc)
  ) CLBLM_R_X35Y123_SLICE_X53Y123_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y127_IOB_X0Y127_I),
.I2(1'b1),
.I3(1'b1),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(1'b1),
.O5(CLBLM_R_X35Y123_SLICE_X53Y123_BO5),
.O6(CLBLM_R_X35Y123_SLICE_X53Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c3c3c3c3c3c)
  ) CLBLM_R_X35Y123_SLICE_X53Y123_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y125_IOB_X0Y126_I),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y123_SLICE_X53Y123_AO5),
.O6(CLBLM_R_X35Y123_SLICE_X53Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X35Y124_SLICE_X52Y124_CARRY4 (
.CI(CLBLM_R_X35Y123_SLICE_X52Y123_D_CY),
.CO({CLBLM_R_X35Y124_SLICE_X52Y124_D_CY, CLBLM_R_X35Y124_SLICE_X52Y124_C_CY, CLBLM_R_X35Y124_SLICE_X52Y124_B_CY, CLBLM_R_X35Y124_SLICE_X52Y124_A_CY}),
.CYINIT(1'b0),
.DI({RIOB33_X105Y113_IOB_X1Y113_I, RIOB33_X105Y111_IOB_X1Y112_I, RIOB33_X105Y111_IOB_X1Y111_I, RIOB33_X105Y109_IOB_X1Y110_I}),
.O({CLBLM_R_X35Y124_SLICE_X52Y124_D_XOR, CLBLM_R_X35Y124_SLICE_X52Y124_C_XOR, CLBLM_R_X35Y124_SLICE_X52Y124_B_XOR, CLBLM_R_X35Y124_SLICE_X52Y124_A_XOR}),
.S({CLBLM_R_X35Y124_SLICE_X52Y124_DO6, CLBLM_R_X35Y124_SLICE_X52Y124_CO6, CLBLM_R_X35Y124_SLICE_X52Y124_BO6, CLBLM_R_X35Y124_SLICE_X52Y124_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0000ff00ff)
  ) CLBLM_R_X35Y124_SLICE_X52Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(1'b1),
.I5(LIOB33_X0Y141_IOB_X0Y141_I),
.O5(CLBLM_R_X35Y124_SLICE_X52Y124_DO5),
.O6(CLBLM_R_X35Y124_SLICE_X52Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf00ff00ff00ff00f)
  ) CLBLM_R_X35Y124_SLICE_X52Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y139_IOB_X0Y140_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y124_SLICE_X52Y124_CO5),
.O6(CLBLM_R_X35Y124_SLICE_X52Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9999999999999999)
  ) CLBLM_R_X35Y124_SLICE_X52Y124_BLUT (
.I0(LIOB33_X0Y139_IOB_X0Y139_I),
.I1(RIOB33_X105Y111_IOB_X1Y111_I),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y124_SLICE_X52Y124_BO5),
.O6(CLBLM_R_X35Y124_SLICE_X52Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf00ff00ff00ff00f)
  ) CLBLM_R_X35Y124_SLICE_X52Y124_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(LIOB33_X0Y137_IOB_X0Y138_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y124_SLICE_X52Y124_AO5),
.O6(CLBLM_R_X35Y124_SLICE_X52Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X35Y124_SLICE_X53Y124_CARRY4 (
.CI(CLBLM_R_X35Y123_SLICE_X53Y123_D_CY),
.CO({CLBLM_R_X35Y124_SLICE_X53Y124_D_CY, CLBLM_R_X35Y124_SLICE_X53Y124_C_CY, CLBLM_R_X35Y124_SLICE_X53Y124_B_CY, CLBLM_R_X35Y124_SLICE_X53Y124_A_CY}),
.CYINIT(1'b0),
.DI({RIOB33_X105Y105_IOB_X1Y105_I, RIOB33_X105Y103_IOB_X1Y104_I, RIOB33_X105Y103_IOB_X1Y103_I, RIOB33_X105Y101_IOB_X1Y102_I}),
.O({CLBLM_R_X35Y124_SLICE_X53Y124_D_XOR, CLBLM_R_X35Y124_SLICE_X53Y124_C_XOR, CLBLM_R_X35Y124_SLICE_X53Y124_B_XOR, CLBLM_R_X35Y124_SLICE_X53Y124_A_XOR}),
.S({CLBLM_R_X35Y124_SLICE_X53Y124_DO6, CLBLM_R_X35Y124_SLICE_X53Y124_CO6, CLBLM_R_X35Y124_SLICE_X53Y124_BO6, CLBLM_R_X35Y124_SLICE_X53Y124_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6666666666666666)
  ) CLBLM_R_X35Y124_SLICE_X53Y124_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y133_IOB_X0Y133_I),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y124_SLICE_X53Y124_DO5),
.O6(CLBLM_R_X35Y124_SLICE_X53Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333333cccccccc)
  ) CLBLM_R_X35Y124_SLICE_X53Y124_CLUT (
.I0(1'b1),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y131_IOB_X0Y132_I),
.O5(CLBLM_R_X35Y124_SLICE_X53Y124_CO5),
.O6(CLBLM_R_X35Y124_SLICE_X53Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6666666666666666)
  ) CLBLM_R_X35Y124_SLICE_X53Y124_BLUT (
.I0(LIOB33_X0Y131_IOB_X0Y131_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y124_SLICE_X53Y124_BO5),
.O6(CLBLM_R_X35Y124_SLICE_X53Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff00ff00ff00ff0)
  ) CLBLM_R_X35Y124_SLICE_X53Y124_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y129_IOB_X0Y130_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y124_SLICE_X53Y124_AO5),
.O6(CLBLM_R_X35Y124_SLICE_X53Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X35Y125_SLICE_X52Y125_CARRY4 (
.CI(CLBLM_R_X35Y124_SLICE_X52Y124_D_CY),
.CO({CLBLM_R_X35Y125_SLICE_X52Y125_D_CY, CLBLM_R_X35Y125_SLICE_X52Y125_C_CY, CLBLM_R_X35Y125_SLICE_X52Y125_B_CY, CLBLM_R_X35Y125_SLICE_X52Y125_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, RIOB33_X105Y115_IOB_X1Y116_I, RIOB33_X105Y115_IOB_X1Y115_I, RIOB33_X105Y113_IOB_X1Y114_I}),
.O({CLBLM_R_X35Y125_SLICE_X52Y125_D_XOR, CLBLM_R_X35Y125_SLICE_X52Y125_C_XOR, CLBLM_R_X35Y125_SLICE_X52Y125_B_XOR, CLBLM_R_X35Y125_SLICE_X52Y125_A_XOR}),
.S({CLBLM_R_X35Y125_SLICE_X52Y125_DO6, CLBLM_R_X35Y125_SLICE_X52Y125_CO6, CLBLM_R_X35Y125_SLICE_X52Y125_BO6, CLBLM_R_X35Y125_SLICE_X52Y125_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f00f0f0f0f)
  ) CLBLM_R_X35Y125_SLICE_X52Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y145_IOB_X0Y145_I),
.I3(1'b1),
.I4(1'b1),
.I5(RIOB33_X105Y117_IOB_X1Y117_I),
.O5(CLBLM_R_X35Y125_SLICE_X52Y125_DO5),
.O6(CLBLM_R_X35Y125_SLICE_X52Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa55aa55aa55aa55)
  ) CLBLM_R_X35Y125_SLICE_X52Y125_CLUT (
.I0(LIOB33_X0Y143_IOB_X0Y144_I),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y115_IOB_X1Y116_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y125_SLICE_X52Y125_CO5),
.O6(CLBLM_R_X35Y125_SLICE_X52Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc33333333)
  ) CLBLM_R_X35Y125_SLICE_X52Y125_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y115_IOB_X1Y115_I),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y143_IOB_X0Y143_I),
.O5(CLBLM_R_X35Y125_SLICE_X52Y125_BO5),
.O6(CLBLM_R_X35Y125_SLICE_X52Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa55aa55aa55aa55)
  ) CLBLM_R_X35Y125_SLICE_X52Y125_ALUT (
.I0(LIOB33_X0Y141_IOB_X0Y142_I),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y113_IOB_X1Y114_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y125_SLICE_X52Y125_AO5),
.O6(CLBLM_R_X35Y125_SLICE_X52Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X35Y125_SLICE_X53Y125_CARRY4 (
.CI(CLBLM_R_X35Y124_SLICE_X53Y124_D_CY),
.CO({CLBLM_R_X35Y125_SLICE_X53Y125_D_CY, CLBLM_R_X35Y125_SLICE_X53Y125_C_CY, CLBLM_R_X35Y125_SLICE_X53Y125_B_CY, CLBLM_R_X35Y125_SLICE_X53Y125_A_CY}),
.CYINIT(1'b0),
.DI({RIOB33_X105Y109_IOB_X1Y109_I, RIOB33_X105Y107_IOB_X1Y108_I, RIOB33_X105Y107_IOB_X1Y107_I, RIOB33_X105Y105_IOB_X1Y106_I}),
.O({CLBLM_R_X35Y125_SLICE_X53Y125_D_XOR, CLBLM_R_X35Y125_SLICE_X53Y125_C_XOR, CLBLM_R_X35Y125_SLICE_X53Y125_B_XOR, CLBLM_R_X35Y125_SLICE_X53Y125_A_XOR}),
.S({CLBLM_R_X35Y125_SLICE_X53Y125_DO6, CLBLM_R_X35Y125_SLICE_X53Y125_CO6, CLBLM_R_X35Y125_SLICE_X53Y125_BO6, CLBLM_R_X35Y125_SLICE_X53Y125_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0ff0f0f0f0)
  ) CLBLM_R_X35Y125_SLICE_X53Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y109_IOB_X1Y109_I),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y137_IOB_X0Y137_I),
.O5(CLBLM_R_X35Y125_SLICE_X53Y125_DO5),
.O6(CLBLM_R_X35Y125_SLICE_X53Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0ff0f00f0ff0f0)
  ) CLBLM_R_X35Y125_SLICE_X53Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(1'b1),
.I4(LIOB33_X0Y135_IOB_X0Y136_I),
.I5(1'b1),
.O5(CLBLM_R_X35Y125_SLICE_X53Y125_CO5),
.O6(CLBLM_R_X35Y125_SLICE_X53Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333333cccccccc)
  ) CLBLM_R_X35Y125_SLICE_X53Y125_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y135_IOB_X0Y135_I),
.O5(CLBLM_R_X35Y125_SLICE_X53Y125_BO5),
.O6(CLBLM_R_X35Y125_SLICE_X53Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33cc33cc33cc33cc)
  ) CLBLM_R_X35Y125_SLICE_X53Y125_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(1'b1),
.I3(LIOB33_X0Y133_IOB_X0Y134_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y125_SLICE_X53Y125_AO5),
.O6(CLBLM_R_X35Y125_SLICE_X53Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h80d0d080c0c0c0c0)
  ) CLBLM_R_X35Y126_SLICE_X52Y126_DLUT (
.I0(LIOB33_X0Y147_IOB_X0Y147_I),
.I1(CLBLM_R_X35Y126_SLICE_X53Y126_C_XOR),
.I2(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(LIOB33_X0Y139_IOB_X0Y140_I),
.I5(LIOB33_X0Y145_IOB_X0Y146_I),
.O5(CLBLM_R_X35Y126_SLICE_X52Y126_DO5),
.O6(CLBLM_R_X35Y126_SLICE_X52Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ba00ff003000)
  ) CLBLM_R_X35Y126_SLICE_X52Y126_CLUT (
.I0(CLBLM_R_X35Y124_SLICE_X52Y124_C_XOR),
.I1(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.I2(CLBLM_R_X35Y126_SLICE_X53Y126_C_XOR),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(CLBLM_R_X35Y126_SLICE_X52Y126_DO6),
.I5(CLBLL_L_X36Y122_SLICE_X55Y122_AO6),
.O5(CLBLM_R_X35Y126_SLICE_X52Y126_CO5),
.O6(CLBLM_R_X35Y126_SLICE_X52Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffef0f8f0)
  ) CLBLM_R_X35Y126_SLICE_X52Y126_BLUT (
.I0(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I1(LIOB33_X0Y139_IOB_X0Y140_I),
.I2(CLBLL_L_X36Y126_SLICE_X54Y126_BO6),
.I3(CLBLL_L_X36Y116_SLICE_X55Y116_AO5),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(CLBLM_R_X35Y126_SLICE_X52Y126_CO6),
.O5(CLBLM_R_X35Y126_SLICE_X52Y126_BO5),
.O6(CLBLM_R_X35Y126_SLICE_X52Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8aa80220aaaa0000)
  ) CLBLM_R_X35Y126_SLICE_X52Y126_ALUT (
.I0(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I1(LIOB33_X0Y147_IOB_X0Y147_I),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(LIOB33_X0Y137_IOB_X0Y138_I),
.I4(CLBLM_R_X35Y126_SLICE_X53Y126_A_XOR),
.I5(LIOB33_X0Y145_IOB_X0Y146_I),
.O5(CLBLM_R_X35Y126_SLICE_X52Y126_AO5),
.O6(CLBLM_R_X35Y126_SLICE_X52Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X35Y126_SLICE_X53Y126_CARRY4 (
.CI(CLBLM_R_X35Y125_SLICE_X53Y125_D_CY),
.CO({CLBLM_R_X35Y126_SLICE_X53Y126_D_CY, CLBLM_R_X35Y126_SLICE_X53Y126_C_CY, CLBLM_R_X35Y126_SLICE_X53Y126_B_CY, CLBLM_R_X35Y126_SLICE_X53Y126_A_CY}),
.CYINIT(1'b0),
.DI({RIOB33_X105Y113_IOB_X1Y113_I, RIOB33_X105Y111_IOB_X1Y112_I, RIOB33_X105Y111_IOB_X1Y111_I, RIOB33_X105Y109_IOB_X1Y110_I}),
.O({CLBLM_R_X35Y126_SLICE_X53Y126_D_XOR, CLBLM_R_X35Y126_SLICE_X53Y126_C_XOR, CLBLM_R_X35Y126_SLICE_X53Y126_B_XOR, CLBLM_R_X35Y126_SLICE_X53Y126_A_XOR}),
.S({CLBLM_R_X35Y126_SLICE_X53Y126_DO6, CLBLM_R_X35Y126_SLICE_X53Y126_CO6, CLBLM_R_X35Y126_SLICE_X53Y126_BO6, CLBLM_R_X35Y126_SLICE_X53Y126_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0ff0f0f0f0)
  ) CLBLM_R_X35Y126_SLICE_X53Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y141_IOB_X0Y141_I),
.O5(CLBLM_R_X35Y126_SLICE_X53Y126_DO5),
.O6(CLBLM_R_X35Y126_SLICE_X53Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555555aaaaaaaa)
  ) CLBLM_R_X35Y126_SLICE_X53Y126_CLUT (
.I0(RIOB33_X105Y111_IOB_X1Y112_I),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y139_IOB_X0Y140_I),
.O5(CLBLM_R_X35Y126_SLICE_X53Y126_CO5),
.O6(CLBLM_R_X35Y126_SLICE_X53Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6666666666666666)
  ) CLBLM_R_X35Y126_SLICE_X53Y126_BLUT (
.I0(LIOB33_X0Y139_IOB_X0Y139_I),
.I1(RIOB33_X105Y111_IOB_X1Y111_I),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y126_SLICE_X53Y126_BO5),
.O6(CLBLM_R_X35Y126_SLICE_X53Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff00ff00ff00ff0)
  ) CLBLM_R_X35Y126_SLICE_X53Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(LIOB33_X0Y137_IOB_X0Y138_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y126_SLICE_X53Y126_AO5),
.O6(CLBLM_R_X35Y126_SLICE_X53Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa55555555)
  ) CLBLM_R_X35Y127_SLICE_X52Y127_DLUT (
.I0(RIOB33_X105Y115_IOB_X1Y115_I),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y143_IOB_X0Y143_I),
.O5(CLBLM_R_X35Y127_SLICE_X52Y127_DO5),
.O6(CLBLM_R_X35Y127_SLICE_X52Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc30fc3022220000)
  ) CLBLM_R_X35Y127_SLICE_X52Y127_CLUT (
.I0(CLBLL_L_X36Y125_SLICE_X55Y125_BO6),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(CLBLL_L_X34Y127_SLICE_X50Y127_BO6),
.I3(CLBLL_L_X34Y126_SLICE_X50Y126_DO6),
.I4(CLBLL_L_X36Y116_SLICE_X54Y116_BO5),
.I5(LIOB33_X0Y145_IOB_X0Y146_I),
.O5(CLBLM_R_X35Y127_SLICE_X52Y127_CO5),
.O6(CLBLM_R_X35Y127_SLICE_X52Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f030fc2222f0f0)
  ) CLBLM_R_X35Y127_SLICE_X52Y127_BLUT (
.I0(CLBLM_R_X35Y125_SLICE_X52Y125_B_XOR),
.I1(LIOB33_X0Y145_IOB_X0Y146_I),
.I2(CLBLM_R_X35Y127_SLICE_X53Y127_B_XOR),
.I3(CLBLM_R_X35Y127_SLICE_X52Y127_DO6),
.I4(LIOB33_X0Y147_IOB_X0Y147_I),
.I5(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.O5(CLBLM_R_X35Y127_SLICE_X52Y127_BO5),
.O6(CLBLM_R_X35Y127_SLICE_X52Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00fe54ea40)
  ) CLBLM_R_X35Y127_SLICE_X52Y127_ALUT (
.I0(LIOB33_X0Y147_IOB_X0Y148_I),
.I1(RIOB33_X105Y115_IOB_X1Y115_I),
.I2(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I3(CLBLM_R_X35Y127_SLICE_X52Y127_BO6),
.I4(LIOB33_X0Y143_IOB_X0Y143_I),
.I5(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.O5(CLBLM_R_X35Y127_SLICE_X52Y127_AO5),
.O6(CLBLM_R_X35Y127_SLICE_X52Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X35Y127_SLICE_X53Y127_CARRY4 (
.CI(CLBLM_R_X35Y126_SLICE_X53Y126_D_CY),
.CO({CLBLM_R_X35Y127_SLICE_X53Y127_D_CY, CLBLM_R_X35Y127_SLICE_X53Y127_C_CY, CLBLM_R_X35Y127_SLICE_X53Y127_B_CY, CLBLM_R_X35Y127_SLICE_X53Y127_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, RIOB33_X105Y115_IOB_X1Y116_I, RIOB33_X105Y115_IOB_X1Y115_I, RIOB33_X105Y113_IOB_X1Y114_I}),
.O({CLBLM_R_X35Y127_SLICE_X53Y127_D_XOR, CLBLM_R_X35Y127_SLICE_X53Y127_C_XOR, CLBLM_R_X35Y127_SLICE_X53Y127_B_XOR, CLBLM_R_X35Y127_SLICE_X53Y127_A_XOR}),
.S({CLBLM_R_X35Y127_SLICE_X53Y127_DO6, CLBLM_R_X35Y127_SLICE_X53Y127_CO6, CLBLM_R_X35Y127_SLICE_X53Y127_BO6, CLBLM_R_X35Y127_SLICE_X53Y127_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333333cccccccc)
  ) CLBLM_R_X35Y127_SLICE_X53Y127_DLUT (
.I0(1'b1),
.I1(RIOB33_X105Y117_IOB_X1Y117_I),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y145_IOB_X0Y145_I),
.O5(CLBLM_R_X35Y127_SLICE_X53Y127_DO5),
.O6(CLBLM_R_X35Y127_SLICE_X53Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333333cccccccc)
  ) CLBLM_R_X35Y127_SLICE_X53Y127_CLUT (
.I0(1'b1),
.I1(RIOB33_X105Y115_IOB_X1Y116_I),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y143_IOB_X0Y144_I),
.O5(CLBLM_R_X35Y127_SLICE_X53Y127_CO5),
.O6(CLBLM_R_X35Y127_SLICE_X53Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333cccc3333cccc)
  ) CLBLM_R_X35Y127_SLICE_X53Y127_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y143_IOB_X0Y143_I),
.I2(1'b1),
.I3(1'b1),
.I4(RIOB33_X105Y115_IOB_X1Y115_I),
.I5(1'b1),
.O5(CLBLM_R_X35Y127_SLICE_X53Y127_BO5),
.O6(CLBLM_R_X35Y127_SLICE_X53Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0ff0f0f0f0)
  ) CLBLM_R_X35Y127_SLICE_X53Y127_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y113_IOB_X1Y114_I),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y141_IOB_X0Y142_I),
.O5(CLBLM_R_X35Y127_SLICE_X53Y127_AO5),
.O6(CLBLM_R_X35Y127_SLICE_X53Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X35Y128_SLICE_X52Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y128_SLICE_X52Y128_DO5),
.O6(CLBLM_R_X35Y128_SLICE_X52Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0f5e4e4a0)
  ) CLBLM_R_X35Y128_SLICE_X52Y128_CLUT (
.I0(LIOB33_X0Y147_IOB_X0Y148_I),
.I1(LIOB33_X0Y141_IOB_X0Y142_I),
.I2(CLBLM_R_X35Y128_SLICE_X53Y128_BO6),
.I3(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I4(RIOB33_X105Y113_IOB_X1Y114_I),
.I5(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.O5(CLBLM_R_X35Y128_SLICE_X52Y128_CO5),
.O6(CLBLM_R_X35Y128_SLICE_X52Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b80000fc300000)
  ) CLBLM_R_X35Y128_SLICE_X52Y128_BLUT (
.I0(CLBLM_R_X35Y127_SLICE_X53Y127_D_XOR),
.I1(LIOB33_X0Y147_IOB_X0Y147_I),
.I2(CLBLM_R_X35Y127_SLICE_X52Y127_CO6),
.I3(RIOB33_X105Y117_IOB_X1Y117_I),
.I4(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I5(LIOB33_X0Y145_IOB_X0Y146_I),
.O5(CLBLM_R_X35Y128_SLICE_X52Y128_BO5),
.O6(CLBLM_R_X35Y128_SLICE_X52Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0f3c0e2c0e2c0c0)
  ) CLBLM_R_X35Y128_SLICE_X52Y128_ALUT (
.I0(LIOB33_X0Y143_IOB_X0Y144_I),
.I1(LIOB33_X0Y147_IOB_X0Y148_I),
.I2(CLBLM_R_X35Y128_SLICE_X53Y128_AO6),
.I3(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.I4(RIOB33_X105Y115_IOB_X1Y116_I),
.I5(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.O5(CLBLM_R_X35Y128_SLICE_X52Y128_AO5),
.O6(CLBLM_R_X35Y128_SLICE_X52Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc3c3c3c3c3c3c3c3)
  ) CLBLM_R_X35Y128_SLICE_X53Y128_DLUT (
.I0(1'b1),
.I1(LIOB33_X0Y141_IOB_X0Y142_I),
.I2(RIOB33_X105Y113_IOB_X1Y114_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y128_SLICE_X53Y128_DO5),
.O6(CLBLM_R_X35Y128_SLICE_X53Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc33cc33cc33cc33)
  ) CLBLM_R_X35Y128_SLICE_X53Y128_CLUT (
.I0(1'b1),
.I1(LIOB33_X0Y143_IOB_X0Y144_I),
.I2(1'b1),
.I3(RIOB33_X105Y115_IOB_X1Y116_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y128_SLICE_X53Y128_CO5),
.O6(CLBLM_R_X35Y128_SLICE_X53Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5ff05000fcf00c0)
  ) CLBLM_R_X35Y128_SLICE_X53Y128_BLUT (
.I0(CLBLM_R_X35Y128_SLICE_X53Y128_DO6),
.I1(CLBLM_R_X35Y125_SLICE_X52Y125_A_XOR),
.I2(LIOB33_X0Y147_IOB_X0Y147_I),
.I3(LIOB33_X0Y145_IOB_X0Y146_I),
.I4(CLBLM_R_X35Y127_SLICE_X53Y127_A_XOR),
.I5(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.O5(CLBLM_R_X35Y128_SLICE_X53Y128_BO5),
.O6(CLBLM_R_X35Y128_SLICE_X53Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha23aa20aae3aae0a)
  ) CLBLM_R_X35Y128_SLICE_X53Y128_ALUT (
.I0(CLBLM_R_X35Y127_SLICE_X53Y127_C_XOR),
.I1(LIOB33_X0Y145_IOB_X0Y146_I),
.I2(LIOB33_X0Y147_IOB_X0Y147_I),
.I3(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I4(CLBLM_R_X35Y125_SLICE_X52Y125_C_XOR),
.I5(CLBLM_R_X35Y128_SLICE_X53Y128_CO6),
.O5(CLBLM_R_X35Y128_SLICE_X53Y128_AO5),
.O6(CLBLM_R_X35Y128_SLICE_X53Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X35Y129_SLICE_X52Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y129_SLICE_X52Y129_DO5),
.O6(CLBLM_R_X35Y129_SLICE_X52Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc3c3c3c3c3c3c3c3)
  ) CLBLM_R_X35Y129_SLICE_X52Y129_CLUT (
.I0(1'b1),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(LIOB33_X0Y141_IOB_X0Y141_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y129_SLICE_X52Y129_CO5),
.O6(CLBLM_R_X35Y129_SLICE_X52Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb1a07070b1a0f8f8)
  ) CLBLM_R_X35Y129_SLICE_X52Y129_BLUT (
.I0(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I1(LIOB33_X0Y145_IOB_X0Y146_I),
.I2(CLBLM_R_X35Y126_SLICE_X53Y126_D_XOR),
.I3(CLBLM_R_X35Y124_SLICE_X52Y124_D_XOR),
.I4(LIOB33_X0Y147_IOB_X0Y147_I),
.I5(CLBLM_R_X35Y129_SLICE_X52Y129_CO6),
.O5(CLBLM_R_X35Y129_SLICE_X52Y129_BO5),
.O6(CLBLM_R_X35Y129_SLICE_X52Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ff00e8e8)
  ) CLBLM_R_X35Y129_SLICE_X52Y129_ALUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(LIOB33_X0Y141_IOB_X0Y141_I),
.I2(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I3(CLBLM_R_X35Y129_SLICE_X52Y129_BO6),
.I4(LIOB33_X0Y147_IOB_X0Y148_I),
.I5(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.O5(CLBLM_R_X35Y129_SLICE_X52Y129_AO5),
.O6(CLBLM_R_X35Y129_SLICE_X52Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X35Y129_SLICE_X53Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X35Y129_SLICE_X53Y129_DO5),
.O6(CLBLM_R_X35Y129_SLICE_X53Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc33333333)
  ) CLBLM_R_X35Y129_SLICE_X53Y129_CLUT (
.I0(1'b1),
.I1(RIOB33_X105Y117_IOB_X1Y117_I),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y145_IOB_X0Y145_I),
.O5(CLBLM_R_X35Y129_SLICE_X53Y129_CO5),
.O6(CLBLM_R_X35Y129_SLICE_X53Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5050554450504400)
  ) CLBLM_R_X35Y129_SLICE_X53Y129_BLUT (
.I0(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I1(LIOB33_X0Y145_IOB_X0Y145_I),
.I2(CLBLM_R_X35Y127_SLICE_X53Y127_D_XOR),
.I3(LIOB33_X0Y145_IOB_X0Y146_I),
.I4(LIOB33_X0Y147_IOB_X0Y147_I),
.I5(RIOB33_X105Y117_IOB_X1Y117_I),
.O5(CLBLM_R_X35Y129_SLICE_X53Y129_BO5),
.O6(CLBLM_R_X35Y129_SLICE_X53Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0e450f0a0e4faf0)
  ) CLBLM_R_X35Y129_SLICE_X53Y129_ALUT (
.I0(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I1(CLBLM_R_X35Y125_SLICE_X52Y125_D_XOR),
.I2(CLBLM_R_X35Y127_SLICE_X53Y127_D_XOR),
.I3(LIOB33_X0Y145_IOB_X0Y146_I),
.I4(LIOB33_X0Y147_IOB_X0Y147_I),
.I5(CLBLM_R_X35Y129_SLICE_X53Y129_CO6),
.O5(CLBLM_R_X35Y129_SLICE_X53Y129_AO5),
.O6(CLBLM_R_X35Y129_SLICE_X53Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y117_SLICE_X56Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y117_SLICE_X56Y117_DO5),
.O6(CLBLM_R_X37Y117_SLICE_X56Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y117_SLICE_X56Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y117_SLICE_X56Y117_CO5),
.O6(CLBLM_R_X37Y117_SLICE_X56Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y117_SLICE_X56Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y117_SLICE_X56Y117_BO5),
.O6(CLBLM_R_X37Y117_SLICE_X56Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe32ce0232320202)
  ) CLBLM_R_X37Y117_SLICE_X56Y117_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y117_IOB_X0Y118_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(RIOB33_X105Y117_IOB_X1Y117_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(1'b1),
.O5(CLBLM_R_X37Y117_SLICE_X56Y117_AO5),
.O6(CLBLM_R_X37Y117_SLICE_X56Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y117_SLICE_X57Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y117_SLICE_X57Y117_DO5),
.O6(CLBLM_R_X37Y117_SLICE_X57Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y117_SLICE_X57Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y117_SLICE_X57Y117_CO5),
.O6(CLBLM_R_X37Y117_SLICE_X57Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y117_SLICE_X57Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y117_SLICE_X57Y117_BO5),
.O6(CLBLM_R_X37Y117_SLICE_X57Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y117_SLICE_X57Y117_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y117_SLICE_X57Y117_AO5),
.O6(CLBLM_R_X37Y117_SLICE_X57Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hddd8ddd888d888d8)
  ) CLBLM_R_X37Y118_SLICE_X56Y118_DLUT (
.I0(LIOB33_X0Y145_IOB_X0Y146_I),
.I1(CLBLM_R_X35Y124_SLICE_X53Y124_A_XOR),
.I2(CLBLM_R_X37Y118_SLICE_X57Y118_BO6),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(1'b1),
.I5(CLBLM_R_X37Y118_SLICE_X56Y118_BO6),
.O5(CLBLM_R_X37Y118_SLICE_X56Y118_DO5),
.O6(CLBLM_R_X37Y118_SLICE_X56Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ccccff00aaaa)
  ) CLBLM_R_X37Y118_SLICE_X56Y118_CLUT (
.I0(CLBLM_R_X37Y117_SLICE_X56Y117_AO6),
.I1(CLBLL_L_X36Y117_SLICE_X55Y117_BO5),
.I2(CLBLL_L_X38Y118_SLICE_X58Y118_AO5),
.I3(CLBLL_L_X36Y118_SLICE_X55Y118_AO5),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLM_R_X37Y118_SLICE_X56Y118_CO5),
.O6(CLBLM_R_X37Y118_SLICE_X56Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8ffb8ccb833b800)
  ) CLBLM_R_X37Y118_SLICE_X56Y118_BLUT (
.I0(CLBLL_L_X36Y117_SLICE_X55Y117_BO5),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(CLBLM_R_X37Y117_SLICE_X56Y117_AO6),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(CLBLM_R_X35Y118_SLICE_X53Y118_AO6),
.I5(CLBLL_L_X36Y118_SLICE_X55Y118_AO5),
.O5(CLBLM_R_X37Y118_SLICE_X56Y118_BO5),
.O6(CLBLM_R_X37Y118_SLICE_X56Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb080b080f0f00000)
  ) CLBLM_R_X37Y118_SLICE_X56Y118_ALUT (
.I0(CLBLM_R_X37Y118_SLICE_X56Y118_DO6),
.I1(LIOB33_X0Y147_IOB_X0Y147_I),
.I2(CLBLL_L_X34Y128_SLICE_X50Y128_AO6),
.I3(CLBLL_L_X36Y118_SLICE_X54Y118_CO6),
.I4(CLBLM_R_X35Y124_SLICE_X53Y124_A_XOR),
.I5(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.O5(CLBLM_R_X37Y118_SLICE_X56Y118_AO5),
.O6(CLBLM_R_X37Y118_SLICE_X56Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee2222fc30fc30)
  ) CLBLM_R_X37Y118_SLICE_X57Y118_DLUT (
.I0(CLBLL_L_X38Y118_SLICE_X58Y118_AO6),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(CLBLL_L_X36Y117_SLICE_X55Y117_AO5),
.I3(CLBLL_L_X36Y116_SLICE_X54Y116_AO5),
.I4(CLBLL_L_X34Y119_SLICE_X51Y119_AO6),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLM_R_X37Y118_SLICE_X57Y118_DO5),
.O6(CLBLM_R_X37Y118_SLICE_X57Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0afa0fcfc0c0c)
  ) CLBLM_R_X37Y118_SLICE_X57Y118_CLUT (
.I0(CLBLL_L_X38Y118_SLICE_X58Y118_AO6),
.I1(CLBLL_L_X36Y115_SLICE_X54Y115_AO6),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(CLBLL_L_X36Y116_SLICE_X54Y116_AO5),
.I4(CLBLL_L_X36Y117_SLICE_X55Y117_AO5),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLM_R_X37Y118_SLICE_X57Y118_CO5),
.O6(CLBLM_R_X37Y118_SLICE_X57Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3c0bbbbf3c08888)
  ) CLBLM_R_X37Y118_SLICE_X57Y118_BLUT (
.I0(CLBLL_L_X36Y117_SLICE_X55Y117_AO5),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(CLBLL_L_X36Y116_SLICE_X54Y116_AO5),
.I3(CLBLL_L_X36Y115_SLICE_X54Y115_AO6),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(CLBLM_R_X37Y118_SLICE_X57Y118_AO5),
.O5(CLBLM_R_X37Y118_SLICE_X57Y118_BO5),
.O6(CLBLM_R_X37Y118_SLICE_X57Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33002222f3c0e2e2)
  ) CLBLM_R_X37Y118_SLICE_X57Y118_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(LIOB33_X0Y117_IOB_X0Y118_I),
.I2(RIOB33_X105Y117_IOB_X1Y117_I),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(1'b1),
.O5(CLBLM_R_X37Y118_SLICE_X57Y118_AO5),
.O6(CLBLM_R_X37Y118_SLICE_X57Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5b1f5b1e4a0e4a0)
  ) CLBLM_R_X37Y119_SLICE_X56Y119_DLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(CLBLM_R_X37Y119_SLICE_X57Y119_BO6),
.I3(CLBLL_L_X38Y118_SLICE_X58Y118_AO5),
.I4(1'b1),
.I5(CLBLL_L_X36Y118_SLICE_X55Y118_AO5),
.O5(CLBLM_R_X37Y119_SLICE_X56Y119_DO5),
.O6(CLBLM_R_X37Y119_SLICE_X56Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5f5f5a0a0a0)
  ) CLBLM_R_X37Y119_SLICE_X56Y119_CLUT (
.I0(LIOB33_X0Y145_IOB_X0Y146_I),
.I1(1'b1),
.I2(CLBLM_R_X35Y124_SLICE_X53Y124_B_XOR),
.I3(CLBLM_R_X37Y118_SLICE_X57Y118_CO6),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(CLBLM_R_X37Y118_SLICE_X56Y118_BO6),
.O5(CLBLM_R_X37Y119_SLICE_X56Y119_CO5),
.O6(CLBLM_R_X37Y119_SLICE_X56Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafcfcaaaa0c0c)
  ) CLBLM_R_X37Y119_SLICE_X56Y119_BLUT (
.I0(CLBLM_R_X35Y123_SLICE_X53Y123_D_XOR),
.I1(CLBLL_L_X36Y118_SLICE_X55Y118_BO6),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(1'b1),
.I4(LIOB33_X0Y145_IOB_X0Y146_I),
.I5(CLBLM_R_X37Y118_SLICE_X57Y118_BO6),
.O5(CLBLM_R_X37Y119_SLICE_X56Y119_BO5),
.O6(CLBLM_R_X37Y119_SLICE_X56Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcb8000074300000)
  ) CLBLM_R_X37Y119_SLICE_X56Y119_ALUT (
.I0(LIOB33_X0Y147_IOB_X0Y147_I),
.I1(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I2(CLBLM_R_X35Y124_SLICE_X53Y124_B_XOR),
.I3(CLBLL_L_X36Y119_SLICE_X54Y119_CO6),
.I4(CLBLL_L_X34Y128_SLICE_X50Y128_AO6),
.I5(CLBLM_R_X37Y119_SLICE_X56Y119_CO6),
.O5(CLBLM_R_X37Y119_SLICE_X56Y119_AO5),
.O6(CLBLM_R_X37Y119_SLICE_X56Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55ff55aa00aa00)
  ) CLBLM_R_X37Y119_SLICE_X57Y119_DLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X37Y119_SLICE_X57Y119_CO6),
.I4(1'b1),
.I5(CLBLL_L_X38Y119_SLICE_X58Y119_AO6),
.O5(CLBLM_R_X37Y119_SLICE_X57Y119_DO5),
.O6(CLBLM_R_X37Y119_SLICE_X57Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000033b800b8)
  ) CLBLM_R_X37Y119_SLICE_X57Y119_CLUT (
.I0(RIOB33_X105Y117_IOB_X1Y117_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(RIOB33_X105Y109_IOB_X1Y109_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(LIOB33_X0Y117_IOB_X0Y118_I),
.O5(CLBLM_R_X37Y119_SLICE_X57Y119_CO5),
.O6(CLBLM_R_X37Y119_SLICE_X57Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefe0202fffc0300)
  ) CLBLM_R_X37Y119_SLICE_X57Y119_BLUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(LIOB33_X0Y117_IOB_X0Y118_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(RIOB33_X105Y109_IOB_X1Y109_I),
.I4(RIOB33_X105Y117_IOB_X1Y117_I),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLM_R_X37Y119_SLICE_X57Y119_BO5),
.O6(CLBLM_R_X37Y119_SLICE_X57Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc480ffffc4800000)
  ) CLBLM_R_X37Y119_SLICE_X57Y119_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(CLBLL_L_X36Y121_SLICE_X54Y121_AO5),
.I2(RIOB33_X105Y115_IOB_X1Y115_I),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(CLBLM_R_X37Y119_SLICE_X57Y119_CO6),
.O5(CLBLM_R_X37Y119_SLICE_X57Y119_AO5),
.O6(CLBLM_R_X37Y119_SLICE_X57Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0dd88f0f0dd88)
  ) CLBLM_R_X37Y120_SLICE_X56Y120_DLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(CLBLM_R_X37Y118_SLICE_X57Y118_DO6),
.I2(CLBLM_R_X35Y124_SLICE_X53Y124_D_XOR),
.I3(CLBLM_R_X37Y118_SLICE_X56Y118_CO6),
.I4(LIOB33_X0Y145_IOB_X0Y146_I),
.I5(1'b1),
.O5(CLBLM_R_X37Y120_SLICE_X56Y120_DO5),
.O6(CLBLM_R_X37Y120_SLICE_X56Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0afa0acacacac)
  ) CLBLM_R_X37Y120_SLICE_X56Y120_CLUT (
.I0(CLBLM_R_X35Y124_SLICE_X53Y124_C_XOR),
.I1(CLBLM_R_X37Y118_SLICE_X57Y118_CO6),
.I2(LIOB33_X0Y145_IOB_X0Y146_I),
.I3(CLBLM_R_X37Y118_SLICE_X56Y118_CO6),
.I4(1'b1),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLM_R_X37Y120_SLICE_X56Y120_CO5),
.O6(CLBLM_R_X37Y120_SLICE_X56Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88c0ccc088c000c0)
  ) CLBLM_R_X37Y120_SLICE_X56Y120_BLUT (
.I0(CLBLM_R_X37Y120_SLICE_X56Y120_DO6),
.I1(CLBLL_L_X34Y128_SLICE_X50Y128_AO6),
.I2(CLBLM_R_X35Y124_SLICE_X53Y124_D_XOR),
.I3(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I4(LIOB33_X0Y147_IOB_X0Y147_I),
.I5(CLBLL_L_X36Y120_SLICE_X55Y120_AO6),
.O5(CLBLM_R_X37Y120_SLICE_X56Y120_BO5),
.O6(CLBLM_R_X37Y120_SLICE_X56Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccc088c000c088c0)
  ) CLBLM_R_X37Y120_SLICE_X56Y120_ALUT (
.I0(CLBLL_L_X36Y120_SLICE_X54Y120_CO6),
.I1(CLBLL_L_X34Y128_SLICE_X50Y128_AO6),
.I2(CLBLM_R_X35Y124_SLICE_X53Y124_C_XOR),
.I3(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I4(LIOB33_X0Y147_IOB_X0Y147_I),
.I5(CLBLM_R_X37Y120_SLICE_X56Y120_CO6),
.O5(CLBLM_R_X37Y120_SLICE_X56Y120_AO5),
.O6(CLBLM_R_X37Y120_SLICE_X56Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y120_SLICE_X57Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y120_SLICE_X57Y120_DO5),
.O6(CLBLM_R_X37Y120_SLICE_X57Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y120_SLICE_X57Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y120_SLICE_X57Y120_CO5),
.O6(CLBLM_R_X37Y120_SLICE_X57Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y120_SLICE_X57Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y120_SLICE_X57Y120_BO5),
.O6(CLBLM_R_X37Y120_SLICE_X57Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y120_SLICE_X57Y120_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y120_SLICE_X57Y120_AO5),
.O6(CLBLM_R_X37Y120_SLICE_X57Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000fef80e08)
  ) CLBLM_R_X37Y121_SLICE_X56Y121_DLUT (
.I0(LIOB33_X0Y129_IOB_X0Y130_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(LIOB33_X0Y147_IOB_X0Y148_I),
.I3(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I4(CLBLM_R_X37Y122_SLICE_X56Y122_CO6),
.I5(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.O5(CLBLM_R_X37Y121_SLICE_X56Y121_DO5),
.O6(CLBLM_R_X37Y121_SLICE_X56Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_R_X37Y121_SLICE_X56Y121_CLUT (
.I0(CLBLM_R_X37Y119_SLICE_X56Y119_AO6),
.I1(CLBLM_R_X37Y118_SLICE_X56Y118_AO6),
.I2(CLBLM_R_X37Y121_SLICE_X57Y121_BO6),
.I3(CLBLL_L_X38Y121_SLICE_X58Y121_BO6),
.I4(CLBLM_R_X37Y121_SLICE_X56Y121_DO6),
.I5(CLBLL_L_X36Y119_SLICE_X55Y119_AO6),
.O5(CLBLM_R_X37Y121_SLICE_X56Y121_CO5),
.O6(CLBLM_R_X37Y121_SLICE_X56Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdf00fd0002002000)
  ) CLBLM_R_X37Y121_SLICE_X56Y121_BLUT (
.I0(LIOB33_X0Y145_IOB_X0Y146_I),
.I1(LIOB33_X0Y147_IOB_X0Y147_I),
.I2(LIOB33_X0Y129_IOB_X0Y130_I),
.I3(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(CLBLM_R_X35Y124_SLICE_X53Y124_A_XOR),
.O5(CLBLM_R_X37Y121_SLICE_X56Y121_BO5),
.O6(CLBLM_R_X37Y121_SLICE_X56Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaa2aaa0aa22aa00)
  ) CLBLM_R_X37Y121_SLICE_X56Y121_ALUT (
.I0(LIOB33_X0Y147_IOB_X0Y148_I),
.I1(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.I2(CLBLL_L_X36Y122_SLICE_X55Y122_AO6),
.I3(CLBLM_R_X37Y121_SLICE_X56Y121_BO6),
.I4(CLBLM_R_X35Y124_SLICE_X53Y124_A_XOR),
.I5(CLBLM_R_X35Y122_SLICE_X52Y122_A_XOR),
.O5(CLBLM_R_X37Y121_SLICE_X56Y121_AO5),
.O6(CLBLM_R_X37Y121_SLICE_X56Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00f0faa55aa55)
  ) CLBLM_R_X37Y121_SLICE_X57Y121_DLUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(1'b1),
.I2(LIOB33_X0Y131_IOB_X0Y131_I),
.I3(LIOB33_X0Y127_IOB_X0Y128_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(1'b1),
.O5(CLBLM_R_X37Y121_SLICE_X57Y121_DO5),
.O6(CLBLM_R_X37Y121_SLICE_X57Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0aaafa0caa0caa)
  ) CLBLM_R_X37Y121_SLICE_X57Y121_CLUT (
.I0(CLBLM_R_X35Y124_SLICE_X53Y124_B_XOR),
.I1(CLBLM_R_X35Y122_SLICE_X52Y122_B_XOR),
.I2(LIOB33_X0Y145_IOB_X0Y146_I),
.I3(LIOB33_X0Y147_IOB_X0Y147_I),
.I4(CLBLM_R_X37Y121_SLICE_X57Y121_DO6),
.I5(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.O5(CLBLM_R_X37Y121_SLICE_X57Y121_CO5),
.O6(CLBLM_R_X37Y121_SLICE_X57Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00e8000000e8)
  ) CLBLM_R_X37Y121_SLICE_X57Y121_BLUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I2(LIOB33_X0Y131_IOB_X0Y131_I),
.I3(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.I4(LIOB33_X0Y147_IOB_X0Y148_I),
.I5(CLBLM_R_X37Y121_SLICE_X57Y121_CO6),
.O5(CLBLM_R_X37Y121_SLICE_X57Y121_BO5),
.O6(CLBLM_R_X37Y121_SLICE_X57Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffafff8fff8fff0)
  ) CLBLM_R_X37Y121_SLICE_X57Y121_ALUT (
.I0(CLBLL_L_X36Y116_SLICE_X55Y116_AO5),
.I1(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I2(CLBLM_R_X37Y121_SLICE_X56Y121_AO6),
.I3(CLBLM_R_X37Y118_SLICE_X56Y118_AO6),
.I4(LIOB33_X0Y129_IOB_X0Y130_I),
.I5(RIOB33_X105Y101_IOB_X1Y102_I),
.O5(CLBLM_R_X37Y121_SLICE_X57Y121_AO5),
.O6(CLBLM_R_X37Y121_SLICE_X57Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa55555555)
  ) CLBLM_R_X37Y122_SLICE_X56Y122_DLUT (
.I0(LIOB33_X0Y129_IOB_X0Y130_I),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(RIOB33_X105Y101_IOB_X1Y102_I),
.O5(CLBLM_R_X37Y122_SLICE_X56Y122_DO5),
.O6(CLBLM_R_X37Y122_SLICE_X56Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haf00ff505d085d08)
  ) CLBLM_R_X37Y122_SLICE_X56Y122_CLUT (
.I0(LIOB33_X0Y147_IOB_X0Y147_I),
.I1(CLBLM_R_X35Y122_SLICE_X52Y122_A_XOR),
.I2(LIOB33_X0Y145_IOB_X0Y146_I),
.I3(CLBLM_R_X35Y124_SLICE_X53Y124_A_XOR),
.I4(CLBLM_R_X37Y122_SLICE_X56Y122_DO6),
.I5(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.O5(CLBLM_R_X37Y122_SLICE_X56Y122_CO5),
.O6(CLBLM_R_X37Y122_SLICE_X56Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c04488c0c0c0c0)
  ) CLBLM_R_X37Y122_SLICE_X56Y122_BLUT (
.I0(LIOB33_X0Y131_IOB_X0Y131_I),
.I1(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I2(CLBLM_R_X35Y124_SLICE_X53Y124_B_XOR),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(LIOB33_X0Y147_IOB_X0Y147_I),
.I5(LIOB33_X0Y145_IOB_X0Y146_I),
.O5(CLBLM_R_X37Y122_SLICE_X56Y122_BO5),
.O6(CLBLM_R_X37Y122_SLICE_X56Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff20000ff220000)
  ) CLBLM_R_X37Y122_SLICE_X56Y122_ALUT (
.I0(CLBLM_R_X35Y124_SLICE_X53Y124_B_XOR),
.I1(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.I2(CLBLL_L_X36Y122_SLICE_X55Y122_AO6),
.I3(CLBLM_R_X37Y122_SLICE_X56Y122_BO6),
.I4(LIOB33_X0Y147_IOB_X0Y148_I),
.I5(CLBLM_R_X35Y122_SLICE_X52Y122_B_XOR),
.O5(CLBLM_R_X37Y122_SLICE_X56Y122_AO5),
.O6(CLBLM_R_X37Y122_SLICE_X56Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y122_SLICE_X57Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y122_SLICE_X57Y122_DO5),
.O6(CLBLM_R_X37Y122_SLICE_X57Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8dd8cccc00000000)
  ) CLBLM_R_X37Y122_SLICE_X57Y122_CLUT (
.I0(LIOB33_X0Y147_IOB_X0Y147_I),
.I1(CLBLM_R_X35Y124_SLICE_X53Y124_D_XOR),
.I2(LIOB33_X0Y133_IOB_X0Y133_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y145_IOB_X0Y146_I),
.I5(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.O5(CLBLM_R_X37Y122_SLICE_X57Y122_CO5),
.O6(CLBLM_R_X37Y122_SLICE_X57Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffd5c000000000)
  ) CLBLM_R_X37Y122_SLICE_X57Y122_BLUT (
.I0(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.I1(CLBLM_R_X35Y122_SLICE_X52Y122_D_XOR),
.I2(CLBLL_L_X36Y122_SLICE_X55Y122_AO6),
.I3(CLBLM_R_X35Y124_SLICE_X53Y124_D_XOR),
.I4(CLBLM_R_X37Y122_SLICE_X57Y122_CO6),
.I5(LIOB33_X0Y147_IOB_X0Y148_I),
.O5(CLBLM_R_X37Y122_SLICE_X57Y122_BO5),
.O6(CLBLM_R_X37Y122_SLICE_X57Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffefff8fff0fff0)
  ) CLBLM_R_X37Y122_SLICE_X57Y122_ALUT (
.I0(LIOB33_X0Y131_IOB_X0Y131_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(CLBLM_R_X37Y122_SLICE_X56Y122_AO6),
.I3(CLBLM_R_X37Y119_SLICE_X56Y119_AO6),
.I4(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I5(CLBLL_L_X36Y116_SLICE_X55Y116_AO5),
.O5(CLBLM_R_X37Y122_SLICE_X57Y122_AO5),
.O6(CLBLM_R_X37Y122_SLICE_X57Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe04ff05fe04fa00)
  ) CLBLM_R_X37Y123_SLICE_X56Y123_DLUT (
.I0(LIOB33_X0Y117_IOB_X0Y118_I),
.I1(RIOB33_X105Y115_IOB_X1Y116_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(RIOB33_X105Y117_IOB_X1Y117_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_R_X37Y123_SLICE_X56Y123_DO5),
.O6(CLBLM_R_X37Y123_SLICE_X56Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff05fe04fa00fe04)
  ) CLBLM_R_X37Y123_SLICE_X56Y123_CLUT (
.I0(LIOB33_X0Y117_IOB_X0Y118_I),
.I1(RIOB33_X105Y111_IOB_X1Y111_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(RIOB33_X105Y117_IOB_X1Y117_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(RIOB33_X105Y115_IOB_X1Y115_I),
.O5(CLBLM_R_X37Y123_SLICE_X56Y123_CO5),
.O6(CLBLM_R_X37Y123_SLICE_X56Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffef8f0f0)
  ) CLBLM_R_X37Y123_SLICE_X56Y123_BLUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I2(CLBLL_L_X36Y123_SLICE_X54Y123_BO6),
.I3(LIOB33_X0Y135_IOB_X0Y135_I),
.I4(CLBLL_L_X36Y116_SLICE_X55Y116_AO5),
.I5(CLBLL_L_X36Y123_SLICE_X55Y123_AO6),
.O5(CLBLM_R_X37Y123_SLICE_X56Y123_BO5),
.O6(CLBLM_R_X37Y123_SLICE_X56Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffa880)
  ) CLBLM_R_X37Y123_SLICE_X56Y123_ALUT (
.I0(CLBLL_L_X36Y116_SLICE_X55Y116_AO5),
.I1(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(LIOB33_X0Y131_IOB_X0Y132_I),
.I4(CLBLL_L_X36Y122_SLICE_X55Y122_CO6),
.I5(CLBLM_R_X37Y120_SLICE_X56Y120_AO6),
.O5(CLBLM_R_X37Y123_SLICE_X56Y123_AO5),
.O6(CLBLM_R_X37Y123_SLICE_X56Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa55aa55cccc3333)
  ) CLBLM_R_X37Y123_SLICE_X57Y123_DLUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(LIOB33_X0Y131_IOB_X0Y132_I),
.I4(LIOB33_X0Y133_IOB_X0Y133_I),
.I5(1'b1),
.O5(CLBLM_R_X37Y123_SLICE_X57Y123_DO5),
.O6(CLBLM_R_X37Y123_SLICE_X57Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc030e2f0c0fce2f0)
  ) CLBLM_R_X37Y123_SLICE_X57Y123_CLUT (
.I0(CLBLM_R_X35Y122_SLICE_X52Y122_D_XOR),
.I1(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I2(CLBLM_R_X35Y124_SLICE_X53Y124_D_XOR),
.I3(LIOB33_X0Y147_IOB_X0Y147_I),
.I4(LIOB33_X0Y145_IOB_X0Y146_I),
.I5(CLBLM_R_X37Y123_SLICE_X57Y123_DO5),
.O5(CLBLM_R_X37Y123_SLICE_X57Y123_CO5),
.O6(CLBLM_R_X37Y123_SLICE_X57Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd1d1c0c070f870f8)
  ) CLBLM_R_X37Y123_SLICE_X57Y123_BLUT (
.I0(LIOB33_X0Y145_IOB_X0Y146_I),
.I1(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I2(CLBLM_R_X35Y124_SLICE_X53Y124_C_XOR),
.I3(CLBLM_R_X37Y123_SLICE_X57Y123_DO6),
.I4(CLBLM_R_X35Y122_SLICE_X52Y122_C_XOR),
.I5(LIOB33_X0Y147_IOB_X0Y147_I),
.O5(CLBLM_R_X37Y123_SLICE_X57Y123_BO5),
.O6(CLBLM_R_X37Y123_SLICE_X57Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffef0fffff8f0)
  ) CLBLM_R_X37Y123_SLICE_X57Y123_ALUT (
.I0(LIOB33_X0Y133_IOB_X0Y133_I),
.I1(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I2(CLBLM_R_X37Y122_SLICE_X57Y122_BO6),
.I3(CLBLL_L_X36Y116_SLICE_X55Y116_AO5),
.I4(CLBLM_R_X37Y120_SLICE_X56Y120_BO6),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X37Y123_SLICE_X57Y123_AO5),
.O6(CLBLM_R_X37Y123_SLICE_X57Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000400)
  ) CLBLM_R_X37Y124_SLICE_X56Y124_DLUT (
.I0(CLBLL_L_X36Y122_SLICE_X54Y122_BO6),
.I1(CLBLM_R_X37Y121_SLICE_X56Y121_CO6),
.I2(CLBLM_R_X35Y119_SLICE_X53Y119_AO6),
.I3(CLBLM_R_X37Y124_SLICE_X56Y124_CO6),
.I4(CLBLM_R_X33Y123_SLICE_X49Y123_AO6),
.I5(CLBLM_R_X33Y121_SLICE_X48Y121_AO6),
.O5(CLBLM_R_X37Y124_SLICE_X56Y124_DO5),
.O6(CLBLM_R_X37Y124_SLICE_X56Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000ff00ab)
  ) CLBLM_R_X37Y124_SLICE_X56Y124_CLUT (
.I0(CLBLM_R_X37Y124_SLICE_X57Y124_BO6),
.I1(CLBLM_R_X37Y124_SLICE_X57Y124_AO6),
.I2(CLBLM_R_X37Y120_SLICE_X56Y120_AO6),
.I3(CLBLL_L_X36Y120_SLICE_X55Y120_BO6),
.I4(CLBLM_R_X37Y120_SLICE_X56Y120_BO6),
.I5(CLBLL_L_X38Y124_SLICE_X58Y124_AO6),
.O5(CLBLM_R_X37Y124_SLICE_X56Y124_CO5),
.O6(CLBLM_R_X37Y124_SLICE_X56Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff007d2800000000)
  ) CLBLM_R_X37Y124_SLICE_X56Y124_BLUT (
.I0(LIOB33_X0Y145_IOB_X0Y146_I),
.I1(LIOB33_X0Y133_IOB_X0Y134_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(CLBLM_R_X35Y125_SLICE_X53Y125_A_XOR),
.I4(LIOB33_X0Y147_IOB_X0Y147_I),
.I5(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.O5(CLBLM_R_X37Y124_SLICE_X56Y124_BO5),
.O6(CLBLM_R_X37Y124_SLICE_X56Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaeaeae00000000)
  ) CLBLM_R_X37Y124_SLICE_X56Y124_ALUT (
.I0(CLBLM_R_X37Y124_SLICE_X56Y124_BO6),
.I1(CLBLM_R_X35Y125_SLICE_X53Y125_A_XOR),
.I2(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.I3(CLBLM_R_X35Y123_SLICE_X52Y123_A_XOR),
.I4(CLBLL_L_X36Y122_SLICE_X55Y122_AO6),
.I5(LIOB33_X0Y147_IOB_X0Y148_I),
.O5(CLBLM_R_X37Y124_SLICE_X56Y124_AO5),
.O6(CLBLM_R_X37Y124_SLICE_X56Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y124_SLICE_X57Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y124_SLICE_X57Y124_DO5),
.O6(CLBLM_R_X37Y124_SLICE_X57Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y124_SLICE_X57Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y124_SLICE_X57Y124_CO5),
.O6(CLBLM_R_X37Y124_SLICE_X57Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00000e080e08)
  ) CLBLM_R_X37Y124_SLICE_X57Y124_BLUT (
.I0(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I1(LIOB33_X0Y133_IOB_X0Y133_I),
.I2(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X37Y123_SLICE_X57Y123_CO6),
.I5(LIOB33_X0Y147_IOB_X0Y148_I),
.O5(CLBLM_R_X37Y124_SLICE_X57Y124_BO5),
.O6(CLBLM_R_X37Y124_SLICE_X57Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa0000fcc0)
  ) CLBLM_R_X37Y124_SLICE_X57Y124_ALUT (
.I0(CLBLM_R_X37Y123_SLICE_X57Y123_BO6),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I3(LIOB33_X0Y131_IOB_X0Y132_I),
.I4(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.I5(LIOB33_X0Y147_IOB_X0Y148_I),
.O5(CLBLM_R_X37Y124_SLICE_X57Y124_AO5),
.O6(CLBLM_R_X37Y124_SLICE_X57Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdf8adf8fd580d080)
  ) CLBLM_R_X37Y125_SLICE_X56Y125_DLUT (
.I0(LIOB33_X0Y147_IOB_X0Y147_I),
.I1(CLBLL_L_X36Y124_SLICE_X54Y124_DO6),
.I2(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I3(CLBLL_L_X36Y123_SLICE_X54Y123_DO6),
.I4(LIOB33_X0Y145_IOB_X0Y146_I),
.I5(CLBLM_R_X35Y125_SLICE_X53Y125_D_XOR),
.O5(CLBLM_R_X37Y125_SLICE_X56Y125_DO5),
.O6(CLBLM_R_X37Y125_SLICE_X56Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2300000020000000)
  ) CLBLM_R_X37Y125_SLICE_X56Y125_CLUT (
.I0(RIOB33_X105Y117_IOB_X1Y117_I),
.I1(LIOB33_X0Y145_IOB_X0Y146_I),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(CLBLL_L_X36Y121_SLICE_X54Y121_AO5),
.I4(CLBLL_L_X36Y116_SLICE_X54Y116_BO5),
.I5(RIOB33_X105Y115_IOB_X1Y116_I),
.O5(CLBLM_R_X37Y125_SLICE_X56Y125_CO5),
.O6(CLBLM_R_X37Y125_SLICE_X56Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000003200000010)
  ) CLBLM_R_X37Y125_SLICE_X56Y125_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(RIOB33_X105Y113_IOB_X1Y114_I),
.I3(LIOB33_X0Y117_IOB_X0Y118_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(RIOB33_X105Y115_IOB_X1Y116_I),
.O5(CLBLM_R_X37Y125_SLICE_X56Y125_BO5),
.O6(CLBLM_R_X37Y125_SLICE_X56Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffefefcfcfcfcfc)
  ) CLBLM_R_X37Y125_SLICE_X56Y125_ALUT (
.I0(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I1(CLBLM_R_X37Y124_SLICE_X56Y124_AO6),
.I2(CLBLL_L_X36Y120_SLICE_X55Y120_BO6),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(LIOB33_X0Y133_IOB_X0Y134_I),
.I5(CLBLL_L_X36Y116_SLICE_X55Y116_AO5),
.O5(CLBLM_R_X37Y125_SLICE_X56Y125_AO5),
.O6(CLBLM_R_X37Y125_SLICE_X56Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hef004f00e0004000)
  ) CLBLM_R_X37Y125_SLICE_X57Y125_DLUT (
.I0(LIOB33_X0Y147_IOB_X0Y147_I),
.I1(CLBLL_L_X36Y123_SLICE_X54Y123_DO6),
.I2(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I3(CLBLL_L_X34Y128_SLICE_X50Y128_AO6),
.I4(CLBLL_L_X36Y124_SLICE_X54Y124_DO6),
.I5(CLBLM_R_X35Y125_SLICE_X53Y125_D_XOR),
.O5(CLBLM_R_X37Y125_SLICE_X57Y125_DO5),
.O6(CLBLM_R_X37Y125_SLICE_X57Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbffb044000000000)
  ) CLBLM_R_X37Y125_SLICE_X57Y125_CLUT (
.I0(LIOB33_X0Y147_IOB_X0Y147_I),
.I1(LIOB33_X0Y145_IOB_X0Y146_I),
.I2(LIOB33_X0Y135_IOB_X0Y136_I),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(CLBLM_R_X35Y125_SLICE_X53Y125_C_XOR),
.I5(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.O5(CLBLM_R_X37Y125_SLICE_X57Y125_CO5),
.O6(CLBLM_R_X37Y125_SLICE_X57Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000c0ea0000)
  ) CLBLM_R_X37Y125_SLICE_X57Y125_BLUT (
.I0(CLBLM_R_X35Y125_SLICE_X53Y125_C_XOR),
.I1(CLBLL_L_X36Y122_SLICE_X55Y122_AO6),
.I2(CLBLM_R_X35Y123_SLICE_X52Y123_C_XOR),
.I3(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.I4(LIOB33_X0Y147_IOB_X0Y148_I),
.I5(CLBLM_R_X37Y125_SLICE_X57Y125_CO6),
.O5(CLBLM_R_X37Y125_SLICE_X57Y125_BO5),
.O6(CLBLM_R_X37Y125_SLICE_X57Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffe8ffffff00)
  ) CLBLM_R_X37Y125_SLICE_X57Y125_ALUT (
.I0(LIOB33_X0Y135_IOB_X0Y136_I),
.I1(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(CLBLM_R_X37Y125_SLICE_X57Y125_BO6),
.I4(CLBLL_L_X36Y124_SLICE_X55Y124_AO6),
.I5(CLBLL_L_X36Y116_SLICE_X55Y116_AO5),
.O5(CLBLM_R_X37Y125_SLICE_X57Y125_AO5),
.O6(CLBLM_R_X37Y125_SLICE_X57Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffc00000030)
  ) CLBLM_R_X37Y126_SLICE_X56Y126_DLUT (
.I0(1'b1),
.I1(LIOB33_X0Y117_IOB_X0Y118_I),
.I2(RIOB33_X105Y113_IOB_X1Y114_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(RIOB33_X105Y117_IOB_X1Y117_I),
.O5(CLBLM_R_X37Y126_SLICE_X56Y126_DO5),
.O6(CLBLM_R_X37Y126_SLICE_X56Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdeccccc00000000)
  ) CLBLM_R_X37Y126_SLICE_X56Y126_CLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(CLBLM_R_X37Y125_SLICE_X56Y125_CO6),
.I2(CLBLL_L_X34Y127_SLICE_X50Y127_AO6),
.I3(CLBLL_L_X34Y126_SLICE_X50Y126_DO6),
.I4(LIOB33_X0Y145_IOB_X0Y146_I),
.I5(CLBLL_L_X36Y122_SLICE_X55Y122_AO5),
.O5(CLBLM_R_X37Y126_SLICE_X56Y126_CO5),
.O6(CLBLM_R_X37Y126_SLICE_X56Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff00ffffba00)
  ) CLBLM_R_X37Y126_SLICE_X56Y126_BLUT (
.I0(CLBLM_R_X37Y127_SLICE_X56Y127_CO6),
.I1(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I2(CLBLM_R_X35Y127_SLICE_X53Y127_C_XOR),
.I3(CLBLL_L_X34Y128_SLICE_X50Y128_AO6),
.I4(CLBLM_R_X35Y128_SLICE_X52Y128_AO6),
.I5(CLBLM_R_X37Y126_SLICE_X56Y126_CO6),
.O5(CLBLM_R_X37Y126_SLICE_X56Y126_BO5),
.O6(CLBLM_R_X37Y126_SLICE_X56Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaff00f0f0aaaa)
  ) CLBLM_R_X37Y126_SLICE_X56Y126_ALUT (
.I0(CLBLM_R_X37Y126_SLICE_X56Y126_DO6),
.I1(1'b1),
.I2(CLBLM_R_X37Y126_SLICE_X57Y126_CO6),
.I3(CLBLM_R_X37Y123_SLICE_X56Y123_DO6),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(1'b1),
.O5(CLBLM_R_X37Y126_SLICE_X56Y126_AO5),
.O6(CLBLM_R_X37Y126_SLICE_X56Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc33333333)
  ) CLBLM_R_X37Y126_SLICE_X57Y126_DLUT (
.I0(1'b1),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y137_IOB_X0Y137_I),
.O5(CLBLM_R_X37Y126_SLICE_X57Y126_DO5),
.O6(CLBLM_R_X37Y126_SLICE_X57Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffa00000500)
  ) CLBLM_R_X37Y126_SLICE_X57Y126_CLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(1'b1),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(RIOB33_X105Y115_IOB_X1Y116_I),
.I4(LIOB33_X0Y117_IOB_X0Y118_I),
.I5(RIOB33_X105Y117_IOB_X1Y117_I),
.O5(CLBLM_R_X37Y126_SLICE_X57Y126_CO5),
.O6(CLBLM_R_X37Y126_SLICE_X57Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcf03cc007f407f40)
  ) CLBLM_R_X37Y126_SLICE_X57Y126_BLUT (
.I0(CLBLM_R_X37Y126_SLICE_X57Y126_DO6),
.I1(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I2(LIOB33_X0Y145_IOB_X0Y146_I),
.I3(CLBLM_R_X35Y125_SLICE_X53Y125_D_XOR),
.I4(CLBLM_R_X35Y123_SLICE_X52Y123_D_XOR),
.I5(LIOB33_X0Y147_IOB_X0Y147_I),
.O5(CLBLM_R_X37Y126_SLICE_X57Y126_BO5),
.O6(CLBLM_R_X37Y126_SLICE_X57Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0054544040)
  ) CLBLM_R_X37Y126_SLICE_X57Y126_ALUT (
.I0(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.I1(CLBLL_L_X34Y127_SLICE_X50Y127_DO6),
.I2(RIOB33_X105Y109_IOB_X1Y109_I),
.I3(CLBLM_R_X37Y126_SLICE_X57Y126_BO6),
.I4(LIOB33_X0Y137_IOB_X0Y137_I),
.I5(LIOB33_X0Y147_IOB_X0Y148_I),
.O5(CLBLM_R_X37Y126_SLICE_X57Y126_AO5),
.O6(CLBLM_R_X37Y126_SLICE_X57Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000055550515)
  ) CLBLM_R_X37Y127_SLICE_X56Y127_DLUT (
.I0(CLBLM_R_X37Y126_SLICE_X57Y126_AO6),
.I1(CLBLM_R_X37Y125_SLICE_X56Y125_DO6),
.I2(CLBLL_L_X34Y129_SLICE_X50Y129_AO6),
.I3(CLBLL_L_X36Y127_SLICE_X55Y127_BO6),
.I4(LIOB33_X0Y147_IOB_X0Y148_I),
.I5(CLBLM_R_X35Y128_SLICE_X52Y128_CO6),
.O5(CLBLM_R_X37Y127_SLICE_X56Y127_DO5),
.O6(CLBLM_R_X37Y127_SLICE_X56Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa30000aca00000)
  ) CLBLM_R_X37Y127_SLICE_X56Y127_CLUT (
.I0(CLBLM_R_X35Y127_SLICE_X53Y127_C_XOR),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(LIOB33_X0Y145_IOB_X0Y146_I),
.I3(RIOB33_X105Y117_IOB_X1Y117_I),
.I4(CLBLL_L_X36Y116_SLICE_X55Y116_AO6),
.I5(CLBLM_R_X37Y127_SLICE_X56Y127_BO6),
.O5(CLBLM_R_X37Y127_SLICE_X56Y127_CO5),
.O6(CLBLM_R_X37Y127_SLICE_X56Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0001fffe0000)
  ) CLBLM_R_X37Y127_SLICE_X56Y127_BLUT (
.I0(LIOB33_X0Y117_IOB_X0Y118_I),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(RIOB33_X105Y117_IOB_X1Y117_I),
.I5(RIOB33_X105Y115_IOB_X1Y116_I),
.O5(CLBLM_R_X37Y127_SLICE_X56Y127_BO5),
.O6(CLBLM_R_X37Y127_SLICE_X56Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000005040100)
  ) CLBLM_R_X37Y127_SLICE_X56Y127_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y118_I),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(RIOB33_X105Y115_IOB_X1Y115_I),
.I4(RIOB33_X105Y117_IOB_X1Y117_I),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X37Y127_SLICE_X56Y127_AO5),
.O6(CLBLM_R_X37Y127_SLICE_X56Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y127_SLICE_X57Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y127_SLICE_X57Y127_DO5),
.O6(CLBLM_R_X37Y127_SLICE_X57Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y127_SLICE_X57Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y127_SLICE_X57Y127_CO5),
.O6(CLBLM_R_X37Y127_SLICE_X57Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y127_SLICE_X57Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y127_SLICE_X57Y127_BO5),
.O6(CLBLM_R_X37Y127_SLICE_X57Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y127_SLICE_X57Y127_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y127_SLICE_X57Y127_AO5),
.O6(CLBLM_R_X37Y127_SLICE_X57Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y128_SLICE_X56Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y128_SLICE_X56Y128_DO5),
.O6(CLBLM_R_X37Y128_SLICE_X56Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y128_SLICE_X56Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y128_SLICE_X56Y128_CO5),
.O6(CLBLM_R_X37Y128_SLICE_X56Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y128_SLICE_X56Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y128_SLICE_X56Y128_BO5),
.O6(CLBLM_R_X37Y128_SLICE_X56Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000002000000000)
  ) CLBLM_R_X37Y128_SLICE_X56Y128_ALUT (
.I0(CLBLL_L_X36Y128_SLICE_X55Y128_CO6),
.I1(CLBLL_L_X36Y127_SLICE_X54Y127_BO6),
.I2(CLBLL_L_X36Y128_SLICE_X55Y128_BO6),
.I3(CLBLM_R_X35Y126_SLICE_X52Y126_BO6),
.I4(CLBLL_L_X36Y127_SLICE_X54Y127_AO6),
.I5(CLBLM_R_X37Y127_SLICE_X56Y127_DO6),
.O5(CLBLM_R_X37Y128_SLICE_X56Y128_AO5),
.O6(CLBLM_R_X37Y128_SLICE_X56Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y128_SLICE_X57Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y128_SLICE_X57Y128_DO5),
.O6(CLBLM_R_X37Y128_SLICE_X57Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y128_SLICE_X57Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y128_SLICE_X57Y128_CO5),
.O6(CLBLM_R_X37Y128_SLICE_X57Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y128_SLICE_X57Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y128_SLICE_X57Y128_BO5),
.O6(CLBLM_R_X37Y128_SLICE_X57Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y128_SLICE_X57Y128_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y128_SLICE_X57Y128_AO5),
.O6(CLBLM_R_X37Y128_SLICE_X57Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12.0"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y65_IOB_X0Y65_OBUF (
.I(CLBLL_L_X34Y115_SLICE_X51Y115_AO6),
.O(result[0])
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y101_IOB_X0Y101_IBUF (
.I(op1[1]),
.O(LIOB33_X0Y101_IOB_X0Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y101_IOB_X0Y102_IBUF (
.I(op1[2]),
.O(LIOB33_X0Y101_IOB_X0Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y103_IOB_X0Y103_IBUF (
.I(op1[3]),
.O(LIOB33_X0Y103_IOB_X0Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y103_IOB_X0Y104_IBUF (
.I(op1[4]),
.O(LIOB33_X0Y103_IOB_X0Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y105_IOB_X0Y105_IBUF (
.I(op1[5]),
.O(LIOB33_X0Y105_IOB_X0Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y105_IOB_X0Y106_IBUF (
.I(op1[6]),
.O(LIOB33_X0Y105_IOB_X0Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y107_IOB_X0Y107_IBUF (
.I(op1[7]),
.O(LIOB33_X0Y107_IOB_X0Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y107_IOB_X0Y108_IBUF (
.I(op1[8]),
.O(LIOB33_X0Y107_IOB_X0Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y109_IOB_X0Y109_IBUF (
.I(op1[9]),
.O(LIOB33_X0Y109_IOB_X0Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y109_IOB_X0Y110_IBUF (
.I(op1[10]),
.O(LIOB33_X0Y109_IOB_X0Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y111_IOB_X0Y111_IBUF (
.I(op1[11]),
.O(LIOB33_X0Y111_IOB_X0Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y111_IOB_X0Y112_IBUF (
.I(op1[12]),
.O(LIOB33_X0Y111_IOB_X0Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y113_IOB_X0Y113_IBUF (
.I(op1[13]),
.O(LIOB33_X0Y113_IOB_X0Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y113_IOB_X0Y114_IBUF (
.I(op2[0]),
.O(LIOB33_X0Y113_IOB_X0Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y115_IOB_X0Y115_IBUF (
.I(op2[1]),
.O(LIOB33_X0Y115_IOB_X0Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y115_IOB_X0Y116_IBUF (
.I(op2[2]),
.O(LIOB33_X0Y115_IOB_X0Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y117_IOB_X0Y117_IBUF (
.I(op2[3]),
.O(LIOB33_X0Y117_IOB_X0Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y117_IOB_X0Y118_IBUF (
.I(op2[4]),
.O(LIOB33_X0Y117_IOB_X0Y118_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y119_IOB_X0Y119_IBUF (
.I(op2[5]),
.O(LIOB33_X0Y119_IOB_X0Y119_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y119_IOB_X0Y120_IBUF (
.I(op2[6]),
.O(LIOB33_X0Y119_IOB_X0Y120_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y121_IOB_X0Y121_IBUF (
.I(op2[7]),
.O(LIOB33_X0Y121_IOB_X0Y121_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y121_IOB_X0Y122_IBUF (
.I(op2[8]),
.O(LIOB33_X0Y121_IOB_X0Y122_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y123_IOB_X0Y123_IBUF (
.I(op2[9]),
.O(LIOB33_X0Y123_IOB_X0Y123_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y123_IOB_X0Y124_IBUF (
.I(op2[10]),
.O(LIOB33_X0Y123_IOB_X0Y124_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y125_IOB_X0Y125_IBUF (
.I(op2[11]),
.O(LIOB33_X0Y125_IOB_X0Y125_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y125_IOB_X0Y126_IBUF (
.I(op2[12]),
.O(LIOB33_X0Y125_IOB_X0Y126_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y127_IOB_X0Y127_IBUF (
.I(op2[13]),
.O(LIOB33_X0Y127_IOB_X0Y127_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y127_IOB_X0Y128_IBUF (
.I(op2[14]),
.O(LIOB33_X0Y127_IOB_X0Y128_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y129_IOB_X0Y129_IBUF (
.I(op2[15]),
.O(LIOB33_X0Y129_IOB_X0Y129_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y129_IOB_X0Y130_IBUF (
.I(op2[16]),
.O(LIOB33_X0Y129_IOB_X0Y130_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y131_IOB_X0Y131_IBUF (
.I(op2[17]),
.O(LIOB33_X0Y131_IOB_X0Y131_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y131_IOB_X0Y132_IBUF (
.I(op2[18]),
.O(LIOB33_X0Y131_IOB_X0Y132_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y133_IOB_X0Y133_IBUF (
.I(op2[19]),
.O(LIOB33_X0Y133_IOB_X0Y133_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y133_IOB_X0Y134_IBUF (
.I(op2[20]),
.O(LIOB33_X0Y133_IOB_X0Y134_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y135_IOB_X0Y135_IBUF (
.I(op2[21]),
.O(LIOB33_X0Y135_IOB_X0Y135_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y135_IOB_X0Y136_IBUF (
.I(op2[22]),
.O(LIOB33_X0Y135_IOB_X0Y136_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y137_IOB_X0Y137_IBUF (
.I(op2[23]),
.O(LIOB33_X0Y137_IOB_X0Y137_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y137_IOB_X0Y138_IBUF (
.I(op2[24]),
.O(LIOB33_X0Y137_IOB_X0Y138_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y139_IOB_X0Y139_IBUF (
.I(op2[25]),
.O(LIOB33_X0Y139_IOB_X0Y139_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y139_IOB_X0Y140_IBUF (
.I(op2[26]),
.O(LIOB33_X0Y139_IOB_X0Y140_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y141_IOB_X0Y141_IBUF (
.I(op2[27]),
.O(LIOB33_X0Y141_IOB_X0Y141_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y141_IOB_X0Y142_IBUF (
.I(op2[28]),
.O(LIOB33_X0Y141_IOB_X0Y142_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y143_IOB_X0Y143_IBUF (
.I(op2[29]),
.O(LIOB33_X0Y143_IOB_X0Y143_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y143_IOB_X0Y144_IBUF (
.I(op2[30]),
.O(LIOB33_X0Y143_IOB_X0Y144_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y145_IOB_X0Y145_IBUF (
.I(op2[31]),
.O(LIOB33_X0Y145_IOB_X0Y145_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y145_IOB_X0Y146_IBUF (
.I(alu_op[0]),
.O(LIOB33_X0Y145_IOB_X0Y146_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y147_IOB_X0Y147_IBUF (
.I(alu_op[1]),
.O(LIOB33_X0Y147_IOB_X0Y147_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y147_IOB_X0Y148_IBUF (
.I(alu_op[2]),
.O(LIOB33_X0Y147_IOB_X0Y148_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_SING_X0Y100_IOB_X0Y100_IBUF (
.I(op1[0]),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_SING_X0Y149_IOB_X0Y149_IBUF (
.I(alu_op[3]),
.O(LIOB33_SING_X0Y149_IOB_X0Y149_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X105Y101_IOB_X1Y101_IBUF (
.I(op1[15]),
.O(RIOB33_X105Y101_IOB_X1Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X105Y101_IOB_X1Y102_IBUF (
.I(op1[16]),
.O(RIOB33_X105Y101_IOB_X1Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X105Y103_IOB_X1Y103_IBUF (
.I(op1[17]),
.O(RIOB33_X105Y103_IOB_X1Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X105Y103_IOB_X1Y104_IBUF (
.I(op1[18]),
.O(RIOB33_X105Y103_IOB_X1Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X105Y105_IOB_X1Y105_IBUF (
.I(op1[19]),
.O(RIOB33_X105Y105_IOB_X1Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X105Y105_IOB_X1Y106_IBUF (
.I(op1[20]),
.O(RIOB33_X105Y105_IOB_X1Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X105Y107_IOB_X1Y107_IBUF (
.I(op1[21]),
.O(RIOB33_X105Y107_IOB_X1Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X105Y107_IOB_X1Y108_IBUF (
.I(op1[22]),
.O(RIOB33_X105Y107_IOB_X1Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X105Y109_IOB_X1Y109_IBUF (
.I(op1[23]),
.O(RIOB33_X105Y109_IOB_X1Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X105Y109_IOB_X1Y110_IBUF (
.I(op1[24]),
.O(RIOB33_X105Y109_IOB_X1Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X105Y111_IOB_X1Y111_IBUF (
.I(op1[25]),
.O(RIOB33_X105Y111_IOB_X1Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X105Y111_IOB_X1Y112_IBUF (
.I(op1[26]),
.O(RIOB33_X105Y111_IOB_X1Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X105Y113_IOB_X1Y113_IBUF (
.I(op1[27]),
.O(RIOB33_X105Y113_IOB_X1Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X105Y113_IOB_X1Y114_IBUF (
.I(op1[28]),
.O(RIOB33_X105Y113_IOB_X1Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X105Y115_IOB_X1Y115_IBUF (
.I(op1[29]),
.O(RIOB33_X105Y115_IOB_X1Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X105Y115_IOB_X1Y116_IBUF (
.I(op1[30]),
.O(RIOB33_X105Y115_IOB_X1Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X105Y117_IOB_X1Y117_IBUF (
.I(op1[31]),
.O(RIOB33_X105Y117_IOB_X1Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12.0"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X105Y117_IOB_X1Y118_OBUF (
.I(CLBLM_R_X35Y117_SLICE_X53Y117_CO6),
.O(result[1])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12.0"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X105Y119_IOB_X1Y119_OBUF (
.I(CLBLM_R_X33Y116_SLICE_X49Y116_AO6),
.O(result[2])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12.0"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X105Y119_IOB_X1Y120_OBUF (
.I(CLBLM_R_X35Y115_SLICE_X53Y115_AO6),
.O(result[3])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12.0"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X105Y121_IOB_X1Y121_OBUF (
.I(CLBLM_R_X35Y115_SLICE_X52Y115_BO6),
.O(result[4])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12.0"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X105Y121_IOB_X1Y122_OBUF (
.I(CLBLM_R_X35Y116_SLICE_X53Y116_BO6),
.O(result[5])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12.0"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X105Y123_IOB_X1Y123_OBUF (
.I(CLBLL_L_X36Y119_SLICE_X55Y119_BO6),
.O(result[6])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12.0"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X105Y123_IOB_X1Y124_OBUF (
.I(CLBLL_L_X34Y120_SLICE_X51Y120_AO6),
.O(result[7])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12.0"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X105Y125_IOB_X1Y125_OBUF (
.I(CLBLM_R_X33Y121_SLICE_X48Y121_AO6),
.O(result[8])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12.0"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X105Y125_IOB_X1Y126_OBUF (
.I(CLBLL_L_X34Y121_SLICE_X51Y121_AO6),
.O(result[9])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12.0"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X105Y127_IOB_X1Y127_OBUF (
.I(CLBLM_R_X33Y123_SLICE_X49Y123_AO6),
.O(result[10])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12.0"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X105Y127_IOB_X1Y128_OBUF (
.I(CLBLL_L_X36Y122_SLICE_X54Y122_BO6),
.O(result[11])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12.0"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X105Y129_IOB_X1Y129_OBUF (
.I(CLBLL_L_X34Y124_SLICE_X50Y124_AO6),
.O(result[12])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12.0"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X105Y129_IOB_X1Y130_OBUF (
.I(CLBLM_R_X35Y119_SLICE_X53Y119_AO6),
.O(result[13])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12.0"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X105Y131_IOB_X1Y131_OBUF (
.I(CLBLL_L_X36Y121_SLICE_X55Y121_BO6),
.O(result[14])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12.0"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X105Y131_IOB_X1Y132_OBUF (
.I(CLBLL_L_X36Y122_SLICE_X55Y122_BO6),
.O(result[15])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12.0"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X105Y133_IOB_X1Y133_OBUF (
.I(CLBLM_R_X37Y121_SLICE_X57Y121_AO6),
.O(result[16])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12.0"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X105Y133_IOB_X1Y134_OBUF (
.I(CLBLM_R_X37Y122_SLICE_X57Y122_AO6),
.O(result[17])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12.0"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X105Y135_IOB_X1Y135_OBUF (
.I(CLBLM_R_X37Y123_SLICE_X56Y123_AO6),
.O(result[18])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12.0"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X105Y135_IOB_X1Y136_OBUF (
.I(CLBLM_R_X37Y123_SLICE_X57Y123_AO6),
.O(result[19])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12.0"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X105Y137_IOB_X1Y137_OBUF (
.I(CLBLM_R_X37Y125_SLICE_X56Y125_AO6),
.O(result[20])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12.0"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X105Y137_IOB_X1Y138_OBUF (
.I(CLBLM_R_X37Y123_SLICE_X56Y123_BO6),
.O(result[21])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12.0"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X105Y139_IOB_X1Y139_OBUF (
.I(CLBLM_R_X37Y125_SLICE_X57Y125_AO6),
.O(result[22])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12.0"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X105Y139_IOB_X1Y140_OBUF (
.I(CLBLL_L_X38Y126_SLICE_X58Y126_AO6),
.O(result[23])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12.0"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X105Y141_IOB_X1Y141_OBUF (
.I(CLBLL_L_X36Y127_SLICE_X54Y127_AO6),
.O(result[24])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12.0"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X105Y141_IOB_X1Y142_OBUF (
.I(CLBLL_L_X36Y127_SLICE_X54Y127_BO6),
.O(result[25])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12.0"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X105Y143_IOB_X1Y143_OBUF (
.I(CLBLM_R_X35Y126_SLICE_X52Y126_BO6),
.O(result[26])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12.0"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X105Y143_IOB_X1Y144_OBUF (
.I(CLBLL_L_X36Y129_SLICE_X55Y129_AO6),
.O(result[27])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12.0"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X105Y145_IOB_X1Y145_OBUF (
.I(CLBLL_L_X36Y129_SLICE_X54Y129_AO6),
.O(result[28])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12.0"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X105Y145_IOB_X1Y146_OBUF (
.I(CLBLL_L_X36Y128_SLICE_X54Y128_AO6),
.O(result[29])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12.0"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X105Y147_IOB_X1Y147_OBUF (
.I(CLBLM_R_X37Y126_SLICE_X56Y126_BO6),
.O(result[30])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12.0"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X105Y147_IOB_X1Y148_OBUF (
.I(CLBLL_L_X36Y129_SLICE_X55Y129_DO6),
.O(result[31])
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_SING_X105Y100_IOB_X1Y100_IBUF (
.I(op1[14]),
.O(RIOB33_SING_X105Y100_IOB_X1Y100_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12.0"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y149_IOB_X1Y149_OBUF (
.I(CLBLL_L_X38Y126_SLICE_X59Y126_AO6),
.O(zero)
  );
  assign CLBLL_L_X34Y114_SLICE_X50Y114_COUT = CLBLL_L_X34Y114_SLICE_X50Y114_D_CY;
  assign CLBLL_L_X34Y114_SLICE_X50Y114_A = CLBLL_L_X34Y114_SLICE_X50Y114_AO6;
  assign CLBLL_L_X34Y114_SLICE_X50Y114_B = CLBLL_L_X34Y114_SLICE_X50Y114_BO6;
  assign CLBLL_L_X34Y114_SLICE_X50Y114_C = CLBLL_L_X34Y114_SLICE_X50Y114_CO6;
  assign CLBLL_L_X34Y114_SLICE_X50Y114_D = CLBLL_L_X34Y114_SLICE_X50Y114_DO6;
  assign CLBLL_L_X34Y114_SLICE_X51Y114_COUT = CLBLL_L_X34Y114_SLICE_X51Y114_D_CY;
  assign CLBLL_L_X34Y114_SLICE_X51Y114_A = CLBLL_L_X34Y114_SLICE_X51Y114_AO6;
  assign CLBLL_L_X34Y114_SLICE_X51Y114_B = CLBLL_L_X34Y114_SLICE_X51Y114_BO6;
  assign CLBLL_L_X34Y114_SLICE_X51Y114_C = CLBLL_L_X34Y114_SLICE_X51Y114_CO6;
  assign CLBLL_L_X34Y114_SLICE_X51Y114_D = CLBLL_L_X34Y114_SLICE_X51Y114_DO6;
  assign CLBLL_L_X34Y115_SLICE_X50Y115_COUT = CLBLL_L_X34Y115_SLICE_X50Y115_D_CY;
  assign CLBLL_L_X34Y115_SLICE_X50Y115_A = CLBLL_L_X34Y115_SLICE_X50Y115_AO6;
  assign CLBLL_L_X34Y115_SLICE_X50Y115_B = CLBLL_L_X34Y115_SLICE_X50Y115_BO6;
  assign CLBLL_L_X34Y115_SLICE_X50Y115_C = CLBLL_L_X34Y115_SLICE_X50Y115_CO6;
  assign CLBLL_L_X34Y115_SLICE_X50Y115_D = CLBLL_L_X34Y115_SLICE_X50Y115_DO6;
  assign CLBLL_L_X34Y115_SLICE_X50Y115_AMUX = CLBLL_L_X34Y115_SLICE_X50Y115_AO6;
  assign CLBLL_L_X34Y115_SLICE_X51Y115_COUT = CLBLL_L_X34Y115_SLICE_X51Y115_D_CY;
  assign CLBLL_L_X34Y115_SLICE_X51Y115_A = CLBLL_L_X34Y115_SLICE_X51Y115_AO6;
  assign CLBLL_L_X34Y115_SLICE_X51Y115_B = CLBLL_L_X34Y115_SLICE_X51Y115_BO6;
  assign CLBLL_L_X34Y115_SLICE_X51Y115_C = CLBLL_L_X34Y115_SLICE_X51Y115_CO6;
  assign CLBLL_L_X34Y115_SLICE_X51Y115_D = CLBLL_L_X34Y115_SLICE_X51Y115_DO6;
  assign CLBLL_L_X34Y116_SLICE_X50Y116_COUT = CLBLL_L_X34Y116_SLICE_X50Y116_D_CY;
  assign CLBLL_L_X34Y116_SLICE_X50Y116_A = CLBLL_L_X34Y116_SLICE_X50Y116_AO6;
  assign CLBLL_L_X34Y116_SLICE_X50Y116_B = CLBLL_L_X34Y116_SLICE_X50Y116_BO6;
  assign CLBLL_L_X34Y116_SLICE_X50Y116_C = CLBLL_L_X34Y116_SLICE_X50Y116_CO6;
  assign CLBLL_L_X34Y116_SLICE_X50Y116_D = CLBLL_L_X34Y116_SLICE_X50Y116_DO6;
  assign CLBLL_L_X34Y116_SLICE_X50Y116_AMUX = CLBLL_L_X34Y116_SLICE_X50Y116_AO5;
  assign CLBLL_L_X34Y116_SLICE_X51Y116_COUT = CLBLL_L_X34Y116_SLICE_X51Y116_D_CY;
  assign CLBLL_L_X34Y116_SLICE_X51Y116_A = CLBLL_L_X34Y116_SLICE_X51Y116_AO6;
  assign CLBLL_L_X34Y116_SLICE_X51Y116_B = CLBLL_L_X34Y116_SLICE_X51Y116_BO6;
  assign CLBLL_L_X34Y116_SLICE_X51Y116_C = CLBLL_L_X34Y116_SLICE_X51Y116_CO6;
  assign CLBLL_L_X34Y116_SLICE_X51Y116_D = CLBLL_L_X34Y116_SLICE_X51Y116_DO6;
  assign CLBLL_L_X34Y116_SLICE_X51Y116_AMUX = CLBLL_L_X34Y116_SLICE_X51Y116_AO5;
  assign CLBLL_L_X34Y117_SLICE_X50Y117_COUT = CLBLL_L_X34Y117_SLICE_X50Y117_D_CY;
  assign CLBLL_L_X34Y117_SLICE_X50Y117_A = CLBLL_L_X34Y117_SLICE_X50Y117_AO6;
  assign CLBLL_L_X34Y117_SLICE_X50Y117_B = CLBLL_L_X34Y117_SLICE_X50Y117_BO6;
  assign CLBLL_L_X34Y117_SLICE_X50Y117_C = CLBLL_L_X34Y117_SLICE_X50Y117_CO6;
  assign CLBLL_L_X34Y117_SLICE_X50Y117_D = CLBLL_L_X34Y117_SLICE_X50Y117_DO6;
  assign CLBLL_L_X34Y117_SLICE_X51Y117_COUT = CLBLL_L_X34Y117_SLICE_X51Y117_D_CY;
  assign CLBLL_L_X34Y117_SLICE_X51Y117_A = CLBLL_L_X34Y117_SLICE_X51Y117_AO6;
  assign CLBLL_L_X34Y117_SLICE_X51Y117_B = CLBLL_L_X34Y117_SLICE_X51Y117_BO6;
  assign CLBLL_L_X34Y117_SLICE_X51Y117_C = CLBLL_L_X34Y117_SLICE_X51Y117_CO6;
  assign CLBLL_L_X34Y117_SLICE_X51Y117_D = CLBLL_L_X34Y117_SLICE_X51Y117_DO6;
  assign CLBLL_L_X34Y117_SLICE_X51Y117_BMUX = CLBLL_L_X34Y117_SLICE_X51Y117_BO6;
  assign CLBLL_L_X34Y118_SLICE_X50Y118_COUT = CLBLL_L_X34Y118_SLICE_X50Y118_D_CY;
  assign CLBLL_L_X34Y118_SLICE_X50Y118_A = CLBLL_L_X34Y118_SLICE_X50Y118_AO6;
  assign CLBLL_L_X34Y118_SLICE_X50Y118_B = CLBLL_L_X34Y118_SLICE_X50Y118_BO6;
  assign CLBLL_L_X34Y118_SLICE_X50Y118_C = CLBLL_L_X34Y118_SLICE_X50Y118_CO6;
  assign CLBLL_L_X34Y118_SLICE_X50Y118_D = CLBLL_L_X34Y118_SLICE_X50Y118_DO6;
  assign CLBLL_L_X34Y118_SLICE_X51Y118_COUT = CLBLL_L_X34Y118_SLICE_X51Y118_D_CY;
  assign CLBLL_L_X34Y118_SLICE_X51Y118_A = CLBLL_L_X34Y118_SLICE_X51Y118_AO6;
  assign CLBLL_L_X34Y118_SLICE_X51Y118_B = CLBLL_L_X34Y118_SLICE_X51Y118_BO6;
  assign CLBLL_L_X34Y118_SLICE_X51Y118_C = CLBLL_L_X34Y118_SLICE_X51Y118_CO6;
  assign CLBLL_L_X34Y118_SLICE_X51Y118_D = CLBLL_L_X34Y118_SLICE_X51Y118_DO6;
  assign CLBLL_L_X34Y119_SLICE_X50Y119_COUT = CLBLL_L_X34Y119_SLICE_X50Y119_D_CY;
  assign CLBLL_L_X34Y119_SLICE_X50Y119_A = CLBLL_L_X34Y119_SLICE_X50Y119_AO6;
  assign CLBLL_L_X34Y119_SLICE_X50Y119_B = CLBLL_L_X34Y119_SLICE_X50Y119_BO6;
  assign CLBLL_L_X34Y119_SLICE_X50Y119_C = CLBLL_L_X34Y119_SLICE_X50Y119_CO6;
  assign CLBLL_L_X34Y119_SLICE_X50Y119_D = CLBLL_L_X34Y119_SLICE_X50Y119_DO6;
  assign CLBLL_L_X34Y119_SLICE_X51Y119_COUT = CLBLL_L_X34Y119_SLICE_X51Y119_D_CY;
  assign CLBLL_L_X34Y119_SLICE_X51Y119_A = CLBLL_L_X34Y119_SLICE_X51Y119_AO6;
  assign CLBLL_L_X34Y119_SLICE_X51Y119_B = CLBLL_L_X34Y119_SLICE_X51Y119_BO6;
  assign CLBLL_L_X34Y119_SLICE_X51Y119_C = CLBLL_L_X34Y119_SLICE_X51Y119_CO6;
  assign CLBLL_L_X34Y119_SLICE_X51Y119_D = CLBLL_L_X34Y119_SLICE_X51Y119_DO6;
  assign CLBLL_L_X34Y119_SLICE_X51Y119_AMUX = CLBLL_L_X34Y119_SLICE_X51Y119_AO5;
  assign CLBLL_L_X34Y119_SLICE_X51Y119_CMUX = CLBLL_L_X34Y119_SLICE_X51Y119_CO6;
  assign CLBLL_L_X34Y120_SLICE_X50Y120_COUT = CLBLL_L_X34Y120_SLICE_X50Y120_D_CY;
  assign CLBLL_L_X34Y120_SLICE_X50Y120_A = CLBLL_L_X34Y120_SLICE_X50Y120_AO6;
  assign CLBLL_L_X34Y120_SLICE_X50Y120_B = CLBLL_L_X34Y120_SLICE_X50Y120_BO6;
  assign CLBLL_L_X34Y120_SLICE_X50Y120_C = CLBLL_L_X34Y120_SLICE_X50Y120_CO6;
  assign CLBLL_L_X34Y120_SLICE_X50Y120_D = CLBLL_L_X34Y120_SLICE_X50Y120_DO6;
  assign CLBLL_L_X34Y120_SLICE_X51Y120_COUT = CLBLL_L_X34Y120_SLICE_X51Y120_D_CY;
  assign CLBLL_L_X34Y120_SLICE_X51Y120_A = CLBLL_L_X34Y120_SLICE_X51Y120_AO6;
  assign CLBLL_L_X34Y120_SLICE_X51Y120_B = CLBLL_L_X34Y120_SLICE_X51Y120_BO6;
  assign CLBLL_L_X34Y120_SLICE_X51Y120_C = CLBLL_L_X34Y120_SLICE_X51Y120_CO6;
  assign CLBLL_L_X34Y120_SLICE_X51Y120_D = CLBLL_L_X34Y120_SLICE_X51Y120_DO6;
  assign CLBLL_L_X34Y121_SLICE_X50Y121_COUT = CLBLL_L_X34Y121_SLICE_X50Y121_D_CY;
  assign CLBLL_L_X34Y121_SLICE_X50Y121_A = CLBLL_L_X34Y121_SLICE_X50Y121_AO6;
  assign CLBLL_L_X34Y121_SLICE_X50Y121_B = CLBLL_L_X34Y121_SLICE_X50Y121_BO6;
  assign CLBLL_L_X34Y121_SLICE_X50Y121_C = CLBLL_L_X34Y121_SLICE_X50Y121_CO6;
  assign CLBLL_L_X34Y121_SLICE_X50Y121_D = CLBLL_L_X34Y121_SLICE_X50Y121_DO6;
  assign CLBLL_L_X34Y121_SLICE_X51Y121_COUT = CLBLL_L_X34Y121_SLICE_X51Y121_D_CY;
  assign CLBLL_L_X34Y121_SLICE_X51Y121_A = CLBLL_L_X34Y121_SLICE_X51Y121_AO6;
  assign CLBLL_L_X34Y121_SLICE_X51Y121_B = CLBLL_L_X34Y121_SLICE_X51Y121_BO6;
  assign CLBLL_L_X34Y121_SLICE_X51Y121_C = CLBLL_L_X34Y121_SLICE_X51Y121_CO6;
  assign CLBLL_L_X34Y121_SLICE_X51Y121_D = CLBLL_L_X34Y121_SLICE_X51Y121_DO6;
  assign CLBLL_L_X34Y122_SLICE_X50Y122_COUT = CLBLL_L_X34Y122_SLICE_X50Y122_D_CY;
  assign CLBLL_L_X34Y122_SLICE_X50Y122_A = CLBLL_L_X34Y122_SLICE_X50Y122_AO6;
  assign CLBLL_L_X34Y122_SLICE_X50Y122_B = CLBLL_L_X34Y122_SLICE_X50Y122_BO6;
  assign CLBLL_L_X34Y122_SLICE_X50Y122_C = CLBLL_L_X34Y122_SLICE_X50Y122_CO6;
  assign CLBLL_L_X34Y122_SLICE_X50Y122_D = CLBLL_L_X34Y122_SLICE_X50Y122_DO6;
  assign CLBLL_L_X34Y122_SLICE_X51Y122_COUT = CLBLL_L_X34Y122_SLICE_X51Y122_D_CY;
  assign CLBLL_L_X34Y122_SLICE_X51Y122_A = CLBLL_L_X34Y122_SLICE_X51Y122_AO6;
  assign CLBLL_L_X34Y122_SLICE_X51Y122_B = CLBLL_L_X34Y122_SLICE_X51Y122_BO6;
  assign CLBLL_L_X34Y122_SLICE_X51Y122_C = CLBLL_L_X34Y122_SLICE_X51Y122_CO6;
  assign CLBLL_L_X34Y122_SLICE_X51Y122_D = CLBLL_L_X34Y122_SLICE_X51Y122_DO6;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_COUT = CLBLL_L_X34Y123_SLICE_X50Y123_D_CY;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_A = CLBLL_L_X34Y123_SLICE_X50Y123_AO6;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_B = CLBLL_L_X34Y123_SLICE_X50Y123_BO6;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_C = CLBLL_L_X34Y123_SLICE_X50Y123_CO6;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_D = CLBLL_L_X34Y123_SLICE_X50Y123_DO6;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_AMUX = CLBLL_L_X34Y123_SLICE_X50Y123_AO5;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_BMUX = CLBLL_L_X34Y123_SLICE_X50Y123_BO5;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_COUT = CLBLL_L_X34Y123_SLICE_X51Y123_D_CY;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_A = CLBLL_L_X34Y123_SLICE_X51Y123_AO6;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_B = CLBLL_L_X34Y123_SLICE_X51Y123_BO6;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_C = CLBLL_L_X34Y123_SLICE_X51Y123_CO6;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_D = CLBLL_L_X34Y123_SLICE_X51Y123_DO6;
  assign CLBLL_L_X34Y124_SLICE_X50Y124_COUT = CLBLL_L_X34Y124_SLICE_X50Y124_D_CY;
  assign CLBLL_L_X34Y124_SLICE_X50Y124_A = CLBLL_L_X34Y124_SLICE_X50Y124_AO6;
  assign CLBLL_L_X34Y124_SLICE_X50Y124_B = CLBLL_L_X34Y124_SLICE_X50Y124_BO6;
  assign CLBLL_L_X34Y124_SLICE_X50Y124_C = CLBLL_L_X34Y124_SLICE_X50Y124_CO6;
  assign CLBLL_L_X34Y124_SLICE_X50Y124_D = CLBLL_L_X34Y124_SLICE_X50Y124_DO6;
  assign CLBLL_L_X34Y124_SLICE_X50Y124_CMUX = CLBLL_L_X34Y124_SLICE_X50Y124_CO6;
  assign CLBLL_L_X34Y124_SLICE_X51Y124_COUT = CLBLL_L_X34Y124_SLICE_X51Y124_D_CY;
  assign CLBLL_L_X34Y124_SLICE_X51Y124_A = CLBLL_L_X34Y124_SLICE_X51Y124_AO6;
  assign CLBLL_L_X34Y124_SLICE_X51Y124_B = CLBLL_L_X34Y124_SLICE_X51Y124_BO6;
  assign CLBLL_L_X34Y124_SLICE_X51Y124_C = CLBLL_L_X34Y124_SLICE_X51Y124_CO6;
  assign CLBLL_L_X34Y124_SLICE_X51Y124_D = CLBLL_L_X34Y124_SLICE_X51Y124_DO6;
  assign CLBLL_L_X34Y125_SLICE_X50Y125_COUT = CLBLL_L_X34Y125_SLICE_X50Y125_D_CY;
  assign CLBLL_L_X34Y125_SLICE_X50Y125_A = CLBLL_L_X34Y125_SLICE_X50Y125_AO6;
  assign CLBLL_L_X34Y125_SLICE_X50Y125_B = CLBLL_L_X34Y125_SLICE_X50Y125_BO6;
  assign CLBLL_L_X34Y125_SLICE_X50Y125_C = CLBLL_L_X34Y125_SLICE_X50Y125_CO6;
  assign CLBLL_L_X34Y125_SLICE_X50Y125_D = CLBLL_L_X34Y125_SLICE_X50Y125_DO6;
  assign CLBLL_L_X34Y125_SLICE_X51Y125_COUT = CLBLL_L_X34Y125_SLICE_X51Y125_D_CY;
  assign CLBLL_L_X34Y125_SLICE_X51Y125_A = CLBLL_L_X34Y125_SLICE_X51Y125_AO6;
  assign CLBLL_L_X34Y125_SLICE_X51Y125_B = CLBLL_L_X34Y125_SLICE_X51Y125_BO6;
  assign CLBLL_L_X34Y125_SLICE_X51Y125_C = CLBLL_L_X34Y125_SLICE_X51Y125_CO6;
  assign CLBLL_L_X34Y125_SLICE_X51Y125_D = CLBLL_L_X34Y125_SLICE_X51Y125_DO6;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_COUT = CLBLL_L_X34Y126_SLICE_X50Y126_D_CY;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_A = CLBLL_L_X34Y126_SLICE_X50Y126_AO6;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_B = CLBLL_L_X34Y126_SLICE_X50Y126_BO6;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_C = CLBLL_L_X34Y126_SLICE_X50Y126_CO6;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_D = CLBLL_L_X34Y126_SLICE_X50Y126_DO6;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_COUT = CLBLL_L_X34Y126_SLICE_X51Y126_D_CY;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_A = CLBLL_L_X34Y126_SLICE_X51Y126_AO6;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_B = CLBLL_L_X34Y126_SLICE_X51Y126_BO6;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_C = CLBLL_L_X34Y126_SLICE_X51Y126_CO6;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_D = CLBLL_L_X34Y126_SLICE_X51Y126_DO6;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_DMUX = CLBLL_L_X34Y126_SLICE_X51Y126_D_CY;
  assign CLBLL_L_X34Y127_SLICE_X50Y127_COUT = CLBLL_L_X34Y127_SLICE_X50Y127_D_CY;
  assign CLBLL_L_X34Y127_SLICE_X50Y127_A = CLBLL_L_X34Y127_SLICE_X50Y127_AO6;
  assign CLBLL_L_X34Y127_SLICE_X50Y127_B = CLBLL_L_X34Y127_SLICE_X50Y127_BO6;
  assign CLBLL_L_X34Y127_SLICE_X50Y127_C = CLBLL_L_X34Y127_SLICE_X50Y127_CO6;
  assign CLBLL_L_X34Y127_SLICE_X50Y127_D = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLL_L_X34Y127_SLICE_X51Y127_COUT = CLBLL_L_X34Y127_SLICE_X51Y127_D_CY;
  assign CLBLL_L_X34Y127_SLICE_X51Y127_A = CLBLL_L_X34Y127_SLICE_X51Y127_AO6;
  assign CLBLL_L_X34Y127_SLICE_X51Y127_B = CLBLL_L_X34Y127_SLICE_X51Y127_BO6;
  assign CLBLL_L_X34Y127_SLICE_X51Y127_C = CLBLL_L_X34Y127_SLICE_X51Y127_CO6;
  assign CLBLL_L_X34Y127_SLICE_X51Y127_D = CLBLL_L_X34Y127_SLICE_X51Y127_DO6;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_COUT = CLBLL_L_X34Y128_SLICE_X50Y128_D_CY;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_A = CLBLL_L_X34Y128_SLICE_X50Y128_AO6;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_B = CLBLL_L_X34Y128_SLICE_X50Y128_BO6;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_C = CLBLL_L_X34Y128_SLICE_X50Y128_CO6;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_D = CLBLL_L_X34Y128_SLICE_X50Y128_DO6;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_COUT = CLBLL_L_X34Y128_SLICE_X51Y128_D_CY;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_A = CLBLL_L_X34Y128_SLICE_X51Y128_AO6;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_B = CLBLL_L_X34Y128_SLICE_X51Y128_BO6;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_C = CLBLL_L_X34Y128_SLICE_X51Y128_CO6;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_D = CLBLL_L_X34Y128_SLICE_X51Y128_DO6;
  assign CLBLL_L_X34Y129_SLICE_X50Y129_COUT = CLBLL_L_X34Y129_SLICE_X50Y129_D_CY;
  assign CLBLL_L_X34Y129_SLICE_X50Y129_A = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLL_L_X34Y129_SLICE_X50Y129_B = CLBLL_L_X34Y129_SLICE_X50Y129_BO6;
  assign CLBLL_L_X34Y129_SLICE_X50Y129_C = CLBLL_L_X34Y129_SLICE_X50Y129_CO6;
  assign CLBLL_L_X34Y129_SLICE_X50Y129_D = CLBLL_L_X34Y129_SLICE_X50Y129_DO6;
  assign CLBLL_L_X34Y129_SLICE_X51Y129_COUT = CLBLL_L_X34Y129_SLICE_X51Y129_D_CY;
  assign CLBLL_L_X34Y129_SLICE_X51Y129_A = CLBLL_L_X34Y129_SLICE_X51Y129_AO6;
  assign CLBLL_L_X34Y129_SLICE_X51Y129_B = CLBLL_L_X34Y129_SLICE_X51Y129_BO6;
  assign CLBLL_L_X34Y129_SLICE_X51Y129_C = CLBLL_L_X34Y129_SLICE_X51Y129_CO6;
  assign CLBLL_L_X34Y129_SLICE_X51Y129_D = CLBLL_L_X34Y129_SLICE_X51Y129_DO6;
  assign CLBLL_L_X36Y115_SLICE_X54Y115_COUT = CLBLL_L_X36Y115_SLICE_X54Y115_D_CY;
  assign CLBLL_L_X36Y115_SLICE_X54Y115_A = CLBLL_L_X36Y115_SLICE_X54Y115_AO6;
  assign CLBLL_L_X36Y115_SLICE_X54Y115_B = CLBLL_L_X36Y115_SLICE_X54Y115_BO6;
  assign CLBLL_L_X36Y115_SLICE_X54Y115_C = CLBLL_L_X36Y115_SLICE_X54Y115_CO6;
  assign CLBLL_L_X36Y115_SLICE_X54Y115_D = CLBLL_L_X36Y115_SLICE_X54Y115_DO6;
  assign CLBLL_L_X36Y115_SLICE_X54Y115_AMUX = CLBLL_L_X36Y115_SLICE_X54Y115_AO5;
  assign CLBLL_L_X36Y115_SLICE_X55Y115_COUT = CLBLL_L_X36Y115_SLICE_X55Y115_D_CY;
  assign CLBLL_L_X36Y115_SLICE_X55Y115_A = CLBLL_L_X36Y115_SLICE_X55Y115_AO6;
  assign CLBLL_L_X36Y115_SLICE_X55Y115_B = CLBLL_L_X36Y115_SLICE_X55Y115_BO6;
  assign CLBLL_L_X36Y115_SLICE_X55Y115_C = CLBLL_L_X36Y115_SLICE_X55Y115_CO6;
  assign CLBLL_L_X36Y115_SLICE_X55Y115_D = CLBLL_L_X36Y115_SLICE_X55Y115_DO6;
  assign CLBLL_L_X36Y116_SLICE_X54Y116_COUT = CLBLL_L_X36Y116_SLICE_X54Y116_D_CY;
  assign CLBLL_L_X36Y116_SLICE_X54Y116_A = CLBLL_L_X36Y116_SLICE_X54Y116_AO6;
  assign CLBLL_L_X36Y116_SLICE_X54Y116_B = CLBLL_L_X36Y116_SLICE_X54Y116_BO6;
  assign CLBLL_L_X36Y116_SLICE_X54Y116_C = CLBLL_L_X36Y116_SLICE_X54Y116_CO6;
  assign CLBLL_L_X36Y116_SLICE_X54Y116_D = CLBLL_L_X36Y116_SLICE_X54Y116_DO6;
  assign CLBLL_L_X36Y116_SLICE_X54Y116_AMUX = CLBLL_L_X36Y116_SLICE_X54Y116_AO5;
  assign CLBLL_L_X36Y116_SLICE_X54Y116_BMUX = CLBLL_L_X36Y116_SLICE_X54Y116_BO5;
  assign CLBLL_L_X36Y116_SLICE_X54Y116_CMUX = CLBLL_L_X36Y116_SLICE_X54Y116_CO5;
  assign CLBLL_L_X36Y116_SLICE_X55Y116_COUT = CLBLL_L_X36Y116_SLICE_X55Y116_D_CY;
  assign CLBLL_L_X36Y116_SLICE_X55Y116_A = CLBLL_L_X36Y116_SLICE_X55Y116_AO6;
  assign CLBLL_L_X36Y116_SLICE_X55Y116_B = CLBLL_L_X36Y116_SLICE_X55Y116_BO6;
  assign CLBLL_L_X36Y116_SLICE_X55Y116_C = CLBLL_L_X36Y116_SLICE_X55Y116_CO6;
  assign CLBLL_L_X36Y116_SLICE_X55Y116_D = CLBLL_L_X36Y116_SLICE_X55Y116_DO6;
  assign CLBLL_L_X36Y116_SLICE_X55Y116_AMUX = CLBLL_L_X36Y116_SLICE_X55Y116_AO5;
  assign CLBLL_L_X36Y117_SLICE_X54Y117_COUT = CLBLL_L_X36Y117_SLICE_X54Y117_D_CY;
  assign CLBLL_L_X36Y117_SLICE_X54Y117_A = CLBLL_L_X36Y117_SLICE_X54Y117_AO6;
  assign CLBLL_L_X36Y117_SLICE_X54Y117_B = CLBLL_L_X36Y117_SLICE_X54Y117_BO6;
  assign CLBLL_L_X36Y117_SLICE_X54Y117_C = CLBLL_L_X36Y117_SLICE_X54Y117_CO6;
  assign CLBLL_L_X36Y117_SLICE_X54Y117_D = CLBLL_L_X36Y117_SLICE_X54Y117_DO6;
  assign CLBLL_L_X36Y117_SLICE_X55Y117_COUT = CLBLL_L_X36Y117_SLICE_X55Y117_D_CY;
  assign CLBLL_L_X36Y117_SLICE_X55Y117_A = CLBLL_L_X36Y117_SLICE_X55Y117_AO6;
  assign CLBLL_L_X36Y117_SLICE_X55Y117_B = CLBLL_L_X36Y117_SLICE_X55Y117_BO6;
  assign CLBLL_L_X36Y117_SLICE_X55Y117_C = CLBLL_L_X36Y117_SLICE_X55Y117_CO6;
  assign CLBLL_L_X36Y117_SLICE_X55Y117_D = CLBLL_L_X36Y117_SLICE_X55Y117_DO6;
  assign CLBLL_L_X36Y117_SLICE_X55Y117_AMUX = CLBLL_L_X36Y117_SLICE_X55Y117_AO5;
  assign CLBLL_L_X36Y117_SLICE_X55Y117_BMUX = CLBLL_L_X36Y117_SLICE_X55Y117_BO5;
  assign CLBLL_L_X36Y118_SLICE_X54Y118_COUT = CLBLL_L_X36Y118_SLICE_X54Y118_D_CY;
  assign CLBLL_L_X36Y118_SLICE_X54Y118_A = CLBLL_L_X36Y118_SLICE_X54Y118_AO6;
  assign CLBLL_L_X36Y118_SLICE_X54Y118_B = CLBLL_L_X36Y118_SLICE_X54Y118_BO6;
  assign CLBLL_L_X36Y118_SLICE_X54Y118_C = CLBLL_L_X36Y118_SLICE_X54Y118_CO6;
  assign CLBLL_L_X36Y118_SLICE_X54Y118_D = CLBLL_L_X36Y118_SLICE_X54Y118_DO6;
  assign CLBLL_L_X36Y118_SLICE_X55Y118_COUT = CLBLL_L_X36Y118_SLICE_X55Y118_D_CY;
  assign CLBLL_L_X36Y118_SLICE_X55Y118_A = CLBLL_L_X36Y118_SLICE_X55Y118_AO6;
  assign CLBLL_L_X36Y118_SLICE_X55Y118_B = CLBLL_L_X36Y118_SLICE_X55Y118_BO6;
  assign CLBLL_L_X36Y118_SLICE_X55Y118_C = CLBLL_L_X36Y118_SLICE_X55Y118_CO6;
  assign CLBLL_L_X36Y118_SLICE_X55Y118_D = CLBLL_L_X36Y118_SLICE_X55Y118_DO6;
  assign CLBLL_L_X36Y118_SLICE_X55Y118_AMUX = CLBLL_L_X36Y118_SLICE_X55Y118_AO5;
  assign CLBLL_L_X36Y118_SLICE_X55Y118_CMUX = CLBLL_L_X36Y118_SLICE_X55Y118_CO6;
  assign CLBLL_L_X36Y119_SLICE_X54Y119_COUT = CLBLL_L_X36Y119_SLICE_X54Y119_D_CY;
  assign CLBLL_L_X36Y119_SLICE_X54Y119_A = CLBLL_L_X36Y119_SLICE_X54Y119_AO6;
  assign CLBLL_L_X36Y119_SLICE_X54Y119_B = CLBLL_L_X36Y119_SLICE_X54Y119_BO6;
  assign CLBLL_L_X36Y119_SLICE_X54Y119_C = CLBLL_L_X36Y119_SLICE_X54Y119_CO6;
  assign CLBLL_L_X36Y119_SLICE_X54Y119_D = CLBLL_L_X36Y119_SLICE_X54Y119_DO6;
  assign CLBLL_L_X36Y119_SLICE_X55Y119_COUT = CLBLL_L_X36Y119_SLICE_X55Y119_D_CY;
  assign CLBLL_L_X36Y119_SLICE_X55Y119_A = CLBLL_L_X36Y119_SLICE_X55Y119_AO6;
  assign CLBLL_L_X36Y119_SLICE_X55Y119_B = CLBLL_L_X36Y119_SLICE_X55Y119_BO6;
  assign CLBLL_L_X36Y119_SLICE_X55Y119_C = CLBLL_L_X36Y119_SLICE_X55Y119_CO6;
  assign CLBLL_L_X36Y119_SLICE_X55Y119_D = CLBLL_L_X36Y119_SLICE_X55Y119_DO6;
  assign CLBLL_L_X36Y120_SLICE_X54Y120_COUT = CLBLL_L_X36Y120_SLICE_X54Y120_D_CY;
  assign CLBLL_L_X36Y120_SLICE_X54Y120_A = CLBLL_L_X36Y120_SLICE_X54Y120_AO6;
  assign CLBLL_L_X36Y120_SLICE_X54Y120_B = CLBLL_L_X36Y120_SLICE_X54Y120_BO6;
  assign CLBLL_L_X36Y120_SLICE_X54Y120_C = CLBLL_L_X36Y120_SLICE_X54Y120_CO6;
  assign CLBLL_L_X36Y120_SLICE_X54Y120_D = CLBLL_L_X36Y120_SLICE_X54Y120_DO6;
  assign CLBLL_L_X36Y120_SLICE_X55Y120_COUT = CLBLL_L_X36Y120_SLICE_X55Y120_D_CY;
  assign CLBLL_L_X36Y120_SLICE_X55Y120_A = CLBLL_L_X36Y120_SLICE_X55Y120_AO6;
  assign CLBLL_L_X36Y120_SLICE_X55Y120_B = CLBLL_L_X36Y120_SLICE_X55Y120_BO6;
  assign CLBLL_L_X36Y120_SLICE_X55Y120_C = CLBLL_L_X36Y120_SLICE_X55Y120_CO6;
  assign CLBLL_L_X36Y120_SLICE_X55Y120_D = CLBLL_L_X36Y120_SLICE_X55Y120_DO6;
  assign CLBLL_L_X36Y121_SLICE_X54Y121_COUT = CLBLL_L_X36Y121_SLICE_X54Y121_D_CY;
  assign CLBLL_L_X36Y121_SLICE_X54Y121_A = CLBLL_L_X36Y121_SLICE_X54Y121_AO6;
  assign CLBLL_L_X36Y121_SLICE_X54Y121_B = CLBLL_L_X36Y121_SLICE_X54Y121_BO6;
  assign CLBLL_L_X36Y121_SLICE_X54Y121_C = CLBLL_L_X36Y121_SLICE_X54Y121_CO6;
  assign CLBLL_L_X36Y121_SLICE_X54Y121_D = CLBLL_L_X36Y121_SLICE_X54Y121_DO6;
  assign CLBLL_L_X36Y121_SLICE_X54Y121_AMUX = CLBLL_L_X36Y121_SLICE_X54Y121_AO5;
  assign CLBLL_L_X36Y121_SLICE_X55Y121_COUT = CLBLL_L_X36Y121_SLICE_X55Y121_D_CY;
  assign CLBLL_L_X36Y121_SLICE_X55Y121_A = CLBLL_L_X36Y121_SLICE_X55Y121_AO6;
  assign CLBLL_L_X36Y121_SLICE_X55Y121_B = CLBLL_L_X36Y121_SLICE_X55Y121_BO6;
  assign CLBLL_L_X36Y121_SLICE_X55Y121_C = CLBLL_L_X36Y121_SLICE_X55Y121_CO6;
  assign CLBLL_L_X36Y121_SLICE_X55Y121_D = CLBLL_L_X36Y121_SLICE_X55Y121_DO6;
  assign CLBLL_L_X36Y121_SLICE_X55Y121_AMUX = CLBLL_L_X36Y121_SLICE_X55Y121_AO5;
  assign CLBLL_L_X36Y122_SLICE_X54Y122_COUT = CLBLL_L_X36Y122_SLICE_X54Y122_D_CY;
  assign CLBLL_L_X36Y122_SLICE_X54Y122_A = CLBLL_L_X36Y122_SLICE_X54Y122_AO6;
  assign CLBLL_L_X36Y122_SLICE_X54Y122_B = CLBLL_L_X36Y122_SLICE_X54Y122_BO6;
  assign CLBLL_L_X36Y122_SLICE_X54Y122_C = CLBLL_L_X36Y122_SLICE_X54Y122_CO6;
  assign CLBLL_L_X36Y122_SLICE_X54Y122_D = CLBLL_L_X36Y122_SLICE_X54Y122_DO6;
  assign CLBLL_L_X36Y122_SLICE_X54Y122_AMUX = CLBLL_L_X36Y122_SLICE_X54Y122_AO5;
  assign CLBLL_L_X36Y122_SLICE_X55Y122_COUT = CLBLL_L_X36Y122_SLICE_X55Y122_D_CY;
  assign CLBLL_L_X36Y122_SLICE_X55Y122_A = CLBLL_L_X36Y122_SLICE_X55Y122_AO6;
  assign CLBLL_L_X36Y122_SLICE_X55Y122_B = CLBLL_L_X36Y122_SLICE_X55Y122_BO6;
  assign CLBLL_L_X36Y122_SLICE_X55Y122_C = CLBLL_L_X36Y122_SLICE_X55Y122_CO6;
  assign CLBLL_L_X36Y122_SLICE_X55Y122_D = CLBLL_L_X36Y122_SLICE_X55Y122_DO6;
  assign CLBLL_L_X36Y122_SLICE_X55Y122_AMUX = CLBLL_L_X36Y122_SLICE_X55Y122_AO5;
  assign CLBLL_L_X36Y123_SLICE_X54Y123_COUT = CLBLL_L_X36Y123_SLICE_X54Y123_D_CY;
  assign CLBLL_L_X36Y123_SLICE_X54Y123_A = CLBLL_L_X36Y123_SLICE_X54Y123_AO6;
  assign CLBLL_L_X36Y123_SLICE_X54Y123_B = CLBLL_L_X36Y123_SLICE_X54Y123_BO6;
  assign CLBLL_L_X36Y123_SLICE_X54Y123_C = CLBLL_L_X36Y123_SLICE_X54Y123_CO6;
  assign CLBLL_L_X36Y123_SLICE_X54Y123_D = CLBLL_L_X36Y123_SLICE_X54Y123_DO6;
  assign CLBLL_L_X36Y123_SLICE_X54Y123_AMUX = CLBLL_L_X36Y123_SLICE_X54Y123_AO5;
  assign CLBLL_L_X36Y123_SLICE_X55Y123_COUT = CLBLL_L_X36Y123_SLICE_X55Y123_D_CY;
  assign CLBLL_L_X36Y123_SLICE_X55Y123_A = CLBLL_L_X36Y123_SLICE_X55Y123_AO6;
  assign CLBLL_L_X36Y123_SLICE_X55Y123_B = CLBLL_L_X36Y123_SLICE_X55Y123_BO6;
  assign CLBLL_L_X36Y123_SLICE_X55Y123_C = CLBLL_L_X36Y123_SLICE_X55Y123_CO6;
  assign CLBLL_L_X36Y123_SLICE_X55Y123_D = CLBLL_L_X36Y123_SLICE_X55Y123_DO6;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_COUT = CLBLL_L_X36Y124_SLICE_X54Y124_D_CY;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_A = CLBLL_L_X36Y124_SLICE_X54Y124_AO6;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_B = CLBLL_L_X36Y124_SLICE_X54Y124_BO6;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_C = CLBLL_L_X36Y124_SLICE_X54Y124_CO6;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_D = CLBLL_L_X36Y124_SLICE_X54Y124_DO6;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_COUT = CLBLL_L_X36Y124_SLICE_X55Y124_D_CY;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_A = CLBLL_L_X36Y124_SLICE_X55Y124_AO6;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_B = CLBLL_L_X36Y124_SLICE_X55Y124_BO6;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_C = CLBLL_L_X36Y124_SLICE_X55Y124_CO6;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_D = CLBLL_L_X36Y124_SLICE_X55Y124_DO6;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_BMUX = CLBLL_L_X36Y124_SLICE_X55Y124_BO6;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_CMUX = CLBLL_L_X36Y124_SLICE_X55Y124_CO6;
  assign CLBLL_L_X36Y125_SLICE_X54Y125_COUT = CLBLL_L_X36Y125_SLICE_X54Y125_D_CY;
  assign CLBLL_L_X36Y125_SLICE_X54Y125_A = CLBLL_L_X36Y125_SLICE_X54Y125_AO6;
  assign CLBLL_L_X36Y125_SLICE_X54Y125_B = CLBLL_L_X36Y125_SLICE_X54Y125_BO6;
  assign CLBLL_L_X36Y125_SLICE_X54Y125_C = CLBLL_L_X36Y125_SLICE_X54Y125_CO6;
  assign CLBLL_L_X36Y125_SLICE_X54Y125_D = CLBLL_L_X36Y125_SLICE_X54Y125_DO6;
  assign CLBLL_L_X36Y125_SLICE_X55Y125_COUT = CLBLL_L_X36Y125_SLICE_X55Y125_D_CY;
  assign CLBLL_L_X36Y125_SLICE_X55Y125_A = CLBLL_L_X36Y125_SLICE_X55Y125_AO6;
  assign CLBLL_L_X36Y125_SLICE_X55Y125_B = CLBLL_L_X36Y125_SLICE_X55Y125_BO6;
  assign CLBLL_L_X36Y125_SLICE_X55Y125_C = CLBLL_L_X36Y125_SLICE_X55Y125_CO6;
  assign CLBLL_L_X36Y125_SLICE_X55Y125_D = CLBLL_L_X36Y125_SLICE_X55Y125_DO6;
  assign CLBLL_L_X36Y125_SLICE_X55Y125_AMUX = CLBLL_L_X36Y125_SLICE_X55Y125_AO5;
  assign CLBLL_L_X36Y125_SLICE_X55Y125_BMUX = CLBLL_L_X36Y125_SLICE_X55Y125_BO5;
  assign CLBLL_L_X36Y125_SLICE_X55Y125_CMUX = CLBLL_L_X36Y125_SLICE_X55Y125_CO6;
  assign CLBLL_L_X36Y126_SLICE_X54Y126_COUT = CLBLL_L_X36Y126_SLICE_X54Y126_D_CY;
  assign CLBLL_L_X36Y126_SLICE_X54Y126_A = CLBLL_L_X36Y126_SLICE_X54Y126_AO6;
  assign CLBLL_L_X36Y126_SLICE_X54Y126_B = CLBLL_L_X36Y126_SLICE_X54Y126_BO6;
  assign CLBLL_L_X36Y126_SLICE_X54Y126_C = CLBLL_L_X36Y126_SLICE_X54Y126_CO6;
  assign CLBLL_L_X36Y126_SLICE_X54Y126_D = CLBLL_L_X36Y126_SLICE_X54Y126_DO6;
  assign CLBLL_L_X36Y126_SLICE_X54Y126_CMUX = CLBLL_L_X36Y126_SLICE_X54Y126_CO6;
  assign CLBLL_L_X36Y126_SLICE_X55Y126_COUT = CLBLL_L_X36Y126_SLICE_X55Y126_D_CY;
  assign CLBLL_L_X36Y126_SLICE_X55Y126_A = CLBLL_L_X36Y126_SLICE_X55Y126_AO6;
  assign CLBLL_L_X36Y126_SLICE_X55Y126_B = CLBLL_L_X36Y126_SLICE_X55Y126_BO6;
  assign CLBLL_L_X36Y126_SLICE_X55Y126_C = CLBLL_L_X36Y126_SLICE_X55Y126_CO6;
  assign CLBLL_L_X36Y126_SLICE_X55Y126_D = CLBLL_L_X36Y126_SLICE_X55Y126_DO6;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_COUT = CLBLL_L_X36Y127_SLICE_X54Y127_D_CY;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_A = CLBLL_L_X36Y127_SLICE_X54Y127_AO6;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_B = CLBLL_L_X36Y127_SLICE_X54Y127_BO6;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_C = CLBLL_L_X36Y127_SLICE_X54Y127_CO6;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_D = CLBLL_L_X36Y127_SLICE_X54Y127_DO6;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_COUT = CLBLL_L_X36Y127_SLICE_X55Y127_D_CY;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_A = CLBLL_L_X36Y127_SLICE_X55Y127_AO6;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_B = CLBLL_L_X36Y127_SLICE_X55Y127_BO6;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_C = CLBLL_L_X36Y127_SLICE_X55Y127_CO6;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_D = CLBLL_L_X36Y127_SLICE_X55Y127_DO6;
  assign CLBLL_L_X36Y128_SLICE_X54Y128_COUT = CLBLL_L_X36Y128_SLICE_X54Y128_D_CY;
  assign CLBLL_L_X36Y128_SLICE_X54Y128_A = CLBLL_L_X36Y128_SLICE_X54Y128_AO6;
  assign CLBLL_L_X36Y128_SLICE_X54Y128_B = CLBLL_L_X36Y128_SLICE_X54Y128_BO6;
  assign CLBLL_L_X36Y128_SLICE_X54Y128_C = CLBLL_L_X36Y128_SLICE_X54Y128_CO6;
  assign CLBLL_L_X36Y128_SLICE_X54Y128_D = CLBLL_L_X36Y128_SLICE_X54Y128_DO6;
  assign CLBLL_L_X36Y128_SLICE_X55Y128_COUT = CLBLL_L_X36Y128_SLICE_X55Y128_D_CY;
  assign CLBLL_L_X36Y128_SLICE_X55Y128_A = CLBLL_L_X36Y128_SLICE_X55Y128_AO6;
  assign CLBLL_L_X36Y128_SLICE_X55Y128_B = CLBLL_L_X36Y128_SLICE_X55Y128_BO6;
  assign CLBLL_L_X36Y128_SLICE_X55Y128_C = CLBLL_L_X36Y128_SLICE_X55Y128_CO6;
  assign CLBLL_L_X36Y128_SLICE_X55Y128_D = CLBLL_L_X36Y128_SLICE_X55Y128_DO6;
  assign CLBLL_L_X36Y129_SLICE_X54Y129_COUT = CLBLL_L_X36Y129_SLICE_X54Y129_D_CY;
  assign CLBLL_L_X36Y129_SLICE_X54Y129_A = CLBLL_L_X36Y129_SLICE_X54Y129_AO6;
  assign CLBLL_L_X36Y129_SLICE_X54Y129_B = CLBLL_L_X36Y129_SLICE_X54Y129_BO6;
  assign CLBLL_L_X36Y129_SLICE_X54Y129_C = CLBLL_L_X36Y129_SLICE_X54Y129_CO6;
  assign CLBLL_L_X36Y129_SLICE_X54Y129_D = CLBLL_L_X36Y129_SLICE_X54Y129_DO6;
  assign CLBLL_L_X36Y129_SLICE_X55Y129_COUT = CLBLL_L_X36Y129_SLICE_X55Y129_D_CY;
  assign CLBLL_L_X36Y129_SLICE_X55Y129_A = CLBLL_L_X36Y129_SLICE_X55Y129_AO6;
  assign CLBLL_L_X36Y129_SLICE_X55Y129_B = CLBLL_L_X36Y129_SLICE_X55Y129_BO6;
  assign CLBLL_L_X36Y129_SLICE_X55Y129_C = CLBLL_L_X36Y129_SLICE_X55Y129_CO6;
  assign CLBLL_L_X36Y129_SLICE_X55Y129_D = CLBLL_L_X36Y129_SLICE_X55Y129_DO6;
  assign CLBLL_L_X38Y118_SLICE_X58Y118_COUT = CLBLL_L_X38Y118_SLICE_X58Y118_D_CY;
  assign CLBLL_L_X38Y118_SLICE_X58Y118_A = CLBLL_L_X38Y118_SLICE_X58Y118_AO6;
  assign CLBLL_L_X38Y118_SLICE_X58Y118_B = CLBLL_L_X38Y118_SLICE_X58Y118_BO6;
  assign CLBLL_L_X38Y118_SLICE_X58Y118_C = CLBLL_L_X38Y118_SLICE_X58Y118_CO6;
  assign CLBLL_L_X38Y118_SLICE_X58Y118_D = CLBLL_L_X38Y118_SLICE_X58Y118_DO6;
  assign CLBLL_L_X38Y118_SLICE_X58Y118_AMUX = CLBLL_L_X38Y118_SLICE_X58Y118_AO5;
  assign CLBLL_L_X38Y118_SLICE_X59Y118_COUT = CLBLL_L_X38Y118_SLICE_X59Y118_D_CY;
  assign CLBLL_L_X38Y118_SLICE_X59Y118_A = CLBLL_L_X38Y118_SLICE_X59Y118_AO6;
  assign CLBLL_L_X38Y118_SLICE_X59Y118_B = CLBLL_L_X38Y118_SLICE_X59Y118_BO6;
  assign CLBLL_L_X38Y118_SLICE_X59Y118_C = CLBLL_L_X38Y118_SLICE_X59Y118_CO6;
  assign CLBLL_L_X38Y118_SLICE_X59Y118_D = CLBLL_L_X38Y118_SLICE_X59Y118_DO6;
  assign CLBLL_L_X38Y119_SLICE_X58Y119_COUT = CLBLL_L_X38Y119_SLICE_X58Y119_D_CY;
  assign CLBLL_L_X38Y119_SLICE_X58Y119_A = CLBLL_L_X38Y119_SLICE_X58Y119_AO6;
  assign CLBLL_L_X38Y119_SLICE_X58Y119_B = CLBLL_L_X38Y119_SLICE_X58Y119_BO6;
  assign CLBLL_L_X38Y119_SLICE_X58Y119_C = CLBLL_L_X38Y119_SLICE_X58Y119_CO6;
  assign CLBLL_L_X38Y119_SLICE_X58Y119_D = CLBLL_L_X38Y119_SLICE_X58Y119_DO6;
  assign CLBLL_L_X38Y119_SLICE_X59Y119_COUT = CLBLL_L_X38Y119_SLICE_X59Y119_D_CY;
  assign CLBLL_L_X38Y119_SLICE_X59Y119_A = CLBLL_L_X38Y119_SLICE_X59Y119_AO6;
  assign CLBLL_L_X38Y119_SLICE_X59Y119_B = CLBLL_L_X38Y119_SLICE_X59Y119_BO6;
  assign CLBLL_L_X38Y119_SLICE_X59Y119_C = CLBLL_L_X38Y119_SLICE_X59Y119_CO6;
  assign CLBLL_L_X38Y119_SLICE_X59Y119_D = CLBLL_L_X38Y119_SLICE_X59Y119_DO6;
  assign CLBLL_L_X38Y121_SLICE_X58Y121_COUT = CLBLL_L_X38Y121_SLICE_X58Y121_D_CY;
  assign CLBLL_L_X38Y121_SLICE_X58Y121_A = CLBLL_L_X38Y121_SLICE_X58Y121_AO6;
  assign CLBLL_L_X38Y121_SLICE_X58Y121_B = CLBLL_L_X38Y121_SLICE_X58Y121_BO6;
  assign CLBLL_L_X38Y121_SLICE_X58Y121_C = CLBLL_L_X38Y121_SLICE_X58Y121_CO6;
  assign CLBLL_L_X38Y121_SLICE_X58Y121_D = CLBLL_L_X38Y121_SLICE_X58Y121_DO6;
  assign CLBLL_L_X38Y121_SLICE_X59Y121_COUT = CLBLL_L_X38Y121_SLICE_X59Y121_D_CY;
  assign CLBLL_L_X38Y121_SLICE_X59Y121_A = CLBLL_L_X38Y121_SLICE_X59Y121_AO6;
  assign CLBLL_L_X38Y121_SLICE_X59Y121_B = CLBLL_L_X38Y121_SLICE_X59Y121_BO6;
  assign CLBLL_L_X38Y121_SLICE_X59Y121_C = CLBLL_L_X38Y121_SLICE_X59Y121_CO6;
  assign CLBLL_L_X38Y121_SLICE_X59Y121_D = CLBLL_L_X38Y121_SLICE_X59Y121_DO6;
  assign CLBLL_L_X38Y123_SLICE_X58Y123_COUT = CLBLL_L_X38Y123_SLICE_X58Y123_D_CY;
  assign CLBLL_L_X38Y123_SLICE_X58Y123_A = CLBLL_L_X38Y123_SLICE_X58Y123_AO6;
  assign CLBLL_L_X38Y123_SLICE_X58Y123_B = CLBLL_L_X38Y123_SLICE_X58Y123_BO6;
  assign CLBLL_L_X38Y123_SLICE_X58Y123_C = CLBLL_L_X38Y123_SLICE_X58Y123_CO6;
  assign CLBLL_L_X38Y123_SLICE_X58Y123_D = CLBLL_L_X38Y123_SLICE_X58Y123_DO6;
  assign CLBLL_L_X38Y123_SLICE_X59Y123_COUT = CLBLL_L_X38Y123_SLICE_X59Y123_D_CY;
  assign CLBLL_L_X38Y123_SLICE_X59Y123_A = CLBLL_L_X38Y123_SLICE_X59Y123_AO6;
  assign CLBLL_L_X38Y123_SLICE_X59Y123_B = CLBLL_L_X38Y123_SLICE_X59Y123_BO6;
  assign CLBLL_L_X38Y123_SLICE_X59Y123_C = CLBLL_L_X38Y123_SLICE_X59Y123_CO6;
  assign CLBLL_L_X38Y123_SLICE_X59Y123_D = CLBLL_L_X38Y123_SLICE_X59Y123_DO6;
  assign CLBLL_L_X38Y124_SLICE_X58Y124_COUT = CLBLL_L_X38Y124_SLICE_X58Y124_D_CY;
  assign CLBLL_L_X38Y124_SLICE_X58Y124_A = CLBLL_L_X38Y124_SLICE_X58Y124_AO6;
  assign CLBLL_L_X38Y124_SLICE_X58Y124_B = CLBLL_L_X38Y124_SLICE_X58Y124_BO6;
  assign CLBLL_L_X38Y124_SLICE_X58Y124_C = CLBLL_L_X38Y124_SLICE_X58Y124_CO6;
  assign CLBLL_L_X38Y124_SLICE_X58Y124_D = CLBLL_L_X38Y124_SLICE_X58Y124_DO6;
  assign CLBLL_L_X38Y124_SLICE_X58Y124_AMUX = CLBLL_L_X38Y124_SLICE_X58Y124_AO6;
  assign CLBLL_L_X38Y124_SLICE_X59Y124_COUT = CLBLL_L_X38Y124_SLICE_X59Y124_D_CY;
  assign CLBLL_L_X38Y124_SLICE_X59Y124_A = CLBLL_L_X38Y124_SLICE_X59Y124_AO6;
  assign CLBLL_L_X38Y124_SLICE_X59Y124_B = CLBLL_L_X38Y124_SLICE_X59Y124_BO6;
  assign CLBLL_L_X38Y124_SLICE_X59Y124_C = CLBLL_L_X38Y124_SLICE_X59Y124_CO6;
  assign CLBLL_L_X38Y124_SLICE_X59Y124_D = CLBLL_L_X38Y124_SLICE_X59Y124_DO6;
  assign CLBLL_L_X38Y126_SLICE_X58Y126_COUT = CLBLL_L_X38Y126_SLICE_X58Y126_D_CY;
  assign CLBLL_L_X38Y126_SLICE_X58Y126_A = CLBLL_L_X38Y126_SLICE_X58Y126_AO6;
  assign CLBLL_L_X38Y126_SLICE_X58Y126_B = CLBLL_L_X38Y126_SLICE_X58Y126_BO6;
  assign CLBLL_L_X38Y126_SLICE_X58Y126_C = CLBLL_L_X38Y126_SLICE_X58Y126_CO6;
  assign CLBLL_L_X38Y126_SLICE_X58Y126_D = CLBLL_L_X38Y126_SLICE_X58Y126_DO6;
  assign CLBLL_L_X38Y126_SLICE_X59Y126_COUT = CLBLL_L_X38Y126_SLICE_X59Y126_D_CY;
  assign CLBLL_L_X38Y126_SLICE_X59Y126_A = CLBLL_L_X38Y126_SLICE_X59Y126_AO6;
  assign CLBLL_L_X38Y126_SLICE_X59Y126_B = CLBLL_L_X38Y126_SLICE_X59Y126_BO6;
  assign CLBLL_L_X38Y126_SLICE_X59Y126_C = CLBLL_L_X38Y126_SLICE_X59Y126_CO6;
  assign CLBLL_L_X38Y126_SLICE_X59Y126_D = CLBLL_L_X38Y126_SLICE_X59Y126_DO6;
  assign CLBLM_L_X32Y116_SLICE_X46Y116_COUT = CLBLM_L_X32Y116_SLICE_X46Y116_D_CY;
  assign CLBLM_L_X32Y116_SLICE_X46Y116_A = CLBLM_L_X32Y116_SLICE_X46Y116_AO6;
  assign CLBLM_L_X32Y116_SLICE_X46Y116_B = CLBLM_L_X32Y116_SLICE_X46Y116_BO6;
  assign CLBLM_L_X32Y116_SLICE_X46Y116_C = CLBLM_L_X32Y116_SLICE_X46Y116_CO6;
  assign CLBLM_L_X32Y116_SLICE_X46Y116_D = CLBLM_L_X32Y116_SLICE_X46Y116_DO6;
  assign CLBLM_L_X32Y116_SLICE_X47Y116_COUT = CLBLM_L_X32Y116_SLICE_X47Y116_D_CY;
  assign CLBLM_L_X32Y116_SLICE_X47Y116_A = CLBLM_L_X32Y116_SLICE_X47Y116_AO6;
  assign CLBLM_L_X32Y116_SLICE_X47Y116_B = CLBLM_L_X32Y116_SLICE_X47Y116_BO6;
  assign CLBLM_L_X32Y116_SLICE_X47Y116_C = CLBLM_L_X32Y116_SLICE_X47Y116_CO6;
  assign CLBLM_L_X32Y116_SLICE_X47Y116_D = CLBLM_L_X32Y116_SLICE_X47Y116_DO6;
  assign CLBLM_L_X32Y117_SLICE_X46Y117_COUT = CLBLM_L_X32Y117_SLICE_X46Y117_D_CY;
  assign CLBLM_L_X32Y117_SLICE_X46Y117_A = CLBLM_L_X32Y117_SLICE_X46Y117_AO6;
  assign CLBLM_L_X32Y117_SLICE_X46Y117_B = CLBLM_L_X32Y117_SLICE_X46Y117_BO6;
  assign CLBLM_L_X32Y117_SLICE_X46Y117_C = CLBLM_L_X32Y117_SLICE_X46Y117_CO6;
  assign CLBLM_L_X32Y117_SLICE_X46Y117_D = CLBLM_L_X32Y117_SLICE_X46Y117_DO6;
  assign CLBLM_L_X32Y117_SLICE_X47Y117_COUT = CLBLM_L_X32Y117_SLICE_X47Y117_D_CY;
  assign CLBLM_L_X32Y117_SLICE_X47Y117_A = CLBLM_L_X32Y117_SLICE_X47Y117_AO6;
  assign CLBLM_L_X32Y117_SLICE_X47Y117_B = CLBLM_L_X32Y117_SLICE_X47Y117_BO6;
  assign CLBLM_L_X32Y117_SLICE_X47Y117_C = CLBLM_L_X32Y117_SLICE_X47Y117_CO6;
  assign CLBLM_L_X32Y117_SLICE_X47Y117_D = CLBLM_L_X32Y117_SLICE_X47Y117_DO6;
  assign CLBLM_L_X32Y123_SLICE_X46Y123_COUT = CLBLM_L_X32Y123_SLICE_X46Y123_D_CY;
  assign CLBLM_L_X32Y123_SLICE_X46Y123_A = CLBLM_L_X32Y123_SLICE_X46Y123_AO6;
  assign CLBLM_L_X32Y123_SLICE_X46Y123_B = CLBLM_L_X32Y123_SLICE_X46Y123_BO6;
  assign CLBLM_L_X32Y123_SLICE_X46Y123_C = CLBLM_L_X32Y123_SLICE_X46Y123_CO6;
  assign CLBLM_L_X32Y123_SLICE_X46Y123_D = CLBLM_L_X32Y123_SLICE_X46Y123_DO6;
  assign CLBLM_L_X32Y123_SLICE_X47Y123_COUT = CLBLM_L_X32Y123_SLICE_X47Y123_D_CY;
  assign CLBLM_L_X32Y123_SLICE_X47Y123_A = CLBLM_L_X32Y123_SLICE_X47Y123_AO6;
  assign CLBLM_L_X32Y123_SLICE_X47Y123_B = CLBLM_L_X32Y123_SLICE_X47Y123_BO6;
  assign CLBLM_L_X32Y123_SLICE_X47Y123_C = CLBLM_L_X32Y123_SLICE_X47Y123_CO6;
  assign CLBLM_L_X32Y123_SLICE_X47Y123_D = CLBLM_L_X32Y123_SLICE_X47Y123_DO6;
  assign CLBLM_L_X32Y123_SLICE_X47Y123_AMUX = CLBLM_L_X32Y123_SLICE_X47Y123_AO5;
  assign CLBLM_R_X33Y115_SLICE_X48Y115_COUT = CLBLM_R_X33Y115_SLICE_X48Y115_D_CY;
  assign CLBLM_R_X33Y115_SLICE_X48Y115_A = CLBLM_R_X33Y115_SLICE_X48Y115_AO6;
  assign CLBLM_R_X33Y115_SLICE_X48Y115_B = CLBLM_R_X33Y115_SLICE_X48Y115_BO6;
  assign CLBLM_R_X33Y115_SLICE_X48Y115_C = CLBLM_R_X33Y115_SLICE_X48Y115_CO6;
  assign CLBLM_R_X33Y115_SLICE_X48Y115_D = CLBLM_R_X33Y115_SLICE_X48Y115_DO6;
  assign CLBLM_R_X33Y115_SLICE_X49Y115_COUT = CLBLM_R_X33Y115_SLICE_X49Y115_D_CY;
  assign CLBLM_R_X33Y115_SLICE_X49Y115_A = CLBLM_R_X33Y115_SLICE_X49Y115_AO6;
  assign CLBLM_R_X33Y115_SLICE_X49Y115_B = CLBLM_R_X33Y115_SLICE_X49Y115_BO6;
  assign CLBLM_R_X33Y115_SLICE_X49Y115_C = CLBLM_R_X33Y115_SLICE_X49Y115_CO6;
  assign CLBLM_R_X33Y115_SLICE_X49Y115_D = CLBLM_R_X33Y115_SLICE_X49Y115_DO6;
  assign CLBLM_R_X33Y115_SLICE_X49Y115_AMUX = CLBLM_R_X33Y115_SLICE_X49Y115_AO5;
  assign CLBLM_R_X33Y116_SLICE_X48Y116_COUT = CLBLM_R_X33Y116_SLICE_X48Y116_D_CY;
  assign CLBLM_R_X33Y116_SLICE_X48Y116_A = CLBLM_R_X33Y116_SLICE_X48Y116_AO6;
  assign CLBLM_R_X33Y116_SLICE_X48Y116_B = CLBLM_R_X33Y116_SLICE_X48Y116_BO6;
  assign CLBLM_R_X33Y116_SLICE_X48Y116_C = CLBLM_R_X33Y116_SLICE_X48Y116_CO6;
  assign CLBLM_R_X33Y116_SLICE_X48Y116_D = CLBLM_R_X33Y116_SLICE_X48Y116_DO6;
  assign CLBLM_R_X33Y116_SLICE_X49Y116_COUT = CLBLM_R_X33Y116_SLICE_X49Y116_D_CY;
  assign CLBLM_R_X33Y116_SLICE_X49Y116_A = CLBLM_R_X33Y116_SLICE_X49Y116_AO6;
  assign CLBLM_R_X33Y116_SLICE_X49Y116_B = CLBLM_R_X33Y116_SLICE_X49Y116_BO6;
  assign CLBLM_R_X33Y116_SLICE_X49Y116_C = CLBLM_R_X33Y116_SLICE_X49Y116_CO6;
  assign CLBLM_R_X33Y116_SLICE_X49Y116_D = CLBLM_R_X33Y116_SLICE_X49Y116_DO6;
  assign CLBLM_R_X33Y116_SLICE_X49Y116_DMUX = CLBLM_R_X33Y116_SLICE_X49Y116_DO6;
  assign CLBLM_R_X33Y117_SLICE_X48Y117_COUT = CLBLM_R_X33Y117_SLICE_X48Y117_D_CY;
  assign CLBLM_R_X33Y117_SLICE_X48Y117_A = CLBLM_R_X33Y117_SLICE_X48Y117_AO6;
  assign CLBLM_R_X33Y117_SLICE_X48Y117_B = CLBLM_R_X33Y117_SLICE_X48Y117_BO6;
  assign CLBLM_R_X33Y117_SLICE_X48Y117_C = CLBLM_R_X33Y117_SLICE_X48Y117_CO6;
  assign CLBLM_R_X33Y117_SLICE_X48Y117_D = CLBLM_R_X33Y117_SLICE_X48Y117_DO6;
  assign CLBLM_R_X33Y117_SLICE_X49Y117_COUT = CLBLM_R_X33Y117_SLICE_X49Y117_D_CY;
  assign CLBLM_R_X33Y117_SLICE_X49Y117_A = CLBLM_R_X33Y117_SLICE_X49Y117_AO6;
  assign CLBLM_R_X33Y117_SLICE_X49Y117_B = CLBLM_R_X33Y117_SLICE_X49Y117_BO6;
  assign CLBLM_R_X33Y117_SLICE_X49Y117_C = CLBLM_R_X33Y117_SLICE_X49Y117_CO6;
  assign CLBLM_R_X33Y117_SLICE_X49Y117_D = CLBLM_R_X33Y117_SLICE_X49Y117_DO6;
  assign CLBLM_R_X33Y118_SLICE_X48Y118_COUT = CLBLM_R_X33Y118_SLICE_X48Y118_D_CY;
  assign CLBLM_R_X33Y118_SLICE_X48Y118_A = CLBLM_R_X33Y118_SLICE_X48Y118_AO6;
  assign CLBLM_R_X33Y118_SLICE_X48Y118_B = CLBLM_R_X33Y118_SLICE_X48Y118_BO6;
  assign CLBLM_R_X33Y118_SLICE_X48Y118_C = CLBLM_R_X33Y118_SLICE_X48Y118_CO6;
  assign CLBLM_R_X33Y118_SLICE_X48Y118_D = CLBLM_R_X33Y118_SLICE_X48Y118_DO6;
  assign CLBLM_R_X33Y118_SLICE_X48Y118_AMUX = CLBLM_R_X33Y118_SLICE_X48Y118_AO5;
  assign CLBLM_R_X33Y118_SLICE_X49Y118_COUT = CLBLM_R_X33Y118_SLICE_X49Y118_D_CY;
  assign CLBLM_R_X33Y118_SLICE_X49Y118_A = CLBLM_R_X33Y118_SLICE_X49Y118_AO6;
  assign CLBLM_R_X33Y118_SLICE_X49Y118_B = CLBLM_R_X33Y118_SLICE_X49Y118_BO6;
  assign CLBLM_R_X33Y118_SLICE_X49Y118_C = CLBLM_R_X33Y118_SLICE_X49Y118_CO6;
  assign CLBLM_R_X33Y118_SLICE_X49Y118_D = CLBLM_R_X33Y118_SLICE_X49Y118_DO6;
  assign CLBLM_R_X33Y119_SLICE_X48Y119_COUT = CLBLM_R_X33Y119_SLICE_X48Y119_D_CY;
  assign CLBLM_R_X33Y119_SLICE_X48Y119_A = CLBLM_R_X33Y119_SLICE_X48Y119_AO6;
  assign CLBLM_R_X33Y119_SLICE_X48Y119_B = CLBLM_R_X33Y119_SLICE_X48Y119_BO6;
  assign CLBLM_R_X33Y119_SLICE_X48Y119_C = CLBLM_R_X33Y119_SLICE_X48Y119_CO6;
  assign CLBLM_R_X33Y119_SLICE_X48Y119_D = CLBLM_R_X33Y119_SLICE_X48Y119_DO6;
  assign CLBLM_R_X33Y119_SLICE_X49Y119_COUT = CLBLM_R_X33Y119_SLICE_X49Y119_D_CY;
  assign CLBLM_R_X33Y119_SLICE_X49Y119_A = CLBLM_R_X33Y119_SLICE_X49Y119_AO6;
  assign CLBLM_R_X33Y119_SLICE_X49Y119_B = CLBLM_R_X33Y119_SLICE_X49Y119_BO6;
  assign CLBLM_R_X33Y119_SLICE_X49Y119_C = CLBLM_R_X33Y119_SLICE_X49Y119_CO6;
  assign CLBLM_R_X33Y119_SLICE_X49Y119_D = CLBLM_R_X33Y119_SLICE_X49Y119_DO6;
  assign CLBLM_R_X33Y119_SLICE_X49Y119_AMUX = CLBLM_R_X33Y119_SLICE_X49Y119_AO6;
  assign CLBLM_R_X33Y119_SLICE_X49Y119_BMUX = CLBLM_R_X33Y119_SLICE_X49Y119_BO6;
  assign CLBLM_R_X33Y121_SLICE_X48Y121_COUT = CLBLM_R_X33Y121_SLICE_X48Y121_D_CY;
  assign CLBLM_R_X33Y121_SLICE_X48Y121_A = CLBLM_R_X33Y121_SLICE_X48Y121_AO6;
  assign CLBLM_R_X33Y121_SLICE_X48Y121_B = CLBLM_R_X33Y121_SLICE_X48Y121_BO6;
  assign CLBLM_R_X33Y121_SLICE_X48Y121_C = CLBLM_R_X33Y121_SLICE_X48Y121_CO6;
  assign CLBLM_R_X33Y121_SLICE_X48Y121_D = CLBLM_R_X33Y121_SLICE_X48Y121_DO6;
  assign CLBLM_R_X33Y121_SLICE_X48Y121_DMUX = CLBLM_R_X33Y121_SLICE_X48Y121_DO6;
  assign CLBLM_R_X33Y121_SLICE_X49Y121_COUT = CLBLM_R_X33Y121_SLICE_X49Y121_D_CY;
  assign CLBLM_R_X33Y121_SLICE_X49Y121_A = CLBLM_R_X33Y121_SLICE_X49Y121_AO6;
  assign CLBLM_R_X33Y121_SLICE_X49Y121_B = CLBLM_R_X33Y121_SLICE_X49Y121_BO6;
  assign CLBLM_R_X33Y121_SLICE_X49Y121_C = CLBLM_R_X33Y121_SLICE_X49Y121_CO6;
  assign CLBLM_R_X33Y121_SLICE_X49Y121_D = CLBLM_R_X33Y121_SLICE_X49Y121_DO6;
  assign CLBLM_R_X33Y122_SLICE_X48Y122_COUT = CLBLM_R_X33Y122_SLICE_X48Y122_D_CY;
  assign CLBLM_R_X33Y122_SLICE_X48Y122_A = CLBLM_R_X33Y122_SLICE_X48Y122_AO6;
  assign CLBLM_R_X33Y122_SLICE_X48Y122_B = CLBLM_R_X33Y122_SLICE_X48Y122_BO6;
  assign CLBLM_R_X33Y122_SLICE_X48Y122_C = CLBLM_R_X33Y122_SLICE_X48Y122_CO6;
  assign CLBLM_R_X33Y122_SLICE_X48Y122_D = CLBLM_R_X33Y122_SLICE_X48Y122_DO6;
  assign CLBLM_R_X33Y122_SLICE_X48Y122_AMUX = CLBLM_R_X33Y122_SLICE_X48Y122_AO5;
  assign CLBLM_R_X33Y122_SLICE_X49Y122_COUT = CLBLM_R_X33Y122_SLICE_X49Y122_D_CY;
  assign CLBLM_R_X33Y122_SLICE_X49Y122_A = CLBLM_R_X33Y122_SLICE_X49Y122_AO6;
  assign CLBLM_R_X33Y122_SLICE_X49Y122_B = CLBLM_R_X33Y122_SLICE_X49Y122_BO6;
  assign CLBLM_R_X33Y122_SLICE_X49Y122_C = CLBLM_R_X33Y122_SLICE_X49Y122_CO6;
  assign CLBLM_R_X33Y122_SLICE_X49Y122_D = CLBLM_R_X33Y122_SLICE_X49Y122_DO6;
  assign CLBLM_R_X33Y123_SLICE_X48Y123_COUT = CLBLM_R_X33Y123_SLICE_X48Y123_D_CY;
  assign CLBLM_R_X33Y123_SLICE_X48Y123_A = CLBLM_R_X33Y123_SLICE_X48Y123_AO6;
  assign CLBLM_R_X33Y123_SLICE_X48Y123_B = CLBLM_R_X33Y123_SLICE_X48Y123_BO6;
  assign CLBLM_R_X33Y123_SLICE_X48Y123_C = CLBLM_R_X33Y123_SLICE_X48Y123_CO6;
  assign CLBLM_R_X33Y123_SLICE_X48Y123_D = CLBLM_R_X33Y123_SLICE_X48Y123_DO6;
  assign CLBLM_R_X33Y123_SLICE_X48Y123_DMUX = CLBLM_R_X33Y123_SLICE_X48Y123_DO6;
  assign CLBLM_R_X33Y123_SLICE_X49Y123_COUT = CLBLM_R_X33Y123_SLICE_X49Y123_D_CY;
  assign CLBLM_R_X33Y123_SLICE_X49Y123_A = CLBLM_R_X33Y123_SLICE_X49Y123_AO6;
  assign CLBLM_R_X33Y123_SLICE_X49Y123_B = CLBLM_R_X33Y123_SLICE_X49Y123_BO6;
  assign CLBLM_R_X33Y123_SLICE_X49Y123_C = CLBLM_R_X33Y123_SLICE_X49Y123_CO6;
  assign CLBLM_R_X33Y123_SLICE_X49Y123_D = CLBLM_R_X33Y123_SLICE_X49Y123_DO6;
  assign CLBLM_R_X33Y124_SLICE_X48Y124_COUT = CLBLM_R_X33Y124_SLICE_X48Y124_D_CY;
  assign CLBLM_R_X33Y124_SLICE_X48Y124_A = CLBLM_R_X33Y124_SLICE_X48Y124_AO6;
  assign CLBLM_R_X33Y124_SLICE_X48Y124_B = CLBLM_R_X33Y124_SLICE_X48Y124_BO6;
  assign CLBLM_R_X33Y124_SLICE_X48Y124_C = CLBLM_R_X33Y124_SLICE_X48Y124_CO6;
  assign CLBLM_R_X33Y124_SLICE_X48Y124_D = CLBLM_R_X33Y124_SLICE_X48Y124_DO6;
  assign CLBLM_R_X33Y124_SLICE_X48Y124_AMUX = CLBLM_R_X33Y124_SLICE_X48Y124_AO5;
  assign CLBLM_R_X33Y124_SLICE_X49Y124_COUT = CLBLM_R_X33Y124_SLICE_X49Y124_D_CY;
  assign CLBLM_R_X33Y124_SLICE_X49Y124_A = CLBLM_R_X33Y124_SLICE_X49Y124_AO6;
  assign CLBLM_R_X33Y124_SLICE_X49Y124_B = CLBLM_R_X33Y124_SLICE_X49Y124_BO6;
  assign CLBLM_R_X33Y124_SLICE_X49Y124_C = CLBLM_R_X33Y124_SLICE_X49Y124_CO6;
  assign CLBLM_R_X33Y124_SLICE_X49Y124_D = CLBLM_R_X33Y124_SLICE_X49Y124_DO6;
  assign CLBLM_R_X33Y124_SLICE_X49Y124_AMUX = CLBLM_R_X33Y124_SLICE_X49Y124_AO5;
  assign CLBLM_R_X33Y125_SLICE_X48Y125_COUT = CLBLM_R_X33Y125_SLICE_X48Y125_D_CY;
  assign CLBLM_R_X33Y125_SLICE_X48Y125_A = CLBLM_R_X33Y125_SLICE_X48Y125_AO6;
  assign CLBLM_R_X33Y125_SLICE_X48Y125_B = CLBLM_R_X33Y125_SLICE_X48Y125_BO6;
  assign CLBLM_R_X33Y125_SLICE_X48Y125_C = CLBLM_R_X33Y125_SLICE_X48Y125_CO6;
  assign CLBLM_R_X33Y125_SLICE_X48Y125_D = CLBLM_R_X33Y125_SLICE_X48Y125_DO6;
  assign CLBLM_R_X33Y125_SLICE_X49Y125_COUT = CLBLM_R_X33Y125_SLICE_X49Y125_D_CY;
  assign CLBLM_R_X33Y125_SLICE_X49Y125_A = CLBLM_R_X33Y125_SLICE_X49Y125_AO6;
  assign CLBLM_R_X33Y125_SLICE_X49Y125_B = CLBLM_R_X33Y125_SLICE_X49Y125_BO6;
  assign CLBLM_R_X33Y125_SLICE_X49Y125_C = CLBLM_R_X33Y125_SLICE_X49Y125_CO6;
  assign CLBLM_R_X33Y125_SLICE_X49Y125_D = CLBLM_R_X33Y125_SLICE_X49Y125_DO6;
  assign CLBLM_R_X33Y125_SLICE_X49Y125_AMUX = CLBLM_R_X33Y125_SLICE_X49Y125_AO5;
  assign CLBLM_R_X33Y125_SLICE_X49Y125_BMUX = CLBLM_R_X33Y125_SLICE_X49Y125_BO5;
  assign CLBLM_R_X35Y114_SLICE_X52Y114_COUT = CLBLM_R_X35Y114_SLICE_X52Y114_D_CY;
  assign CLBLM_R_X35Y114_SLICE_X52Y114_A = CLBLM_R_X35Y114_SLICE_X52Y114_AO6;
  assign CLBLM_R_X35Y114_SLICE_X52Y114_B = CLBLM_R_X35Y114_SLICE_X52Y114_BO6;
  assign CLBLM_R_X35Y114_SLICE_X52Y114_C = CLBLM_R_X35Y114_SLICE_X52Y114_CO6;
  assign CLBLM_R_X35Y114_SLICE_X52Y114_D = CLBLM_R_X35Y114_SLICE_X52Y114_DO6;
  assign CLBLM_R_X35Y114_SLICE_X53Y114_COUT = CLBLM_R_X35Y114_SLICE_X53Y114_D_CY;
  assign CLBLM_R_X35Y114_SLICE_X53Y114_A = CLBLM_R_X35Y114_SLICE_X53Y114_AO6;
  assign CLBLM_R_X35Y114_SLICE_X53Y114_B = CLBLM_R_X35Y114_SLICE_X53Y114_BO6;
  assign CLBLM_R_X35Y114_SLICE_X53Y114_C = CLBLM_R_X35Y114_SLICE_X53Y114_CO6;
  assign CLBLM_R_X35Y114_SLICE_X53Y114_D = CLBLM_R_X35Y114_SLICE_X53Y114_DO6;
  assign CLBLM_R_X35Y115_SLICE_X52Y115_COUT = CLBLM_R_X35Y115_SLICE_X52Y115_D_CY;
  assign CLBLM_R_X35Y115_SLICE_X52Y115_A = CLBLM_R_X35Y115_SLICE_X52Y115_AO6;
  assign CLBLM_R_X35Y115_SLICE_X52Y115_B = CLBLM_R_X35Y115_SLICE_X52Y115_BO6;
  assign CLBLM_R_X35Y115_SLICE_X52Y115_C = CLBLM_R_X35Y115_SLICE_X52Y115_CO6;
  assign CLBLM_R_X35Y115_SLICE_X52Y115_D = CLBLM_R_X35Y115_SLICE_X52Y115_DO6;
  assign CLBLM_R_X35Y115_SLICE_X52Y115_AMUX = CLBLM_R_X35Y115_SLICE_X52Y115_AO5;
  assign CLBLM_R_X35Y115_SLICE_X53Y115_COUT = CLBLM_R_X35Y115_SLICE_X53Y115_D_CY;
  assign CLBLM_R_X35Y115_SLICE_X53Y115_A = CLBLM_R_X35Y115_SLICE_X53Y115_AO6;
  assign CLBLM_R_X35Y115_SLICE_X53Y115_B = CLBLM_R_X35Y115_SLICE_X53Y115_BO6;
  assign CLBLM_R_X35Y115_SLICE_X53Y115_C = CLBLM_R_X35Y115_SLICE_X53Y115_CO6;
  assign CLBLM_R_X35Y115_SLICE_X53Y115_D = CLBLM_R_X35Y115_SLICE_X53Y115_DO6;
  assign CLBLM_R_X35Y115_SLICE_X53Y115_CMUX = CLBLM_R_X35Y115_SLICE_X53Y115_CO6;
  assign CLBLM_R_X35Y116_SLICE_X52Y116_COUT = CLBLM_R_X35Y116_SLICE_X52Y116_D_CY;
  assign CLBLM_R_X35Y116_SLICE_X52Y116_A = CLBLM_R_X35Y116_SLICE_X52Y116_AO6;
  assign CLBLM_R_X35Y116_SLICE_X52Y116_B = CLBLM_R_X35Y116_SLICE_X52Y116_BO6;
  assign CLBLM_R_X35Y116_SLICE_X52Y116_C = CLBLM_R_X35Y116_SLICE_X52Y116_CO6;
  assign CLBLM_R_X35Y116_SLICE_X52Y116_D = CLBLM_R_X35Y116_SLICE_X52Y116_DO6;
  assign CLBLM_R_X35Y116_SLICE_X52Y116_AMUX = CLBLM_R_X35Y116_SLICE_X52Y116_AO6;
  assign CLBLM_R_X35Y116_SLICE_X53Y116_COUT = CLBLM_R_X35Y116_SLICE_X53Y116_D_CY;
  assign CLBLM_R_X35Y116_SLICE_X53Y116_A = CLBLM_R_X35Y116_SLICE_X53Y116_AO6;
  assign CLBLM_R_X35Y116_SLICE_X53Y116_B = CLBLM_R_X35Y116_SLICE_X53Y116_BO6;
  assign CLBLM_R_X35Y116_SLICE_X53Y116_C = CLBLM_R_X35Y116_SLICE_X53Y116_CO6;
  assign CLBLM_R_X35Y116_SLICE_X53Y116_D = CLBLM_R_X35Y116_SLICE_X53Y116_DO6;
  assign CLBLM_R_X35Y117_SLICE_X52Y117_COUT = CLBLM_R_X35Y117_SLICE_X52Y117_D_CY;
  assign CLBLM_R_X35Y117_SLICE_X52Y117_A = CLBLM_R_X35Y117_SLICE_X52Y117_AO6;
  assign CLBLM_R_X35Y117_SLICE_X52Y117_B = CLBLM_R_X35Y117_SLICE_X52Y117_BO6;
  assign CLBLM_R_X35Y117_SLICE_X52Y117_C = CLBLM_R_X35Y117_SLICE_X52Y117_CO6;
  assign CLBLM_R_X35Y117_SLICE_X52Y117_D = CLBLM_R_X35Y117_SLICE_X52Y117_DO6;
  assign CLBLM_R_X35Y117_SLICE_X52Y117_AMUX = CLBLM_R_X35Y117_SLICE_X52Y117_AO6;
  assign CLBLM_R_X35Y117_SLICE_X53Y117_COUT = CLBLM_R_X35Y117_SLICE_X53Y117_D_CY;
  assign CLBLM_R_X35Y117_SLICE_X53Y117_A = CLBLM_R_X35Y117_SLICE_X53Y117_AO6;
  assign CLBLM_R_X35Y117_SLICE_X53Y117_B = CLBLM_R_X35Y117_SLICE_X53Y117_BO6;
  assign CLBLM_R_X35Y117_SLICE_X53Y117_C = CLBLM_R_X35Y117_SLICE_X53Y117_CO6;
  assign CLBLM_R_X35Y117_SLICE_X53Y117_D = CLBLM_R_X35Y117_SLICE_X53Y117_DO6;
  assign CLBLM_R_X35Y117_SLICE_X53Y117_BMUX = CLBLM_R_X35Y117_SLICE_X53Y117_BO6;
  assign CLBLM_R_X35Y118_SLICE_X52Y118_COUT = CLBLM_R_X35Y118_SLICE_X52Y118_D_CY;
  assign CLBLM_R_X35Y118_SLICE_X52Y118_A = CLBLM_R_X35Y118_SLICE_X52Y118_AO6;
  assign CLBLM_R_X35Y118_SLICE_X52Y118_B = CLBLM_R_X35Y118_SLICE_X52Y118_BO6;
  assign CLBLM_R_X35Y118_SLICE_X52Y118_C = CLBLM_R_X35Y118_SLICE_X52Y118_CO6;
  assign CLBLM_R_X35Y118_SLICE_X52Y118_D = CLBLM_R_X35Y118_SLICE_X52Y118_DO6;
  assign CLBLM_R_X35Y118_SLICE_X52Y118_AMUX = CLBLM_R_X35Y118_SLICE_X52Y118_A_XOR;
  assign CLBLM_R_X35Y118_SLICE_X52Y118_BMUX = CLBLM_R_X35Y118_SLICE_X52Y118_B_XOR;
  assign CLBLM_R_X35Y118_SLICE_X52Y118_CMUX = CLBLM_R_X35Y118_SLICE_X52Y118_C_XOR;
  assign CLBLM_R_X35Y118_SLICE_X52Y118_DMUX = CLBLM_R_X35Y118_SLICE_X52Y118_D_XOR;
  assign CLBLM_R_X35Y118_SLICE_X53Y118_COUT = CLBLM_R_X35Y118_SLICE_X53Y118_D_CY;
  assign CLBLM_R_X35Y118_SLICE_X53Y118_A = CLBLM_R_X35Y118_SLICE_X53Y118_AO6;
  assign CLBLM_R_X35Y118_SLICE_X53Y118_B = CLBLM_R_X35Y118_SLICE_X53Y118_BO6;
  assign CLBLM_R_X35Y118_SLICE_X53Y118_C = CLBLM_R_X35Y118_SLICE_X53Y118_CO6;
  assign CLBLM_R_X35Y118_SLICE_X53Y118_D = CLBLM_R_X35Y118_SLICE_X53Y118_DO6;
  assign CLBLM_R_X35Y118_SLICE_X53Y118_AMUX = CLBLM_R_X35Y118_SLICE_X53Y118_AO5;
  assign CLBLM_R_X35Y118_SLICE_X53Y118_BMUX = CLBLM_R_X35Y118_SLICE_X53Y118_BO5;
  assign CLBLM_R_X35Y119_SLICE_X52Y119_COUT = CLBLM_R_X35Y119_SLICE_X52Y119_D_CY;
  assign CLBLM_R_X35Y119_SLICE_X52Y119_A = CLBLM_R_X35Y119_SLICE_X52Y119_AO6;
  assign CLBLM_R_X35Y119_SLICE_X52Y119_B = CLBLM_R_X35Y119_SLICE_X52Y119_BO6;
  assign CLBLM_R_X35Y119_SLICE_X52Y119_C = CLBLM_R_X35Y119_SLICE_X52Y119_CO6;
  assign CLBLM_R_X35Y119_SLICE_X52Y119_D = CLBLM_R_X35Y119_SLICE_X52Y119_DO6;
  assign CLBLM_R_X35Y119_SLICE_X52Y119_AMUX = CLBLM_R_X35Y119_SLICE_X52Y119_A_XOR;
  assign CLBLM_R_X35Y119_SLICE_X52Y119_BMUX = CLBLM_R_X35Y119_SLICE_X52Y119_B_XOR;
  assign CLBLM_R_X35Y119_SLICE_X52Y119_CMUX = CLBLM_R_X35Y119_SLICE_X52Y119_C_XOR;
  assign CLBLM_R_X35Y119_SLICE_X52Y119_DMUX = CLBLM_R_X35Y119_SLICE_X52Y119_D_XOR;
  assign CLBLM_R_X35Y119_SLICE_X53Y119_COUT = CLBLM_R_X35Y119_SLICE_X53Y119_D_CY;
  assign CLBLM_R_X35Y119_SLICE_X53Y119_A = CLBLM_R_X35Y119_SLICE_X53Y119_AO6;
  assign CLBLM_R_X35Y119_SLICE_X53Y119_B = CLBLM_R_X35Y119_SLICE_X53Y119_BO6;
  assign CLBLM_R_X35Y119_SLICE_X53Y119_C = CLBLM_R_X35Y119_SLICE_X53Y119_CO6;
  assign CLBLM_R_X35Y119_SLICE_X53Y119_D = CLBLM_R_X35Y119_SLICE_X53Y119_DO6;
  assign CLBLM_R_X35Y120_SLICE_X52Y120_COUT = CLBLM_R_X35Y120_SLICE_X52Y120_D_CY;
  assign CLBLM_R_X35Y120_SLICE_X52Y120_A = CLBLM_R_X35Y120_SLICE_X52Y120_AO6;
  assign CLBLM_R_X35Y120_SLICE_X52Y120_B = CLBLM_R_X35Y120_SLICE_X52Y120_BO6;
  assign CLBLM_R_X35Y120_SLICE_X52Y120_C = CLBLM_R_X35Y120_SLICE_X52Y120_CO6;
  assign CLBLM_R_X35Y120_SLICE_X52Y120_D = CLBLM_R_X35Y120_SLICE_X52Y120_DO6;
  assign CLBLM_R_X35Y120_SLICE_X52Y120_AMUX = CLBLM_R_X35Y120_SLICE_X52Y120_A_XOR;
  assign CLBLM_R_X35Y120_SLICE_X52Y120_BMUX = CLBLM_R_X35Y120_SLICE_X52Y120_B_XOR;
  assign CLBLM_R_X35Y120_SLICE_X52Y120_CMUX = CLBLM_R_X35Y120_SLICE_X52Y120_C_XOR;
  assign CLBLM_R_X35Y120_SLICE_X52Y120_DMUX = CLBLM_R_X35Y120_SLICE_X52Y120_D_XOR;
  assign CLBLM_R_X35Y120_SLICE_X53Y120_COUT = CLBLM_R_X35Y120_SLICE_X53Y120_D_CY;
  assign CLBLM_R_X35Y120_SLICE_X53Y120_A = CLBLM_R_X35Y120_SLICE_X53Y120_AO6;
  assign CLBLM_R_X35Y120_SLICE_X53Y120_B = CLBLM_R_X35Y120_SLICE_X53Y120_BO6;
  assign CLBLM_R_X35Y120_SLICE_X53Y120_C = CLBLM_R_X35Y120_SLICE_X53Y120_CO6;
  assign CLBLM_R_X35Y120_SLICE_X53Y120_D = CLBLM_R_X35Y120_SLICE_X53Y120_DO6;
  assign CLBLM_R_X35Y120_SLICE_X53Y120_AMUX = CLBLM_R_X35Y120_SLICE_X53Y120_A_XOR;
  assign CLBLM_R_X35Y120_SLICE_X53Y120_BMUX = CLBLM_R_X35Y120_SLICE_X53Y120_B_XOR;
  assign CLBLM_R_X35Y120_SLICE_X53Y120_CMUX = CLBLM_R_X35Y120_SLICE_X53Y120_C_XOR;
  assign CLBLM_R_X35Y120_SLICE_X53Y120_DMUX = CLBLM_R_X35Y120_SLICE_X53Y120_D_XOR;
  assign CLBLM_R_X35Y121_SLICE_X52Y121_COUT = CLBLM_R_X35Y121_SLICE_X52Y121_D_CY;
  assign CLBLM_R_X35Y121_SLICE_X52Y121_A = CLBLM_R_X35Y121_SLICE_X52Y121_AO6;
  assign CLBLM_R_X35Y121_SLICE_X52Y121_B = CLBLM_R_X35Y121_SLICE_X52Y121_BO6;
  assign CLBLM_R_X35Y121_SLICE_X52Y121_C = CLBLM_R_X35Y121_SLICE_X52Y121_CO6;
  assign CLBLM_R_X35Y121_SLICE_X52Y121_D = CLBLM_R_X35Y121_SLICE_X52Y121_DO6;
  assign CLBLM_R_X35Y121_SLICE_X52Y121_AMUX = CLBLM_R_X35Y121_SLICE_X52Y121_A_XOR;
  assign CLBLM_R_X35Y121_SLICE_X52Y121_BMUX = CLBLM_R_X35Y121_SLICE_X52Y121_B_XOR;
  assign CLBLM_R_X35Y121_SLICE_X52Y121_CMUX = CLBLM_R_X35Y121_SLICE_X52Y121_C_XOR;
  assign CLBLM_R_X35Y121_SLICE_X52Y121_DMUX = CLBLM_R_X35Y121_SLICE_X52Y121_D_XOR;
  assign CLBLM_R_X35Y121_SLICE_X53Y121_COUT = CLBLM_R_X35Y121_SLICE_X53Y121_D_CY;
  assign CLBLM_R_X35Y121_SLICE_X53Y121_A = CLBLM_R_X35Y121_SLICE_X53Y121_AO6;
  assign CLBLM_R_X35Y121_SLICE_X53Y121_B = CLBLM_R_X35Y121_SLICE_X53Y121_BO6;
  assign CLBLM_R_X35Y121_SLICE_X53Y121_C = CLBLM_R_X35Y121_SLICE_X53Y121_CO6;
  assign CLBLM_R_X35Y121_SLICE_X53Y121_D = CLBLM_R_X35Y121_SLICE_X53Y121_DO6;
  assign CLBLM_R_X35Y121_SLICE_X53Y121_AMUX = CLBLM_R_X35Y121_SLICE_X53Y121_A_XOR;
  assign CLBLM_R_X35Y121_SLICE_X53Y121_BMUX = CLBLM_R_X35Y121_SLICE_X53Y121_B_XOR;
  assign CLBLM_R_X35Y121_SLICE_X53Y121_CMUX = CLBLM_R_X35Y121_SLICE_X53Y121_C_XOR;
  assign CLBLM_R_X35Y121_SLICE_X53Y121_DMUX = CLBLM_R_X35Y121_SLICE_X53Y121_D_XOR;
  assign CLBLM_R_X35Y122_SLICE_X52Y122_COUT = CLBLM_R_X35Y122_SLICE_X52Y122_D_CY;
  assign CLBLM_R_X35Y122_SLICE_X52Y122_A = CLBLM_R_X35Y122_SLICE_X52Y122_AO6;
  assign CLBLM_R_X35Y122_SLICE_X52Y122_B = CLBLM_R_X35Y122_SLICE_X52Y122_BO6;
  assign CLBLM_R_X35Y122_SLICE_X52Y122_C = CLBLM_R_X35Y122_SLICE_X52Y122_CO6;
  assign CLBLM_R_X35Y122_SLICE_X52Y122_D = CLBLM_R_X35Y122_SLICE_X52Y122_DO6;
  assign CLBLM_R_X35Y122_SLICE_X52Y122_AMUX = CLBLM_R_X35Y122_SLICE_X52Y122_A_XOR;
  assign CLBLM_R_X35Y122_SLICE_X52Y122_BMUX = CLBLM_R_X35Y122_SLICE_X52Y122_B_XOR;
  assign CLBLM_R_X35Y122_SLICE_X52Y122_CMUX = CLBLM_R_X35Y122_SLICE_X52Y122_C_XOR;
  assign CLBLM_R_X35Y122_SLICE_X52Y122_DMUX = CLBLM_R_X35Y122_SLICE_X52Y122_D_XOR;
  assign CLBLM_R_X35Y122_SLICE_X53Y122_COUT = CLBLM_R_X35Y122_SLICE_X53Y122_D_CY;
  assign CLBLM_R_X35Y122_SLICE_X53Y122_A = CLBLM_R_X35Y122_SLICE_X53Y122_AO6;
  assign CLBLM_R_X35Y122_SLICE_X53Y122_B = CLBLM_R_X35Y122_SLICE_X53Y122_BO6;
  assign CLBLM_R_X35Y122_SLICE_X53Y122_C = CLBLM_R_X35Y122_SLICE_X53Y122_CO6;
  assign CLBLM_R_X35Y122_SLICE_X53Y122_D = CLBLM_R_X35Y122_SLICE_X53Y122_DO6;
  assign CLBLM_R_X35Y122_SLICE_X53Y122_AMUX = CLBLM_R_X35Y122_SLICE_X53Y122_A_XOR;
  assign CLBLM_R_X35Y122_SLICE_X53Y122_BMUX = CLBLM_R_X35Y122_SLICE_X53Y122_B_XOR;
  assign CLBLM_R_X35Y122_SLICE_X53Y122_CMUX = CLBLM_R_X35Y122_SLICE_X53Y122_C_XOR;
  assign CLBLM_R_X35Y122_SLICE_X53Y122_DMUX = CLBLM_R_X35Y122_SLICE_X53Y122_D_XOR;
  assign CLBLM_R_X35Y123_SLICE_X52Y123_COUT = CLBLM_R_X35Y123_SLICE_X52Y123_D_CY;
  assign CLBLM_R_X35Y123_SLICE_X52Y123_A = CLBLM_R_X35Y123_SLICE_X52Y123_AO6;
  assign CLBLM_R_X35Y123_SLICE_X52Y123_B = CLBLM_R_X35Y123_SLICE_X52Y123_BO6;
  assign CLBLM_R_X35Y123_SLICE_X52Y123_C = CLBLM_R_X35Y123_SLICE_X52Y123_CO6;
  assign CLBLM_R_X35Y123_SLICE_X52Y123_D = CLBLM_R_X35Y123_SLICE_X52Y123_DO6;
  assign CLBLM_R_X35Y123_SLICE_X52Y123_AMUX = CLBLM_R_X35Y123_SLICE_X52Y123_A_XOR;
  assign CLBLM_R_X35Y123_SLICE_X52Y123_BMUX = CLBLM_R_X35Y123_SLICE_X52Y123_B_XOR;
  assign CLBLM_R_X35Y123_SLICE_X52Y123_CMUX = CLBLM_R_X35Y123_SLICE_X52Y123_C_XOR;
  assign CLBLM_R_X35Y123_SLICE_X52Y123_DMUX = CLBLM_R_X35Y123_SLICE_X52Y123_D_XOR;
  assign CLBLM_R_X35Y123_SLICE_X53Y123_COUT = CLBLM_R_X35Y123_SLICE_X53Y123_D_CY;
  assign CLBLM_R_X35Y123_SLICE_X53Y123_A = CLBLM_R_X35Y123_SLICE_X53Y123_AO6;
  assign CLBLM_R_X35Y123_SLICE_X53Y123_B = CLBLM_R_X35Y123_SLICE_X53Y123_BO6;
  assign CLBLM_R_X35Y123_SLICE_X53Y123_C = CLBLM_R_X35Y123_SLICE_X53Y123_CO6;
  assign CLBLM_R_X35Y123_SLICE_X53Y123_D = CLBLM_R_X35Y123_SLICE_X53Y123_DO6;
  assign CLBLM_R_X35Y123_SLICE_X53Y123_AMUX = CLBLM_R_X35Y123_SLICE_X53Y123_A_XOR;
  assign CLBLM_R_X35Y123_SLICE_X53Y123_BMUX = CLBLM_R_X35Y123_SLICE_X53Y123_B_XOR;
  assign CLBLM_R_X35Y123_SLICE_X53Y123_CMUX = CLBLM_R_X35Y123_SLICE_X53Y123_C_XOR;
  assign CLBLM_R_X35Y123_SLICE_X53Y123_DMUX = CLBLM_R_X35Y123_SLICE_X53Y123_D_XOR;
  assign CLBLM_R_X35Y124_SLICE_X52Y124_COUT = CLBLM_R_X35Y124_SLICE_X52Y124_D_CY;
  assign CLBLM_R_X35Y124_SLICE_X52Y124_A = CLBLM_R_X35Y124_SLICE_X52Y124_AO6;
  assign CLBLM_R_X35Y124_SLICE_X52Y124_B = CLBLM_R_X35Y124_SLICE_X52Y124_BO6;
  assign CLBLM_R_X35Y124_SLICE_X52Y124_C = CLBLM_R_X35Y124_SLICE_X52Y124_CO6;
  assign CLBLM_R_X35Y124_SLICE_X52Y124_D = CLBLM_R_X35Y124_SLICE_X52Y124_DO6;
  assign CLBLM_R_X35Y124_SLICE_X52Y124_AMUX = CLBLM_R_X35Y124_SLICE_X52Y124_A_XOR;
  assign CLBLM_R_X35Y124_SLICE_X52Y124_BMUX = CLBLM_R_X35Y124_SLICE_X52Y124_B_XOR;
  assign CLBLM_R_X35Y124_SLICE_X52Y124_CMUX = CLBLM_R_X35Y124_SLICE_X52Y124_C_XOR;
  assign CLBLM_R_X35Y124_SLICE_X52Y124_DMUX = CLBLM_R_X35Y124_SLICE_X52Y124_D_XOR;
  assign CLBLM_R_X35Y124_SLICE_X53Y124_COUT = CLBLM_R_X35Y124_SLICE_X53Y124_D_CY;
  assign CLBLM_R_X35Y124_SLICE_X53Y124_A = CLBLM_R_X35Y124_SLICE_X53Y124_AO6;
  assign CLBLM_R_X35Y124_SLICE_X53Y124_B = CLBLM_R_X35Y124_SLICE_X53Y124_BO6;
  assign CLBLM_R_X35Y124_SLICE_X53Y124_C = CLBLM_R_X35Y124_SLICE_X53Y124_CO6;
  assign CLBLM_R_X35Y124_SLICE_X53Y124_D = CLBLM_R_X35Y124_SLICE_X53Y124_DO6;
  assign CLBLM_R_X35Y124_SLICE_X53Y124_AMUX = CLBLM_R_X35Y124_SLICE_X53Y124_A_XOR;
  assign CLBLM_R_X35Y124_SLICE_X53Y124_BMUX = CLBLM_R_X35Y124_SLICE_X53Y124_B_XOR;
  assign CLBLM_R_X35Y124_SLICE_X53Y124_CMUX = CLBLM_R_X35Y124_SLICE_X53Y124_C_XOR;
  assign CLBLM_R_X35Y124_SLICE_X53Y124_DMUX = CLBLM_R_X35Y124_SLICE_X53Y124_D_XOR;
  assign CLBLM_R_X35Y125_SLICE_X52Y125_COUT = CLBLM_R_X35Y125_SLICE_X52Y125_D_CY;
  assign CLBLM_R_X35Y125_SLICE_X52Y125_A = CLBLM_R_X35Y125_SLICE_X52Y125_AO6;
  assign CLBLM_R_X35Y125_SLICE_X52Y125_B = CLBLM_R_X35Y125_SLICE_X52Y125_BO6;
  assign CLBLM_R_X35Y125_SLICE_X52Y125_C = CLBLM_R_X35Y125_SLICE_X52Y125_CO6;
  assign CLBLM_R_X35Y125_SLICE_X52Y125_D = CLBLM_R_X35Y125_SLICE_X52Y125_DO6;
  assign CLBLM_R_X35Y125_SLICE_X52Y125_AMUX = CLBLM_R_X35Y125_SLICE_X52Y125_A_XOR;
  assign CLBLM_R_X35Y125_SLICE_X52Y125_BMUX = CLBLM_R_X35Y125_SLICE_X52Y125_B_XOR;
  assign CLBLM_R_X35Y125_SLICE_X52Y125_CMUX = CLBLM_R_X35Y125_SLICE_X52Y125_C_XOR;
  assign CLBLM_R_X35Y125_SLICE_X52Y125_DMUX = CLBLM_R_X35Y125_SLICE_X52Y125_D_XOR;
  assign CLBLM_R_X35Y125_SLICE_X53Y125_COUT = CLBLM_R_X35Y125_SLICE_X53Y125_D_CY;
  assign CLBLM_R_X35Y125_SLICE_X53Y125_A = CLBLM_R_X35Y125_SLICE_X53Y125_AO6;
  assign CLBLM_R_X35Y125_SLICE_X53Y125_B = CLBLM_R_X35Y125_SLICE_X53Y125_BO6;
  assign CLBLM_R_X35Y125_SLICE_X53Y125_C = CLBLM_R_X35Y125_SLICE_X53Y125_CO6;
  assign CLBLM_R_X35Y125_SLICE_X53Y125_D = CLBLM_R_X35Y125_SLICE_X53Y125_DO6;
  assign CLBLM_R_X35Y125_SLICE_X53Y125_AMUX = CLBLM_R_X35Y125_SLICE_X53Y125_A_XOR;
  assign CLBLM_R_X35Y125_SLICE_X53Y125_BMUX = CLBLM_R_X35Y125_SLICE_X53Y125_B_XOR;
  assign CLBLM_R_X35Y125_SLICE_X53Y125_CMUX = CLBLM_R_X35Y125_SLICE_X53Y125_C_XOR;
  assign CLBLM_R_X35Y125_SLICE_X53Y125_DMUX = CLBLM_R_X35Y125_SLICE_X53Y125_D_XOR;
  assign CLBLM_R_X35Y126_SLICE_X52Y126_COUT = CLBLM_R_X35Y126_SLICE_X52Y126_D_CY;
  assign CLBLM_R_X35Y126_SLICE_X52Y126_A = CLBLM_R_X35Y126_SLICE_X52Y126_AO6;
  assign CLBLM_R_X35Y126_SLICE_X52Y126_B = CLBLM_R_X35Y126_SLICE_X52Y126_BO6;
  assign CLBLM_R_X35Y126_SLICE_X52Y126_C = CLBLM_R_X35Y126_SLICE_X52Y126_CO6;
  assign CLBLM_R_X35Y126_SLICE_X52Y126_D = CLBLM_R_X35Y126_SLICE_X52Y126_DO6;
  assign CLBLM_R_X35Y126_SLICE_X53Y126_COUT = CLBLM_R_X35Y126_SLICE_X53Y126_D_CY;
  assign CLBLM_R_X35Y126_SLICE_X53Y126_A = CLBLM_R_X35Y126_SLICE_X53Y126_AO6;
  assign CLBLM_R_X35Y126_SLICE_X53Y126_B = CLBLM_R_X35Y126_SLICE_X53Y126_BO6;
  assign CLBLM_R_X35Y126_SLICE_X53Y126_C = CLBLM_R_X35Y126_SLICE_X53Y126_CO6;
  assign CLBLM_R_X35Y126_SLICE_X53Y126_D = CLBLM_R_X35Y126_SLICE_X53Y126_DO6;
  assign CLBLM_R_X35Y126_SLICE_X53Y126_AMUX = CLBLM_R_X35Y126_SLICE_X53Y126_A_XOR;
  assign CLBLM_R_X35Y126_SLICE_X53Y126_BMUX = CLBLM_R_X35Y126_SLICE_X53Y126_B_XOR;
  assign CLBLM_R_X35Y126_SLICE_X53Y126_CMUX = CLBLM_R_X35Y126_SLICE_X53Y126_C_XOR;
  assign CLBLM_R_X35Y126_SLICE_X53Y126_DMUX = CLBLM_R_X35Y126_SLICE_X53Y126_D_XOR;
  assign CLBLM_R_X35Y127_SLICE_X52Y127_COUT = CLBLM_R_X35Y127_SLICE_X52Y127_D_CY;
  assign CLBLM_R_X35Y127_SLICE_X52Y127_A = CLBLM_R_X35Y127_SLICE_X52Y127_AO6;
  assign CLBLM_R_X35Y127_SLICE_X52Y127_B = CLBLM_R_X35Y127_SLICE_X52Y127_BO6;
  assign CLBLM_R_X35Y127_SLICE_X52Y127_C = CLBLM_R_X35Y127_SLICE_X52Y127_CO6;
  assign CLBLM_R_X35Y127_SLICE_X52Y127_D = CLBLM_R_X35Y127_SLICE_X52Y127_DO6;
  assign CLBLM_R_X35Y127_SLICE_X52Y127_DMUX = CLBLM_R_X35Y127_SLICE_X52Y127_DO6;
  assign CLBLM_R_X35Y127_SLICE_X53Y127_COUT = CLBLM_R_X35Y127_SLICE_X53Y127_D_CY;
  assign CLBLM_R_X35Y127_SLICE_X53Y127_A = CLBLM_R_X35Y127_SLICE_X53Y127_AO6;
  assign CLBLM_R_X35Y127_SLICE_X53Y127_B = CLBLM_R_X35Y127_SLICE_X53Y127_BO6;
  assign CLBLM_R_X35Y127_SLICE_X53Y127_C = CLBLM_R_X35Y127_SLICE_X53Y127_CO6;
  assign CLBLM_R_X35Y127_SLICE_X53Y127_D = CLBLM_R_X35Y127_SLICE_X53Y127_DO6;
  assign CLBLM_R_X35Y127_SLICE_X53Y127_AMUX = CLBLM_R_X35Y127_SLICE_X53Y127_A_XOR;
  assign CLBLM_R_X35Y127_SLICE_X53Y127_BMUX = CLBLM_R_X35Y127_SLICE_X53Y127_B_XOR;
  assign CLBLM_R_X35Y127_SLICE_X53Y127_CMUX = CLBLM_R_X35Y127_SLICE_X53Y127_C_XOR;
  assign CLBLM_R_X35Y127_SLICE_X53Y127_DMUX = CLBLM_R_X35Y127_SLICE_X53Y127_D_XOR;
  assign CLBLM_R_X35Y128_SLICE_X52Y128_COUT = CLBLM_R_X35Y128_SLICE_X52Y128_D_CY;
  assign CLBLM_R_X35Y128_SLICE_X52Y128_A = CLBLM_R_X35Y128_SLICE_X52Y128_AO6;
  assign CLBLM_R_X35Y128_SLICE_X52Y128_B = CLBLM_R_X35Y128_SLICE_X52Y128_BO6;
  assign CLBLM_R_X35Y128_SLICE_X52Y128_C = CLBLM_R_X35Y128_SLICE_X52Y128_CO6;
  assign CLBLM_R_X35Y128_SLICE_X52Y128_D = CLBLM_R_X35Y128_SLICE_X52Y128_DO6;
  assign CLBLM_R_X35Y128_SLICE_X52Y128_BMUX = CLBLM_R_X35Y128_SLICE_X52Y128_BO6;
  assign CLBLM_R_X35Y128_SLICE_X53Y128_COUT = CLBLM_R_X35Y128_SLICE_X53Y128_D_CY;
  assign CLBLM_R_X35Y128_SLICE_X53Y128_A = CLBLM_R_X35Y128_SLICE_X53Y128_AO6;
  assign CLBLM_R_X35Y128_SLICE_X53Y128_B = CLBLM_R_X35Y128_SLICE_X53Y128_BO6;
  assign CLBLM_R_X35Y128_SLICE_X53Y128_C = CLBLM_R_X35Y128_SLICE_X53Y128_CO6;
  assign CLBLM_R_X35Y128_SLICE_X53Y128_D = CLBLM_R_X35Y128_SLICE_X53Y128_DO6;
  assign CLBLM_R_X35Y128_SLICE_X53Y128_BMUX = CLBLM_R_X35Y128_SLICE_X53Y128_BO6;
  assign CLBLM_R_X35Y129_SLICE_X52Y129_COUT = CLBLM_R_X35Y129_SLICE_X52Y129_D_CY;
  assign CLBLM_R_X35Y129_SLICE_X52Y129_A = CLBLM_R_X35Y129_SLICE_X52Y129_AO6;
  assign CLBLM_R_X35Y129_SLICE_X52Y129_B = CLBLM_R_X35Y129_SLICE_X52Y129_BO6;
  assign CLBLM_R_X35Y129_SLICE_X52Y129_C = CLBLM_R_X35Y129_SLICE_X52Y129_CO6;
  assign CLBLM_R_X35Y129_SLICE_X52Y129_D = CLBLM_R_X35Y129_SLICE_X52Y129_DO6;
  assign CLBLM_R_X35Y129_SLICE_X53Y129_COUT = CLBLM_R_X35Y129_SLICE_X53Y129_D_CY;
  assign CLBLM_R_X35Y129_SLICE_X53Y129_A = CLBLM_R_X35Y129_SLICE_X53Y129_AO6;
  assign CLBLM_R_X35Y129_SLICE_X53Y129_B = CLBLM_R_X35Y129_SLICE_X53Y129_BO6;
  assign CLBLM_R_X35Y129_SLICE_X53Y129_C = CLBLM_R_X35Y129_SLICE_X53Y129_CO6;
  assign CLBLM_R_X35Y129_SLICE_X53Y129_D = CLBLM_R_X35Y129_SLICE_X53Y129_DO6;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_COUT = CLBLM_R_X37Y117_SLICE_X56Y117_D_CY;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_A = CLBLM_R_X37Y117_SLICE_X56Y117_AO6;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_B = CLBLM_R_X37Y117_SLICE_X56Y117_BO6;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_C = CLBLM_R_X37Y117_SLICE_X56Y117_CO6;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_D = CLBLM_R_X37Y117_SLICE_X56Y117_DO6;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_AMUX = CLBLM_R_X37Y117_SLICE_X56Y117_AO5;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_COUT = CLBLM_R_X37Y117_SLICE_X57Y117_D_CY;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_A = CLBLM_R_X37Y117_SLICE_X57Y117_AO6;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_B = CLBLM_R_X37Y117_SLICE_X57Y117_BO6;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_C = CLBLM_R_X37Y117_SLICE_X57Y117_CO6;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_D = CLBLM_R_X37Y117_SLICE_X57Y117_DO6;
  assign CLBLM_R_X37Y118_SLICE_X56Y118_COUT = CLBLM_R_X37Y118_SLICE_X56Y118_D_CY;
  assign CLBLM_R_X37Y118_SLICE_X56Y118_A = CLBLM_R_X37Y118_SLICE_X56Y118_AO6;
  assign CLBLM_R_X37Y118_SLICE_X56Y118_B = CLBLM_R_X37Y118_SLICE_X56Y118_BO6;
  assign CLBLM_R_X37Y118_SLICE_X56Y118_C = CLBLM_R_X37Y118_SLICE_X56Y118_CO6;
  assign CLBLM_R_X37Y118_SLICE_X56Y118_D = CLBLM_R_X37Y118_SLICE_X56Y118_DO6;
  assign CLBLM_R_X37Y118_SLICE_X57Y118_COUT = CLBLM_R_X37Y118_SLICE_X57Y118_D_CY;
  assign CLBLM_R_X37Y118_SLICE_X57Y118_A = CLBLM_R_X37Y118_SLICE_X57Y118_AO6;
  assign CLBLM_R_X37Y118_SLICE_X57Y118_B = CLBLM_R_X37Y118_SLICE_X57Y118_BO6;
  assign CLBLM_R_X37Y118_SLICE_X57Y118_C = CLBLM_R_X37Y118_SLICE_X57Y118_CO6;
  assign CLBLM_R_X37Y118_SLICE_X57Y118_D = CLBLM_R_X37Y118_SLICE_X57Y118_DO6;
  assign CLBLM_R_X37Y118_SLICE_X57Y118_AMUX = CLBLM_R_X37Y118_SLICE_X57Y118_AO5;
  assign CLBLM_R_X37Y118_SLICE_X57Y118_BMUX = CLBLM_R_X37Y118_SLICE_X57Y118_BO6;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_COUT = CLBLM_R_X37Y119_SLICE_X56Y119_D_CY;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_A = CLBLM_R_X37Y119_SLICE_X56Y119_AO6;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_B = CLBLM_R_X37Y119_SLICE_X56Y119_BO6;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_C = CLBLM_R_X37Y119_SLICE_X56Y119_CO6;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_D = CLBLM_R_X37Y119_SLICE_X56Y119_DO6;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_COUT = CLBLM_R_X37Y119_SLICE_X57Y119_D_CY;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_A = CLBLM_R_X37Y119_SLICE_X57Y119_AO6;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_B = CLBLM_R_X37Y119_SLICE_X57Y119_BO6;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_C = CLBLM_R_X37Y119_SLICE_X57Y119_CO6;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_D = CLBLM_R_X37Y119_SLICE_X57Y119_DO6;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_BMUX = CLBLM_R_X37Y119_SLICE_X57Y119_BO6;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_COUT = CLBLM_R_X37Y120_SLICE_X56Y120_D_CY;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_A = CLBLM_R_X37Y120_SLICE_X56Y120_AO6;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_B = CLBLM_R_X37Y120_SLICE_X56Y120_BO6;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_C = CLBLM_R_X37Y120_SLICE_X56Y120_CO6;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_D = CLBLM_R_X37Y120_SLICE_X56Y120_DO6;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_COUT = CLBLM_R_X37Y120_SLICE_X57Y120_D_CY;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_A = CLBLM_R_X37Y120_SLICE_X57Y120_AO6;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_B = CLBLM_R_X37Y120_SLICE_X57Y120_BO6;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_C = CLBLM_R_X37Y120_SLICE_X57Y120_CO6;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_D = CLBLM_R_X37Y120_SLICE_X57Y120_DO6;
  assign CLBLM_R_X37Y121_SLICE_X56Y121_COUT = CLBLM_R_X37Y121_SLICE_X56Y121_D_CY;
  assign CLBLM_R_X37Y121_SLICE_X56Y121_A = CLBLM_R_X37Y121_SLICE_X56Y121_AO6;
  assign CLBLM_R_X37Y121_SLICE_X56Y121_B = CLBLM_R_X37Y121_SLICE_X56Y121_BO6;
  assign CLBLM_R_X37Y121_SLICE_X56Y121_C = CLBLM_R_X37Y121_SLICE_X56Y121_CO6;
  assign CLBLM_R_X37Y121_SLICE_X56Y121_D = CLBLM_R_X37Y121_SLICE_X56Y121_DO6;
  assign CLBLM_R_X37Y121_SLICE_X57Y121_COUT = CLBLM_R_X37Y121_SLICE_X57Y121_D_CY;
  assign CLBLM_R_X37Y121_SLICE_X57Y121_A = CLBLM_R_X37Y121_SLICE_X57Y121_AO6;
  assign CLBLM_R_X37Y121_SLICE_X57Y121_B = CLBLM_R_X37Y121_SLICE_X57Y121_BO6;
  assign CLBLM_R_X37Y121_SLICE_X57Y121_C = CLBLM_R_X37Y121_SLICE_X57Y121_CO6;
  assign CLBLM_R_X37Y121_SLICE_X57Y121_D = CLBLM_R_X37Y121_SLICE_X57Y121_DO6;
  assign CLBLM_R_X37Y121_SLICE_X57Y121_BMUX = CLBLM_R_X37Y121_SLICE_X57Y121_BO6;
  assign CLBLM_R_X37Y121_SLICE_X57Y121_DMUX = CLBLM_R_X37Y121_SLICE_X57Y121_DO5;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_COUT = CLBLM_R_X37Y122_SLICE_X56Y122_D_CY;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_A = CLBLM_R_X37Y122_SLICE_X56Y122_AO6;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_B = CLBLM_R_X37Y122_SLICE_X56Y122_BO6;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_C = CLBLM_R_X37Y122_SLICE_X56Y122_CO6;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_D = CLBLM_R_X37Y122_SLICE_X56Y122_DO6;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_COUT = CLBLM_R_X37Y122_SLICE_X57Y122_D_CY;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_A = CLBLM_R_X37Y122_SLICE_X57Y122_AO6;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_B = CLBLM_R_X37Y122_SLICE_X57Y122_BO6;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_C = CLBLM_R_X37Y122_SLICE_X57Y122_CO6;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_D = CLBLM_R_X37Y122_SLICE_X57Y122_DO6;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_CMUX = CLBLM_R_X37Y122_SLICE_X57Y122_CO6;
  assign CLBLM_R_X37Y123_SLICE_X56Y123_COUT = CLBLM_R_X37Y123_SLICE_X56Y123_D_CY;
  assign CLBLM_R_X37Y123_SLICE_X56Y123_A = CLBLM_R_X37Y123_SLICE_X56Y123_AO6;
  assign CLBLM_R_X37Y123_SLICE_X56Y123_B = CLBLM_R_X37Y123_SLICE_X56Y123_BO6;
  assign CLBLM_R_X37Y123_SLICE_X56Y123_C = CLBLM_R_X37Y123_SLICE_X56Y123_CO6;
  assign CLBLM_R_X37Y123_SLICE_X56Y123_D = CLBLM_R_X37Y123_SLICE_X56Y123_DO6;
  assign CLBLM_R_X37Y123_SLICE_X56Y123_CMUX = CLBLM_R_X37Y123_SLICE_X56Y123_CO6;
  assign CLBLM_R_X37Y123_SLICE_X56Y123_DMUX = CLBLM_R_X37Y123_SLICE_X56Y123_DO6;
  assign CLBLM_R_X37Y123_SLICE_X57Y123_COUT = CLBLM_R_X37Y123_SLICE_X57Y123_D_CY;
  assign CLBLM_R_X37Y123_SLICE_X57Y123_A = CLBLM_R_X37Y123_SLICE_X57Y123_AO6;
  assign CLBLM_R_X37Y123_SLICE_X57Y123_B = CLBLM_R_X37Y123_SLICE_X57Y123_BO6;
  assign CLBLM_R_X37Y123_SLICE_X57Y123_C = CLBLM_R_X37Y123_SLICE_X57Y123_CO6;
  assign CLBLM_R_X37Y123_SLICE_X57Y123_D = CLBLM_R_X37Y123_SLICE_X57Y123_DO6;
  assign CLBLM_R_X37Y123_SLICE_X57Y123_BMUX = CLBLM_R_X37Y123_SLICE_X57Y123_BO6;
  assign CLBLM_R_X37Y123_SLICE_X57Y123_DMUX = CLBLM_R_X37Y123_SLICE_X57Y123_DO5;
  assign CLBLM_R_X37Y124_SLICE_X56Y124_COUT = CLBLM_R_X37Y124_SLICE_X56Y124_D_CY;
  assign CLBLM_R_X37Y124_SLICE_X56Y124_A = CLBLM_R_X37Y124_SLICE_X56Y124_AO6;
  assign CLBLM_R_X37Y124_SLICE_X56Y124_B = CLBLM_R_X37Y124_SLICE_X56Y124_BO6;
  assign CLBLM_R_X37Y124_SLICE_X56Y124_C = CLBLM_R_X37Y124_SLICE_X56Y124_CO6;
  assign CLBLM_R_X37Y124_SLICE_X56Y124_D = CLBLM_R_X37Y124_SLICE_X56Y124_DO6;
  assign CLBLM_R_X37Y124_SLICE_X56Y124_BMUX = CLBLM_R_X37Y124_SLICE_X56Y124_BO6;
  assign CLBLM_R_X37Y124_SLICE_X57Y124_COUT = CLBLM_R_X37Y124_SLICE_X57Y124_D_CY;
  assign CLBLM_R_X37Y124_SLICE_X57Y124_A = CLBLM_R_X37Y124_SLICE_X57Y124_AO6;
  assign CLBLM_R_X37Y124_SLICE_X57Y124_B = CLBLM_R_X37Y124_SLICE_X57Y124_BO6;
  assign CLBLM_R_X37Y124_SLICE_X57Y124_C = CLBLM_R_X37Y124_SLICE_X57Y124_CO6;
  assign CLBLM_R_X37Y124_SLICE_X57Y124_D = CLBLM_R_X37Y124_SLICE_X57Y124_DO6;
  assign CLBLM_R_X37Y125_SLICE_X56Y125_COUT = CLBLM_R_X37Y125_SLICE_X56Y125_D_CY;
  assign CLBLM_R_X37Y125_SLICE_X56Y125_A = CLBLM_R_X37Y125_SLICE_X56Y125_AO6;
  assign CLBLM_R_X37Y125_SLICE_X56Y125_B = CLBLM_R_X37Y125_SLICE_X56Y125_BO6;
  assign CLBLM_R_X37Y125_SLICE_X56Y125_C = CLBLM_R_X37Y125_SLICE_X56Y125_CO6;
  assign CLBLM_R_X37Y125_SLICE_X56Y125_D = CLBLM_R_X37Y125_SLICE_X56Y125_DO6;
  assign CLBLM_R_X37Y125_SLICE_X57Y125_COUT = CLBLM_R_X37Y125_SLICE_X57Y125_D_CY;
  assign CLBLM_R_X37Y125_SLICE_X57Y125_A = CLBLM_R_X37Y125_SLICE_X57Y125_AO6;
  assign CLBLM_R_X37Y125_SLICE_X57Y125_B = CLBLM_R_X37Y125_SLICE_X57Y125_BO6;
  assign CLBLM_R_X37Y125_SLICE_X57Y125_C = CLBLM_R_X37Y125_SLICE_X57Y125_CO6;
  assign CLBLM_R_X37Y125_SLICE_X57Y125_D = CLBLM_R_X37Y125_SLICE_X57Y125_DO6;
  assign CLBLM_R_X37Y126_SLICE_X56Y126_COUT = CLBLM_R_X37Y126_SLICE_X56Y126_D_CY;
  assign CLBLM_R_X37Y126_SLICE_X56Y126_A = CLBLM_R_X37Y126_SLICE_X56Y126_AO6;
  assign CLBLM_R_X37Y126_SLICE_X56Y126_B = CLBLM_R_X37Y126_SLICE_X56Y126_BO6;
  assign CLBLM_R_X37Y126_SLICE_X56Y126_C = CLBLM_R_X37Y126_SLICE_X56Y126_CO6;
  assign CLBLM_R_X37Y126_SLICE_X56Y126_D = CLBLM_R_X37Y126_SLICE_X56Y126_DO6;
  assign CLBLM_R_X37Y126_SLICE_X56Y126_AMUX = CLBLM_R_X37Y126_SLICE_X56Y126_AO5;
  assign CLBLM_R_X37Y126_SLICE_X57Y126_COUT = CLBLM_R_X37Y126_SLICE_X57Y126_D_CY;
  assign CLBLM_R_X37Y126_SLICE_X57Y126_A = CLBLM_R_X37Y126_SLICE_X57Y126_AO6;
  assign CLBLM_R_X37Y126_SLICE_X57Y126_B = CLBLM_R_X37Y126_SLICE_X57Y126_BO6;
  assign CLBLM_R_X37Y126_SLICE_X57Y126_C = CLBLM_R_X37Y126_SLICE_X57Y126_CO6;
  assign CLBLM_R_X37Y126_SLICE_X57Y126_D = CLBLM_R_X37Y126_SLICE_X57Y126_DO6;
  assign CLBLM_R_X37Y126_SLICE_X57Y126_CMUX = CLBLM_R_X37Y126_SLICE_X57Y126_CO6;
  assign CLBLM_R_X37Y127_SLICE_X56Y127_COUT = CLBLM_R_X37Y127_SLICE_X56Y127_D_CY;
  assign CLBLM_R_X37Y127_SLICE_X56Y127_A = CLBLM_R_X37Y127_SLICE_X56Y127_AO6;
  assign CLBLM_R_X37Y127_SLICE_X56Y127_B = CLBLM_R_X37Y127_SLICE_X56Y127_BO6;
  assign CLBLM_R_X37Y127_SLICE_X56Y127_C = CLBLM_R_X37Y127_SLICE_X56Y127_CO6;
  assign CLBLM_R_X37Y127_SLICE_X56Y127_D = CLBLM_R_X37Y127_SLICE_X56Y127_DO6;
  assign CLBLM_R_X37Y127_SLICE_X57Y127_COUT = CLBLM_R_X37Y127_SLICE_X57Y127_D_CY;
  assign CLBLM_R_X37Y127_SLICE_X57Y127_A = CLBLM_R_X37Y127_SLICE_X57Y127_AO6;
  assign CLBLM_R_X37Y127_SLICE_X57Y127_B = CLBLM_R_X37Y127_SLICE_X57Y127_BO6;
  assign CLBLM_R_X37Y127_SLICE_X57Y127_C = CLBLM_R_X37Y127_SLICE_X57Y127_CO6;
  assign CLBLM_R_X37Y127_SLICE_X57Y127_D = CLBLM_R_X37Y127_SLICE_X57Y127_DO6;
  assign CLBLM_R_X37Y128_SLICE_X56Y128_COUT = CLBLM_R_X37Y128_SLICE_X56Y128_D_CY;
  assign CLBLM_R_X37Y128_SLICE_X56Y128_A = CLBLM_R_X37Y128_SLICE_X56Y128_AO6;
  assign CLBLM_R_X37Y128_SLICE_X56Y128_B = CLBLM_R_X37Y128_SLICE_X56Y128_BO6;
  assign CLBLM_R_X37Y128_SLICE_X56Y128_C = CLBLM_R_X37Y128_SLICE_X56Y128_CO6;
  assign CLBLM_R_X37Y128_SLICE_X56Y128_D = CLBLM_R_X37Y128_SLICE_X56Y128_DO6;
  assign CLBLM_R_X37Y128_SLICE_X57Y128_COUT = CLBLM_R_X37Y128_SLICE_X57Y128_D_CY;
  assign CLBLM_R_X37Y128_SLICE_X57Y128_A = CLBLM_R_X37Y128_SLICE_X57Y128_AO6;
  assign CLBLM_R_X37Y128_SLICE_X57Y128_B = CLBLM_R_X37Y128_SLICE_X57Y128_BO6;
  assign CLBLM_R_X37Y128_SLICE_X57Y128_C = CLBLM_R_X37Y128_SLICE_X57Y128_CO6;
  assign CLBLM_R_X37Y128_SLICE_X57Y128_D = CLBLM_R_X37Y128_SLICE_X57Y128_DO6;
  assign LIOI3_X0Y65_OLOGIC_X0Y65_OQ = CLBLL_L_X34Y115_SLICE_X51Y115_AO6;
  assign LIOI3_X0Y65_OLOGIC_X0Y65_TQ = 1'b1;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_O = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_O = LIOB33_X0Y101_IOB_X0Y101_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_O = LIOB33_X0Y103_IOB_X0Y104_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_O = LIOB33_X0Y103_IOB_X0Y103_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_O = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_O = LIOB33_X0Y105_IOB_X0Y105_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y110_O = LIOB33_X0Y109_IOB_X0Y110_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_O = LIOB33_X0Y109_IOB_X0Y109_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_O = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y111_O = LIOB33_X0Y111_IOB_X0Y111_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y116_O = LIOB33_X0Y115_IOB_X0Y116_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y115_O = LIOB33_X0Y115_IOB_X0Y115_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y118_O = LIOB33_X0Y117_IOB_X0Y118_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y117_O = LIOB33_X0Y117_IOB_X0Y117_I;
  assign LIOI3_X0Y121_ILOGIC_X0Y122_O = LIOB33_X0Y121_IOB_X0Y122_I;
  assign LIOI3_X0Y121_ILOGIC_X0Y121_O = LIOB33_X0Y121_IOB_X0Y121_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y124_O = LIOB33_X0Y123_IOB_X0Y124_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y123_O = LIOB33_X0Y123_IOB_X0Y123_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y126_O = LIOB33_X0Y125_IOB_X0Y126_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y125_O = LIOB33_X0Y125_IOB_X0Y125_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y128_O = LIOB33_X0Y127_IOB_X0Y128_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y127_O = LIOB33_X0Y127_IOB_X0Y127_I;
  assign LIOI3_X0Y129_ILOGIC_X0Y130_O = LIOB33_X0Y129_IOB_X0Y130_I;
  assign LIOI3_X0Y129_ILOGIC_X0Y129_O = LIOB33_X0Y129_IOB_X0Y129_I;
  assign LIOI3_X0Y133_ILOGIC_X0Y134_O = LIOB33_X0Y133_IOB_X0Y134_I;
  assign LIOI3_X0Y133_ILOGIC_X0Y133_O = LIOB33_X0Y133_IOB_X0Y133_I;
  assign LIOI3_X0Y135_ILOGIC_X0Y136_O = LIOB33_X0Y135_IOB_X0Y136_I;
  assign LIOI3_X0Y135_ILOGIC_X0Y135_O = LIOB33_X0Y135_IOB_X0Y135_I;
  assign LIOI3_X0Y139_ILOGIC_X0Y140_O = LIOB33_X0Y139_IOB_X0Y140_I;
  assign LIOI3_X0Y139_ILOGIC_X0Y139_O = LIOB33_X0Y139_IOB_X0Y139_I;
  assign LIOI3_X0Y141_ILOGIC_X0Y142_O = LIOB33_X0Y141_IOB_X0Y142_I;
  assign LIOI3_X0Y141_ILOGIC_X0Y141_O = LIOB33_X0Y141_IOB_X0Y141_I;
  assign LIOI3_X0Y145_ILOGIC_X0Y146_O = LIOB33_X0Y145_IOB_X0Y146_I;
  assign LIOI3_X0Y145_ILOGIC_X0Y145_O = LIOB33_X0Y145_IOB_X0Y145_I;
  assign LIOI3_X0Y147_ILOGIC_X0Y148_O = LIOB33_X0Y147_IOB_X0Y148_I;
  assign LIOI3_X0Y147_ILOGIC_X0Y147_O = LIOB33_X0Y147_IOB_X0Y147_I;
  assign LIOI3_SING_X0Y100_ILOGIC_X0Y100_O = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOI3_SING_X0Y149_ILOGIC_X0Y149_O = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O = LIOB33_X0Y107_IOB_X0Y107_I;
  assign LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y120_O = LIOB33_X0Y119_IOB_X0Y120_I;
  assign LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y119_O = LIOB33_X0Y119_IOB_X0Y119_I;
  assign LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y132_O = LIOB33_X0Y131_IOB_X0Y132_I;
  assign LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y131_O = LIOB33_X0Y131_IOB_X0Y131_I;
  assign LIOI3_TBYTESRC_X0Y143_ILOGIC_X0Y144_O = LIOB33_X0Y143_IOB_X0Y144_I;
  assign LIOI3_TBYTESRC_X0Y143_ILOGIC_X0Y143_O = LIOB33_X0Y143_IOB_X0Y143_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_O = LIOB33_X0Y113_IOB_X0Y114_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_O = LIOB33_X0Y113_IOB_X0Y113_I;
  assign LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y138_O = LIOB33_X0Y137_IOB_X0Y138_I;
  assign LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_O = LIOB33_X0Y137_IOB_X0Y137_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_O = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign RIOI3_X105Y117_OLOGIC_X1Y118_OQ = CLBLM_R_X35Y117_SLICE_X53Y117_CO6;
  assign RIOI3_X105Y117_OLOGIC_X1Y118_TQ = 1'b1;
  assign RIOI3_X105Y121_OLOGIC_X1Y122_OQ = CLBLM_R_X35Y116_SLICE_X53Y116_BO6;
  assign RIOI3_X105Y121_OLOGIC_X1Y122_TQ = 1'b1;
  assign RIOI3_X105Y121_OLOGIC_X1Y121_OQ = CLBLM_R_X35Y115_SLICE_X52Y115_BO6;
  assign RIOI3_X105Y121_OLOGIC_X1Y121_TQ = 1'b1;
  assign RIOI3_X105Y123_OLOGIC_X1Y124_OQ = CLBLL_L_X34Y120_SLICE_X51Y120_AO6;
  assign RIOI3_X105Y123_OLOGIC_X1Y124_TQ = 1'b1;
  assign RIOI3_X105Y123_OLOGIC_X1Y123_OQ = CLBLL_L_X36Y119_SLICE_X55Y119_BO6;
  assign RIOI3_X105Y123_OLOGIC_X1Y123_TQ = 1'b1;
  assign RIOI3_X105Y125_OLOGIC_X1Y126_OQ = CLBLL_L_X34Y121_SLICE_X51Y121_AO6;
  assign RIOI3_X105Y125_OLOGIC_X1Y126_TQ = 1'b1;
  assign RIOI3_X105Y125_OLOGIC_X1Y125_OQ = CLBLM_R_X33Y121_SLICE_X48Y121_AO6;
  assign RIOI3_X105Y125_OLOGIC_X1Y125_TQ = 1'b1;
  assign RIOI3_X105Y127_OLOGIC_X1Y128_OQ = CLBLL_L_X36Y122_SLICE_X54Y122_BO6;
  assign RIOI3_X105Y127_OLOGIC_X1Y128_TQ = 1'b1;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_OQ = CLBLM_R_X33Y123_SLICE_X49Y123_AO6;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_TQ = 1'b1;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_OQ = CLBLM_R_X35Y119_SLICE_X53Y119_AO6;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_TQ = 1'b1;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_OQ = CLBLL_L_X34Y124_SLICE_X50Y124_AO6;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_TQ = 1'b1;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_OQ = CLBLM_R_X37Y122_SLICE_X57Y122_AO6;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_TQ = 1'b1;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_OQ = CLBLM_R_X37Y121_SLICE_X57Y121_AO6;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_TQ = 1'b1;
  assign RIOI3_X105Y135_OLOGIC_X1Y136_OQ = CLBLM_R_X37Y123_SLICE_X57Y123_AO6;
  assign RIOI3_X105Y135_OLOGIC_X1Y136_TQ = 1'b1;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_OQ = CLBLM_R_X37Y123_SLICE_X56Y123_AO6;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_TQ = 1'b1;
  assign RIOI3_X105Y139_OLOGIC_X1Y140_OQ = CLBLL_L_X38Y126_SLICE_X58Y126_AO6;
  assign RIOI3_X105Y139_OLOGIC_X1Y140_TQ = 1'b1;
  assign RIOI3_X105Y139_OLOGIC_X1Y139_OQ = CLBLM_R_X37Y125_SLICE_X57Y125_AO6;
  assign RIOI3_X105Y139_OLOGIC_X1Y139_TQ = 1'b1;
  assign RIOI3_X105Y141_OLOGIC_X1Y142_OQ = CLBLL_L_X36Y127_SLICE_X54Y127_BO6;
  assign RIOI3_X105Y141_OLOGIC_X1Y142_TQ = 1'b1;
  assign RIOI3_X105Y141_OLOGIC_X1Y141_OQ = CLBLL_L_X36Y127_SLICE_X54Y127_AO6;
  assign RIOI3_X105Y141_OLOGIC_X1Y141_TQ = 1'b1;
  assign RIOI3_X105Y145_OLOGIC_X1Y146_OQ = CLBLL_L_X36Y128_SLICE_X54Y128_AO6;
  assign RIOI3_X105Y145_OLOGIC_X1Y146_TQ = 1'b1;
  assign RIOI3_X105Y145_OLOGIC_X1Y145_OQ = CLBLL_L_X36Y129_SLICE_X54Y129_AO6;
  assign RIOI3_X105Y145_OLOGIC_X1Y145_TQ = 1'b1;
  assign RIOI3_X105Y147_OLOGIC_X1Y148_OQ = CLBLL_L_X36Y129_SLICE_X55Y129_DO6;
  assign RIOI3_X105Y147_OLOGIC_X1Y148_TQ = 1'b1;
  assign RIOI3_X105Y147_OLOGIC_X1Y147_OQ = CLBLM_R_X37Y126_SLICE_X56Y126_BO6;
  assign RIOI3_X105Y147_OLOGIC_X1Y147_TQ = 1'b1;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_SING_X105Y149_OLOGIC_X1Y149_OQ = CLBLL_L_X38Y126_SLICE_X59Y126_AO6;
  assign RIOI3_SING_X105Y149_OLOGIC_X1Y149_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_OQ = CLBLM_R_X35Y115_SLICE_X53Y115_AO6;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_OQ = CLBLM_R_X33Y116_SLICE_X49Y116_AO6;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_OQ = CLBLL_L_X36Y122_SLICE_X55Y122_BO6;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_OQ = CLBLL_L_X36Y121_SLICE_X55Y121_BO6;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_OQ = CLBLL_L_X36Y129_SLICE_X55Y129_AO6;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_OQ = CLBLM_R_X35Y126_SLICE_X52Y126_BO6;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O = RIOB33_X105Y113_IOB_X1Y114_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_OQ = CLBLM_R_X37Y123_SLICE_X56Y123_BO6;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_OQ = CLBLM_R_X37Y125_SLICE_X56Y125_AO6;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_TQ = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_C1 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_C2 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_C3 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_C4 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_C5 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_C6 = 1'b1;
  assign RIOB33_X105Y137_IOB_X1Y137_O = CLBLM_R_X37Y125_SLICE_X56Y125_AO6;
  assign CLBLM_R_X35Y124_SLICE_X53Y124_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X34Y125_SLICE_X51Y125_A1 = 1'b1;
  assign CLBLL_L_X34Y125_SLICE_X51Y125_A2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X34Y125_SLICE_X51Y125_A3 = LIOB33_X0Y129_IOB_X0Y130_I;
  assign CLBLL_L_X34Y125_SLICE_X51Y125_A4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X34Y125_SLICE_X51Y125_A5 = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLL_L_X34Y125_SLICE_X51Y125_A6 = 1'b1;
  assign CLBLM_R_X35Y129_SLICE_X53Y129_C6 = LIOB33_X0Y145_IOB_X0Y145_I;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_D1 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_D2 = 1'b1;
  assign CLBLL_L_X34Y125_SLICE_X51Y125_B1 = LIOB33_X0Y133_IOB_X0Y133_I;
  assign CLBLL_L_X34Y125_SLICE_X51Y125_B2 = LIOB33_X0Y131_IOB_X0Y132_I;
  assign CLBLL_L_X34Y125_SLICE_X51Y125_B3 = 1'b1;
  assign CLBLL_L_X34Y125_SLICE_X51Y125_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X34Y125_SLICE_X51Y125_B5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X34Y125_SLICE_X51Y125_B6 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_D5 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_D6 = 1'b1;
  assign CLBLL_L_X34Y125_SLICE_X51Y125_C1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X34Y125_SLICE_X51Y125_C2 = 1'b1;
  assign CLBLL_L_X34Y125_SLICE_X51Y125_C3 = LIOB33_X0Y135_IOB_X0Y135_I;
  assign CLBLL_L_X34Y125_SLICE_X51Y125_C4 = LIOB33_X0Y133_IOB_X0Y134_I;
  assign CLBLL_L_X34Y125_SLICE_X51Y125_C5 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X34Y125_SLICE_X51Y125_C6 = 1'b1;
  assign LIOI3_X0Y139_ILOGIC_X0Y139_D = LIOB33_X0Y139_IOB_X0Y139_I;
  assign CLBLL_L_X34Y125_SLICE_X51Y125_CIN = CLBLL_L_X34Y124_SLICE_X51Y124_D_CY;
  assign CLBLM_R_X33Y125_SLICE_X49Y125_D6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X34Y125_SLICE_X51Y125_D1 = LIOB33_X0Y137_IOB_X0Y137_I;
  assign CLBLL_L_X34Y125_SLICE_X51Y125_D2 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X34Y125_SLICE_X51Y125_D3 = LIOB33_X0Y135_IOB_X0Y136_I;
  assign CLBLL_L_X34Y125_SLICE_X51Y125_D4 = 1'b1;
  assign CLBLL_L_X34Y125_SLICE_X51Y125_D5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X34Y125_SLICE_X51Y125_D6 = 1'b1;
  assign CLBLL_L_X38Y119_SLICE_X58Y119_A1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X38Y119_SLICE_X58Y119_A2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X38Y119_SLICE_X58Y119_A3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X38Y119_SLICE_X58Y119_A4 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X38Y119_SLICE_X58Y119_A5 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X38Y119_SLICE_X58Y119_A6 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X38Y119_SLICE_X58Y119_B1 = 1'b1;
  assign CLBLL_L_X38Y119_SLICE_X58Y119_B2 = 1'b1;
  assign CLBLL_L_X38Y119_SLICE_X58Y119_B3 = 1'b1;
  assign CLBLL_L_X38Y119_SLICE_X58Y119_B4 = 1'b1;
  assign CLBLL_L_X38Y119_SLICE_X58Y119_B5 = 1'b1;
  assign CLBLL_L_X38Y119_SLICE_X58Y119_B6 = 1'b1;
  assign CLBLL_L_X38Y119_SLICE_X58Y119_C1 = 1'b1;
  assign CLBLL_L_X38Y119_SLICE_X58Y119_C2 = 1'b1;
  assign CLBLL_L_X38Y119_SLICE_X58Y119_C3 = 1'b1;
  assign CLBLL_L_X38Y119_SLICE_X58Y119_C4 = 1'b1;
  assign CLBLL_L_X38Y119_SLICE_X58Y119_C5 = 1'b1;
  assign CLBLL_L_X38Y119_SLICE_X58Y119_C6 = 1'b1;
  assign RIOI3_X105Y139_OLOGIC_X1Y140_D1 = CLBLL_L_X38Y126_SLICE_X58Y126_AO6;
  assign CLBLL_L_X38Y119_SLICE_X58Y119_D1 = 1'b1;
  assign CLBLL_L_X38Y119_SLICE_X58Y119_D2 = 1'b1;
  assign CLBLL_L_X38Y119_SLICE_X58Y119_D3 = 1'b1;
  assign CLBLL_L_X38Y119_SLICE_X58Y119_D4 = 1'b1;
  assign CLBLL_L_X38Y119_SLICE_X58Y119_D5 = 1'b1;
  assign CLBLL_L_X38Y119_SLICE_X58Y119_D6 = 1'b1;
  assign RIOI3_X105Y139_OLOGIC_X1Y140_T1 = 1'b1;
  assign LIOI3_X0Y65_OLOGIC_X0Y65_D1 = CLBLL_L_X34Y115_SLICE_X51Y115_AO6;
  assign RIOI3_X105Y139_OLOGIC_X1Y139_D1 = CLBLM_R_X37Y125_SLICE_X57Y125_AO6;
  assign LIOI3_X0Y65_OLOGIC_X0Y65_T1 = 1'b1;
  assign RIOI3_X105Y139_OLOGIC_X1Y139_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_D1 = CLBLM_R_X37Y123_SLICE_X56Y123_BO6;
  assign CLBLL_L_X38Y119_SLICE_X59Y119_A1 = 1'b1;
  assign CLBLL_L_X38Y119_SLICE_X59Y119_A2 = 1'b1;
  assign CLBLL_L_X38Y119_SLICE_X59Y119_A3 = 1'b1;
  assign CLBLL_L_X38Y119_SLICE_X59Y119_A4 = 1'b1;
  assign CLBLL_L_X38Y119_SLICE_X59Y119_A5 = 1'b1;
  assign CLBLL_L_X38Y119_SLICE_X59Y119_A6 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_T1 = 1'b1;
  assign CLBLL_L_X38Y119_SLICE_X59Y119_B1 = 1'b1;
  assign CLBLL_L_X38Y119_SLICE_X59Y119_B2 = 1'b1;
  assign CLBLL_L_X38Y119_SLICE_X59Y119_B3 = 1'b1;
  assign CLBLL_L_X38Y119_SLICE_X59Y119_B4 = 1'b1;
  assign CLBLL_L_X38Y119_SLICE_X59Y119_B5 = 1'b1;
  assign CLBLL_L_X38Y119_SLICE_X59Y119_B6 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_D1 = CLBLM_R_X37Y125_SLICE_X56Y125_AO6;
  assign CLBLL_L_X38Y119_SLICE_X59Y119_C1 = 1'b1;
  assign CLBLL_L_X38Y119_SLICE_X59Y119_C2 = 1'b1;
  assign CLBLL_L_X38Y119_SLICE_X59Y119_C3 = 1'b1;
  assign CLBLL_L_X38Y119_SLICE_X59Y119_C4 = 1'b1;
  assign CLBLL_L_X38Y119_SLICE_X59Y119_C5 = 1'b1;
  assign CLBLL_L_X38Y119_SLICE_X59Y119_C6 = 1'b1;
  assign CLBLM_R_X35Y128_SLICE_X53Y128_C2 = LIOB33_X0Y143_IOB_X0Y144_I;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_T1 = 1'b1;
  assign CLBLL_L_X38Y119_SLICE_X59Y119_D1 = 1'b1;
  assign CLBLL_L_X38Y119_SLICE_X59Y119_D2 = 1'b1;
  assign CLBLL_L_X38Y119_SLICE_X59Y119_D3 = 1'b1;
  assign CLBLL_L_X38Y119_SLICE_X59Y119_D4 = 1'b1;
  assign CLBLL_L_X38Y119_SLICE_X59Y119_D5 = 1'b1;
  assign CLBLL_L_X38Y119_SLICE_X59Y119_D6 = 1'b1;
  assign CLBLL_L_X36Y123_SLICE_X55Y123_B1 = CLBLL_L_X36Y116_SLICE_X54Y116_DO6;
  assign CLBLL_L_X36Y123_SLICE_X55Y123_B2 = CLBLM_R_X37Y119_SLICE_X57Y119_DO6;
  assign CLBLM_R_X35Y128_SLICE_X53Y128_C3 = 1'b1;
  assign CLBLL_L_X36Y123_SLICE_X55Y123_B3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X36Y123_SLICE_X55Y123_B4 = CLBLM_R_X33Y123_SLICE_X48Y123_CO6;
  assign CLBLL_L_X36Y123_SLICE_X55Y123_B5 = CLBLM_R_X33Y122_SLICE_X48Y122_BO6;
  assign CLBLL_L_X36Y123_SLICE_X55Y123_B6 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X35Y128_SLICE_X53Y128_C4 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X37Y118_SLICE_X57Y118_A1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X37Y118_SLICE_X57Y118_A2 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X37Y118_SLICE_X57Y118_A3 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X37Y118_SLICE_X57Y118_A4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X37Y118_SLICE_X57Y118_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X37Y118_SLICE_X57Y118_A6 = 1'b1;
  assign RIOB33_X105Y117_IOB_X1Y118_O = CLBLM_R_X35Y117_SLICE_X53Y117_CO6;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_A1 = CLBLL_L_X34Y123_SLICE_X50Y123_BO5;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_A2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_A3 = CLBLM_R_X33Y125_SLICE_X49Y125_BO5;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_A4 = CLBLM_R_X33Y122_SLICE_X48Y122_AO5;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_A5 = CLBLL_L_X34Y125_SLICE_X50Y125_BO6;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_A6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X35Y128_SLICE_X53Y128_C5 = 1'b1;
  assign CLBLM_R_X37Y118_SLICE_X57Y118_B1 = CLBLL_L_X36Y117_SLICE_X55Y117_AO5;
  assign CLBLM_R_X37Y118_SLICE_X57Y118_B2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_B1 = CLBLL_L_X34Y123_SLICE_X50Y123_BO5;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_B2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_B3 = CLBLM_R_X33Y125_SLICE_X49Y125_BO5;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_B4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_B5 = CLBLL_L_X34Y125_SLICE_X50Y125_BO6;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_B6 = CLBLM_R_X33Y125_SLICE_X49Y125_CO6;
  assign CLBLM_R_X37Y118_SLICE_X57Y118_B6 = CLBLM_R_X37Y118_SLICE_X57Y118_AO5;
  assign CLBLM_R_X37Y118_SLICE_X57Y118_C1 = CLBLL_L_X38Y118_SLICE_X58Y118_AO6;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_C1 = CLBLM_R_X33Y124_SLICE_X49Y124_DO6;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_C2 = CLBLL_L_X34Y123_SLICE_X50Y123_AO5;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_C3 = CLBLM_R_X33Y125_SLICE_X49Y125_DO6;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_C4 = CLBLL_L_X34Y125_SLICE_X50Y125_DO6;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_C5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_C6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X37Y118_SLICE_X57Y118_C6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X37Y118_SLICE_X57Y118_D1 = CLBLL_L_X38Y118_SLICE_X58Y118_AO6;
  assign CLBLM_R_X37Y118_SLICE_X57Y118_D2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X35Y128_SLICE_X53Y128_C6 = 1'b1;
  assign CLBLM_R_X37Y118_SLICE_X57Y118_D3 = CLBLL_L_X36Y117_SLICE_X55Y117_AO5;
  assign CLBLM_R_X37Y118_SLICE_X57Y118_D4 = CLBLL_L_X36Y116_SLICE_X54Y116_AO5;
  assign CLBLM_R_X33Y125_SLICE_X48Y125_D3 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_D1 = CLBLM_R_X33Y124_SLICE_X49Y124_DO6;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_D2 = CLBLL_L_X34Y122_SLICE_X51Y122_CO6;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_D3 = CLBLM_R_X33Y125_SLICE_X49Y125_DO6;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_D4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_D5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X34Y126_SLICE_X50Y126_D6 = CLBLL_L_X34Y125_SLICE_X50Y125_DO6;
  assign CLBLM_R_X33Y125_SLICE_X48Y125_D4 = 1'b1;
  assign CLBLM_R_X37Y118_SLICE_X56Y118_A1 = CLBLM_R_X37Y118_SLICE_X56Y118_DO6;
  assign CLBLM_R_X33Y125_SLICE_X48Y125_D5 = 1'b1;
  assign CLBLM_R_X37Y118_SLICE_X56Y118_A2 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_R_X37Y118_SLICE_X56Y118_A3 = CLBLL_L_X34Y128_SLICE_X50Y128_AO6;
  assign CLBLM_R_X37Y118_SLICE_X56Y118_A4 = CLBLL_L_X36Y118_SLICE_X54Y118_CO6;
  assign CLBLM_R_X37Y118_SLICE_X56Y118_A5 = CLBLM_R_X35Y124_SLICE_X53Y124_A_XOR;
  assign CLBLM_R_X33Y125_SLICE_X48Y125_D6 = 1'b1;
  assign CLBLM_R_X37Y118_SLICE_X56Y118_A6 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLM_R_X37Y118_SLICE_X56Y118_B1 = CLBLL_L_X36Y117_SLICE_X55Y117_BO5;
  assign CLBLM_R_X37Y118_SLICE_X56Y118_B2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X37Y118_SLICE_X56Y118_B3 = CLBLM_R_X37Y117_SLICE_X56Y117_AO6;
  assign CLBLM_R_X37Y118_SLICE_X56Y118_B4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X37Y118_SLICE_X56Y118_B5 = CLBLM_R_X35Y118_SLICE_X53Y118_AO6;
  assign CLBLM_R_X37Y118_SLICE_X56Y118_B6 = CLBLL_L_X36Y118_SLICE_X55Y118_AO5;
  assign CLBLM_R_X37Y118_SLICE_X56Y118_C1 = CLBLM_R_X37Y117_SLICE_X56Y117_AO6;
  assign CLBLM_R_X37Y118_SLICE_X56Y118_C2 = CLBLL_L_X36Y117_SLICE_X55Y117_BO5;
  assign CLBLM_R_X37Y118_SLICE_X56Y118_C3 = CLBLL_L_X38Y118_SLICE_X58Y118_AO5;
  assign CLBLM_R_X37Y118_SLICE_X56Y118_C4 = CLBLL_L_X36Y118_SLICE_X55Y118_AO5;
  assign CLBLM_R_X37Y118_SLICE_X56Y118_C5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X37Y118_SLICE_X56Y118_C6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_A1 = LIOB33_X0Y137_IOB_X0Y138_I;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_A2 = LIOB33_X0Y139_IOB_X0Y139_I;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_A3 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_A4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_A5 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_A6 = 1'b1;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_D = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X37Y118_SLICE_X56Y118_D1 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X37Y118_SLICE_X56Y118_D2 = CLBLM_R_X35Y124_SLICE_X53Y124_A_XOR;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_B1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_B2 = LIOB33_X0Y139_IOB_X0Y140_I;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_B3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_B4 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_B5 = LIOB33_X0Y141_IOB_X0Y141_I;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_B6 = 1'b1;
  assign CLBLM_R_X37Y118_SLICE_X56Y118_D3 = CLBLM_R_X37Y118_SLICE_X57Y118_BO6;
  assign CLBLM_R_X37Y118_SLICE_X56Y118_D4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X37Y118_SLICE_X56Y118_D5 = 1'b1;
  assign CLBLM_R_X37Y118_SLICE_X56Y118_D6 = CLBLM_R_X37Y118_SLICE_X56Y118_BO6;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_C1 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_C2 = LIOB33_X0Y143_IOB_X0Y143_I;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_C3 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_C4 = LIOB33_X0Y141_IOB_X0Y142_I;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_C5 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_C6 = 1'b1;
  assign CLBLM_R_X35Y125_SLICE_X53Y125_CX = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_CIN = CLBLL_L_X34Y125_SLICE_X51Y125_D_CY;
  assign LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y119_D = LIOB33_X0Y119_IOB_X0Y119_I;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_D1 = LIOB33_X0Y143_IOB_X0Y144_I;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_D2 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_D3 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_D4 = LIOB33_X0Y145_IOB_X0Y145_I;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_D5 = 1'b1;
  assign CLBLL_L_X34Y126_SLICE_X51Y126_D6 = 1'b1;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_D = RIOB33_X105Y109_IOB_X1Y109_I;
  assign LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y120_D = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLM_R_X35Y127_SLICE_X53Y127_A3 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X35Y127_SLICE_X53Y127_A4 = 1'b1;
  assign CLBLM_R_X35Y127_SLICE_X53Y127_A5 = 1'b1;
  assign CLBLM_R_X35Y127_SLICE_X53Y127_A6 = LIOB33_X0Y141_IOB_X0Y142_I;
  assign RIOB33_X105Y119_IOB_X1Y120_O = CLBLM_R_X35Y115_SLICE_X53Y115_AO6;
  assign RIOB33_X105Y119_IOB_X1Y119_O = CLBLM_R_X33Y116_SLICE_X49Y116_AO6;
  assign CLBLM_R_X35Y127_SLICE_X53Y127_AX = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X35Y127_SLICE_X53Y127_B3 = 1'b1;
  assign CLBLM_R_X33Y115_SLICE_X49Y115_D2 = CLBLM_R_X35Y121_SLICE_X53Y121_A_XOR;
  assign CLBLM_R_X35Y127_SLICE_X53Y127_B4 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_A1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X34Y127_SLICE_X50Y127_A1 = CLBLL_L_X34Y123_SLICE_X50Y123_BO5;
  assign CLBLL_L_X34Y127_SLICE_X50Y127_A2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X34Y127_SLICE_X50Y127_A3 = CLBLL_L_X34Y125_SLICE_X50Y125_BO6;
  assign CLBLL_L_X34Y127_SLICE_X50Y127_A4 = CLBLM_R_X33Y125_SLICE_X49Y125_CO6;
  assign CLBLL_L_X34Y127_SLICE_X50Y127_A5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X34Y127_SLICE_X50Y127_A6 = CLBLL_L_X34Y125_SLICE_X50Y125_CO6;
  assign CLBLM_R_X35Y127_SLICE_X53Y127_B5 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X35Y127_SLICE_X53Y127_B6 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_A4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X34Y127_SLICE_X50Y127_B1 = CLBLL_L_X34Y125_SLICE_X50Y125_CO6;
  assign CLBLL_L_X34Y127_SLICE_X50Y127_B2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X34Y127_SLICE_X50Y127_B3 = CLBLL_L_X34Y125_SLICE_X50Y125_BO6;
  assign CLBLL_L_X34Y127_SLICE_X50Y127_B4 = CLBLM_R_X33Y125_SLICE_X49Y125_CO6;
  assign CLBLL_L_X34Y127_SLICE_X50Y127_B5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X34Y127_SLICE_X50Y127_B6 = CLBLL_L_X34Y127_SLICE_X50Y127_CO6;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_B1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_B2 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_B4 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X34Y127_SLICE_X50Y127_C1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X34Y127_SLICE_X50Y127_C2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X34Y127_SLICE_X50Y127_C3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X34Y127_SLICE_X50Y127_C4 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X34Y127_SLICE_X50Y127_C5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X34Y127_SLICE_X50Y127_C6 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X35Y127_SLICE_X53Y127_BX = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_C2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_C3 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_C4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_C5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_C6 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X35Y127_SLICE_X53Y127_C1 = 1'b1;
  assign CLBLL_L_X34Y127_SLICE_X50Y127_D1 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X34Y127_SLICE_X50Y127_D2 = 1'b1;
  assign CLBLL_L_X34Y127_SLICE_X50Y127_D3 = 1'b1;
  assign CLBLL_L_X34Y127_SLICE_X50Y127_D4 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLL_L_X34Y127_SLICE_X50Y127_D5 = 1'b1;
  assign CLBLL_L_X34Y127_SLICE_X50Y127_D6 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_R_X35Y127_SLICE_X53Y127_C2 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X35Y127_SLICE_X53Y127_C3 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_D4 = CLBLM_R_X37Y119_SLICE_X57Y119_CO6;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_A1 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_A2 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLM_R_X35Y127_SLICE_X53Y127_C4 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_A3 = CLBLM_R_X35Y124_SLICE_X53Y124_B_XOR;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_A4 = CLBLL_L_X36Y119_SLICE_X54Y119_CO6;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_A5 = CLBLL_L_X34Y128_SLICE_X50Y128_AO6;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_A6 = CLBLM_R_X37Y119_SLICE_X56Y119_CO6;
  assign CLBLM_R_X35Y127_SLICE_X53Y127_C5 = 1'b1;
  assign RIOB33_X105Y137_IOB_X1Y138_O = CLBLM_R_X37Y123_SLICE_X56Y123_BO6;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_B1 = CLBLM_R_X35Y123_SLICE_X53Y123_D_XOR;
  assign CLBLM_R_X35Y127_SLICE_X53Y127_C6 = LIOB33_X0Y143_IOB_X0Y144_I;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_B2 = CLBLL_L_X36Y118_SLICE_X55Y118_BO6;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_B3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_B4 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_B5 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_B6 = CLBLM_R_X37Y118_SLICE_X57Y118_BO6;
  assign CLBLM_R_X35Y127_SLICE_X53Y127_CIN = CLBLM_R_X35Y126_SLICE_X53Y126_D_CY;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_C1 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_C2 = 1'b1;
  assign CLBLL_L_X34Y127_SLICE_X51Y127_A1 = 1'b1;
  assign CLBLL_L_X34Y127_SLICE_X51Y127_A2 = 1'b1;
  assign CLBLL_L_X34Y127_SLICE_X51Y127_A3 = 1'b1;
  assign CLBLL_L_X34Y127_SLICE_X51Y127_A4 = 1'b1;
  assign CLBLL_L_X34Y127_SLICE_X51Y127_A5 = 1'b1;
  assign CLBLL_L_X34Y127_SLICE_X51Y127_A6 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_C3 = CLBLM_R_X35Y124_SLICE_X53Y124_B_XOR;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_C4 = CLBLM_R_X37Y118_SLICE_X57Y118_CO6;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_C5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X34Y127_SLICE_X51Y127_B1 = 1'b1;
  assign CLBLL_L_X34Y127_SLICE_X51Y127_B2 = 1'b1;
  assign CLBLL_L_X34Y127_SLICE_X51Y127_B3 = 1'b1;
  assign CLBLL_L_X34Y127_SLICE_X51Y127_B4 = 1'b1;
  assign CLBLL_L_X34Y127_SLICE_X51Y127_B5 = 1'b1;
  assign CLBLL_L_X34Y127_SLICE_X51Y127_B6 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_D1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_D2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X34Y127_SLICE_X51Y127_C1 = 1'b1;
  assign CLBLL_L_X34Y127_SLICE_X51Y127_C2 = 1'b1;
  assign CLBLL_L_X34Y127_SLICE_X51Y127_C3 = 1'b1;
  assign CLBLL_L_X34Y127_SLICE_X51Y127_C4 = 1'b1;
  assign CLBLL_L_X34Y127_SLICE_X51Y127_C5 = 1'b1;
  assign CLBLL_L_X34Y127_SLICE_X51Y127_C6 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_D5 = 1'b1;
  assign CLBLM_R_X35Y127_SLICE_X53Y127_CX = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X34Y127_SLICE_X51Y127_D1 = 1'b1;
  assign CLBLL_L_X34Y127_SLICE_X51Y127_D2 = 1'b1;
  assign CLBLL_L_X34Y127_SLICE_X51Y127_D3 = 1'b1;
  assign CLBLL_L_X34Y127_SLICE_X51Y127_D4 = 1'b1;
  assign CLBLL_L_X34Y127_SLICE_X51Y127_D5 = 1'b1;
  assign CLBLL_L_X34Y127_SLICE_X51Y127_D6 = 1'b1;
  assign CLBLM_R_X35Y127_SLICE_X53Y127_D1 = 1'b1;
  assign CLBLM_R_X35Y127_SLICE_X53Y127_D2 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X37Y127_SLICE_X57Y127_A6 = 1'b1;
  assign CLBLM_R_X35Y127_SLICE_X53Y127_D3 = 1'b1;
  assign CLBLM_R_X35Y127_SLICE_X53Y127_D4 = 1'b1;
  assign CLBLM_R_X35Y127_SLICE_X53Y127_D5 = 1'b1;
  assign CLBLM_R_X35Y127_SLICE_X53Y127_D6 = LIOB33_X0Y145_IOB_X0Y145_I;
  assign CLBLM_R_X37Y127_SLICE_X57Y127_B1 = 1'b1;
  assign CLBLL_L_X38Y121_SLICE_X58Y121_A1 = CLBLL_L_X38Y121_SLICE_X58Y121_DO6;
  assign CLBLL_L_X38Y121_SLICE_X58Y121_A2 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLL_L_X38Y121_SLICE_X58Y121_A3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X38Y121_SLICE_X58Y121_A4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X38Y121_SLICE_X58Y121_A5 = CLBLL_L_X36Y121_SLICE_X54Y121_AO5;
  assign CLBLL_L_X38Y121_SLICE_X58Y121_A6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X35Y127_SLICE_X53Y127_DX = 1'b0;
  assign CLBLM_R_X37Y127_SLICE_X57Y127_B2 = 1'b1;
  assign CLBLM_R_X37Y127_SLICE_X57Y127_B3 = 1'b1;
  assign CLBLL_L_X38Y121_SLICE_X58Y121_B1 = LIOB33_X0Y127_IOB_X0Y128_I;
  assign CLBLL_L_X38Y121_SLICE_X58Y121_B2 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLL_L_X38Y121_SLICE_X58Y121_B3 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X38Y121_SLICE_X58Y121_B4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X38Y121_SLICE_X58Y121_B5 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLL_L_X38Y121_SLICE_X58Y121_B6 = CLBLL_L_X38Y121_SLICE_X58Y121_CO6;
  assign CLBLM_R_X37Y127_SLICE_X57Y127_B4 = 1'b1;
  assign CLBLM_R_X37Y127_SLICE_X57Y127_B5 = 1'b1;
  assign CLBLL_L_X38Y121_SLICE_X58Y121_C1 = CLBLM_R_X35Y123_SLICE_X53Y123_C_XOR;
  assign CLBLL_L_X38Y121_SLICE_X58Y121_C2 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLL_L_X38Y121_SLICE_X58Y121_C3 = CLBLM_R_X37Y121_SLICE_X57Y121_DO5;
  assign CLBLL_L_X38Y121_SLICE_X58Y121_C4 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X38Y121_SLICE_X58Y121_C5 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X38Y121_SLICE_X58Y121_C6 = CLBLM_R_X35Y121_SLICE_X52Y121_C_XOR;
  assign CLBLM_R_X37Y127_SLICE_X57Y127_B6 = 1'b1;
  assign CLBLM_R_X37Y128_SLICE_X56Y128_A3 = CLBLL_L_X36Y128_SLICE_X55Y128_BO6;
  assign CLBLL_L_X38Y121_SLICE_X58Y121_D1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X38Y121_SLICE_X58Y121_D2 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X38Y121_SLICE_X58Y121_D3 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X38Y121_SLICE_X58Y121_D4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X38Y121_SLICE_X58Y121_D5 = 1'b1;
  assign CLBLL_L_X38Y121_SLICE_X58Y121_D6 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X35Y127_SLICE_X52Y127_A3 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLM_R_X35Y127_SLICE_X52Y127_A4 = CLBLM_R_X35Y127_SLICE_X52Y127_BO6;
  assign CLBLM_R_X35Y127_SLICE_X52Y127_A5 = LIOB33_X0Y143_IOB_X0Y143_I;
  assign CLBLM_R_X37Y127_SLICE_X57Y127_C2 = 1'b1;
  assign CLBLM_R_X35Y127_SLICE_X52Y127_A6 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLM_R_X37Y127_SLICE_X57Y127_C3 = 1'b1;
  assign CLBLM_R_X37Y127_SLICE_X57Y127_C4 = 1'b1;
  assign CLBLM_R_X37Y127_SLICE_X57Y127_C5 = 1'b1;
  assign CLBLL_L_X38Y121_SLICE_X59Y121_A1 = 1'b1;
  assign CLBLL_L_X38Y121_SLICE_X59Y121_A2 = 1'b1;
  assign CLBLL_L_X38Y121_SLICE_X59Y121_A3 = 1'b1;
  assign CLBLL_L_X38Y121_SLICE_X59Y121_A4 = 1'b1;
  assign CLBLL_L_X38Y121_SLICE_X59Y121_A5 = 1'b1;
  assign CLBLL_L_X38Y121_SLICE_X59Y121_A6 = 1'b1;
  assign CLBLM_R_X37Y127_SLICE_X57Y127_C6 = 1'b1;
  assign CLBLL_L_X38Y121_SLICE_X59Y121_B1 = 1'b1;
  assign CLBLL_L_X38Y121_SLICE_X59Y121_B2 = 1'b1;
  assign CLBLL_L_X38Y121_SLICE_X59Y121_B3 = 1'b1;
  assign CLBLL_L_X38Y121_SLICE_X59Y121_B4 = 1'b1;
  assign CLBLL_L_X38Y121_SLICE_X59Y121_B5 = 1'b1;
  assign CLBLL_L_X38Y121_SLICE_X59Y121_B6 = 1'b1;
  assign CLBLM_R_X35Y127_SLICE_X52Y127_B1 = CLBLM_R_X35Y125_SLICE_X52Y125_B_XOR;
  assign CLBLM_R_X35Y127_SLICE_X52Y127_B2 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X38Y121_SLICE_X59Y121_C1 = 1'b1;
  assign CLBLL_L_X38Y121_SLICE_X59Y121_C2 = 1'b1;
  assign CLBLL_L_X38Y121_SLICE_X59Y121_C3 = 1'b1;
  assign CLBLL_L_X38Y121_SLICE_X59Y121_C4 = 1'b1;
  assign CLBLL_L_X38Y121_SLICE_X59Y121_C5 = 1'b1;
  assign CLBLL_L_X38Y121_SLICE_X59Y121_C6 = 1'b1;
  assign CLBLM_R_X35Y127_SLICE_X52Y127_B3 = CLBLM_R_X35Y127_SLICE_X53Y127_B_XOR;
  assign CLBLM_R_X35Y127_SLICE_X52Y127_B4 = CLBLM_R_X35Y127_SLICE_X52Y127_DO6;
  assign CLBLM_R_X35Y127_SLICE_X52Y127_B5 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X38Y121_SLICE_X59Y121_D1 = 1'b1;
  assign CLBLL_L_X38Y121_SLICE_X59Y121_D2 = 1'b1;
  assign CLBLL_L_X38Y121_SLICE_X59Y121_D3 = 1'b1;
  assign CLBLL_L_X38Y121_SLICE_X59Y121_D4 = 1'b1;
  assign CLBLL_L_X38Y121_SLICE_X59Y121_D5 = 1'b1;
  assign CLBLL_L_X38Y121_SLICE_X59Y121_D6 = 1'b1;
  assign CLBLM_R_X35Y127_SLICE_X52Y127_B6 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign RIOB33_X105Y121_IOB_X1Y121_O = CLBLM_R_X35Y115_SLICE_X52Y115_BO6;
  assign RIOB33_X105Y121_IOB_X1Y122_O = CLBLM_R_X35Y116_SLICE_X53Y116_BO6;
  assign CLBLM_R_X37Y127_SLICE_X57Y127_D1 = 1'b1;
  assign CLBLM_R_X37Y127_SLICE_X57Y127_D2 = 1'b1;
  assign CLBLM_R_X37Y127_SLICE_X57Y127_D3 = 1'b1;
  assign CLBLM_R_X37Y127_SLICE_X57Y127_D4 = 1'b1;
  assign CLBLM_R_X35Y127_SLICE_X52Y127_C1 = CLBLL_L_X36Y125_SLICE_X55Y125_BO6;
  assign CLBLM_R_X37Y127_SLICE_X57Y127_D5 = 1'b1;
  assign CLBLM_R_X35Y127_SLICE_X52Y127_C2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X37Y127_SLICE_X57Y127_D6 = 1'b1;
  assign CLBLM_R_X35Y127_SLICE_X52Y127_C3 = CLBLL_L_X34Y127_SLICE_X50Y127_BO6;
  assign RIOI3_X105Y141_OLOGIC_X1Y142_D1 = CLBLL_L_X36Y127_SLICE_X54Y127_BO6;
  assign CLBLM_R_X35Y127_SLICE_X52Y127_C4 = CLBLL_L_X34Y126_SLICE_X50Y126_DO6;
  assign CLBLM_R_X35Y127_SLICE_X52Y127_C5 = CLBLL_L_X36Y116_SLICE_X54Y116_BO5;
  assign RIOI3_X105Y141_OLOGIC_X1Y142_T1 = 1'b1;
  assign CLBLM_R_X35Y127_SLICE_X52Y127_C6 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_A1 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_A2 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_A3 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_A4 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_A5 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_A6 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_A1 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_A2 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_A3 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_B1 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_B2 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_B3 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_B4 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_B5 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_B6 = 1'b1;
  assign CLBLM_R_X35Y114_SLICE_X53Y114_A1 = 1'b1;
  assign CLBLM_R_X35Y114_SLICE_X53Y114_A2 = 1'b1;
  assign CLBLM_R_X35Y114_SLICE_X53Y114_A3 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_C1 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_C2 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_C3 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_C4 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_C5 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_C6 = 1'b1;
  assign CLBLM_R_X35Y114_SLICE_X53Y114_B1 = 1'b1;
  assign CLBLM_R_X35Y114_SLICE_X53Y114_B2 = 1'b1;
  assign CLBLM_R_X35Y114_SLICE_X53Y114_B3 = 1'b1;
  assign CLBLM_R_X35Y114_SLICE_X53Y114_B4 = 1'b1;
  assign CLBLM_R_X35Y114_SLICE_X53Y114_B5 = 1'b1;
  assign CLBLM_R_X35Y114_SLICE_X53Y114_B6 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_D1 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_D2 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_D3 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_D4 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_D5 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X50Y128_D6 = 1'b1;
  assign CLBLM_R_X35Y114_SLICE_X53Y114_C1 = 1'b1;
  assign CLBLM_R_X35Y114_SLICE_X53Y114_C2 = 1'b1;
  assign CLBLM_R_X35Y114_SLICE_X53Y114_C3 = 1'b1;
  assign CLBLM_R_X35Y114_SLICE_X53Y114_C4 = 1'b1;
  assign CLBLM_R_X35Y114_SLICE_X53Y114_C5 = 1'b1;
  assign CLBLM_R_X35Y114_SLICE_X53Y114_C6 = 1'b1;
  assign CLBLM_R_X35Y114_SLICE_X53Y114_D1 = 1'b1;
  assign CLBLM_R_X35Y114_SLICE_X53Y114_D2 = 1'b1;
  assign CLBLM_R_X35Y114_SLICE_X53Y114_D3 = 1'b1;
  assign CLBLM_R_X35Y114_SLICE_X53Y114_D4 = 1'b1;
  assign CLBLM_R_X35Y114_SLICE_X53Y114_D5 = 1'b1;
  assign CLBLM_R_X35Y114_SLICE_X53Y114_D6 = 1'b1;
  assign CLBLM_R_X35Y127_SLICE_X52Y127_D1 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_A1 = CLBLL_L_X36Y120_SLICE_X54Y120_CO6;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_A2 = CLBLL_L_X34Y128_SLICE_X50Y128_AO6;
  assign CLBLM_R_X35Y127_SLICE_X52Y127_D2 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_A3 = CLBLM_R_X35Y124_SLICE_X53Y124_C_XOR;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_A4 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLM_R_X35Y114_SLICE_X52Y114_A1 = LIOB33_X0Y119_IOB_X0Y119_I;
  assign CLBLM_R_X35Y114_SLICE_X52Y114_A2 = 1'b1;
  assign CLBLM_R_X35Y114_SLICE_X52Y114_A3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X35Y114_SLICE_X52Y114_A4 = 1'b1;
  assign CLBLM_R_X35Y114_SLICE_X52Y114_A5 = 1'b1;
  assign CLBLM_R_X35Y114_SLICE_X52Y114_A6 = 1'b1;
  assign CLBLM_R_X35Y127_SLICE_X52Y127_D3 = 1'b1;
  assign CLBLM_R_X35Y127_SLICE_X52Y127_D4 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_A1 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_A2 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_A3 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_A4 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_A5 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_A6 = 1'b1;
  assign CLBLM_R_X35Y114_SLICE_X52Y114_B1 = 1'b1;
  assign CLBLM_R_X35Y114_SLICE_X52Y114_B2 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_B1 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_B2 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_B3 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_B4 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_B5 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_B6 = 1'b1;
  assign CLBLM_R_X35Y114_SLICE_X52Y114_B5 = 1'b1;
  assign CLBLM_R_X35Y114_SLICE_X52Y114_B6 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_C1 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_C2 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_C3 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_C4 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_C5 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_C6 = 1'b1;
  assign CLBLM_R_X35Y114_SLICE_X52Y114_C4 = 1'b1;
  assign CLBLM_R_X35Y114_SLICE_X52Y114_C5 = 1'b1;
  assign CLBLM_R_X35Y114_SLICE_X52Y114_C6 = 1'b1;
  assign CLBLM_R_X35Y114_SLICE_X52Y114_D1 = 1'b1;
  assign CLBLM_R_X35Y114_SLICE_X52Y114_D2 = 1'b1;
  assign CLBLM_R_X35Y114_SLICE_X52Y114_D3 = 1'b1;
  assign CLBLM_R_X35Y114_SLICE_X52Y114_D4 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_D1 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_D2 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_D3 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_D4 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_D5 = 1'b1;
  assign CLBLL_L_X34Y128_SLICE_X51Y128_D6 = 1'b1;
  assign CLBLM_R_X35Y114_SLICE_X52Y114_D5 = 1'b1;
  assign CLBLM_R_X35Y114_SLICE_X52Y114_D6 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_B3 = CLBLL_L_X36Y122_SLICE_X55Y122_AO6;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_B4 = CLBLM_R_X35Y124_SLICE_X53Y124_D_XOR;
  assign CLBLM_R_X37Y123_SLICE_X56Y123_B6 = CLBLL_L_X36Y123_SLICE_X55Y123_AO6;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_B5 = CLBLM_R_X37Y122_SLICE_X57Y122_CO6;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_B6 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign RIOI3_SING_X105Y149_OLOGIC_X1Y149_D1 = CLBLL_L_X38Y126_SLICE_X59Y126_AO6;
  assign CLBLM_R_X37Y127_SLICE_X56Y127_C1 = CLBLM_R_X35Y127_SLICE_X53Y127_C_XOR;
  assign CLBLM_R_X37Y127_SLICE_X56Y127_C2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X37Y127_SLICE_X56Y127_C3 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X37Y127_SLICE_X56Y127_C4 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_C1 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_R_X37Y127_SLICE_X56Y127_C5 = CLBLL_L_X36Y116_SLICE_X55Y116_AO6;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_C2 = CLBLM_R_X35Y124_SLICE_X53Y124_D_XOR;
  assign CLBLM_R_X37Y127_SLICE_X56Y127_C6 = CLBLM_R_X37Y127_SLICE_X56Y127_BO6;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_C3 = LIOB33_X0Y133_IOB_X0Y133_I;
  assign CLBLM_R_X35Y125_SLICE_X53Y125_C4 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y128_D = LIOB33_X0Y127_IOB_X0Y128_I;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_C5 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y127_D = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_C6 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign RIOB33_X105Y135_IOB_X1Y135_O = CLBLM_R_X37Y123_SLICE_X56Y123_AO6;
  assign RIOI3_SING_X105Y149_OLOGIC_X1Y149_T1 = 1'b1;
  assign CLBLM_R_X35Y125_SLICE_X53Y125_C5 = LIOB33_X0Y135_IOB_X0Y136_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_D = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_D = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_D1 = CLBLM_R_X33Y123_SLICE_X49Y123_AO6;
  assign CLBLM_R_X35Y125_SLICE_X53Y125_C6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y132_D = LIOB33_X0Y131_IOB_X0Y132_I;
  assign LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y131_D = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLM_R_X37Y127_SLICE_X56Y127_D2 = CLBLM_R_X37Y125_SLICE_X56Y125_DO6;
  assign CLBLM_R_X35Y123_SLICE_X53Y123_CX = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOB33_X105Y123_IOB_X1Y124_O = CLBLL_L_X34Y120_SLICE_X51Y120_AO6;
  assign RIOB33_X105Y123_IOB_X1Y123_O = CLBLL_L_X36Y119_SLICE_X55Y119_BO6;
  assign CLBLM_R_X37Y127_SLICE_X56Y127_D4 = CLBLL_L_X36Y127_SLICE_X55Y127_BO6;
  assign CLBLM_R_X37Y127_SLICE_X56Y127_D5 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_D3 = 1'b1;
  assign CLBLM_R_X37Y128_SLICE_X56Y128_A6 = CLBLM_R_X37Y127_SLICE_X56Y127_DO6;
  assign CLBLM_R_X37Y127_SLICE_X56Y127_D6 = CLBLM_R_X35Y128_SLICE_X52Y128_CO6;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_D4 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_D5 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_D6 = 1'b1;
  assign CLBLM_R_X37Y123_SLICE_X57Y123_A1 = LIOB33_X0Y133_IOB_X0Y133_I;
  assign CLBLM_R_X35Y125_SLICE_X53Y125_CIN = CLBLM_R_X35Y124_SLICE_X53Y124_D_CY;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_T1 = 1'b1;
  assign CLBLM_R_X37Y118_SLICE_X57Y118_B3 = CLBLL_L_X36Y116_SLICE_X54Y116_AO5;
  assign CLBLL_L_X34Y129_SLICE_X50Y129_A1 = 1'b1;
  assign CLBLL_L_X34Y129_SLICE_X50Y129_A2 = 1'b1;
  assign CLBLL_L_X34Y129_SLICE_X50Y129_A3 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X34Y129_SLICE_X50Y129_A4 = 1'b1;
  assign CLBLL_L_X34Y129_SLICE_X50Y129_A5 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLL_L_X34Y129_SLICE_X50Y129_A6 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_A6 = CLBLM_R_X35Y122_SLICE_X52Y122_B_XOR;
  assign CLBLM_R_X37Y121_SLICE_X57Y121_A1 = CLBLL_L_X36Y116_SLICE_X55Y116_AO5;
  assign CLBLM_R_X37Y121_SLICE_X57Y121_A2 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLL_L_X34Y129_SLICE_X50Y129_B1 = 1'b1;
  assign CLBLL_L_X34Y129_SLICE_X50Y129_B2 = 1'b1;
  assign CLBLL_L_X34Y129_SLICE_X50Y129_B3 = 1'b1;
  assign CLBLL_L_X34Y129_SLICE_X50Y129_B4 = 1'b1;
  assign CLBLL_L_X34Y129_SLICE_X50Y129_B5 = 1'b1;
  assign CLBLL_L_X34Y129_SLICE_X50Y129_B6 = 1'b1;
  assign CLBLM_R_X37Y121_SLICE_X57Y121_A3 = CLBLM_R_X37Y121_SLICE_X56Y121_AO6;
  assign CLBLM_R_X37Y121_SLICE_X57Y121_A4 = CLBLM_R_X37Y118_SLICE_X56Y118_AO6;
  assign CLBLM_R_X35Y115_SLICE_X53Y115_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X34Y129_SLICE_X50Y129_C1 = 1'b1;
  assign CLBLL_L_X34Y129_SLICE_X50Y129_C2 = 1'b1;
  assign CLBLL_L_X34Y129_SLICE_X50Y129_C3 = 1'b1;
  assign CLBLL_L_X34Y129_SLICE_X50Y129_C4 = 1'b1;
  assign CLBLL_L_X34Y129_SLICE_X50Y129_C5 = 1'b1;
  assign CLBLL_L_X34Y129_SLICE_X50Y129_C6 = 1'b1;
  assign CLBLM_R_X35Y115_SLICE_X53Y115_A2 = CLBLM_R_X33Y116_SLICE_X48Y116_CO6;
  assign CLBLM_R_X35Y115_SLICE_X53Y115_A3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X35Y115_SLICE_X53Y115_A4 = CLBLM_R_X35Y115_SLICE_X53Y115_BO6;
  assign CLBLM_R_X35Y115_SLICE_X53Y115_A5 = CLBLL_L_X36Y116_SLICE_X55Y116_AO5;
  assign CLBLM_R_X35Y115_SLICE_X53Y115_A6 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLM_R_X35Y115_SLICE_X53Y115_B1 = CLBLM_R_X35Y120_SLICE_X53Y120_D_XOR;
  assign CLBLM_R_X35Y115_SLICE_X53Y115_B2 = CLBLM_R_X35Y118_SLICE_X52Y118_D_XOR;
  assign CLBLL_L_X34Y129_SLICE_X50Y129_D1 = 1'b1;
  assign CLBLL_L_X34Y129_SLICE_X50Y129_D2 = 1'b1;
  assign CLBLL_L_X34Y129_SLICE_X50Y129_D3 = 1'b1;
  assign CLBLL_L_X34Y129_SLICE_X50Y129_D4 = 1'b1;
  assign CLBLL_L_X34Y129_SLICE_X50Y129_D5 = 1'b1;
  assign CLBLL_L_X34Y129_SLICE_X50Y129_D6 = 1'b1;
  assign CLBLM_R_X35Y115_SLICE_X53Y115_B4 = CLBLL_L_X36Y122_SLICE_X55Y122_AO6;
  assign CLBLM_R_X35Y115_SLICE_X53Y115_B5 = CLBLM_R_X35Y115_SLICE_X53Y115_CO6;
  assign CLBLM_R_X35Y115_SLICE_X53Y115_C1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X35Y115_SLICE_X53Y115_C2 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_R_X35Y115_SLICE_X53Y115_C3 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X35Y115_SLICE_X53Y115_C4 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLM_R_X35Y115_SLICE_X53Y115_C5 = CLBLM_R_X35Y120_SLICE_X53Y120_D_XOR;
  assign CLBLM_R_X35Y115_SLICE_X53Y115_C6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X37Y121_SLICE_X57Y121_D3 = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLM_R_X35Y115_SLICE_X53Y115_D1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X35Y115_SLICE_X53Y115_D2 = CLBLM_R_X35Y116_SLICE_X53Y116_CO6;
  assign CLBLM_R_X35Y115_SLICE_X53Y115_D3 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLM_R_X35Y115_SLICE_X53Y115_D4 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLM_R_X35Y115_SLICE_X53Y115_D5 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X35Y115_SLICE_X53Y115_D6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_B1 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_B2 = 1'b1;
  assign CLBLM_R_X37Y121_SLICE_X56Y121_A1 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X37Y121_SLICE_X56Y121_A2 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLM_R_X37Y121_SLICE_X56Y121_A3 = CLBLL_L_X36Y122_SLICE_X55Y122_AO6;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_B3 = 1'b1;
  assign CLBLM_R_X35Y115_SLICE_X52Y115_A1 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X35Y115_SLICE_X52Y115_A2 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X35Y115_SLICE_X52Y115_A3 = CLBLM_R_X35Y120_SLICE_X53Y120_A_XOR;
  assign CLBLL_L_X34Y129_SLICE_X51Y129_A1 = 1'b1;
  assign CLBLL_L_X34Y129_SLICE_X51Y129_A2 = 1'b1;
  assign CLBLL_L_X34Y129_SLICE_X51Y129_A3 = 1'b1;
  assign CLBLL_L_X34Y129_SLICE_X51Y129_A4 = 1'b1;
  assign CLBLL_L_X34Y129_SLICE_X51Y129_A5 = 1'b1;
  assign CLBLL_L_X34Y129_SLICE_X51Y129_A6 = 1'b1;
  assign CLBLM_R_X35Y115_SLICE_X52Y115_A4 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_R_X35Y115_SLICE_X52Y115_A5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X35Y115_SLICE_X52Y115_A6 = 1'b1;
  assign CLBLL_L_X34Y129_SLICE_X51Y129_B1 = 1'b1;
  assign CLBLL_L_X34Y129_SLICE_X51Y129_B2 = 1'b1;
  assign CLBLL_L_X34Y129_SLICE_X51Y129_B3 = 1'b1;
  assign CLBLL_L_X34Y129_SLICE_X51Y129_B4 = 1'b1;
  assign CLBLL_L_X34Y129_SLICE_X51Y129_B5 = 1'b1;
  assign CLBLL_L_X34Y129_SLICE_X51Y129_B6 = 1'b1;
  assign CLBLM_R_X35Y115_SLICE_X52Y115_B1 = CLBLL_L_X36Y116_SLICE_X55Y116_AO5;
  assign CLBLM_R_X35Y115_SLICE_X52Y115_B2 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X35Y115_SLICE_X52Y115_B3 = CLBLL_L_X34Y115_SLICE_X51Y115_BO6;
  assign CLBLL_L_X34Y129_SLICE_X51Y129_C1 = 1'b1;
  assign CLBLL_L_X34Y129_SLICE_X51Y129_C2 = 1'b1;
  assign CLBLL_L_X34Y129_SLICE_X51Y129_C3 = 1'b1;
  assign CLBLL_L_X34Y129_SLICE_X51Y129_C4 = 1'b1;
  assign CLBLL_L_X34Y129_SLICE_X51Y129_C5 = 1'b1;
  assign CLBLL_L_X34Y129_SLICE_X51Y129_C6 = 1'b1;
  assign CLBLM_R_X35Y115_SLICE_X52Y115_C1 = CLBLL_L_X34Y115_SLICE_X51Y115_CO6;
  assign CLBLM_R_X35Y115_SLICE_X52Y115_C2 = CLBLL_L_X34Y115_SLICE_X50Y115_BO6;
  assign CLBLM_R_X35Y115_SLICE_X52Y115_C3 = CLBLM_R_X35Y115_SLICE_X53Y115_DO6;
  assign CLBLM_R_X35Y115_SLICE_X52Y115_C4 = CLBLL_L_X34Y116_SLICE_X51Y116_CO6;
  assign CLBLM_R_X35Y115_SLICE_X52Y115_C5 = CLBLM_R_X35Y115_SLICE_X52Y115_DO6;
  assign CLBLM_R_X35Y115_SLICE_X52Y115_C6 = CLBLM_R_X33Y116_SLICE_X48Y116_CO6;
  assign CLBLL_L_X34Y129_SLICE_X51Y129_D1 = 1'b1;
  assign CLBLL_L_X34Y129_SLICE_X51Y129_D2 = 1'b1;
  assign CLBLL_L_X34Y129_SLICE_X51Y129_D3 = 1'b1;
  assign CLBLL_L_X34Y129_SLICE_X51Y129_D4 = 1'b1;
  assign CLBLL_L_X34Y129_SLICE_X51Y129_D5 = 1'b1;
  assign CLBLL_L_X34Y129_SLICE_X51Y129_D6 = 1'b1;
  assign CLBLM_R_X35Y115_SLICE_X52Y115_D1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X35Y115_SLICE_X52Y115_D2 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X35Y115_SLICE_X52Y115_D3 = CLBLM_R_X35Y116_SLICE_X52Y116_DO6;
  assign CLBLM_R_X35Y115_SLICE_X52Y115_D4 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLM_R_X35Y115_SLICE_X52Y115_D5 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLM_R_X35Y115_SLICE_X52Y115_D6 = LIOB33_X0Y119_IOB_X0Y119_I;
  assign CLBLM_R_X35Y117_SLICE_X52Y117_A6 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X35Y124_SLICE_X53Y124_C4 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_C3 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_C6 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_C5 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_C6 = 1'b1;
  assign CLBLM_R_X35Y124_SLICE_X53Y124_C5 = 1'b1;
  assign CLBLL_L_X38Y123_SLICE_X58Y123_A1 = 1'b1;
  assign CLBLL_L_X38Y123_SLICE_X58Y123_A2 = 1'b1;
  assign CLBLL_L_X38Y123_SLICE_X58Y123_A3 = 1'b1;
  assign CLBLL_L_X38Y123_SLICE_X58Y123_A4 = 1'b1;
  assign CLBLL_L_X38Y123_SLICE_X58Y123_A5 = 1'b1;
  assign CLBLL_L_X38Y123_SLICE_X58Y123_A6 = 1'b1;
  assign CLBLM_R_X35Y117_SLICE_X52Y117_B1 = CLBLL_L_X36Y121_SLICE_X55Y121_AO5;
  assign CLBLM_R_X35Y117_SLICE_X52Y117_B2 = CLBLM_R_X35Y117_SLICE_X53Y117_BO6;
  assign CLBLL_L_X38Y123_SLICE_X58Y123_B1 = 1'b1;
  assign CLBLL_L_X38Y123_SLICE_X58Y123_B2 = 1'b1;
  assign CLBLL_L_X38Y123_SLICE_X58Y123_B3 = 1'b1;
  assign CLBLL_L_X38Y123_SLICE_X58Y123_B4 = 1'b1;
  assign CLBLL_L_X38Y123_SLICE_X58Y123_B5 = 1'b1;
  assign CLBLL_L_X38Y123_SLICE_X58Y123_B6 = 1'b1;
  assign CLBLM_R_X35Y117_SLICE_X52Y117_B3 = CLBLM_R_X35Y116_SLICE_X53Y116_AO6;
  assign CLBLM_R_X35Y117_SLICE_X52Y117_B4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X35Y125_SLICE_X53Y125_D1 = 1'b1;
  assign CLBLL_L_X38Y123_SLICE_X58Y123_C1 = 1'b1;
  assign CLBLL_L_X38Y123_SLICE_X58Y123_C2 = 1'b1;
  assign CLBLL_L_X38Y123_SLICE_X58Y123_C3 = 1'b1;
  assign CLBLL_L_X38Y123_SLICE_X58Y123_C4 = 1'b1;
  assign CLBLL_L_X38Y123_SLICE_X58Y123_C5 = 1'b1;
  assign CLBLL_L_X38Y123_SLICE_X58Y123_C6 = 1'b1;
  assign CLBLM_R_X35Y117_SLICE_X52Y117_B5 = CLBLM_R_X35Y118_SLICE_X53Y118_AO6;
  assign CLBLM_R_X35Y124_SLICE_X53Y124_C6 = LIOB33_X0Y131_IOB_X0Y132_I;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_D1 = LIOB33_X0Y129_IOB_X0Y130_I;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_D2 = 1'b1;
  assign CLBLL_L_X38Y123_SLICE_X58Y123_D1 = 1'b1;
  assign CLBLL_L_X38Y123_SLICE_X58Y123_D2 = 1'b1;
  assign CLBLL_L_X38Y123_SLICE_X58Y123_D3 = 1'b1;
  assign CLBLL_L_X38Y123_SLICE_X58Y123_D4 = 1'b1;
  assign CLBLL_L_X38Y123_SLICE_X58Y123_D5 = 1'b1;
  assign CLBLL_L_X38Y123_SLICE_X58Y123_D6 = 1'b1;
  assign CLBLM_R_X35Y125_SLICE_X53Y125_D2 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_D3 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_D4 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_D5 = 1'b1;
  assign CLBLM_R_X37Y123_SLICE_X57Y123_A3 = CLBLM_R_X37Y122_SLICE_X57Y122_BO6;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_D6 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOB33_X105Y125_IOB_X1Y126_O = CLBLL_L_X34Y121_SLICE_X51Y121_AO6;
  assign RIOB33_X105Y125_IOB_X1Y125_O = CLBLM_R_X33Y121_SLICE_X48Y121_AO6;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X37Y125_SLICE_X57Y125_A5 = CLBLL_L_X36Y124_SLICE_X55Y124_AO6;
  assign CLBLL_L_X38Y123_SLICE_X59Y123_A1 = CLBLL_L_X34Y121_SLICE_X51Y121_AO6;
  assign CLBLL_L_X38Y123_SLICE_X59Y123_A2 = CLBLM_R_X33Y121_SLICE_X48Y121_AO6;
  assign CLBLL_L_X38Y123_SLICE_X59Y123_A3 = CLBLM_R_X33Y123_SLICE_X49Y123_AO6;
  assign CLBLL_L_X38Y123_SLICE_X59Y123_A4 = CLBLL_L_X34Y120_SLICE_X51Y120_AO6;
  assign CLBLL_L_X38Y123_SLICE_X59Y123_A5 = CLBLL_L_X36Y122_SLICE_X54Y122_BO6;
  assign CLBLL_L_X38Y123_SLICE_X59Y123_A6 = CLBLL_L_X36Y119_SLICE_X55Y119_BO6;
  assign CLBLM_R_X35Y124_SLICE_X53Y124_CIN = CLBLM_R_X35Y123_SLICE_X53Y123_D_CY;
  assign CLBLL_L_X38Y123_SLICE_X59Y123_B1 = 1'b1;
  assign CLBLL_L_X38Y123_SLICE_X59Y123_B2 = 1'b1;
  assign CLBLL_L_X38Y123_SLICE_X59Y123_B3 = 1'b1;
  assign CLBLL_L_X38Y123_SLICE_X59Y123_B4 = 1'b1;
  assign CLBLL_L_X38Y123_SLICE_X59Y123_B5 = 1'b1;
  assign CLBLL_L_X38Y123_SLICE_X59Y123_B6 = 1'b1;
  assign CLBLM_R_X35Y117_SLICE_X52Y117_C6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X38Y123_SLICE_X59Y123_C1 = 1'b1;
  assign CLBLL_L_X38Y123_SLICE_X59Y123_C2 = 1'b1;
  assign CLBLL_L_X38Y123_SLICE_X59Y123_C3 = 1'b1;
  assign CLBLL_L_X38Y123_SLICE_X59Y123_C4 = 1'b1;
  assign CLBLL_L_X38Y123_SLICE_X59Y123_C5 = 1'b1;
  assign CLBLL_L_X38Y123_SLICE_X59Y123_C6 = 1'b1;
  assign CLBLM_R_X37Y125_SLICE_X57Y125_A6 = CLBLL_L_X36Y116_SLICE_X55Y116_AO5;
  assign CLBLM_R_X35Y122_SLICE_X53Y122_C6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X38Y123_SLICE_X59Y123_D1 = 1'b1;
  assign CLBLL_L_X38Y123_SLICE_X59Y123_D2 = 1'b1;
  assign CLBLL_L_X38Y123_SLICE_X59Y123_D3 = 1'b1;
  assign CLBLL_L_X38Y123_SLICE_X59Y123_D4 = 1'b1;
  assign CLBLL_L_X38Y123_SLICE_X59Y123_D5 = 1'b1;
  assign CLBLL_L_X38Y123_SLICE_X59Y123_D6 = 1'b1;
  assign CLBLM_R_X35Y123_SLICE_X53Y123_D2 = LIOB33_X0Y129_IOB_X0Y129_I;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_B2 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_B3 = 1'b1;
  assign CLBLL_L_X36Y115_SLICE_X54Y115_A1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X36Y115_SLICE_X54Y115_A2 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLL_L_X36Y115_SLICE_X54Y115_A3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X36Y115_SLICE_X54Y115_A4 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X36Y115_SLICE_X54Y115_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X36Y115_SLICE_X54Y115_A6 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_B4 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_B5 = 1'b1;
  assign CLBLL_L_X36Y115_SLICE_X54Y115_B1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X36Y115_SLICE_X54Y115_B2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X36Y115_SLICE_X54Y115_B3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X36Y115_SLICE_X54Y115_B4 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X36Y115_SLICE_X54Y115_B5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X36Y115_SLICE_X54Y115_B6 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_B6 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_A3 = CLBLM_R_X37Y122_SLICE_X56Y122_AO6;
  assign CLBLM_R_X35Y116_SLICE_X53Y116_A1 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X36Y115_SLICE_X54Y115_C1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X36Y115_SLICE_X54Y115_C2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X36Y115_SLICE_X54Y115_C3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X36Y115_SLICE_X54Y115_C4 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X36Y115_SLICE_X54Y115_C5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X36Y115_SLICE_X54Y115_C6 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X35Y116_SLICE_X53Y116_A2 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X35Y116_SLICE_X53Y116_A3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X35Y116_SLICE_X53Y116_A4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X35Y116_SLICE_X53Y116_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X35Y116_SLICE_X53Y116_A6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X35Y116_SLICE_X53Y116_B1 = CLBLL_L_X36Y116_SLICE_X55Y116_AO5;
  assign CLBLM_R_X35Y116_SLICE_X53Y116_B2 = CLBLM_R_X35Y116_SLICE_X52Y116_BO6;
  assign CLBLL_L_X36Y115_SLICE_X54Y115_D1 = 1'b1;
  assign CLBLL_L_X36Y115_SLICE_X54Y115_D2 = 1'b1;
  assign CLBLL_L_X36Y115_SLICE_X54Y115_D3 = 1'b1;
  assign CLBLL_L_X36Y115_SLICE_X54Y115_D4 = 1'b1;
  assign CLBLL_L_X36Y115_SLICE_X54Y115_D5 = 1'b1;
  assign CLBLL_L_X36Y115_SLICE_X54Y115_D6 = 1'b1;
  assign CLBLM_R_X35Y116_SLICE_X53Y116_C1 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_R_X35Y116_SLICE_X53Y116_C2 = CLBLM_R_X35Y118_SLICE_X52Y118_D_XOR;
  assign CLBLM_R_X35Y116_SLICE_X53Y116_C3 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X35Y116_SLICE_X53Y116_C4 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLM_R_X35Y116_SLICE_X53Y116_C5 = CLBLM_R_X35Y118_SLICE_X53Y118_BO5;
  assign CLBLM_R_X35Y116_SLICE_X53Y116_C6 = CLBLM_R_X35Y120_SLICE_X53Y120_D_XOR;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_D1 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_D2 = 1'b1;
  assign CLBLM_R_X35Y129_SLICE_X52Y129_D1 = 1'b1;
  assign CLBLM_R_X35Y116_SLICE_X53Y116_D1 = CLBLM_R_X35Y115_SLICE_X52Y115_CO6;
  assign CLBLM_R_X35Y116_SLICE_X53Y116_D2 = CLBLM_R_X33Y115_SLICE_X49Y115_BO6;
  assign CLBLM_R_X35Y116_SLICE_X53Y116_D3 = CLBLL_L_X34Y120_SLICE_X51Y120_AO6;
  assign CLBLM_R_X35Y116_SLICE_X53Y116_D4 = CLBLM_R_X35Y117_SLICE_X53Y117_CO6;
  assign CLBLM_R_X35Y116_SLICE_X53Y116_D5 = CLBLL_L_X34Y115_SLICE_X51Y115_AO6;
  assign CLBLM_R_X35Y116_SLICE_X53Y116_D6 = CLBLM_R_X35Y116_SLICE_X53Y116_BO6;
  assign CLBLM_R_X35Y124_SLICE_X53Y124_CX = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_A1 = CLBLM_R_X35Y124_SLICE_X53Y124_B_XOR;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_A2 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_A3 = CLBLL_L_X36Y122_SLICE_X55Y122_AO6;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_A4 = CLBLM_R_X37Y122_SLICE_X56Y122_BO6;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_A5 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X35Y116_SLICE_X52Y116_A1 = CLBLL_L_X36Y116_SLICE_X54Y116_BO5;
  assign CLBLM_R_X35Y116_SLICE_X52Y116_A2 = CLBLL_L_X36Y122_SLICE_X55Y122_AO5;
  assign CLBLM_R_X35Y116_SLICE_X52Y116_A3 = CLBLM_R_X35Y115_SLICE_X52Y115_AO6;
  assign CLBLM_R_X35Y116_SLICE_X52Y116_A4 = CLBLM_R_X33Y115_SLICE_X49Y115_AO5;
  assign CLBLL_L_X36Y115_SLICE_X55Y115_A1 = 1'b1;
  assign CLBLL_L_X36Y115_SLICE_X55Y115_A2 = 1'b1;
  assign CLBLL_L_X36Y115_SLICE_X55Y115_A3 = 1'b1;
  assign CLBLL_L_X36Y115_SLICE_X55Y115_A4 = 1'b1;
  assign CLBLL_L_X36Y115_SLICE_X55Y115_A5 = 1'b1;
  assign CLBLL_L_X36Y115_SLICE_X55Y115_A6 = 1'b1;
  assign CLBLM_R_X35Y116_SLICE_X52Y116_A5 = CLBLL_L_X34Y116_SLICE_X51Y116_BO6;
  assign CLBLM_R_X35Y116_SLICE_X52Y116_A6 = CLBLL_L_X34Y116_SLICE_X50Y116_DO6;
  assign CLBLL_L_X36Y115_SLICE_X55Y115_B1 = 1'b1;
  assign CLBLL_L_X36Y115_SLICE_X55Y115_B2 = 1'b1;
  assign CLBLL_L_X36Y115_SLICE_X55Y115_B3 = 1'b1;
  assign CLBLL_L_X36Y115_SLICE_X55Y115_B4 = 1'b1;
  assign CLBLL_L_X36Y115_SLICE_X55Y115_B5 = 1'b1;
  assign CLBLL_L_X36Y115_SLICE_X55Y115_B6 = 1'b1;
  assign CLBLM_R_X35Y116_SLICE_X52Y116_B1 = CLBLM_R_X35Y119_SLICE_X52Y119_B_XOR;
  assign CLBLM_R_X35Y116_SLICE_X52Y116_B2 = CLBLM_R_X35Y121_SLICE_X53Y121_B_XOR;
  assign CLBLM_R_X35Y116_SLICE_X52Y116_B4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X36Y115_SLICE_X55Y115_C1 = 1'b1;
  assign CLBLL_L_X36Y115_SLICE_X55Y115_C2 = 1'b1;
  assign CLBLL_L_X36Y115_SLICE_X55Y115_C3 = 1'b1;
  assign CLBLL_L_X36Y115_SLICE_X55Y115_C4 = 1'b1;
  assign CLBLL_L_X36Y115_SLICE_X55Y115_C5 = 1'b1;
  assign CLBLL_L_X36Y115_SLICE_X55Y115_C6 = 1'b1;
  assign CLBLM_R_X35Y116_SLICE_X52Y116_C1 = LIOB33_X0Y119_IOB_X0Y119_I;
  assign CLBLM_R_X35Y116_SLICE_X52Y116_C2 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_R_X35Y116_SLICE_X52Y116_C3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X35Y116_SLICE_X52Y116_C4 = CLBLM_R_X35Y121_SLICE_X53Y121_B_XOR;
  assign CLBLM_R_X35Y116_SLICE_X52Y116_C5 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X35Y116_SLICE_X52Y116_C6 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLM_R_X35Y116_SLICE_X52Y116_D1 = CLBLM_R_X35Y114_SLICE_X52Y114_AO6;
  assign CLBLL_L_X36Y115_SLICE_X55Y115_D1 = 1'b1;
  assign CLBLL_L_X36Y115_SLICE_X55Y115_D2 = 1'b1;
  assign CLBLL_L_X36Y115_SLICE_X55Y115_D3 = 1'b1;
  assign CLBLL_L_X36Y115_SLICE_X55Y115_D4 = 1'b1;
  assign CLBLL_L_X36Y115_SLICE_X55Y115_D5 = 1'b1;
  assign CLBLL_L_X36Y115_SLICE_X55Y115_D6 = 1'b1;
  assign CLBLM_R_X35Y116_SLICE_X52Y116_D2 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_R_X35Y116_SLICE_X52Y116_D3 = CLBLM_R_X35Y119_SLICE_X52Y119_B_XOR;
  assign CLBLM_R_X35Y116_SLICE_X52Y116_D4 = CLBLM_R_X35Y121_SLICE_X53Y121_B_XOR;
  assign CLBLM_R_X35Y116_SLICE_X52Y116_D5 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X35Y116_SLICE_X52Y116_D6 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign RIOI3_X105Y145_OLOGIC_X1Y146_T1 = 1'b1;
  assign CLBLM_R_X35Y123_SLICE_X53Y123_C6 = 1'b1;
  assign RIOI3_X105Y145_OLOGIC_X1Y145_D1 = CLBLL_L_X36Y129_SLICE_X54Y129_AO6;
  assign CLBLM_R_X35Y129_SLICE_X52Y129_D4 = 1'b1;
  assign CLBLM_R_X35Y124_SLICE_X53Y124_D2 = LIOB33_X0Y133_IOB_X0Y133_I;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_D3 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_D4 = 1'b1;
  assign CLBLL_L_X38Y124_SLICE_X58Y124_A1 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLL_L_X38Y124_SLICE_X58Y124_A2 = LIOB33_X0Y133_IOB_X0Y134_I;
  assign CLBLL_L_X38Y124_SLICE_X58Y124_A3 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X38Y124_SLICE_X58Y124_A4 = CLBLL_L_X38Y124_SLICE_X58Y124_BO6;
  assign CLBLL_L_X38Y124_SLICE_X58Y124_A5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X38Y124_SLICE_X58Y124_A6 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign RIOI3_X105Y145_OLOGIC_X1Y145_T1 = 1'b1;
  assign CLBLL_L_X38Y124_SLICE_X58Y124_B1 = CLBLM_R_X35Y123_SLICE_X52Y123_A_XOR;
  assign CLBLL_L_X38Y124_SLICE_X58Y124_B2 = CLBLM_R_X35Y125_SLICE_X53Y125_A_XOR;
  assign CLBLL_L_X38Y124_SLICE_X58Y124_B3 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLL_L_X38Y124_SLICE_X58Y124_B4 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X38Y124_SLICE_X58Y124_B5 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X38Y124_SLICE_X58Y124_B6 = CLBLL_L_X38Y124_SLICE_X58Y124_CO6;
  assign CLBLL_L_X38Y124_SLICE_X58Y124_C1 = 1'b1;
  assign CLBLL_L_X38Y124_SLICE_X58Y124_C2 = 1'b1;
  assign CLBLL_L_X38Y124_SLICE_X58Y124_C3 = LIOB33_X0Y133_IOB_X0Y134_I;
  assign CLBLL_L_X38Y124_SLICE_X58Y124_C4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X38Y124_SLICE_X58Y124_C5 = 1'b1;
  assign CLBLL_L_X38Y124_SLICE_X58Y124_C6 = 1'b1;
  assign RIOB33_X105Y127_IOB_X1Y128_O = CLBLL_L_X36Y122_SLICE_X54Y122_BO6;
  assign RIOB33_X105Y127_IOB_X1Y127_O = CLBLM_R_X33Y123_SLICE_X49Y123_AO6;
  assign CLBLL_L_X38Y124_SLICE_X58Y124_D1 = 1'b1;
  assign CLBLL_L_X38Y124_SLICE_X58Y124_D2 = 1'b1;
  assign CLBLL_L_X38Y124_SLICE_X58Y124_D3 = 1'b1;
  assign CLBLL_L_X38Y124_SLICE_X58Y124_D4 = 1'b1;
  assign CLBLL_L_X38Y124_SLICE_X58Y124_D5 = 1'b1;
  assign CLBLL_L_X38Y124_SLICE_X58Y124_D6 = 1'b1;
  assign CLBLM_R_X35Y129_SLICE_X52Y129_D6 = 1'b1;
  assign CLBLM_R_X35Y124_SLICE_X53Y124_D4 = 1'b1;
  assign CLBLM_R_X37Y124_SLICE_X57Y124_A6 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X37Y128_SLICE_X56Y128_A1 = CLBLL_L_X36Y128_SLICE_X55Y128_CO6;
  assign CLBLM_R_X35Y124_SLICE_X53Y124_D5 = 1'b1;
  assign CLBLL_L_X38Y124_SLICE_X59Y124_A1 = 1'b1;
  assign CLBLL_L_X38Y124_SLICE_X59Y124_A2 = 1'b1;
  assign CLBLL_L_X38Y124_SLICE_X59Y124_A3 = 1'b1;
  assign CLBLL_L_X38Y124_SLICE_X59Y124_A4 = 1'b1;
  assign CLBLL_L_X38Y124_SLICE_X59Y124_A5 = 1'b1;
  assign CLBLL_L_X38Y124_SLICE_X59Y124_A6 = 1'b1;
  assign CLBLL_L_X38Y124_SLICE_X59Y124_B1 = 1'b1;
  assign CLBLL_L_X38Y124_SLICE_X59Y124_B2 = 1'b1;
  assign CLBLL_L_X38Y124_SLICE_X59Y124_B3 = 1'b1;
  assign CLBLL_L_X38Y124_SLICE_X59Y124_B4 = 1'b1;
  assign CLBLL_L_X38Y124_SLICE_X59Y124_B5 = 1'b1;
  assign CLBLL_L_X38Y124_SLICE_X59Y124_B6 = 1'b1;
  assign CLBLM_R_X37Y128_SLICE_X56Y128_A2 = CLBLL_L_X36Y127_SLICE_X54Y127_BO6;
  assign CLBLL_L_X38Y124_SLICE_X59Y124_C1 = 1'b1;
  assign CLBLL_L_X38Y124_SLICE_X59Y124_C2 = 1'b1;
  assign CLBLL_L_X38Y124_SLICE_X59Y124_C3 = 1'b1;
  assign CLBLL_L_X38Y124_SLICE_X59Y124_C4 = 1'b1;
  assign CLBLL_L_X38Y124_SLICE_X59Y124_C5 = 1'b1;
  assign CLBLL_L_X38Y124_SLICE_X59Y124_C6 = 1'b1;
  assign LIOI3_X0Y125_ILOGIC_X0Y126_D = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLM_L_X32Y123_SLICE_X47Y123_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X32Y123_SLICE_X47Y123_A2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X32Y123_SLICE_X47Y123_A3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X32Y123_SLICE_X47Y123_A4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X32Y123_SLICE_X47Y123_A5 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X38Y124_SLICE_X59Y124_D1 = 1'b1;
  assign CLBLL_L_X38Y124_SLICE_X59Y124_D2 = 1'b1;
  assign CLBLL_L_X38Y124_SLICE_X59Y124_D3 = 1'b1;
  assign CLBLL_L_X38Y124_SLICE_X59Y124_D4 = 1'b1;
  assign CLBLM_L_X32Y123_SLICE_X47Y123_A6 = 1'b1;
  assign CLBLM_L_X32Y123_SLICE_X47Y123_B2 = CLBLL_L_X34Y123_SLICE_X50Y123_BO6;
  assign CLBLM_L_X32Y123_SLICE_X47Y123_B4 = CLBLM_R_X33Y125_SLICE_X49Y125_BO6;
  assign CLBLM_L_X32Y123_SLICE_X47Y123_B6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_L_X32Y123_SLICE_X47Y123_B1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X38Y124_SLICE_X59Y124_D5 = 1'b1;
  assign CLBLL_L_X38Y124_SLICE_X59Y124_D6 = 1'b1;
  assign CLBLM_L_X32Y123_SLICE_X47Y123_C1 = CLBLM_R_X33Y122_SLICE_X48Y122_AO6;
  assign CLBLM_L_X32Y123_SLICE_X47Y123_C2 = CLBLL_L_X34Y123_SLICE_X50Y123_BO6;
  assign CLBLM_L_X32Y123_SLICE_X47Y123_C3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_L_X32Y123_SLICE_X47Y123_C4 = CLBLM_L_X32Y123_SLICE_X47Y123_AO5;
  assign CLBLM_L_X32Y123_SLICE_X47Y123_C5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X32Y123_SLICE_X47Y123_C6 = CLBLM_R_X33Y125_SLICE_X49Y125_BO6;
  assign LIOI3_X0Y125_ILOGIC_X0Y125_D = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLM_L_X32Y123_SLICE_X47Y123_D1 = CLBLM_R_X33Y125_SLICE_X49Y125_BO6;
  assign CLBLM_L_X32Y123_SLICE_X47Y123_D2 = CLBLL_L_X34Y123_SLICE_X50Y123_BO6;
  assign CLBLM_L_X32Y123_SLICE_X47Y123_D3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_L_X32Y123_SLICE_X47Y123_D4 = CLBLM_L_X32Y123_SLICE_X47Y123_AO5;
  assign CLBLM_L_X32Y123_SLICE_X47Y123_D5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X32Y123_SLICE_X47Y123_D6 = CLBLM_R_X33Y122_SLICE_X48Y122_AO5;
  assign CLBLM_R_X37Y128_SLICE_X56Y128_A4 = CLBLM_R_X35Y126_SLICE_X52Y126_BO6;
  assign LIOI3_X0Y129_ILOGIC_X0Y130_D = LIOB33_X0Y129_IOB_X0Y130_I;
  assign CLBLM_L_X32Y123_SLICE_X46Y123_A1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X32Y123_SLICE_X46Y123_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X32Y123_SLICE_X46Y123_A3 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_L_X32Y123_SLICE_X46Y123_A4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X32Y123_SLICE_X46Y123_A5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X32Y123_SLICE_X46Y123_A6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_D = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y129_ILOGIC_X0Y129_D = LIOB33_X0Y129_IOB_X0Y129_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_D = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X32Y123_SLICE_X46Y123_B1 = 1'b1;
  assign CLBLM_L_X32Y123_SLICE_X46Y123_B2 = 1'b1;
  assign CLBLM_L_X32Y123_SLICE_X46Y123_B3 = 1'b1;
  assign CLBLM_L_X32Y123_SLICE_X46Y123_B4 = 1'b1;
  assign CLBLM_L_X32Y123_SLICE_X46Y123_B5 = 1'b1;
  assign CLBLM_L_X32Y123_SLICE_X46Y123_B6 = 1'b1;
  assign CLBLM_R_X37Y128_SLICE_X56Y128_A5 = CLBLL_L_X36Y127_SLICE_X54Y127_AO6;
  assign CLBLM_L_X32Y123_SLICE_X46Y123_C1 = 1'b1;
  assign CLBLM_L_X32Y123_SLICE_X46Y123_C2 = 1'b1;
  assign CLBLM_L_X32Y123_SLICE_X46Y123_C3 = 1'b1;
  assign CLBLL_L_X36Y116_SLICE_X54Y116_A1 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLL_L_X36Y116_SLICE_X54Y116_A2 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X36Y116_SLICE_X54Y116_A3 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X36Y116_SLICE_X54Y116_A4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X36Y116_SLICE_X54Y116_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X36Y116_SLICE_X54Y116_A6 = 1'b1;
  assign CLBLM_L_X32Y123_SLICE_X46Y123_C4 = 1'b1;
  assign CLBLM_L_X32Y123_SLICE_X46Y123_C6 = 1'b1;
  assign CLBLM_L_X32Y123_SLICE_X46Y123_C5 = 1'b1;
  assign CLBLL_L_X36Y116_SLICE_X54Y116_B1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X36Y116_SLICE_X54Y116_B2 = CLBLL_L_X36Y115_SLICE_X54Y115_AO5;
  assign CLBLL_L_X36Y116_SLICE_X54Y116_B3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_L_X32Y123_SLICE_X46Y123_D1 = 1'b1;
  assign CLBLL_L_X36Y116_SLICE_X54Y116_B4 = CLBLL_L_X36Y115_SLICE_X54Y115_BO6;
  assign CLBLL_L_X36Y116_SLICE_X54Y116_B5 = CLBLL_L_X36Y116_SLICE_X54Y116_AO6;
  assign CLBLL_L_X36Y116_SLICE_X54Y116_B6 = 1'b1;
  assign CLBLM_L_X32Y123_SLICE_X46Y123_D2 = 1'b1;
  assign CLBLL_L_X36Y116_SLICE_X54Y116_C1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X36Y116_SLICE_X54Y116_C2 = CLBLL_L_X36Y115_SLICE_X54Y115_CO6;
  assign CLBLL_L_X36Y116_SLICE_X54Y116_C3 = CLBLL_L_X36Y115_SLICE_X54Y115_BO6;
  assign CLBLL_L_X36Y116_SLICE_X54Y116_C4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X36Y116_SLICE_X54Y116_C5 = 1'b1;
  assign CLBLL_L_X36Y116_SLICE_X54Y116_C6 = 1'b1;
  assign CLBLM_L_X32Y123_SLICE_X46Y123_D6 = 1'b1;
  assign CLBLM_R_X35Y117_SLICE_X53Y117_A1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X35Y117_SLICE_X53Y117_A2 = CLBLL_L_X36Y116_SLICE_X55Y116_BO6;
  assign CLBLM_R_X35Y117_SLICE_X53Y117_A3 = CLBLM_R_X37Y118_SLICE_X57Y118_AO6;
  assign CLBLM_R_X35Y117_SLICE_X53Y117_A4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X35Y117_SLICE_X53Y117_A5 = CLBLL_L_X36Y115_SLICE_X54Y115_AO5;
  assign CLBLM_R_X35Y117_SLICE_X53Y117_A6 = CLBLL_L_X34Y117_SLICE_X51Y117_DO6;
  assign CLBLL_L_X36Y116_SLICE_X54Y116_D1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X36Y116_SLICE_X54Y116_D2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X36Y116_SLICE_X54Y116_D3 = CLBLL_L_X36Y121_SLICE_X54Y121_AO5;
  assign CLBLL_L_X36Y116_SLICE_X54Y116_D4 = CLBLL_L_X36Y115_SLICE_X54Y115_CO6;
  assign CLBLL_L_X36Y116_SLICE_X54Y116_D5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X36Y116_SLICE_X54Y116_D6 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X35Y117_SLICE_X53Y117_B1 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X35Y117_SLICE_X53Y117_B2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X35Y117_SLICE_X53Y117_B3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X35Y117_SLICE_X53Y117_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X35Y117_SLICE_X53Y117_B5 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X35Y117_SLICE_X53Y117_B6 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X35Y117_SLICE_X53Y117_C1 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLM_R_X35Y117_SLICE_X53Y117_C2 = CLBLL_L_X34Y128_SLICE_X50Y128_AO6;
  assign CLBLM_R_X35Y117_SLICE_X53Y117_C3 = CLBLM_R_X35Y120_SLICE_X53Y120_B_XOR;
  assign CLBLM_R_X35Y117_SLICE_X53Y117_C4 = CLBLM_R_X35Y116_SLICE_X52Y116_AO6;
  assign CLBLM_R_X35Y117_SLICE_X53Y117_C5 = CLBLM_R_X35Y117_SLICE_X53Y117_DO6;
  assign CLBLM_R_X35Y117_SLICE_X53Y117_C6 = CLBLL_L_X36Y117_SLICE_X54Y117_CO6;
  assign CLBLM_R_X37Y123_SLICE_X57Y123_D1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X37Y123_SLICE_X57Y123_D3 = 1'b1;
  assign CLBLM_R_X35Y117_SLICE_X53Y117_D1 = CLBLL_L_X34Y116_SLICE_X50Y116_DO6;
  assign CLBLM_R_X35Y117_SLICE_X53Y117_D2 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X35Y117_SLICE_X53Y117_D3 = CLBLM_R_X35Y120_SLICE_X53Y120_B_XOR;
  assign CLBLM_R_X35Y117_SLICE_X53Y117_D4 = CLBLL_L_X34Y117_SLICE_X50Y117_BO6;
  assign CLBLM_R_X35Y117_SLICE_X53Y117_D5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X35Y117_SLICE_X53Y117_D6 = CLBLL_L_X36Y116_SLICE_X55Y116_AO6;
  assign CLBLM_R_X35Y123_SLICE_X53Y123_D1 = 1'b1;
  assign CLBLM_R_X37Y123_SLICE_X56Y123_A1 = CLBLL_L_X36Y116_SLICE_X55Y116_AO5;
  assign CLBLM_R_X37Y123_SLICE_X56Y123_A2 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLM_R_X37Y123_SLICE_X56Y123_A3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X37Y123_SLICE_X56Y123_A4 = LIOB33_X0Y131_IOB_X0Y132_I;
  assign CLBLL_L_X36Y116_SLICE_X55Y116_A1 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X36Y116_SLICE_X55Y116_A2 = 1'b1;
  assign CLBLL_L_X36Y116_SLICE_X55Y116_A3 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLL_L_X36Y116_SLICE_X55Y116_A4 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X36Y116_SLICE_X55Y116_A5 = 1'b1;
  assign CLBLL_L_X36Y116_SLICE_X55Y116_A6 = 1'b1;
  assign CLBLM_R_X35Y117_SLICE_X52Y117_A1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X35Y117_SLICE_X52Y117_A2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X35Y117_SLICE_X52Y117_A3 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLL_L_X36Y116_SLICE_X55Y116_B1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X36Y116_SLICE_X55Y116_B2 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X36Y116_SLICE_X55Y116_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X36Y116_SLICE_X55Y116_B4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X36Y116_SLICE_X55Y116_B5 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X36Y116_SLICE_X55Y116_B6 = 1'b1;
  assign CLBLM_R_X33Y121_SLICE_X49Y121_D5 = 1'b1;
  assign CLBLM_R_X33Y121_SLICE_X49Y121_D6 = 1'b1;
  assign CLBLL_L_X36Y116_SLICE_X55Y116_C1 = 1'b1;
  assign CLBLL_L_X36Y116_SLICE_X55Y116_C2 = 1'b1;
  assign CLBLL_L_X36Y116_SLICE_X55Y116_C3 = 1'b1;
  assign CLBLL_L_X36Y116_SLICE_X55Y116_C4 = 1'b1;
  assign CLBLL_L_X36Y116_SLICE_X55Y116_C5 = 1'b1;
  assign CLBLL_L_X36Y116_SLICE_X55Y116_C6 = 1'b1;
  assign CLBLM_R_X35Y117_SLICE_X52Y117_B6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X35Y117_SLICE_X52Y117_C1 = CLBLM_R_X35Y116_SLICE_X53Y116_AO6;
  assign CLBLM_R_X35Y117_SLICE_X52Y117_C2 = CLBLM_R_X35Y117_SLICE_X52Y117_AO6;
  assign CLBLM_R_X35Y117_SLICE_X52Y117_C3 = CLBLM_R_X35Y117_SLICE_X53Y117_BO6;
  assign CLBLM_R_X35Y117_SLICE_X52Y117_C4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X35Y117_SLICE_X52Y117_C5 = CLBLL_L_X34Y115_SLICE_X50Y115_DO6;
  assign CLBLL_L_X36Y116_SLICE_X55Y116_D1 = 1'b1;
  assign CLBLL_L_X36Y116_SLICE_X55Y116_D2 = 1'b1;
  assign CLBLL_L_X36Y116_SLICE_X55Y116_D3 = 1'b1;
  assign CLBLL_L_X36Y116_SLICE_X55Y116_D4 = 1'b1;
  assign CLBLL_L_X36Y116_SLICE_X55Y116_D5 = 1'b1;
  assign CLBLL_L_X36Y116_SLICE_X55Y116_D6 = 1'b1;
  assign CLBLM_R_X35Y117_SLICE_X52Y117_D2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X35Y117_SLICE_X52Y117_D3 = CLBLM_R_X35Y117_SLICE_X53Y117_BO6;
  assign CLBLM_R_X35Y117_SLICE_X52Y117_D4 = CLBLL_L_X34Y115_SLICE_X50Y115_DO6;
  assign CLBLM_R_X35Y117_SLICE_X52Y117_D5 = CLBLL_L_X36Y121_SLICE_X55Y121_AO5;
  assign CLBLM_R_X35Y117_SLICE_X52Y117_D6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X35Y117_SLICE_X52Y117_D1 = CLBLM_R_X35Y116_SLICE_X53Y116_AO6;
  assign CLBLM_R_X35Y123_SLICE_X53Y123_D3 = 1'b1;
  assign CLBLM_R_X37Y123_SLICE_X57Y123_A5 = CLBLM_R_X37Y120_SLICE_X56Y120_BO6;
  assign CLBLM_R_X35Y122_SLICE_X53Y122_CIN = CLBLM_R_X35Y121_SLICE_X53Y121_D_CY;
  assign CLBLM_R_X35Y123_SLICE_X53Y123_D4 = 1'b1;
  assign RIOB33_X105Y129_IOB_X1Y130_O = CLBLM_R_X35Y119_SLICE_X53Y119_AO6;
  assign RIOB33_X105Y129_IOB_X1Y129_O = CLBLL_L_X34Y124_SLICE_X50Y124_AO6;
  assign CLBLM_R_X37Y123_SLICE_X57Y123_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X37Y127_SLICE_X56Y127_A1 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X35Y123_SLICE_X53Y123_D5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X37Y128_SLICE_X56Y128_B1 = 1'b1;
  assign CLBLM_R_X37Y127_SLICE_X56Y127_A2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X37Y127_SLICE_X56Y127_A3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X37Y128_SLICE_X56Y128_B3 = 1'b1;
  assign CLBLM_R_X37Y127_SLICE_X56Y127_A4 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X37Y127_SLICE_X56Y127_A5 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign RIOB33_X105Y133_IOB_X1Y134_O = CLBLM_R_X37Y122_SLICE_X57Y122_AO6;
  assign CLBLM_R_X37Y127_SLICE_X56Y127_A6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X35Y128_SLICE_X53Y128_A5 = CLBLM_R_X35Y125_SLICE_X52Y125_C_XOR;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_A1 = LIOB33_X0Y131_IOB_X0Y131_I;
  assign RIOB33_X105Y133_IOB_X1Y133_O = CLBLM_R_X37Y121_SLICE_X57Y121_AO6;
  assign CLBLM_R_X35Y128_SLICE_X53Y128_A6 = CLBLM_R_X35Y128_SLICE_X53Y128_CO6;
  assign CLBLL_L_X36Y117_SLICE_X54Y117_A1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X36Y117_SLICE_X54Y117_A2 = CLBLM_R_X37Y118_SLICE_X57Y118_AO6;
  assign CLBLL_L_X36Y117_SLICE_X54Y117_A3 = CLBLL_L_X36Y117_SLICE_X55Y117_AO6;
  assign CLBLL_L_X36Y117_SLICE_X54Y117_A4 = CLBLL_L_X36Y115_SLICE_X54Y115_AO5;
  assign CLBLL_L_X36Y117_SLICE_X54Y117_A5 = CLBLL_L_X36Y116_SLICE_X55Y116_BO6;
  assign CLBLL_L_X36Y117_SLICE_X54Y117_A6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_A2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X36Y117_SLICE_X54Y117_B1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X36Y117_SLICE_X54Y117_B2 = CLBLM_R_X37Y118_SLICE_X57Y118_AO6;
  assign CLBLL_L_X36Y117_SLICE_X54Y117_B3 = CLBLL_L_X36Y117_SLICE_X55Y117_AO6;
  assign CLBLL_L_X36Y117_SLICE_X54Y117_B4 = CLBLL_L_X36Y115_SLICE_X54Y115_AO5;
  assign CLBLL_L_X36Y117_SLICE_X54Y117_B5 = CLBLL_L_X36Y116_SLICE_X54Y116_AO6;
  assign CLBLL_L_X36Y117_SLICE_X54Y117_B6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X37Y124_SLICE_X57Y124_A1 = CLBLM_R_X37Y123_SLICE_X57Y123_BO6;
  assign CLBLM_R_X37Y124_SLICE_X57Y124_A2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X37Y124_SLICE_X57Y124_A3 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLL_L_X36Y117_SLICE_X54Y117_C1 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLL_L_X36Y117_SLICE_X54Y117_C2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X36Y117_SLICE_X54Y117_C3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X36Y117_SLICE_X54Y117_C4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X36Y117_SLICE_X54Y117_C5 = CLBLL_L_X36Y117_SLICE_X54Y117_DO6;
  assign CLBLL_L_X36Y117_SLICE_X54Y117_C6 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLM_R_X37Y124_SLICE_X57Y124_A4 = LIOB33_X0Y131_IOB_X0Y132_I;
  assign CLBLM_R_X37Y124_SLICE_X57Y124_A5 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLM_R_X35Y118_SLICE_X53Y118_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X35Y118_SLICE_X53Y118_A2 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X35Y118_SLICE_X53Y118_A3 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X35Y118_SLICE_X53Y118_A4 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X35Y118_SLICE_X53Y118_A5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X35Y118_SLICE_X53Y118_A6 = 1'b1;
  assign CLBLL_L_X36Y117_SLICE_X54Y117_D1 = CLBLM_R_X35Y120_SLICE_X53Y120_B_XOR;
  assign CLBLL_L_X36Y117_SLICE_X54Y117_D2 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLL_L_X36Y117_SLICE_X54Y117_D3 = CLBLM_R_X35Y118_SLICE_X52Y118_B_XOR;
  assign CLBLL_L_X36Y117_SLICE_X54Y117_D4 = CLBLL_L_X36Y116_SLICE_X54Y116_CO5;
  assign CLBLL_L_X36Y117_SLICE_X54Y117_D5 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X36Y117_SLICE_X54Y117_D6 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_R_X35Y118_SLICE_X53Y118_B1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X35Y118_SLICE_X53Y118_B2 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X35Y118_SLICE_X53Y118_B3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X35Y118_SLICE_X53Y118_B4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X35Y118_SLICE_X53Y118_B5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X35Y118_SLICE_X53Y118_B6 = 1'b1;
  assign CLBLM_R_X35Y118_SLICE_X53Y118_C1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X35Y118_SLICE_X53Y118_C2 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X35Y118_SLICE_X53Y118_C3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X35Y118_SLICE_X53Y118_C4 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X35Y118_SLICE_X53Y118_C5 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X35Y118_SLICE_X53Y118_C6 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_A4 = CLBLM_R_X37Y119_SLICE_X56Y119_AO6;
  assign CLBLM_R_X37Y124_SLICE_X57Y124_D6 = 1'b1;
  assign CLBLM_R_X37Y124_SLICE_X57Y124_D1 = 1'b1;
  assign CLBLM_R_X35Y128_SLICE_X53Y128_C1 = 1'b1;
  assign CLBLM_R_X35Y118_SLICE_X53Y118_D1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X35Y118_SLICE_X53Y118_D2 = CLBLL_L_X36Y117_SLICE_X55Y117_AO5;
  assign CLBLM_R_X35Y118_SLICE_X53Y118_D3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X35Y118_SLICE_X53Y118_D4 = CLBLM_R_X35Y118_SLICE_X53Y118_CO6;
  assign CLBLM_R_X35Y118_SLICE_X53Y118_D5 = CLBLM_R_X37Y118_SLICE_X57Y118_AO5;
  assign CLBLM_R_X35Y118_SLICE_X53Y118_D6 = CLBLL_L_X36Y115_SLICE_X54Y115_AO6;
  assign CLBLM_R_X35Y122_SLICE_X53Y122_D3 = 1'b1;
  assign CLBLL_L_X36Y117_SLICE_X55Y117_A1 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLL_L_X36Y117_SLICE_X55Y117_A2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X36Y117_SLICE_X55Y117_A3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X36Y117_SLICE_X55Y117_A4 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X36Y117_SLICE_X55Y117_A5 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X36Y117_SLICE_X55Y117_A6 = 1'b1;
  assign CLBLM_R_X35Y118_SLICE_X52Y118_A1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X35Y118_SLICE_X52Y118_A2 = 1'b1;
  assign CLBLM_R_X35Y118_SLICE_X52Y118_A3 = 1'b1;
  assign CLBLL_L_X36Y117_SLICE_X55Y117_B1 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLL_L_X36Y117_SLICE_X55Y117_B2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X36Y117_SLICE_X55Y117_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X36Y117_SLICE_X55Y117_B4 = 1'b1;
  assign CLBLL_L_X36Y117_SLICE_X55Y117_B5 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X36Y117_SLICE_X55Y117_B6 = 1'b1;
  assign CLBLM_R_X35Y118_SLICE_X52Y118_A4 = 1'b1;
  assign CLBLM_R_X35Y118_SLICE_X52Y118_A5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X35Y118_SLICE_X52Y118_A6 = 1'b1;
  assign CLBLL_L_X36Y117_SLICE_X55Y117_C1 = CLBLM_R_X37Y117_SLICE_X56Y117_AO6;
  assign CLBLL_L_X36Y117_SLICE_X55Y117_C2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X36Y117_SLICE_X55Y117_C3 = CLBLL_L_X36Y121_SLICE_X55Y121_AO5;
  assign CLBLL_L_X36Y117_SLICE_X55Y117_C4 = CLBLM_R_X35Y117_SLICE_X53Y117_BO6;
  assign CLBLL_L_X36Y117_SLICE_X55Y117_C5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X36Y117_SLICE_X55Y117_C6 = CLBLM_R_X35Y118_SLICE_X53Y118_AO6;
  assign CLBLM_R_X35Y118_SLICE_X52Y118_B1 = 1'b1;
  assign CLBLM_R_X35Y118_SLICE_X52Y118_B2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X35Y118_SLICE_X52Y118_B3 = 1'b1;
  assign CLBLM_R_X35Y118_SLICE_X52Y118_B4 = 1'b1;
  assign CLBLM_R_X35Y118_SLICE_X52Y118_B5 = 1'b1;
  assign CLBLM_R_X35Y118_SLICE_X52Y118_B6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X35Y118_SLICE_X52Y118_BX = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X35Y118_SLICE_X52Y118_C1 = 1'b1;
  assign CLBLL_L_X36Y117_SLICE_X55Y117_D1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X36Y117_SLICE_X55Y117_D2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X36Y117_SLICE_X55Y117_D3 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X36Y117_SLICE_X55Y117_D4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X36Y117_SLICE_X55Y117_D5 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLL_L_X36Y117_SLICE_X55Y117_D6 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X35Y118_SLICE_X52Y118_C5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X35Y118_SLICE_X52Y118_C6 = 1'b1;
  assign CLBLM_R_X35Y118_SLICE_X52Y118_CX = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X35Y118_SLICE_X52Y118_D1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X35Y118_SLICE_X52Y118_D2 = 1'b1;
  assign CLBLM_R_X35Y118_SLICE_X52Y118_D3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X35Y118_SLICE_X52Y118_D4 = 1'b1;
  assign CLBLM_R_X35Y118_SLICE_X52Y118_D5 = 1'b1;
  assign CLBLM_R_X35Y118_SLICE_X52Y118_D6 = 1'b1;
  assign CLBLM_R_X35Y122_SLICE_X53Y122_D5 = 1'b1;
  assign RIOB33_X105Y131_IOB_X1Y131_O = CLBLL_L_X36Y121_SLICE_X55Y121_BO6;
  assign CLBLM_R_X35Y118_SLICE_X52Y118_DX = LIOB33_X0Y103_IOB_X0Y103_I;
  assign RIOB33_X105Y131_IOB_X1Y132_O = CLBLL_L_X36Y122_SLICE_X55Y122_BO6;
  assign CLBLM_R_X37Y127_SLICE_X56Y127_B1 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X38Y126_SLICE_X58Y126_A1 = CLBLL_L_X36Y116_SLICE_X55Y116_AO5;
  assign CLBLL_L_X38Y126_SLICE_X58Y126_A2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X38Y126_SLICE_X58Y126_A3 = CLBLM_R_X37Y125_SLICE_X57Y125_DO6;
  assign CLBLL_L_X38Y126_SLICE_X58Y126_A4 = CLBLL_L_X38Y126_SLICE_X58Y126_BO6;
  assign CLBLL_L_X38Y126_SLICE_X58Y126_A5 = LIOB33_X0Y137_IOB_X0Y137_I;
  assign CLBLL_L_X38Y126_SLICE_X58Y126_A6 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLM_R_X35Y122_SLICE_X53Y122_D6 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLM_R_X37Y128_SLICE_X57Y128_A6 = 1'b1;
  assign CLBLL_L_X38Y126_SLICE_X58Y126_B1 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X38Y126_SLICE_X58Y126_B2 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLL_L_X38Y126_SLICE_X58Y126_B3 = CLBLM_R_X35Y125_SLICE_X53Y125_D_XOR;
  assign CLBLL_L_X38Y126_SLICE_X58Y126_B4 = CLBLM_R_X35Y123_SLICE_X52Y123_D_XOR;
  assign CLBLL_L_X38Y126_SLICE_X58Y126_B5 = CLBLL_L_X36Y122_SLICE_X55Y122_AO6;
  assign CLBLL_L_X38Y126_SLICE_X58Y126_B6 = CLBLL_L_X38Y126_SLICE_X58Y126_CO6;
  assign CLBLM_R_X37Y127_SLICE_X56Y127_B2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X38Y126_SLICE_X58Y126_C1 = CLBLM_R_X35Y125_SLICE_X53Y125_D_XOR;
  assign CLBLL_L_X38Y126_SLICE_X58Y126_C2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X38Y126_SLICE_X58Y126_C3 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLL_L_X38Y126_SLICE_X58Y126_C4 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X38Y126_SLICE_X58Y126_C5 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X38Y126_SLICE_X58Y126_C6 = LIOB33_X0Y137_IOB_X0Y137_I;
  assign CLBLM_R_X37Y128_SLICE_X57Y128_B1 = 1'b1;
  assign CLBLL_L_X38Y126_SLICE_X58Y126_D1 = 1'b1;
  assign CLBLL_L_X38Y126_SLICE_X58Y126_D2 = 1'b1;
  assign CLBLL_L_X38Y126_SLICE_X58Y126_D3 = 1'b1;
  assign CLBLL_L_X38Y126_SLICE_X58Y126_D4 = 1'b1;
  assign CLBLL_L_X38Y126_SLICE_X58Y126_D5 = 1'b1;
  assign CLBLL_L_X38Y126_SLICE_X58Y126_D6 = 1'b1;
  assign CLBLM_R_X37Y127_SLICE_X56Y127_B3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X37Y128_SLICE_X57Y128_B2 = 1'b1;
  assign CLBLM_R_X37Y128_SLICE_X57Y128_B4 = 1'b1;
  assign CLBLM_R_X37Y128_SLICE_X57Y128_B5 = 1'b1;
  assign CLBLM_R_X37Y128_SLICE_X57Y128_B6 = 1'b1;
  assign CLBLM_R_X37Y127_SLICE_X56Y127_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign RIOB33_X105Y135_IOB_X1Y136_O = CLBLM_R_X37Y123_SLICE_X57Y123_AO6;
  assign CLBLL_L_X38Y126_SLICE_X59Y126_A1 = CLBLM_R_X35Y116_SLICE_X53Y116_DO6;
  assign CLBLL_L_X38Y126_SLICE_X59Y126_A2 = CLBLM_R_X37Y124_SLICE_X56Y124_DO6;
  assign CLBLL_L_X38Y126_SLICE_X59Y126_A3 = CLBLM_R_X37Y128_SLICE_X56Y128_AO6;
  assign CLBLL_L_X38Y126_SLICE_X59Y126_A4 = CLBLL_L_X38Y126_SLICE_X59Y126_BO6;
  assign CLBLL_L_X38Y126_SLICE_X59Y126_A5 = CLBLL_L_X38Y123_SLICE_X59Y123_AO6;
  assign CLBLL_L_X38Y126_SLICE_X59Y126_A6 = CLBLL_L_X38Y126_SLICE_X59Y126_CO6;
  assign CLBLM_R_X35Y128_SLICE_X52Y128_A3 = CLBLM_R_X35Y128_SLICE_X53Y128_AO6;
  assign CLBLM_R_X35Y128_SLICE_X52Y128_A4 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLL_L_X38Y126_SLICE_X59Y126_B1 = CLBLM_R_X37Y123_SLICE_X57Y123_AO6;
  assign CLBLL_L_X38Y126_SLICE_X59Y126_B2 = CLBLM_R_X37Y125_SLICE_X56Y125_AO6;
  assign CLBLL_L_X38Y126_SLICE_X59Y126_B3 = CLBLM_R_X37Y125_SLICE_X57Y125_AO6;
  assign CLBLL_L_X38Y126_SLICE_X59Y126_B4 = CLBLL_L_X38Y126_SLICE_X58Y126_AO6;
  assign CLBLL_L_X38Y126_SLICE_X59Y126_B5 = CLBLM_R_X37Y123_SLICE_X56Y123_BO6;
  assign CLBLL_L_X38Y126_SLICE_X59Y126_B6 = CLBLM_R_X37Y126_SLICE_X56Y126_BO6;
  assign CLBLM_R_X35Y122_SLICE_X53Y122_DX = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X35Y128_SLICE_X52Y128_A5 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X35Y128_SLICE_X52Y128_A6 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLL_L_X38Y126_SLICE_X59Y126_C1 = CLBLM_R_X37Y122_SLICE_X57Y122_AO6;
  assign CLBLL_L_X38Y126_SLICE_X59Y126_C2 = CLBLL_L_X36Y122_SLICE_X55Y122_BO6;
  assign CLBLL_L_X38Y126_SLICE_X59Y126_C3 = CLBLM_R_X37Y121_SLICE_X57Y121_AO6;
  assign CLBLL_L_X38Y126_SLICE_X59Y126_C4 = CLBLM_R_X35Y119_SLICE_X53Y119_AO6;
  assign CLBLL_L_X38Y126_SLICE_X59Y126_C5 = CLBLL_L_X34Y124_SLICE_X50Y124_AO6;
  assign CLBLL_L_X38Y126_SLICE_X59Y126_C6 = CLBLL_L_X36Y121_SLICE_X55Y121_BO6;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_B1 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLM_R_X37Y127_SLICE_X56Y127_B5 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X37Y128_SLICE_X57Y128_C4 = 1'b1;
  assign RIOI3_X105Y117_OLOGIC_X1Y118_D1 = CLBLM_R_X35Y117_SLICE_X53Y117_CO6;
  assign RIOI3_X105Y147_OLOGIC_X1Y148_T1 = 1'b1;
  assign CLBLM_R_X37Y128_SLICE_X57Y128_C5 = 1'b1;
  assign CLBLL_L_X38Y126_SLICE_X59Y126_D1 = 1'b1;
  assign CLBLL_L_X38Y126_SLICE_X59Y126_D2 = 1'b1;
  assign CLBLL_L_X38Y126_SLICE_X59Y126_D3 = 1'b1;
  assign CLBLL_L_X38Y126_SLICE_X59Y126_D4 = 1'b1;
  assign CLBLL_L_X38Y126_SLICE_X59Y126_D5 = 1'b1;
  assign CLBLL_L_X38Y126_SLICE_X59Y126_D6 = 1'b1;
  assign CLBLM_R_X37Y128_SLICE_X57Y128_C6 = 1'b1;
  assign RIOI3_X105Y117_OLOGIC_X1Y118_T1 = 1'b1;
  assign CLBLM_R_X37Y127_SLICE_X56Y127_B6 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y147_OLOGIC_X1Y147_D1 = CLBLM_R_X37Y126_SLICE_X56Y126_BO6;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_B2 = CLBLM_R_X35Y122_SLICE_X52Y122_D_XOR;
  assign RIOI3_X105Y147_OLOGIC_X1Y147_T1 = 1'b1;
  assign CLBLM_R_X35Y128_SLICE_X52Y128_B3 = CLBLM_R_X35Y127_SLICE_X52Y127_CO6;
  assign CLBLM_R_X35Y128_SLICE_X52Y128_B4 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X35Y128_SLICE_X52Y128_B5 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLM_R_X35Y128_SLICE_X52Y128_B6 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X37Y128_SLICE_X57Y128_D1 = 1'b1;
  assign CLBLM_R_X37Y128_SLICE_X57Y128_D2 = 1'b1;
  assign CLBLM_R_X37Y128_SLICE_X57Y128_D3 = 1'b1;
  assign CLBLL_L_X36Y118_SLICE_X54Y118_A1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X36Y118_SLICE_X54Y118_A2 = CLBLM_R_X35Y118_SLICE_X53Y118_AO5;
  assign CLBLL_L_X36Y118_SLICE_X54Y118_A3 = CLBLL_L_X36Y118_SLICE_X55Y118_AO6;
  assign CLBLL_L_X36Y118_SLICE_X54Y118_A4 = CLBLL_L_X36Y121_SLICE_X55Y121_AO6;
  assign CLBLL_L_X36Y118_SLICE_X54Y118_A5 = CLBLM_R_X37Y117_SLICE_X56Y117_AO5;
  assign CLBLL_L_X36Y118_SLICE_X54Y118_A6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X37Y128_SLICE_X57Y128_D4 = 1'b1;
  assign CLBLM_R_X37Y128_SLICE_X57Y128_D5 = 1'b1;
  assign CLBLM_R_X35Y123_SLICE_X53Y123_BX = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X36Y118_SLICE_X54Y118_B1 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X36Y118_SLICE_X54Y118_B2 = CLBLL_L_X36Y117_SLICE_X54Y117_BO6;
  assign CLBLL_L_X36Y118_SLICE_X54Y118_B3 = CLBLM_L_X32Y123_SLICE_X47Y123_BO6;
  assign CLBLL_L_X36Y118_SLICE_X54Y118_B4 = CLBLM_R_X33Y124_SLICE_X49Y124_BO6;
  assign CLBLL_L_X36Y118_SLICE_X54Y118_B5 = CLBLL_L_X36Y118_SLICE_X54Y118_AO6;
  assign CLBLL_L_X36Y118_SLICE_X54Y118_B6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X37Y128_SLICE_X57Y128_D6 = 1'b1;
  assign RIOI3_X105Y127_OLOGIC_X1Y128_D1 = CLBLL_L_X36Y122_SLICE_X54Y122_BO6;
  assign CLBLM_R_X35Y123_SLICE_X53Y123_C1 = 1'b1;
  assign CLBLL_L_X36Y118_SLICE_X54Y118_C1 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X36Y118_SLICE_X54Y118_C2 = CLBLM_L_X32Y123_SLICE_X47Y123_BO6;
  assign CLBLL_L_X36Y118_SLICE_X54Y118_C3 = CLBLM_R_X33Y124_SLICE_X49Y124_CO6;
  assign CLBLL_L_X36Y118_SLICE_X54Y118_C4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X36Y118_SLICE_X54Y118_C5 = CLBLL_L_X36Y118_SLICE_X54Y118_DO6;
  assign CLBLL_L_X36Y118_SLICE_X54Y118_C6 = CLBLL_L_X36Y117_SLICE_X54Y117_BO6;
  assign CLBLM_L_X32Y117_SLICE_X47Y117_C1 = 1'b1;
  assign CLBLM_R_X35Y123_SLICE_X53Y123_C2 = 1'b1;
  assign CLBLM_R_X37Y125_SLICE_X57Y125_A1 = LIOB33_X0Y135_IOB_X0Y136_I;
  assign CLBLM_R_X35Y123_SLICE_X53Y123_C3 = LIOB33_X0Y127_IOB_X0Y128_I;
  assign CLBLM_R_X37Y125_SLICE_X57Y125_A2 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLM_R_X37Y125_SLICE_X57Y125_A3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X37Y125_SLICE_X57Y125_A4 = CLBLM_R_X37Y125_SLICE_X57Y125_BO6;
  assign CLBLM_R_X35Y119_SLICE_X53Y119_A1 = CLBLL_L_X36Y116_SLICE_X55Y116_AO5;
  assign CLBLL_L_X36Y118_SLICE_X54Y118_D1 = CLBLL_L_X36Y117_SLICE_X55Y117_BO6;
  assign CLBLL_L_X36Y118_SLICE_X54Y118_D2 = CLBLL_L_X36Y118_SLICE_X55Y118_AO6;
  assign CLBLL_L_X36Y118_SLICE_X54Y118_D3 = CLBLM_R_X35Y118_SLICE_X53Y118_AO5;
  assign CLBLL_L_X36Y118_SLICE_X54Y118_D4 = CLBLM_R_X37Y117_SLICE_X56Y117_AO5;
  assign CLBLL_L_X36Y118_SLICE_X54Y118_D5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X36Y118_SLICE_X54Y118_D6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X35Y119_SLICE_X53Y119_A2 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLM_R_X35Y119_SLICE_X53Y119_A3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X35Y119_SLICE_X53Y119_A4 = CLBLM_R_X35Y119_SLICE_X53Y119_BO6;
  assign CLBLM_R_X35Y119_SLICE_X53Y119_A5 = CLBLL_L_X36Y120_SLICE_X54Y120_AO6;
  assign CLBLM_R_X35Y119_SLICE_X53Y119_A6 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLM_R_X35Y119_SLICE_X53Y119_B1 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLM_R_X35Y119_SLICE_X53Y119_B2 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X35Y119_SLICE_X53Y119_B3 = CLBLM_R_X35Y123_SLICE_X53Y123_B_XOR;
  assign CLBLM_R_X35Y119_SLICE_X53Y119_B4 = CLBLM_R_X35Y121_SLICE_X52Y121_B_XOR;
  assign CLBLM_R_X35Y119_SLICE_X53Y119_B5 = CLBLL_L_X36Y122_SLICE_X55Y122_AO6;
  assign CLBLM_R_X35Y119_SLICE_X53Y119_B6 = CLBLM_R_X35Y119_SLICE_X53Y119_CO6;
  assign CLBLM_R_X35Y119_SLICE_X53Y119_C1 = CLBLM_R_X35Y123_SLICE_X53Y123_B_XOR;
  assign CLBLM_R_X35Y119_SLICE_X53Y119_C2 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_R_X35Y119_SLICE_X53Y119_C3 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X35Y119_SLICE_X53Y119_C4 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLM_R_X35Y119_SLICE_X53Y119_C5 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLM_R_X35Y119_SLICE_X53Y119_C6 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X35Y123_SLICE_X53Y123_CIN = CLBLM_R_X35Y122_SLICE_X53Y122_D_CY;
  assign CLBLM_R_X37Y125_SLICE_X57Y125_D1 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_R_X37Y125_SLICE_X57Y125_D2 = CLBLL_L_X36Y123_SLICE_X54Y123_DO6;
  assign CLBLM_R_X37Y125_SLICE_X57Y125_D3 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLM_R_X37Y125_SLICE_X57Y125_D4 = CLBLL_L_X34Y128_SLICE_X50Y128_AO6;
  assign CLBLM_R_X35Y119_SLICE_X53Y119_D1 = CLBLM_R_X35Y121_SLICE_X53Y121_C_XOR;
  assign CLBLM_R_X35Y119_SLICE_X53Y119_D2 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLL_L_X36Y118_SLICE_X55Y118_A1 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLL_L_X36Y118_SLICE_X55Y118_A2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X36Y118_SLICE_X55Y118_A3 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X36Y118_SLICE_X55Y118_A4 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X36Y118_SLICE_X55Y118_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X36Y118_SLICE_X55Y118_A6 = 1'b1;
  assign CLBLM_R_X35Y119_SLICE_X53Y119_D3 = CLBLL_L_X34Y120_SLICE_X51Y120_DO6;
  assign CLBLM_R_X35Y119_SLICE_X53Y119_D4 = CLBLM_R_X33Y119_SLICE_X49Y119_AO6;
  assign CLBLM_R_X35Y119_SLICE_X53Y119_D5 = CLBLL_L_X34Y128_SLICE_X50Y128_AO6;
  assign CLBLL_L_X36Y118_SLICE_X55Y118_B1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X36Y118_SLICE_X55Y118_B2 = CLBLM_R_X35Y118_SLICE_X53Y118_AO6;
  assign CLBLL_L_X36Y118_SLICE_X55Y118_B3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X36Y118_SLICE_X55Y118_B4 = CLBLL_L_X36Y118_SLICE_X55Y118_AO5;
  assign CLBLL_L_X36Y118_SLICE_X55Y118_B5 = CLBLM_R_X37Y117_SLICE_X56Y117_AO6;
  assign CLBLL_L_X36Y118_SLICE_X55Y118_B6 = CLBLL_L_X36Y121_SLICE_X55Y121_AO5;
  assign CLBLM_R_X35Y119_SLICE_X52Y119_A1 = 1'b1;
  assign CLBLM_R_X35Y119_SLICE_X52Y119_A2 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X35Y119_SLICE_X52Y119_A3 = 1'b1;
  assign CLBLL_L_X36Y118_SLICE_X55Y118_C1 = CLBLL_L_X38Y119_SLICE_X58Y119_AO6;
  assign CLBLL_L_X36Y118_SLICE_X55Y118_C2 = CLBLM_R_X37Y117_SLICE_X56Y117_AO5;
  assign CLBLL_L_X36Y118_SLICE_X55Y118_C3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X36Y118_SLICE_X55Y118_C4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X36Y118_SLICE_X55Y118_C5 = 1'b1;
  assign CLBLL_L_X36Y118_SLICE_X55Y118_C6 = CLBLL_L_X36Y117_SLICE_X55Y117_BO6;
  assign CLBLM_R_X35Y119_SLICE_X52Y119_AX = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X35Y119_SLICE_X52Y119_B1 = 1'b1;
  assign CLBLM_R_X35Y119_SLICE_X52Y119_B2 = LIOB33_X0Y119_IOB_X0Y119_I;
  assign CLBLM_R_X35Y119_SLICE_X52Y119_B3 = 1'b1;
  assign CLBLM_R_X35Y119_SLICE_X52Y119_B4 = 1'b1;
  assign CLBLM_R_X35Y119_SLICE_X52Y119_B5 = 1'b1;
  assign CLBLM_R_X35Y119_SLICE_X52Y119_B6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X35Y119_SLICE_X52Y119_BX = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X36Y118_SLICE_X55Y118_D1 = CLBLL_L_X34Y119_SLICE_X51Y119_AO6;
  assign CLBLL_L_X36Y118_SLICE_X55Y118_D2 = 1'b1;
  assign CLBLL_L_X36Y118_SLICE_X55Y118_D3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X36Y118_SLICE_X55Y118_D4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X36Y118_SLICE_X55Y118_D5 = CLBLL_L_X36Y117_SLICE_X55Y117_DO6;
  assign CLBLL_L_X36Y118_SLICE_X55Y118_D6 = CLBLL_L_X36Y116_SLICE_X54Y116_AO5;
  assign CLBLM_R_X35Y119_SLICE_X52Y119_C1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X35Y119_SLICE_X52Y119_C2 = 1'b1;
  assign CLBLM_R_X35Y119_SLICE_X52Y119_C3 = 1'b1;
  assign CLBLM_R_X35Y119_SLICE_X52Y119_C4 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLM_R_X35Y119_SLICE_X52Y119_C5 = 1'b1;
  assign CLBLM_R_X35Y119_SLICE_X52Y119_C6 = 1'b1;
  assign CLBLM_R_X35Y119_SLICE_X52Y119_CIN = CLBLM_R_X35Y118_SLICE_X52Y118_D_CY;
  assign CLBLM_R_X35Y119_SLICE_X52Y119_CX = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X35Y119_SLICE_X52Y119_D1 = 1'b1;
  assign CLBLM_R_X35Y119_SLICE_X52Y119_D2 = 1'b1;
  assign CLBLM_R_X35Y119_SLICE_X52Y119_D3 = 1'b1;
  assign CLBLM_R_X35Y119_SLICE_X52Y119_D4 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLM_R_X35Y119_SLICE_X52Y119_D5 = 1'b1;
  assign CLBLM_R_X35Y119_SLICE_X52Y119_D6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X35Y123_SLICE_X53Y123_D6 = 1'b1;
  assign CLBLM_R_X37Y123_SLICE_X57Y123_B1 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X35Y119_SLICE_X52Y119_DX = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X37Y128_SLICE_X56Y128_B4 = 1'b1;
  assign CLBLM_R_X37Y128_SLICE_X56Y128_B5 = 1'b1;
  assign CLBLM_R_X37Y128_SLICE_X56Y128_B6 = 1'b1;
  assign CLBLM_R_X37Y123_SLICE_X57Y123_B2 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_D = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X35Y123_SLICE_X53Y123_DX = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X37Y123_SLICE_X57Y123_B3 = CLBLM_R_X35Y124_SLICE_X53Y124_C_XOR;
  assign CLBLM_R_X37Y123_SLICE_X57Y123_B4 = CLBLM_R_X37Y123_SLICE_X57Y123_DO6;
  assign CLBLM_R_X37Y123_SLICE_X57Y123_B5 = CLBLM_R_X35Y122_SLICE_X52Y122_C_XOR;
  assign CLBLM_R_X37Y123_SLICE_X57Y123_B6 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign RIOI3_X105Y147_OLOGIC_X1Y148_D1 = CLBLL_L_X36Y129_SLICE_X55Y129_DO6;
  assign CLBLM_R_X37Y128_SLICE_X56Y128_C1 = 1'b1;
  assign CLBLM_R_X35Y123_SLICE_X52Y123_A2 = 1'b1;
  assign CLBLM_R_X37Y128_SLICE_X56Y128_C2 = 1'b1;
  assign CLBLM_R_X35Y123_SLICE_X52Y123_A3 = 1'b1;
  assign CLBLM_R_X37Y128_SLICE_X56Y128_C3 = 1'b1;
  assign CLBLM_R_X35Y123_SLICE_X52Y123_A4 = LIOB33_X0Y133_IOB_X0Y134_I;
  assign CLBLM_R_X37Y128_SLICE_X56Y128_C4 = 1'b1;
  assign CLBLM_R_X37Y123_SLICE_X57Y123_C1 = CLBLM_R_X35Y122_SLICE_X52Y122_D_XOR;
  assign CLBLM_R_X35Y123_SLICE_X52Y123_A5 = 1'b1;
  assign CLBLM_R_X37Y128_SLICE_X56Y128_C5 = 1'b1;
  assign CLBLM_R_X37Y123_SLICE_X57Y123_C2 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLM_R_X35Y123_SLICE_X52Y123_A6 = 1'b1;
  assign CLBLM_R_X37Y128_SLICE_X56Y128_C6 = 1'b1;
  assign CLBLM_R_X37Y123_SLICE_X57Y123_C3 = CLBLM_R_X35Y124_SLICE_X53Y124_D_XOR;
  assign CLBLM_R_X35Y120_SLICE_X53Y120_CX = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X37Y123_SLICE_X57Y123_C4 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_R_X37Y123_SLICE_X57Y123_C5 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X37Y125_SLICE_X56Y125_A6 = CLBLL_L_X36Y116_SLICE_X55Y116_AO5;
  assign CLBLM_R_X37Y123_SLICE_X57Y123_C6 = CLBLM_R_X37Y123_SLICE_X57Y123_DO5;
  assign CLBLM_R_X35Y123_SLICE_X52Y123_AX = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X35Y123_SLICE_X52Y123_B1 = 1'b1;
  assign CLBLM_R_X35Y123_SLICE_X52Y123_B2 = 1'b1;
  assign CLBLM_R_X35Y123_SLICE_X52Y123_B6 = LIOB33_X0Y135_IOB_X0Y135_I;
  assign CLBLM_R_X35Y120_SLICE_X53Y120_D1 = 1'b1;
  assign CLBLM_R_X37Y128_SLICE_X56Y128_D2 = 1'b1;
  assign CLBLM_R_X37Y128_SLICE_X56Y128_D4 = 1'b1;
  assign CLBLM_R_X37Y123_SLICE_X57Y123_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X37Y128_SLICE_X56Y128_D5 = 1'b1;
  assign CLBLM_R_X37Y128_SLICE_X56Y128_D6 = 1'b1;
  assign CLBLM_R_X35Y120_SLICE_X53Y120_D2 = 1'b1;
  assign CLBLM_R_X37Y123_SLICE_X57Y123_D4 = LIOB33_X0Y131_IOB_X0Y132_I;
  assign CLBLM_R_X35Y123_SLICE_X52Y123_C1 = 1'b1;
  assign CLBLM_R_X37Y123_SLICE_X57Y123_D5 = LIOB33_X0Y133_IOB_X0Y133_I;
  assign CLBLM_R_X35Y123_SLICE_X52Y123_C2 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_A4 = 1'b1;
  assign CLBLM_R_X37Y123_SLICE_X57Y123_D6 = 1'b1;
  assign CLBLM_R_X35Y120_SLICE_X53Y120_D3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X35Y123_SLICE_X52Y123_C6 = LIOB33_X0Y135_IOB_X0Y136_I;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_A5 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_B5 = 1'b1;
  assign CLBLL_L_X36Y119_SLICE_X54Y119_A1 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X36Y119_SLICE_X54Y119_A2 = CLBLM_R_X33Y124_SLICE_X49Y124_BO6;
  assign CLBLL_L_X36Y119_SLICE_X54Y119_A3 = CLBLL_L_X36Y118_SLICE_X54Y118_AO6;
  assign CLBLL_L_X36Y119_SLICE_X54Y119_A4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X36Y119_SLICE_X54Y119_A5 = CLBLL_L_X36Y117_SLICE_X54Y117_AO6;
  assign CLBLL_L_X36Y119_SLICE_X54Y119_A6 = CLBLL_L_X34Y123_SLICE_X50Y123_DO6;
  assign CLBLL_L_X36Y119_SLICE_X54Y119_B1 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X36Y119_SLICE_X54Y119_B2 = CLBLL_L_X34Y128_SLICE_X50Y128_AO6;
  assign CLBLL_L_X36Y119_SLICE_X54Y119_B3 = CLBLM_R_X35Y123_SLICE_X53Y123_D_XOR;
  assign CLBLL_L_X36Y119_SLICE_X54Y119_B4 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLL_L_X36Y119_SLICE_X54Y119_B5 = CLBLL_L_X36Y118_SLICE_X54Y118_BO6;
  assign CLBLL_L_X36Y119_SLICE_X54Y119_B6 = CLBLM_R_X37Y119_SLICE_X56Y119_BO6;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_A6 = 1'b1;
  assign CLBLL_L_X36Y119_SLICE_X54Y119_C1 = CLBLL_L_X36Y116_SLICE_X54Y116_BO6;
  assign CLBLL_L_X36Y119_SLICE_X54Y119_C2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X36Y119_SLICE_X54Y119_C3 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X36Y119_SLICE_X54Y119_C4 = CLBLM_L_X32Y123_SLICE_X47Y123_CO6;
  assign CLBLL_L_X36Y119_SLICE_X54Y119_C5 = CLBLM_R_X33Y124_SLICE_X49Y124_CO6;
  assign CLBLL_L_X36Y119_SLICE_X54Y119_C6 = CLBLL_L_X36Y118_SLICE_X54Y118_DO6;
  assign CLBLM_R_X37Y126_SLICE_X57Y126_A1 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLM_R_X37Y126_SLICE_X57Y126_A2 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLM_R_X37Y123_SLICE_X56Y123_A5 = CLBLL_L_X36Y122_SLICE_X55Y122_CO6;
  assign CLBLM_R_X37Y126_SLICE_X57Y126_A3 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X37Y126_SLICE_X57Y126_A4 = CLBLM_R_X37Y126_SLICE_X57Y126_BO6;
  assign CLBLM_R_X37Y126_SLICE_X57Y126_A5 = LIOB33_X0Y137_IOB_X0Y137_I;
  assign CLBLM_R_X37Y126_SLICE_X57Y126_A6 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X37Y123_SLICE_X56Y123_A6 = CLBLM_R_X37Y120_SLICE_X56Y120_AO6;
  assign CLBLL_L_X36Y119_SLICE_X54Y119_D1 = CLBLM_R_X35Y123_SLICE_X53Y123_C_XOR;
  assign CLBLL_L_X36Y119_SLICE_X54Y119_D2 = CLBLM_R_X35Y118_SLICE_X53Y118_DO6;
  assign CLBLL_L_X36Y119_SLICE_X54Y119_D3 = 1'b1;
  assign CLBLL_L_X36Y119_SLICE_X54Y119_D4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X36Y119_SLICE_X54Y119_D5 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X36Y119_SLICE_X54Y119_D6 = CLBLL_L_X36Y118_SLICE_X55Y118_BO6;
  assign CLBLM_R_X35Y120_SLICE_X53Y120_A1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X35Y120_SLICE_X53Y120_A2 = 1'b1;
  assign CLBLM_R_X35Y120_SLICE_X53Y120_A3 = 1'b1;
  assign CLBLM_R_X35Y120_SLICE_X53Y120_A4 = 1'b1;
  assign CLBLM_R_X35Y120_SLICE_X53Y120_A5 = 1'b1;
  assign CLBLM_R_X35Y120_SLICE_X53Y120_A6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X35Y120_SLICE_X53Y120_AX = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X35Y120_SLICE_X53Y120_B1 = 1'b1;
  assign CLBLM_R_X35Y120_SLICE_X53Y120_B2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X35Y120_SLICE_X53Y120_B3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X35Y120_SLICE_X53Y120_B4 = 1'b1;
  assign CLBLM_R_X35Y120_SLICE_X53Y120_B5 = 1'b1;
  assign CLBLM_R_X35Y120_SLICE_X53Y120_B6 = 1'b1;
  assign CLBLM_R_X35Y120_SLICE_X53Y120_BX = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X37Y126_SLICE_X57Y126_C3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X35Y120_SLICE_X53Y120_C1 = 1'b1;
  assign CLBLM_R_X35Y120_SLICE_X53Y120_C2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X35Y120_SLICE_X53Y120_C3 = 1'b1;
  assign CLBLM_R_X35Y120_SLICE_X53Y120_C4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X35Y120_SLICE_X53Y120_C5 = 1'b1;
  assign CLBLM_R_X35Y120_SLICE_X53Y120_C6 = 1'b1;
  assign CLBLM_R_X37Y123_SLICE_X56Y123_B1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X37Y125_SLICE_X56Y125_B2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X37Y126_SLICE_X57Y126_D1 = 1'b1;
  assign CLBLM_R_X37Y123_SLICE_X56Y123_B2 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLM_R_X37Y126_SLICE_X57Y126_D2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X36Y119_SLICE_X55Y119_A1 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLL_L_X36Y119_SLICE_X55Y119_A2 = CLBLL_L_X34Y128_SLICE_X50Y128_AO6;
  assign CLBLL_L_X36Y119_SLICE_X55Y119_A3 = CLBLL_L_X36Y119_SLICE_X54Y119_AO6;
  assign CLBLL_L_X36Y119_SLICE_X55Y119_A4 = CLBLM_R_X35Y123_SLICE_X53Y123_C_XOR;
  assign CLBLL_L_X36Y119_SLICE_X55Y119_A5 = CLBLL_L_X36Y119_SLICE_X54Y119_DO6;
  assign CLBLL_L_X36Y119_SLICE_X55Y119_A6 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_R_X35Y120_SLICE_X53Y120_D4 = 1'b1;
  assign CLBLM_R_X35Y120_SLICE_X53Y120_D5 = 1'b1;
  assign CLBLM_R_X35Y120_SLICE_X53Y120_D6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X36Y119_SLICE_X55Y119_B1 = CLBLL_L_X36Y116_SLICE_X55Y116_AO5;
  assign CLBLL_L_X36Y119_SLICE_X55Y119_B2 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLL_L_X36Y119_SLICE_X55Y119_B3 = CLBLM_R_X35Y119_SLICE_X53Y119_DO6;
  assign CLBLL_L_X36Y119_SLICE_X55Y119_B4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X36Y119_SLICE_X55Y119_B5 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X36Y119_SLICE_X55Y119_B6 = CLBLL_L_X36Y119_SLICE_X55Y119_CO6;
  assign CLBLM_R_X35Y120_SLICE_X52Y120_A1 = 1'b1;
  assign CLBLM_R_X35Y120_SLICE_X52Y120_A2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X35Y120_SLICE_X52Y120_A3 = 1'b1;
  assign CLBLL_L_X36Y119_SLICE_X55Y119_C1 = CLBLL_L_X36Y122_SLICE_X55Y122_AO6;
  assign CLBLL_L_X36Y119_SLICE_X55Y119_C2 = CLBLM_R_X35Y119_SLICE_X52Y119_C_XOR;
  assign CLBLL_L_X36Y119_SLICE_X55Y119_C3 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLL_L_X36Y119_SLICE_X55Y119_C4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X36Y119_SLICE_X55Y119_C5 = CLBLL_L_X36Y119_SLICE_X55Y119_DO6;
  assign CLBLL_L_X36Y119_SLICE_X55Y119_C6 = CLBLM_R_X35Y121_SLICE_X53Y121_C_XOR;
  assign CLBLM_R_X35Y120_SLICE_X52Y120_A4 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLM_R_X35Y120_SLICE_X52Y120_A5 = 1'b1;
  assign CLBLM_R_X35Y120_SLICE_X52Y120_A6 = 1'b1;
  assign CLBLM_R_X35Y120_SLICE_X52Y120_AX = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X35Y120_SLICE_X52Y120_B1 = 1'b1;
  assign CLBLM_R_X35Y120_SLICE_X52Y120_B2 = 1'b1;
  assign CLBLM_R_X35Y120_SLICE_X52Y120_B3 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_L_X36Y119_SLICE_X55Y119_D1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X36Y119_SLICE_X55Y119_D2 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X36Y119_SLICE_X55Y119_D3 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X36Y119_SLICE_X55Y119_D4 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X36Y119_SLICE_X55Y119_D5 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLL_L_X36Y119_SLICE_X55Y119_D6 = CLBLM_R_X35Y121_SLICE_X53Y121_C_XOR;
  assign CLBLM_R_X35Y120_SLICE_X52Y120_B6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X35Y120_SLICE_X52Y120_BX = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X35Y120_SLICE_X52Y120_C1 = 1'b1;
  assign CLBLM_R_X35Y120_SLICE_X52Y120_C2 = 1'b1;
  assign CLBLM_R_X35Y120_SLICE_X52Y120_C3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X35Y120_SLICE_X52Y120_C4 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLM_R_X35Y120_SLICE_X52Y120_C5 = 1'b1;
  assign CLBLM_R_X35Y120_SLICE_X52Y120_C6 = 1'b1;
  assign CLBLM_R_X35Y120_SLICE_X52Y120_CIN = CLBLM_R_X35Y119_SLICE_X52Y119_D_CY;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_B6 = 1'b1;
  assign CLBLM_R_X35Y120_SLICE_X52Y120_CX = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X37Y123_SLICE_X56Y123_C1 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X35Y120_SLICE_X52Y120_D1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X35Y120_SLICE_X52Y120_D2 = 1'b1;
  assign CLBLM_R_X35Y120_SLICE_X52Y120_D3 = 1'b1;
  assign CLBLM_R_X35Y120_SLICE_X52Y120_D4 = 1'b1;
  assign CLBLM_R_X35Y120_SLICE_X52Y120_D5 = 1'b1;
  assign CLBLM_R_X35Y120_SLICE_X52Y120_D6 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLM_R_X37Y123_SLICE_X56Y123_C2 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X37Y123_SLICE_X56Y123_C3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X35Y120_SLICE_X52Y120_DX = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X37Y123_SLICE_X56Y123_C4 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X35Y120_SLICE_X53Y120_DX = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X37Y123_SLICE_X56Y123_C5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X37Y118_SLICE_X57Y118_C2 = CLBLL_L_X36Y115_SLICE_X54Y115_AO6;
  assign CLBLM_R_X37Y125_SLICE_X56Y125_B5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X37Y123_SLICE_X56Y123_C6 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X37Y118_SLICE_X57Y118_C3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X37Y118_SLICE_X57Y118_C4 = CLBLL_L_X36Y116_SLICE_X54Y116_AO5;
  assign CLBLM_R_X37Y118_SLICE_X57Y118_C5 = CLBLL_L_X36Y117_SLICE_X55Y117_AO5;
  assign CLBLM_R_X37Y124_SLICE_X56Y124_A6 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X35Y118_SLICE_X52Y118_AX = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X37Y125_SLICE_X56Y125_B6 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_B2 = 1'b1;
  assign CLBLM_R_X35Y127_SLICE_X52Y127_D5 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_A2 = CLBLL_L_X36Y121_SLICE_X54Y121_AO5;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_B3 = 1'b1;
  assign CLBLM_R_X37Y123_SLICE_X56Y123_D1 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X37Y123_SLICE_X56Y123_D2 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X37Y123_SLICE_X56Y123_D3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_A3 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X37Y123_SLICE_X56Y123_D4 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_B4 = 1'b1;
  assign CLBLM_R_X37Y123_SLICE_X56Y123_D5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X37Y123_SLICE_X56Y123_D6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X37Y118_SLICE_X57Y118_D5 = CLBLL_L_X34Y119_SLICE_X51Y119_AO6;
  assign CLBLM_R_X35Y118_SLICE_X52Y118_C2 = 1'b1;
  assign CLBLM_R_X37Y118_SLICE_X57Y118_D6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X35Y118_SLICE_X52Y118_C3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X35Y118_SLICE_X52Y118_C4 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_A5 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y138_D = LIOB33_X0Y137_IOB_X0Y138_I;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_A5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_D = LIOB33_X0Y137_IOB_X0Y137_I;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_A6 = CLBLM_R_X37Y119_SLICE_X57Y119_CO6;
  assign CLBLM_R_X35Y127_SLICE_X52Y127_D6 = LIOB33_X0Y143_IOB_X0Y143_I;
  assign CLBLM_R_X37Y124_SLICE_X56Y124_B1 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X36Y120_SLICE_X54Y120_A1 = CLBLL_L_X36Y120_SLICE_X54Y120_DO6;
  assign CLBLL_L_X36Y120_SLICE_X54Y120_A2 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLL_L_X36Y120_SLICE_X54Y120_A3 = CLBLM_R_X35Y123_SLICE_X53Y123_B_XOR;
  assign CLBLL_L_X36Y120_SLICE_X54Y120_A4 = CLBLL_L_X36Y120_SLICE_X54Y120_BO6;
  assign CLBLL_L_X36Y120_SLICE_X54Y120_A5 = CLBLL_L_X34Y128_SLICE_X50Y128_AO6;
  assign CLBLL_L_X36Y120_SLICE_X54Y120_A6 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_R_X35Y122_SLICE_X53Y122_D4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X36Y120_SLICE_X54Y120_B1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X36Y120_SLICE_X54Y120_B2 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X36Y120_SLICE_X54Y120_B3 = CLBLL_L_X36Y117_SLICE_X54Y117_AO6;
  assign CLBLL_L_X36Y120_SLICE_X54Y120_B4 = CLBLL_L_X34Y119_SLICE_X51Y119_BO6;
  assign CLBLL_L_X36Y120_SLICE_X54Y120_B5 = CLBLM_R_X33Y123_SLICE_X49Y123_DO6;
  assign CLBLL_L_X36Y120_SLICE_X54Y120_B6 = CLBLL_L_X34Y123_SLICE_X50Y123_DO6;
  assign CLBLL_L_X36Y120_SLICE_X54Y120_C1 = CLBLL_L_X36Y118_SLICE_X55Y118_CO6;
  assign CLBLL_L_X36Y120_SLICE_X54Y120_C2 = CLBLL_L_X36Y116_SLICE_X54Y116_BO6;
  assign CLBLL_L_X36Y120_SLICE_X54Y120_C3 = CLBLM_R_X33Y123_SLICE_X48Y123_BO6;
  assign CLBLL_L_X36Y120_SLICE_X54Y120_C4 = CLBLM_L_X32Y123_SLICE_X47Y123_CO6;
  assign CLBLL_L_X36Y120_SLICE_X54Y120_C5 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X36Y120_SLICE_X54Y120_C6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X37Y124_SLICE_X56Y124_B2 = LIOB33_X0Y133_IOB_X0Y134_I;
  assign CLBLM_R_X37Y125_SLICE_X56Y125_C2 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X37Y127_SLICE_X57Y127_A1 = 1'b1;
  assign CLBLM_R_X37Y127_SLICE_X57Y127_A2 = 1'b1;
  assign CLBLM_R_X37Y127_SLICE_X57Y127_A3 = 1'b1;
  assign CLBLL_L_X36Y120_SLICE_X54Y120_D1 = CLBLM_R_X35Y123_SLICE_X53Y123_B_XOR;
  assign CLBLL_L_X36Y120_SLICE_X54Y120_D2 = 1'b1;
  assign CLBLL_L_X36Y120_SLICE_X54Y120_D3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X36Y120_SLICE_X54Y120_D4 = CLBLM_R_X35Y118_SLICE_X53Y118_DO6;
  assign CLBLL_L_X36Y120_SLICE_X54Y120_D5 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X36Y120_SLICE_X54Y120_D6 = CLBLL_L_X36Y117_SLICE_X55Y117_CO6;
  assign CLBLM_R_X37Y127_SLICE_X57Y127_A4 = 1'b1;
  assign CLBLM_R_X37Y127_SLICE_X57Y127_A5 = 1'b1;
  assign CLBLM_R_X35Y121_SLICE_X53Y121_A1 = 1'b1;
  assign CLBLM_R_X35Y121_SLICE_X53Y121_A2 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X35Y121_SLICE_X53Y121_A3 = 1'b1;
  assign CLBLM_R_X35Y121_SLICE_X53Y121_A4 = 1'b1;
  assign CLBLM_R_X35Y121_SLICE_X53Y121_A5 = 1'b1;
  assign CLBLM_R_X35Y121_SLICE_X53Y121_A6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X35Y121_SLICE_X53Y121_AX = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X37Y124_SLICE_X56Y124_B3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X35Y121_SLICE_X53Y121_B1 = 1'b1;
  assign CLBLM_R_X35Y121_SLICE_X53Y121_B2 = LIOB33_X0Y119_IOB_X0Y119_I;
  assign CLBLM_R_X35Y121_SLICE_X53Y121_B3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X35Y121_SLICE_X53Y121_B4 = 1'b1;
  assign CLBLM_R_X35Y121_SLICE_X53Y121_B5 = 1'b1;
  assign CLBLM_R_X35Y121_SLICE_X53Y121_B6 = 1'b1;
  assign CLBLM_R_X37Y125_SLICE_X56Y125_C3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X37Y127_SLICE_X57Y127_C1 = 1'b1;
  assign CLBLM_R_X35Y121_SLICE_X53Y121_BX = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X37Y122_SLICE_X57Y122_A6 = CLBLL_L_X36Y116_SLICE_X55Y116_AO5;
  assign CLBLM_R_X35Y121_SLICE_X53Y121_C1 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLM_R_X35Y121_SLICE_X53Y121_C2 = 1'b1;
  assign CLBLM_R_X35Y121_SLICE_X53Y121_C3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X35Y121_SLICE_X53Y121_C4 = 1'b1;
  assign CLBLM_R_X35Y121_SLICE_X53Y121_C5 = 1'b1;
  assign CLBLM_R_X35Y121_SLICE_X53Y121_C6 = 1'b1;
  assign CLBLL_L_X36Y120_SLICE_X55Y120_A1 = CLBLM_R_X33Y123_SLICE_X48Y123_BO6;
  assign CLBLL_L_X36Y120_SLICE_X55Y120_A2 = CLBLM_L_X32Y123_SLICE_X47Y123_DO6;
  assign CLBLL_L_X36Y120_SLICE_X55Y120_A3 = CLBLL_L_X36Y116_SLICE_X54Y116_CO6;
  assign CLBLL_L_X36Y120_SLICE_X55Y120_A4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X36Y120_SLICE_X55Y120_A5 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X36Y120_SLICE_X55Y120_A6 = CLBLL_L_X36Y118_SLICE_X55Y118_CO6;
  assign CLBLM_R_X35Y121_SLICE_X53Y121_CIN = CLBLM_R_X35Y120_SLICE_X53Y120_D_CY;
  assign CLBLM_R_X35Y121_SLICE_X53Y121_CX = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X35Y121_SLICE_X53Y121_D1 = 1'b1;
  assign CLBLL_L_X36Y120_SLICE_X55Y120_B1 = CLBLL_L_X36Y120_SLICE_X55Y120_DO6;
  assign CLBLL_L_X36Y120_SLICE_X55Y120_B2 = CLBLM_R_X35Y125_SLICE_X53Y125_A_XOR;
  assign CLBLL_L_X36Y120_SLICE_X55Y120_B3 = CLBLL_L_X34Y128_SLICE_X50Y128_AO6;
  assign CLBLL_L_X36Y120_SLICE_X55Y120_B4 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X36Y120_SLICE_X55Y120_B5 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLL_L_X36Y120_SLICE_X55Y120_B6 = CLBLL_L_X36Y120_SLICE_X55Y120_CO6;
  assign CLBLM_R_X35Y121_SLICE_X53Y121_D2 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLM_R_X35Y121_SLICE_X53Y121_D3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X35Y121_SLICE_X53Y121_D4 = 1'b1;
  assign CLBLL_L_X36Y120_SLICE_X55Y120_C1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X36Y120_SLICE_X55Y120_C2 = CLBLL_L_X36Y116_SLICE_X54Y116_CO6;
  assign CLBLL_L_X36Y120_SLICE_X55Y120_C3 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X36Y120_SLICE_X55Y120_C4 = CLBLM_R_X33Y123_SLICE_X48Y123_CO6;
  assign CLBLL_L_X36Y120_SLICE_X55Y120_C5 = CLBLM_R_X37Y119_SLICE_X57Y119_DO6;
  assign CLBLL_L_X36Y120_SLICE_X55Y120_C6 = CLBLM_L_X32Y123_SLICE_X47Y123_DO6;
  assign CLBLM_R_X35Y121_SLICE_X52Y121_A1 = 1'b1;
  assign CLBLM_R_X35Y121_SLICE_X52Y121_A2 = 1'b1;
  assign CLBLM_R_X35Y121_SLICE_X52Y121_A3 = 1'b1;
  assign CLBLM_R_X35Y121_SLICE_X52Y121_A4 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLM_R_X35Y121_SLICE_X52Y121_A5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X35Y121_SLICE_X52Y121_A6 = 1'b1;
  assign CLBLM_R_X35Y121_SLICE_X52Y121_AX = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X35Y121_SLICE_X52Y121_B1 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLL_L_X36Y120_SLICE_X55Y120_D1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X36Y120_SLICE_X55Y120_D2 = CLBLM_R_X35Y125_SLICE_X53Y125_A_XOR;
  assign CLBLL_L_X36Y120_SLICE_X55Y120_D3 = CLBLM_R_X37Y118_SLICE_X57Y118_DO6;
  assign CLBLL_L_X36Y120_SLICE_X55Y120_D4 = CLBLM_R_X37Y119_SLICE_X56Y119_DO6;
  assign CLBLL_L_X36Y120_SLICE_X55Y120_D5 = 1'b1;
  assign CLBLL_L_X36Y120_SLICE_X55Y120_D6 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X35Y121_SLICE_X52Y121_B2 = 1'b1;
  assign CLBLM_R_X35Y121_SLICE_X52Y121_B3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X35Y121_SLICE_X52Y121_B4 = 1'b1;
  assign CLBLM_R_X35Y121_SLICE_X52Y121_B5 = 1'b1;
  assign CLBLM_R_X35Y121_SLICE_X52Y121_B6 = 1'b1;
  assign CLBLM_R_X35Y121_SLICE_X52Y121_BX = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X35Y121_SLICE_X52Y121_C1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X35Y121_SLICE_X52Y121_C2 = 1'b1;
  assign CLBLM_R_X35Y121_SLICE_X52Y121_C3 = 1'b1;
  assign CLBLM_R_X35Y121_SLICE_X52Y121_C4 = 1'b1;
  assign CLBLM_R_X35Y121_SLICE_X52Y121_C5 = LIOB33_X0Y127_IOB_X0Y128_I;
  assign CLBLM_R_X35Y121_SLICE_X52Y121_C6 = 1'b1;
  assign CLBLM_R_X35Y121_SLICE_X52Y121_CIN = CLBLM_R_X35Y120_SLICE_X52Y120_D_CY;
  assign CLBLM_R_X37Y124_SLICE_X56Y124_B6 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLM_R_X37Y127_SLICE_X56Y127_D1 = CLBLM_R_X37Y126_SLICE_X57Y126_AO6;
  assign CLBLM_R_X35Y121_SLICE_X52Y121_CX = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X37Y127_SLICE_X56Y127_D3 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLM_R_X35Y121_SLICE_X52Y121_D1 = 1'b1;
  assign CLBLM_R_X35Y121_SLICE_X52Y121_D2 = 1'b1;
  assign CLBLM_R_X35Y121_SLICE_X52Y121_D3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X35Y121_SLICE_X52Y121_D4 = LIOB33_X0Y129_IOB_X0Y129_I;
  assign CLBLM_R_X35Y121_SLICE_X52Y121_D5 = 1'b1;
  assign CLBLM_R_X35Y121_SLICE_X52Y121_D6 = 1'b1;
  assign CLBLM_R_X37Y125_SLICE_X56Y125_C6 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X35Y121_SLICE_X52Y121_DX = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_B5 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign LIOI3_X0Y135_ILOGIC_X0Y136_D = LIOB33_X0Y135_IOB_X0Y136_I;
  assign LIOI3_X0Y135_ILOGIC_X0Y135_D = LIOB33_X0Y135_IOB_X0Y135_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_D = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_B6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_D = LIOB33_X0Y105_IOB_X0Y105_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_D = LIOB33_X0Y113_IOB_X0Y114_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_D = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X37Y124_SLICE_X56Y124_C1 = CLBLM_R_X37Y124_SLICE_X57Y124_BO6;
  assign CLBLM_R_X37Y124_SLICE_X56Y124_C2 = CLBLM_R_X37Y124_SLICE_X57Y124_AO6;
  assign CLBLL_L_X36Y121_SLICE_X54Y121_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X36Y121_SLICE_X54Y121_A2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X36Y121_SLICE_X54Y121_A3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X36Y121_SLICE_X54Y121_A4 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X36Y121_SLICE_X54Y121_A5 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X36Y121_SLICE_X54Y121_A6 = 1'b1;
  assign CLBLM_R_X37Y123_SLICE_X56Y123_B3 = CLBLL_L_X36Y123_SLICE_X54Y123_BO6;
  assign CLBLL_L_X36Y121_SLICE_X54Y121_B1 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLL_L_X36Y121_SLICE_X54Y121_B2 = CLBLM_R_X35Y120_SLICE_X52Y120_D_XOR;
  assign CLBLL_L_X36Y121_SLICE_X54Y121_B3 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X36Y121_SLICE_X54Y121_B4 = CLBLM_R_X35Y122_SLICE_X53Y122_D_XOR;
  assign CLBLL_L_X36Y121_SLICE_X54Y121_B5 = CLBLL_L_X36Y122_SLICE_X55Y122_AO6;
  assign CLBLL_L_X36Y121_SLICE_X54Y121_B6 = CLBLL_L_X36Y121_SLICE_X54Y121_CO6;
  assign CLBLL_L_X36Y125_SLICE_X55Y125_C1 = CLBLL_L_X34Y125_SLICE_X50Y125_AO6;
  assign CLBLM_R_X37Y124_SLICE_X56Y124_C3 = CLBLM_R_X37Y120_SLICE_X56Y120_AO6;
  assign CLBLL_L_X36Y125_SLICE_X55Y125_C2 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X36Y121_SLICE_X54Y121_C1 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLL_L_X36Y121_SLICE_X54Y121_C2 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLL_L_X36Y121_SLICE_X54Y121_C3 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X36Y121_SLICE_X54Y121_C4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X36Y121_SLICE_X54Y121_C5 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X36Y121_SLICE_X54Y121_C6 = CLBLM_R_X35Y122_SLICE_X53Y122_D_XOR;
  assign CLBLM_R_X37Y123_SLICE_X56Y123_B4 = LIOB33_X0Y135_IOB_X0Y135_I;
  assign CLBLL_L_X36Y125_SLICE_X55Y125_C5 = CLBLL_L_X36Y124_SLICE_X55Y124_BO6;
  assign CLBLL_L_X36Y121_SLICE_X54Y121_D1 = CLBLL_L_X36Y121_SLICE_X54Y121_AO6;
  assign CLBLL_L_X36Y121_SLICE_X54Y121_D2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X36Y121_SLICE_X54Y121_D3 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X36Y121_SLICE_X54Y121_D4 = CLBLL_L_X36Y121_SLICE_X54Y121_AO5;
  assign CLBLL_L_X36Y121_SLICE_X54Y121_D5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X36Y121_SLICE_X54Y121_D6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X37Y128_SLICE_X57Y128_A1 = 1'b1;
  assign CLBLM_R_X37Y128_SLICE_X57Y128_A2 = 1'b1;
  assign CLBLM_R_X33Y122_SLICE_X49Y122_C5 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X37Y128_SLICE_X57Y128_A3 = 1'b1;
  assign CLBLM_R_X37Y128_SLICE_X57Y128_A4 = 1'b1;
  assign CLBLM_R_X37Y128_SLICE_X57Y128_A5 = 1'b1;
  assign CLBLM_R_X33Y122_SLICE_X49Y122_C6 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X35Y122_SLICE_X53Y122_A1 = 1'b1;
  assign CLBLM_R_X35Y122_SLICE_X53Y122_A2 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLM_R_X35Y122_SLICE_X53Y122_A3 = 1'b1;
  assign CLBLM_R_X35Y122_SLICE_X53Y122_A4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X35Y122_SLICE_X53Y122_A5 = 1'b1;
  assign CLBLM_R_X35Y122_SLICE_X53Y122_A6 = 1'b1;
  assign CLBLM_R_X37Y123_SLICE_X56Y123_B5 = CLBLL_L_X36Y116_SLICE_X55Y116_AO5;
  assign CLBLM_R_X35Y122_SLICE_X53Y122_AX = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X37Y128_SLICE_X57Y128_B3 = 1'b1;
  assign CLBLM_R_X35Y122_SLICE_X53Y122_B1 = 1'b1;
  assign CLBLM_R_X35Y122_SLICE_X53Y122_B2 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLM_R_X35Y122_SLICE_X53Y122_B3 = 1'b1;
  assign CLBLM_R_X35Y122_SLICE_X53Y122_B4 = 1'b1;
  assign CLBLM_R_X35Y122_SLICE_X53Y122_B5 = 1'b1;
  assign CLBLM_R_X35Y122_SLICE_X53Y122_B6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X37Y128_SLICE_X57Y128_C1 = 1'b1;
  assign CLBLM_R_X37Y128_SLICE_X57Y128_C2 = 1'b1;
  assign CLBLM_R_X35Y122_SLICE_X53Y122_BX = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X37Y128_SLICE_X57Y128_C3 = 1'b1;
  assign CLBLM_R_X35Y122_SLICE_X53Y122_C1 = 1'b1;
  assign CLBLM_R_X35Y122_SLICE_X53Y122_C2 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_L_X36Y121_SLICE_X55Y121_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X36Y121_SLICE_X55Y121_A2 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLL_L_X36Y121_SLICE_X55Y121_A3 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X36Y121_SLICE_X55Y121_A4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X36Y121_SLICE_X55Y121_A5 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X36Y121_SLICE_X55Y121_A6 = 1'b1;
  assign CLBLM_R_X35Y122_SLICE_X53Y122_C3 = 1'b1;
  assign CLBLM_R_X35Y122_SLICE_X53Y122_C4 = 1'b1;
  assign CLBLM_R_X35Y122_SLICE_X53Y122_C5 = 1'b1;
  assign CLBLL_L_X36Y121_SLICE_X55Y121_B1 = LIOB33_X0Y127_IOB_X0Y128_I;
  assign CLBLL_L_X36Y121_SLICE_X55Y121_B2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X36Y121_SLICE_X55Y121_B3 = CLBLL_L_X36Y119_SLICE_X55Y119_AO6;
  assign CLBLL_L_X36Y121_SLICE_X55Y121_B4 = CLBLL_L_X36Y116_SLICE_X55Y116_AO5;
  assign CLBLL_L_X36Y121_SLICE_X55Y121_B5 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLL_L_X36Y121_SLICE_X55Y121_B6 = CLBLL_L_X36Y121_SLICE_X55Y121_CO6;
  assign CLBLM_R_X35Y122_SLICE_X53Y122_CX = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X35Y122_SLICE_X53Y122_D1 = 1'b1;
  assign CLBLM_R_X35Y122_SLICE_X53Y122_D2 = 1'b1;
  assign CLBLL_L_X36Y121_SLICE_X55Y121_C1 = CLBLM_R_X35Y123_SLICE_X53Y123_C_XOR;
  assign CLBLL_L_X36Y121_SLICE_X55Y121_C2 = CLBLL_L_X36Y122_SLICE_X55Y122_AO6;
  assign CLBLL_L_X36Y121_SLICE_X55Y121_C3 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLL_L_X36Y121_SLICE_X55Y121_C4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X36Y121_SLICE_X55Y121_C5 = CLBLL_L_X36Y121_SLICE_X55Y121_DO6;
  assign CLBLL_L_X36Y121_SLICE_X55Y121_C6 = CLBLM_R_X35Y121_SLICE_X52Y121_C_XOR;
  assign CLBLM_R_X35Y122_SLICE_X52Y122_A1 = 1'b1;
  assign CLBLM_R_X35Y122_SLICE_X52Y122_A2 = 1'b1;
  assign CLBLM_R_X35Y122_SLICE_X52Y122_A3 = LIOB33_X0Y129_IOB_X0Y130_I;
  assign CLBLM_R_X35Y122_SLICE_X52Y122_A4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X35Y122_SLICE_X52Y122_A5 = 1'b1;
  assign CLBLM_R_X35Y122_SLICE_X52Y122_A6 = 1'b1;
  assign CLBLM_R_X37Y128_SLICE_X56Y128_B2 = 1'b1;
  assign CLBLM_R_X33Y122_SLICE_X49Y122_D2 = CLBLM_R_X35Y117_SLICE_X52Y117_BO6;
  assign CLBLL_L_X36Y121_SLICE_X55Y121_D1 = CLBLM_R_X35Y123_SLICE_X53Y123_C_XOR;
  assign CLBLL_L_X36Y121_SLICE_X55Y121_D2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X36Y121_SLICE_X55Y121_D3 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLL_L_X36Y121_SLICE_X55Y121_D4 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X36Y121_SLICE_X55Y121_D5 = LIOB33_X0Y127_IOB_X0Y128_I;
  assign CLBLL_L_X36Y121_SLICE_X55Y121_D6 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_R_X33Y122_SLICE_X49Y122_D3 = 1'b1;
  assign CLBLM_R_X35Y122_SLICE_X52Y122_AX = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X33Y122_SLICE_X49Y122_D4 = CLBLL_L_X34Y118_SLICE_X50Y118_AO6;
  assign CLBLM_R_X35Y122_SLICE_X52Y122_B1 = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLM_R_X35Y122_SLICE_X52Y122_B2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X35Y122_SLICE_X52Y122_B3 = 1'b1;
  assign CLBLM_R_X33Y122_SLICE_X49Y122_D5 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X35Y122_SLICE_X52Y122_B4 = 1'b1;
  assign CLBLM_R_X35Y122_SLICE_X52Y122_B5 = 1'b1;
  assign CLBLM_R_X35Y122_SLICE_X52Y122_B6 = 1'b1;
  assign CLBLM_R_X35Y122_SLICE_X52Y122_BX = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X35Y122_SLICE_X52Y122_C1 = 1'b1;
  assign CLBLM_R_X33Y122_SLICE_X49Y122_D6 = CLBLM_R_X35Y122_SLICE_X53Y122_C_XOR;
  assign CLBLM_R_X35Y122_SLICE_X52Y122_C2 = 1'b1;
  assign CLBLM_R_X35Y122_SLICE_X52Y122_C3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X35Y122_SLICE_X52Y122_C4 = 1'b1;
  assign CLBLM_R_X35Y122_SLICE_X52Y122_C5 = 1'b1;
  assign CLBLM_R_X35Y122_SLICE_X52Y122_C6 = LIOB33_X0Y131_IOB_X0Y132_I;
  assign CLBLM_R_X35Y122_SLICE_X52Y122_CIN = CLBLM_R_X35Y121_SLICE_X52Y121_D_CY;
  assign CLBLM_R_X37Y128_SLICE_X56Y128_D1 = 1'b1;
  assign CLBLM_R_X35Y122_SLICE_X52Y122_CX = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X37Y128_SLICE_X56Y128_D3 = 1'b1;
  assign CLBLM_R_X35Y122_SLICE_X52Y122_D1 = LIOB33_X0Y133_IOB_X0Y133_I;
  assign CLBLM_R_X35Y122_SLICE_X52Y122_D2 = 1'b1;
  assign CLBLM_R_X35Y122_SLICE_X52Y122_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X35Y122_SLICE_X52Y122_D4 = 1'b1;
  assign CLBLM_R_X35Y122_SLICE_X52Y122_D5 = 1'b1;
  assign CLBLM_R_X35Y122_SLICE_X52Y122_D6 = 1'b1;
  assign CLBLM_R_X37Y118_SLICE_X57Y118_B4 = CLBLL_L_X36Y115_SLICE_X54Y115_AO6;
  assign CLBLM_R_X35Y122_SLICE_X52Y122_DX = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_A4 = 1'b1;
  assign CLBLM_R_X37Y118_SLICE_X57Y118_B5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_A5 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_A6 = 1'b1;
  assign CLBLM_R_X33Y117_SLICE_X49Y117_A5 = CLBLL_L_X34Y117_SLICE_X51Y117_BO6;
  assign CLBLM_R_X33Y117_SLICE_X49Y117_A6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_B1 = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_B2 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_B3 = CLBLM_R_X35Y124_SLICE_X53Y124_B_XOR;
  assign CLBLM_R_X33Y117_SLICE_X49Y117_C1 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign RIOB33_X105Y141_IOB_X1Y142_O = CLBLL_L_X36Y127_SLICE_X54Y127_BO6;
  assign CLBLM_R_X33Y117_SLICE_X49Y117_C2 = CLBLM_R_X33Y118_SLICE_X49Y118_CO6;
  assign RIOB33_X105Y141_IOB_X1Y141_O = CLBLL_L_X36Y127_SLICE_X54Y127_AO6;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_B4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X33Y117_SLICE_X49Y117_C3 = CLBLM_R_X33Y117_SLICE_X48Y117_DO6;
  assign CLBLM_R_X33Y117_SLICE_X49Y117_C4 = CLBLL_L_X34Y118_SLICE_X50Y118_CO6;
  assign CLBLL_L_X36Y122_SLICE_X54Y122_A1 = CLBLM_R_X33Y122_SLICE_X49Y122_CO6;
  assign CLBLL_L_X36Y122_SLICE_X54Y122_A2 = CLBLM_R_X37Y123_SLICE_X56Y123_CO6;
  assign CLBLL_L_X36Y122_SLICE_X54Y122_A3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X36Y122_SLICE_X54Y122_A4 = CLBLM_L_X32Y123_SLICE_X46Y123_AO6;
  assign CLBLL_L_X36Y122_SLICE_X54Y122_A5 = CLBLM_R_X37Y119_SLICE_X57Y119_BO6;
  assign CLBLL_L_X36Y122_SLICE_X54Y122_A6 = 1'b1;
  assign CLBLM_R_X35Y129_SLICE_X53Y129_A3 = CLBLM_R_X35Y127_SLICE_X53Y127_D_XOR;
  assign CLBLL_L_X36Y122_SLICE_X54Y122_B1 = CLBLL_L_X36Y116_SLICE_X55Y116_AO5;
  assign CLBLL_L_X36Y122_SLICE_X54Y122_B2 = CLBLL_L_X34Y122_SLICE_X50Y122_BO6;
  assign CLBLL_L_X36Y122_SLICE_X54Y122_B3 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLL_L_X36Y122_SLICE_X54Y122_B4 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLL_L_X36Y122_SLICE_X54Y122_B5 = CLBLL_L_X36Y121_SLICE_X54Y121_BO6;
  assign CLBLL_L_X36Y122_SLICE_X54Y122_B6 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X35Y129_SLICE_X53Y129_A4 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X35Y129_SLICE_X53Y129_A5 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_B5 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X36Y122_SLICE_X54Y122_C1 = CLBLM_R_X35Y123_SLICE_X53Y123_D_XOR;
  assign CLBLL_L_X36Y122_SLICE_X54Y122_C2 = CLBLM_R_X35Y121_SLICE_X52Y121_D_XOR;
  assign CLBLL_L_X36Y122_SLICE_X54Y122_C3 = CLBLL_L_X36Y122_SLICE_X55Y122_AO6;
  assign CLBLL_L_X36Y122_SLICE_X54Y122_C4 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLL_L_X36Y122_SLICE_X54Y122_C5 = CLBLL_L_X36Y122_SLICE_X54Y122_DO6;
  assign CLBLL_L_X36Y122_SLICE_X54Y122_C6 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X36Y122_SLICE_X54Y122_D1 = CLBLM_R_X35Y123_SLICE_X53Y123_D_XOR;
  assign CLBLL_L_X36Y122_SLICE_X54Y122_D2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X36Y122_SLICE_X54Y122_D3 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X36Y122_SLICE_X54Y122_D4 = LIOB33_X0Y129_IOB_X0Y129_I;
  assign CLBLL_L_X36Y122_SLICE_X54Y122_D5 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLL_L_X36Y122_SLICE_X54Y122_D6 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_B6 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X35Y129_SLICE_X53Y129_B1 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLM_R_X35Y129_SLICE_X53Y129_B2 = LIOB33_X0Y145_IOB_X0Y145_I;
  assign CLBLM_R_X35Y123_SLICE_X53Y123_A1 = 1'b1;
  assign CLBLM_R_X35Y123_SLICE_X53Y123_A2 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLM_R_X35Y123_SLICE_X53Y123_A3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X35Y123_SLICE_X53Y123_A4 = 1'b1;
  assign CLBLM_R_X35Y123_SLICE_X53Y123_A5 = 1'b1;
  assign CLBLM_R_X35Y123_SLICE_X53Y123_A6 = 1'b1;
  assign CLBLM_R_X35Y129_SLICE_X53Y129_B3 = CLBLM_R_X35Y127_SLICE_X53Y127_D_XOR;
  assign CLBLM_R_X35Y129_SLICE_X53Y129_B4 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X35Y123_SLICE_X53Y123_AX = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X35Y123_SLICE_X53Y123_B1 = 1'b1;
  assign CLBLM_R_X35Y123_SLICE_X53Y123_B2 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLM_R_X35Y123_SLICE_X53Y123_B3 = 1'b1;
  assign CLBLM_R_X35Y123_SLICE_X53Y123_B4 = 1'b1;
  assign CLBLM_R_X35Y123_SLICE_X53Y123_B5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X35Y123_SLICE_X53Y123_B6 = 1'b1;
  assign CLBLM_R_X33Y115_SLICE_X49Y115_A1 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X33Y115_SLICE_X49Y115_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X33Y115_SLICE_X49Y115_A3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X33Y115_SLICE_X49Y115_A4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X33Y115_SLICE_X49Y115_A5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X33Y115_SLICE_X49Y115_A6 = 1'b1;
  assign CLBLL_L_X36Y122_SLICE_X55Y122_A4 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X36Y122_SLICE_X55Y122_A5 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLL_L_X36Y122_SLICE_X55Y122_A6 = 1'b1;
  assign CLBLM_R_X33Y115_SLICE_X49Y115_B1 = CLBLM_R_X33Y115_SLICE_X49Y115_DO6;
  assign CLBLM_R_X33Y115_SLICE_X49Y115_B2 = CLBLL_L_X34Y115_SLICE_X51Y115_CO6;
  assign CLBLM_R_X33Y115_SLICE_X49Y115_B3 = CLBLM_R_X33Y115_SLICE_X48Y115_AO6;
  assign CLBLM_R_X33Y115_SLICE_X49Y115_B4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X33Y115_SLICE_X49Y115_B5 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLM_R_X33Y115_SLICE_X49Y115_B6 = CLBLM_R_X33Y115_SLICE_X49Y115_CO6;
  assign CLBLL_L_X36Y122_SLICE_X55Y122_B1 = CLBLL_L_X36Y116_SLICE_X55Y116_AO5;
  assign CLBLM_R_X33Y115_SLICE_X49Y115_C1 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLM_R_X33Y115_SLICE_X49Y115_C2 = CLBLM_R_X33Y116_SLICE_X49Y116_CO6;
  assign CLBLM_R_X33Y115_SLICE_X49Y115_C3 = CLBLM_R_X35Y120_SLICE_X53Y120_C_XOR;
  assign CLBLM_R_X33Y115_SLICE_X49Y115_C4 = CLBLM_R_X33Y116_SLICE_X49Y116_DO6;
  assign CLBLM_R_X33Y115_SLICE_X49Y115_C5 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X33Y115_SLICE_X49Y115_C6 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X36Y122_SLICE_X55Y122_C1 = CLBLL_L_X36Y122_SLICE_X55Y122_AO6;
  assign CLBLL_L_X36Y122_SLICE_X55Y122_C2 = CLBLM_R_X35Y122_SLICE_X52Y122_C_XOR;
  assign CLBLL_L_X36Y122_SLICE_X55Y122_C3 = CLBLM_R_X35Y124_SLICE_X53Y124_C_XOR;
  assign CLBLL_L_X36Y122_SLICE_X55Y122_C4 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLL_L_X36Y122_SLICE_X55Y122_C5 = CLBLL_L_X36Y122_SLICE_X55Y122_DO6;
  assign CLBLL_L_X36Y122_SLICE_X55Y122_C6 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X35Y123_SLICE_X52Y123_A1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X33Y115_SLICE_X49Y115_D1 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLL_L_X36Y122_SLICE_X55Y122_D1 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLL_L_X36Y122_SLICE_X55Y122_D2 = LIOB33_X0Y131_IOB_X0Y132_I;
  assign CLBLL_L_X36Y122_SLICE_X55Y122_D3 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X33Y115_SLICE_X49Y115_D5 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X33Y115_SLICE_X49Y115_D6 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X36Y122_SLICE_X55Y122_D4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X36Y122_SLICE_X55Y122_D5 = CLBLM_R_X35Y124_SLICE_X53Y124_C_XOR;
  assign CLBLL_L_X36Y122_SLICE_X55Y122_D6 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_R_X33Y115_SLICE_X49Y115_D3 = CLBLL_L_X34Y116_SLICE_X50Y116_AO5;
  assign CLBLM_R_X33Y115_SLICE_X49Y115_D4 = CLBLM_R_X33Y117_SLICE_X48Y117_CO6;
  assign CLBLM_R_X33Y115_SLICE_X48Y115_A1 = CLBLM_R_X33Y118_SLICE_X48Y118_CO6;
  assign CLBLM_R_X33Y115_SLICE_X48Y115_A2 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLM_R_X33Y115_SLICE_X48Y115_A3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X33Y115_SLICE_X48Y115_A4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X33Y115_SLICE_X48Y115_A5 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLM_R_X33Y115_SLICE_X48Y115_A6 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X35Y123_SLICE_X52Y123_B3 = 1'b1;
  assign CLBLM_R_X35Y123_SLICE_X52Y123_B4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X35Y123_SLICE_X52Y123_B5 = 1'b1;
  assign CLBLM_R_X35Y123_SLICE_X52Y123_BX = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X33Y115_SLICE_X48Y115_B1 = 1'b1;
  assign CLBLM_R_X33Y115_SLICE_X48Y115_B2 = 1'b1;
  assign CLBLM_R_X33Y115_SLICE_X48Y115_B3 = 1'b1;
  assign CLBLM_R_X33Y115_SLICE_X48Y115_B4 = 1'b1;
  assign CLBLM_R_X33Y115_SLICE_X48Y115_B5 = 1'b1;
  assign CLBLM_R_X33Y115_SLICE_X48Y115_B6 = 1'b1;
  assign CLBLM_R_X35Y123_SLICE_X52Y123_C3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X35Y123_SLICE_X52Y123_C4 = 1'b1;
  assign CLBLM_R_X35Y123_SLICE_X52Y123_C5 = 1'b1;
  assign CLBLM_R_X35Y123_SLICE_X52Y123_CIN = CLBLM_R_X35Y122_SLICE_X52Y122_D_CY;
  assign CLBLM_R_X33Y115_SLICE_X48Y115_C1 = 1'b1;
  assign CLBLM_R_X33Y115_SLICE_X48Y115_C2 = 1'b1;
  assign CLBLM_R_X33Y115_SLICE_X48Y115_C3 = 1'b1;
  assign CLBLM_R_X33Y115_SLICE_X48Y115_C4 = 1'b1;
  assign CLBLM_R_X33Y115_SLICE_X48Y115_C5 = 1'b1;
  assign CLBLM_R_X33Y115_SLICE_X48Y115_C6 = 1'b1;
  assign CLBLM_R_X35Y123_SLICE_X52Y123_CX = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X35Y123_SLICE_X52Y123_D1 = 1'b1;
  assign CLBLM_R_X35Y123_SLICE_X52Y123_D2 = LIOB33_X0Y137_IOB_X0Y137_I;
  assign CLBLM_R_X35Y123_SLICE_X52Y123_D3 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X35Y123_SLICE_X52Y123_D4 = 1'b1;
  assign CLBLM_R_X35Y123_SLICE_X52Y123_D5 = 1'b1;
  assign CLBLM_R_X35Y123_SLICE_X52Y123_D6 = 1'b1;
  assign CLBLM_R_X35Y123_SLICE_X52Y123_DX = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X33Y115_SLICE_X48Y115_D1 = 1'b1;
  assign CLBLM_R_X33Y115_SLICE_X48Y115_D2 = 1'b1;
  assign CLBLM_R_X33Y115_SLICE_X48Y115_D3 = 1'b1;
  assign CLBLM_R_X33Y115_SLICE_X48Y115_D4 = 1'b1;
  assign CLBLM_R_X33Y115_SLICE_X48Y115_D5 = 1'b1;
  assign CLBLM_R_X33Y115_SLICE_X48Y115_D6 = 1'b1;
  assign CLBLM_R_X35Y129_SLICE_X53Y129_D1 = 1'b1;
  assign RIOI3_X105Y123_OLOGIC_X1Y124_D1 = CLBLL_L_X34Y120_SLICE_X51Y120_AO6;
  assign CLBLM_R_X35Y129_SLICE_X53Y129_D2 = 1'b1;
  assign CLBLM_R_X35Y129_SLICE_X53Y129_D3 = 1'b1;
  assign RIOI3_X105Y123_OLOGIC_X1Y124_T1 = 1'b1;
  assign CLBLM_R_X35Y129_SLICE_X53Y129_D4 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_C1 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_R_X35Y129_SLICE_X53Y129_D5 = 1'b1;
  assign RIOI3_X105Y123_OLOGIC_X1Y123_D1 = CLBLL_L_X36Y119_SLICE_X55Y119_BO6;
  assign CLBLM_R_X35Y129_SLICE_X53Y129_D6 = 1'b1;
  assign CLBLM_R_X35Y117_SLICE_X52Y117_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign RIOI3_X105Y123_OLOGIC_X1Y123_T1 = 1'b1;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_C2 = CLBLM_R_X35Y122_SLICE_X52Y122_A_XOR;
  assign CLBLM_R_X35Y117_SLICE_X52Y117_A5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X35Y129_SLICE_X52Y129_A1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_C3 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X35Y129_SLICE_X52Y129_A2 = LIOB33_X0Y141_IOB_X0Y141_I;
  assign CLBLM_R_X35Y129_SLICE_X52Y129_A3 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLM_R_X35Y129_SLICE_X52Y129_A4 = CLBLM_R_X35Y129_SLICE_X52Y129_BO6;
  assign CLBLM_R_X35Y129_SLICE_X52Y129_A5 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X35Y129_SLICE_X52Y129_A6 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_C4 = CLBLM_R_X35Y124_SLICE_X53Y124_A_XOR;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_C1 = 1'b1;
  assign RIOB33_X105Y143_IOB_X1Y144_O = CLBLL_L_X36Y129_SLICE_X55Y129_AO6;
  assign RIOB33_X105Y143_IOB_X1Y143_O = CLBLM_R_X35Y126_SLICE_X52Y126_BO6;
  assign CLBLM_R_X37Y122_SLICE_X56Y122_C5 = CLBLM_R_X37Y122_SLICE_X56Y122_DO6;
  assign CLBLM_R_X35Y129_SLICE_X52Y129_B1 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLM_R_X35Y129_SLICE_X52Y129_B2 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X35Y129_SLICE_X52Y129_B3 = CLBLM_R_X35Y126_SLICE_X53Y126_D_XOR;
  assign CLBLM_R_X35Y129_SLICE_X52Y129_B4 = CLBLM_R_X35Y124_SLICE_X52Y124_D_XOR;
  assign CLBLL_L_X36Y123_SLICE_X54Y123_A1 = CLBLL_L_X36Y117_SLICE_X55Y117_DO6;
  assign CLBLL_L_X36Y123_SLICE_X54Y123_A2 = CLBLL_L_X34Y123_SLICE_X50Y123_CO6;
  assign CLBLL_L_X36Y123_SLICE_X54Y123_A3 = CLBLM_R_X37Y123_SLICE_X56Y123_DO6;
  assign CLBLL_L_X36Y123_SLICE_X54Y123_A4 = CLBLM_R_X33Y123_SLICE_X48Y123_AO6;
  assign CLBLL_L_X36Y123_SLICE_X54Y123_A5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X36Y123_SLICE_X54Y123_A6 = 1'b1;
  assign CLBLM_R_X35Y129_SLICE_X52Y129_B5 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_R_X35Y129_SLICE_X52Y129_B6 = CLBLM_R_X35Y129_SLICE_X52Y129_CO6;
  assign CLBLL_L_X36Y123_SLICE_X54Y123_B1 = CLBLM_R_X35Y125_SLICE_X53Y125_B_XOR;
  assign CLBLL_L_X36Y123_SLICE_X54Y123_B2 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLL_L_X36Y123_SLICE_X54Y123_B3 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X36Y123_SLICE_X54Y123_B4 = CLBLM_R_X35Y123_SLICE_X52Y123_B_XOR;
  assign CLBLL_L_X36Y123_SLICE_X54Y123_B5 = CLBLL_L_X36Y122_SLICE_X55Y122_AO6;
  assign CLBLL_L_X36Y123_SLICE_X54Y123_B6 = CLBLL_L_X36Y123_SLICE_X54Y123_CO6;
  assign CLBLM_R_X35Y124_SLICE_X53Y124_B3 = 1'b1;
  assign CLBLM_R_X35Y124_SLICE_X53Y124_B4 = 1'b1;
  assign CLBLL_L_X36Y123_SLICE_X54Y123_C1 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLL_L_X36Y123_SLICE_X54Y123_C2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X36Y123_SLICE_X54Y123_C3 = CLBLM_R_X35Y125_SLICE_X53Y125_B_XOR;
  assign CLBLL_L_X36Y123_SLICE_X54Y123_C4 = LIOB33_X0Y135_IOB_X0Y135_I;
  assign CLBLL_L_X36Y123_SLICE_X54Y123_C5 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X36Y123_SLICE_X54Y123_C6 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_R_X35Y124_SLICE_X53Y124_B5 = 1'b1;
  assign CLBLM_R_X35Y124_SLICE_X53Y124_B6 = 1'b1;
  assign LIOI3_X0Y139_ILOGIC_X0Y140_D = LIOB33_X0Y139_IOB_X0Y140_I;
  assign CLBLL_L_X36Y123_SLICE_X54Y123_D1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X36Y123_SLICE_X54Y123_D2 = CLBLL_L_X36Y121_SLICE_X54Y121_DO6;
  assign CLBLL_L_X36Y123_SLICE_X54Y123_D3 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X36Y123_SLICE_X54Y123_D4 = CLBLM_R_X33Y123_SLICE_X48Y123_DO6;
  assign CLBLL_L_X36Y123_SLICE_X54Y123_D5 = CLBLM_R_X37Y119_SLICE_X57Y119_AO6;
  assign CLBLL_L_X36Y123_SLICE_X54Y123_D6 = CLBLM_R_X33Y124_SLICE_X48Y124_BO6;
  assign CLBLM_R_X35Y129_SLICE_X52Y129_C1 = 1'b1;
  assign CLBLM_R_X35Y129_SLICE_X52Y129_C2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X35Y124_SLICE_X53Y124_BX = RIOB33_X105Y103_IOB_X1Y103_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y110_D = LIOB33_X0Y109_IOB_X0Y110_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_D = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X35Y129_SLICE_X52Y129_C3 = LIOB33_X0Y141_IOB_X0Y141_I;
  assign CLBLM_R_X35Y129_SLICE_X52Y129_C4 = 1'b1;
  assign CLBLM_R_X35Y124_SLICE_X53Y124_C1 = 1'b1;
  assign CLBLM_R_X35Y129_SLICE_X52Y129_C5 = 1'b1;
  assign CLBLM_R_X35Y124_SLICE_X53Y124_A1 = 1'b1;
  assign CLBLM_R_X35Y124_SLICE_X53Y124_A2 = 1'b1;
  assign CLBLM_R_X35Y124_SLICE_X53Y124_A3 = LIOB33_X0Y129_IOB_X0Y130_I;
  assign CLBLM_R_X35Y124_SLICE_X53Y124_A4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X35Y124_SLICE_X53Y124_A5 = 1'b1;
  assign CLBLM_R_X35Y124_SLICE_X53Y124_A6 = 1'b1;
  assign CLBLM_R_X35Y124_SLICE_X53Y124_C2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X35Y124_SLICE_X53Y124_C3 = 1'b1;
  assign CLBLM_R_X35Y124_SLICE_X53Y124_AX = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X35Y129_SLICE_X52Y129_C6 = 1'b1;
  assign CLBLM_R_X35Y124_SLICE_X53Y124_B1 = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLM_R_X35Y124_SLICE_X53Y124_B2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X36Y123_SLICE_X55Y123_A1 = CLBLL_L_X36Y123_SLICE_X55Y123_DO6;
  assign CLBLL_L_X36Y123_SLICE_X55Y123_A2 = CLBLL_L_X34Y128_SLICE_X50Y128_AO6;
  assign CLBLL_L_X36Y123_SLICE_X55Y123_A3 = CLBLM_R_X35Y125_SLICE_X53Y125_B_XOR;
  assign CLBLL_L_X36Y123_SLICE_X55Y123_A4 = CLBLL_L_X36Y123_SLICE_X55Y123_BO6;
  assign CLBLL_L_X36Y123_SLICE_X55Y123_A5 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X36Y123_SLICE_X55Y123_A6 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLM_R_X33Y116_SLICE_X49Y116_A1 = CLBLL_L_X36Y116_SLICE_X55Y116_AO5;
  assign CLBLM_R_X33Y116_SLICE_X49Y116_A2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X33Y116_SLICE_X49Y116_A3 = CLBLM_R_X33Y116_SLICE_X48Y116_AO6;
  assign CLBLM_R_X33Y116_SLICE_X49Y116_A4 = CLBLM_R_X33Y116_SLICE_X49Y116_BO6;
  assign CLBLM_R_X33Y116_SLICE_X49Y116_A5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X33Y116_SLICE_X49Y116_A6 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLM_R_X33Y116_SLICE_X49Y116_B1 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_R_X33Y116_SLICE_X49Y116_B2 = CLBLM_R_X33Y116_SLICE_X49Y116_CO6;
  assign CLBLM_R_X33Y116_SLICE_X49Y116_B3 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLM_R_X33Y116_SLICE_X49Y116_B4 = CLBLM_R_X33Y116_SLICE_X49Y116_DO6;
  assign CLBLM_R_X33Y116_SLICE_X49Y116_B5 = CLBLM_R_X35Y120_SLICE_X53Y120_C_XOR;
  assign CLBLM_R_X33Y116_SLICE_X49Y116_B6 = CLBLL_L_X34Y128_SLICE_X50Y128_AO6;
  assign CLBLL_L_X36Y123_SLICE_X55Y123_C1 = CLBLM_R_X37Y119_SLICE_X57Y119_AO6;
  assign CLBLL_L_X36Y123_SLICE_X55Y123_C2 = CLBLM_R_X33Y123_SLICE_X48Y123_DO6;
  assign CLBLL_L_X36Y123_SLICE_X55Y123_C3 = CLBLM_R_X33Y122_SLICE_X48Y122_BO6;
  assign CLBLL_L_X36Y123_SLICE_X55Y123_C4 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X36Y123_SLICE_X55Y123_C5 = CLBLL_L_X36Y116_SLICE_X54Y116_DO6;
  assign CLBLM_R_X33Y116_SLICE_X49Y116_C1 = CLBLM_R_X33Y115_SLICE_X49Y115_AO6;
  assign CLBLM_R_X33Y116_SLICE_X49Y116_C2 = CLBLM_R_X33Y117_SLICE_X49Y117_AO6;
  assign CLBLM_R_X33Y116_SLICE_X49Y116_C3 = CLBLL_L_X34Y118_SLICE_X50Y118_BO6;
  assign CLBLM_R_X33Y116_SLICE_X49Y116_C4 = CLBLM_L_X32Y116_SLICE_X47Y116_AO6;
  assign CLBLM_R_X33Y116_SLICE_X49Y116_C5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X33Y116_SLICE_X49Y116_C6 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X36Y123_SLICE_X55Y123_C6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X35Y124_SLICE_X53Y124_D3 = 1'b1;
  assign CLBLL_L_X36Y123_SLICE_X55Y123_D1 = 1'b1;
  assign CLBLL_L_X36Y123_SLICE_X55Y123_D2 = CLBLM_R_X37Y119_SLICE_X56Y119_DO6;
  assign CLBLL_L_X36Y123_SLICE_X55Y123_D3 = CLBLL_L_X36Y118_SLICE_X55Y118_DO6;
  assign CLBLL_L_X36Y123_SLICE_X55Y123_D4 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X36Y123_SLICE_X55Y123_D5 = CLBLM_R_X35Y125_SLICE_X53Y125_B_XOR;
  assign CLBLM_R_X33Y116_SLICE_X49Y116_D1 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X33Y116_SLICE_X49Y116_D2 = CLBLL_L_X34Y117_SLICE_X50Y117_CO6;
  assign CLBLM_R_X33Y116_SLICE_X49Y116_D5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X36Y123_SLICE_X55Y123_D6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X33Y116_SLICE_X49Y116_D3 = CLBLM_R_X35Y120_SLICE_X53Y120_C_XOR;
  assign CLBLM_R_X33Y116_SLICE_X49Y116_D4 = 1'b1;
  assign CLBLM_R_X33Y116_SLICE_X49Y116_D6 = CLBLL_L_X34Y117_SLICE_X50Y117_BO6;
  assign CLBLM_R_X35Y124_SLICE_X52Y124_B1 = LIOB33_X0Y139_IOB_X0Y139_I;
  assign CLBLM_R_X35Y124_SLICE_X52Y124_B2 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X33Y116_SLICE_X48Y116_A1 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLM_R_X33Y116_SLICE_X48Y116_A2 = CLBLM_R_X35Y120_SLICE_X53Y120_C_XOR;
  assign CLBLM_R_X33Y116_SLICE_X48Y116_A3 = CLBLM_R_X35Y118_SLICE_X52Y118_C_XOR;
  assign CLBLM_R_X33Y116_SLICE_X48Y116_A4 = CLBLM_R_X33Y116_SLICE_X48Y116_BO6;
  assign CLBLM_R_X33Y116_SLICE_X48Y116_A5 = CLBLL_L_X36Y122_SLICE_X55Y122_AO6;
  assign CLBLM_R_X33Y116_SLICE_X48Y116_A6 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X35Y124_SLICE_X52Y124_B3 = 1'b1;
  assign CLBLM_R_X35Y124_SLICE_X52Y124_B4 = 1'b1;
  assign CLBLM_R_X35Y124_SLICE_X52Y124_B5 = 1'b1;
  assign CLBLM_R_X35Y124_SLICE_X52Y124_BX = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X33Y116_SLICE_X48Y116_B1 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_R_X33Y116_SLICE_X48Y116_B2 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X33Y116_SLICE_X48Y116_B3 = CLBLM_R_X35Y120_SLICE_X53Y120_C_XOR;
  assign CLBLM_R_X33Y116_SLICE_X48Y116_B4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X33Y116_SLICE_X48Y116_B5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X33Y116_SLICE_X48Y116_B6 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLM_R_X35Y124_SLICE_X52Y124_C3 = LIOB33_X0Y139_IOB_X0Y140_I;
  assign CLBLM_R_X35Y124_SLICE_X52Y124_C4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X35Y124_SLICE_X52Y124_C5 = 1'b1;
  assign CLBLM_R_X35Y124_SLICE_X52Y124_CIN = CLBLM_R_X35Y123_SLICE_X52Y123_D_CY;
  assign CLBLM_R_X33Y116_SLICE_X48Y116_C1 = CLBLL_L_X34Y128_SLICE_X50Y128_AO6;
  assign CLBLM_R_X33Y116_SLICE_X48Y116_C2 = CLBLM_R_X33Y117_SLICE_X48Y117_BO6;
  assign CLBLM_R_X33Y116_SLICE_X48Y116_C3 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_R_X33Y116_SLICE_X48Y116_C4 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLM_R_X33Y116_SLICE_X48Y116_C5 = CLBLM_R_X33Y116_SLICE_X48Y116_DO6;
  assign CLBLM_R_X33Y116_SLICE_X48Y116_C6 = CLBLM_R_X35Y120_SLICE_X53Y120_D_XOR;
  assign CLBLM_R_X35Y124_SLICE_X52Y124_CX = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X35Y124_SLICE_X52Y124_D1 = 1'b1;
  assign CLBLM_R_X35Y124_SLICE_X52Y124_D2 = 1'b1;
  assign CLBLM_R_X35Y124_SLICE_X52Y124_D3 = 1'b1;
  assign CLBLM_R_X35Y124_SLICE_X52Y124_D4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X35Y124_SLICE_X52Y124_D5 = 1'b1;
  assign CLBLM_R_X35Y124_SLICE_X52Y124_D6 = LIOB33_X0Y141_IOB_X0Y141_I;
  assign CLBLM_R_X35Y124_SLICE_X52Y124_DX = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X35Y124_SLICE_X53Y124_D6 = 1'b1;
  assign CLBLM_R_X33Y116_SLICE_X48Y116_D1 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X33Y116_SLICE_X48Y116_D2 = CLBLL_L_X34Y117_SLICE_X51Y117_CO6;
  assign CLBLM_R_X33Y116_SLICE_X48Y116_D3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X33Y116_SLICE_X48Y116_D4 = CLBLL_L_X34Y117_SLICE_X50Y117_CO6;
  assign CLBLM_R_X33Y116_SLICE_X48Y116_D5 = 1'b1;
  assign CLBLM_R_X33Y116_SLICE_X48Y116_D6 = CLBLM_R_X35Y120_SLICE_X53Y120_D_XOR;
  assign CLBLM_R_X37Y124_SLICE_X57Y124_B1 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLM_R_X37Y124_SLICE_X57Y124_B2 = LIOB33_X0Y133_IOB_X0Y133_I;
  assign CLBLM_R_X35Y124_SLICE_X53Y124_DX = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X37Y124_SLICE_X57Y124_B3 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLM_R_X37Y124_SLICE_X57Y124_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X37Y124_SLICE_X57Y124_B5 = CLBLM_R_X37Y123_SLICE_X57Y123_CO6;
  assign CLBLM_R_X37Y124_SLICE_X57Y124_B6 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign RIOB33_SING_X105Y149_IOB_X1Y149_O = CLBLL_L_X38Y126_SLICE_X59Y126_AO6;
  assign CLBLM_R_X35Y124_SLICE_X52Y124_A1 = 1'b1;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_T1 = 1'b1;
  assign CLBLM_R_X35Y124_SLICE_X52Y124_A2 = 1'b1;
  assign CLBLM_R_X35Y124_SLICE_X52Y124_A3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X35Y124_SLICE_X52Y124_A4 = LIOB33_X0Y137_IOB_X0Y138_I;
  assign CLBLM_R_X37Y124_SLICE_X57Y124_C1 = 1'b1;
  assign CLBLM_R_X35Y124_SLICE_X52Y124_A5 = 1'b1;
  assign CLBLM_R_X37Y124_SLICE_X57Y124_C2 = 1'b1;
  assign CLBLM_R_X35Y124_SLICE_X52Y124_A6 = 1'b1;
  assign CLBLM_R_X37Y124_SLICE_X57Y124_C3 = 1'b1;
  assign CLBLM_R_X37Y124_SLICE_X57Y124_C4 = 1'b1;
  assign CLBLM_R_X37Y124_SLICE_X57Y124_C5 = 1'b1;
  assign CLBLM_R_X37Y124_SLICE_X57Y124_C6 = 1'b1;
  assign CLBLM_R_X35Y124_SLICE_X52Y124_AX = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOB33_X105Y145_IOB_X1Y146_O = CLBLL_L_X36Y128_SLICE_X54Y128_AO6;
  assign RIOB33_X105Y145_IOB_X1Y145_O = CLBLL_L_X36Y129_SLICE_X54Y129_AO6;
  assign CLBLM_R_X35Y124_SLICE_X52Y124_B6 = 1'b1;
  assign CLBLM_R_X37Y124_SLICE_X57Y124_D2 = 1'b1;
  assign CLBLM_R_X37Y124_SLICE_X57Y124_D3 = 1'b1;
  assign CLBLM_R_X37Y124_SLICE_X57Y124_D4 = 1'b1;
  assign CLBLM_R_X35Y124_SLICE_X52Y124_C1 = 1'b1;
  assign CLBLM_R_X37Y124_SLICE_X57Y124_D5 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_A1 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_A2 = CLBLL_L_X38Y121_SLICE_X58Y121_AO6;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_A3 = CLBLL_L_X34Y124_SLICE_X50Y124_DO6;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_A4 = CLBLL_L_X36Y121_SLICE_X54Y121_DO6;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_A5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_A6 = CLBLM_R_X33Y124_SLICE_X48Y124_BO6;
  assign CLBLM_R_X35Y124_SLICE_X52Y124_C2 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_T1 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_B1 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_B2 = CLBLL_L_X38Y121_SLICE_X58Y121_AO6;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_B3 = CLBLL_L_X34Y126_SLICE_X50Y126_AO6;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_B4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_B5 = CLBLL_L_X34Y124_SLICE_X50Y124_DO6;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_B6 = CLBLL_L_X36Y124_SLICE_X54Y124_CO6;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_C1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_C2 = CLBLL_L_X36Y121_SLICE_X54Y121_AO5;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_C3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_C4 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_C5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_C6 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X35Y124_SLICE_X52Y124_C6 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_D1 = CLBLL_L_X36Y122_SLICE_X54Y122_AO6;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_D2 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_D3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_D4 = CLBLL_L_X36Y123_SLICE_X54Y123_AO5;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_D5 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_D6 = CLBLM_R_X35Y125_SLICE_X53Y125_D_XOR;
  assign CLBLM_R_X37Y124_SLICE_X56Y124_A1 = CLBLM_R_X37Y124_SLICE_X56Y124_BO6;
  assign CLBLM_R_X37Y124_SLICE_X56Y124_A2 = CLBLM_R_X35Y125_SLICE_X53Y125_A_XOR;
  assign CLBLM_R_X37Y124_SLICE_X56Y124_A3 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLM_R_X37Y124_SLICE_X56Y124_A4 = CLBLM_R_X35Y123_SLICE_X52Y123_A_XOR;
  assign CLBLM_R_X35Y125_SLICE_X53Y125_A1 = 1'b1;
  assign CLBLM_R_X35Y125_SLICE_X53Y125_A2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X35Y125_SLICE_X53Y125_A3 = 1'b1;
  assign CLBLM_R_X35Y125_SLICE_X53Y125_A4 = LIOB33_X0Y133_IOB_X0Y134_I;
  assign CLBLM_R_X35Y125_SLICE_X53Y125_A5 = 1'b1;
  assign CLBLM_R_X35Y125_SLICE_X53Y125_A6 = 1'b1;
  assign CLBLM_R_X37Y124_SLICE_X56Y124_A5 = CLBLL_L_X36Y122_SLICE_X55Y122_AO6;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_A1 = CLBLM_R_X35Y125_SLICE_X53Y125_C_XOR;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_A2 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_A3 = CLBLL_L_X34Y128_SLICE_X50Y128_AO6;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_A4 = CLBLL_L_X36Y123_SLICE_X55Y123_CO6;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_A5 = CLBLL_L_X36Y124_SLICE_X55Y124_CO6;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_A6 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLM_R_X35Y125_SLICE_X53Y125_AX = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X35Y125_SLICE_X53Y125_B1 = 1'b1;
  assign CLBLM_R_X33Y117_SLICE_X49Y117_A1 = CLBLM_R_X33Y117_SLICE_X49Y117_DO6;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_B1 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_B2 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_B3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_B4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_B5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_B6 = CLBLL_L_X36Y121_SLICE_X54Y121_AO5;
  assign CLBLM_R_X33Y117_SLICE_X49Y117_A2 = CLBLL_L_X34Y114_SLICE_X51Y114_CO6;
  assign CLBLM_R_X33Y117_SLICE_X49Y117_A3 = CLBLM_R_X33Y117_SLICE_X48Y117_AO6;
  assign CLBLM_R_X33Y117_SLICE_X49Y117_A4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_C1 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_C2 = CLBLL_L_X36Y118_SLICE_X55Y118_DO6;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_C3 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_C4 = CLBLL_L_X36Y122_SLICE_X54Y122_AO6;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_C5 = CLBLM_R_X35Y125_SLICE_X53Y125_C_XOR;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_C6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X33Y117_SLICE_X49Y117_B1 = CLBLM_R_X33Y117_SLICE_X49Y117_DO6;
  assign CLBLM_R_X33Y117_SLICE_X49Y117_B2 = CLBLL_L_X34Y114_SLICE_X51Y114_CO6;
  assign CLBLM_R_X33Y117_SLICE_X49Y117_B3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X33Y117_SLICE_X49Y117_B4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X33Y117_SLICE_X49Y117_B5 = CLBLL_L_X34Y117_SLICE_X51Y117_BO6;
  assign CLBLM_R_X33Y117_SLICE_X49Y117_B6 = CLBLM_R_X33Y118_SLICE_X48Y118_DO6;
  assign CLBLM_R_X33Y117_SLICE_X49Y117_C5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_D1 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_D2 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_D3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_D4 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_D5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_D6 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X33Y117_SLICE_X49Y117_C6 = CLBLM_R_X33Y119_SLICE_X49Y119_BO6;
  assign CLBLM_R_X33Y117_SLICE_X49Y117_D1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X33Y117_SLICE_X49Y117_D2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X33Y117_SLICE_X49Y117_D3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X33Y117_SLICE_X49Y117_D4 = 1'b1;
  assign CLBLM_R_X33Y117_SLICE_X49Y117_D5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X33Y117_SLICE_X49Y117_D6 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X35Y119_SLICE_X53Y119_D6 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_R_X35Y125_SLICE_X52Y125_A2 = 1'b1;
  assign CLBLM_R_X35Y125_SLICE_X52Y125_A4 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X35Y125_SLICE_X52Y125_A5 = 1'b1;
  assign CLBLM_R_X35Y125_SLICE_X52Y125_A6 = 1'b1;
  assign CLBLM_R_X35Y125_SLICE_X52Y125_AX = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X33Y117_SLICE_X48Y117_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X33Y117_SLICE_X48Y117_A2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X33Y117_SLICE_X48Y117_A3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X33Y117_SLICE_X48Y117_A4 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X33Y117_SLICE_X48Y117_A5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X33Y117_SLICE_X48Y117_A6 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X35Y125_SLICE_X52Y125_B4 = 1'b1;
  assign CLBLM_R_X35Y125_SLICE_X52Y125_B5 = 1'b1;
  assign CLBLM_R_X35Y125_SLICE_X52Y125_BX = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X33Y117_SLICE_X48Y117_B1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X33Y117_SLICE_X48Y117_B2 = CLBLM_R_X33Y117_SLICE_X49Y117_BO6;
  assign CLBLM_R_X33Y117_SLICE_X48Y117_B3 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X33Y117_SLICE_X48Y117_B4 = CLBLL_L_X34Y118_SLICE_X50Y118_BO6;
  assign CLBLM_R_X33Y117_SLICE_X48Y117_B5 = CLBLM_L_X32Y116_SLICE_X47Y116_AO6;
  assign CLBLM_R_X33Y117_SLICE_X48Y117_B6 = CLBLM_L_X32Y117_SLICE_X47Y117_AO6;
  assign CLBLM_R_X35Y125_SLICE_X52Y125_C3 = 1'b1;
  assign CLBLM_R_X35Y125_SLICE_X52Y125_C4 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X35Y125_SLICE_X52Y125_C5 = 1'b1;
  assign CLBLM_R_X35Y125_SLICE_X52Y125_CIN = CLBLM_R_X35Y124_SLICE_X52Y124_D_CY;
  assign CLBLM_R_X33Y117_SLICE_X48Y117_C1 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X33Y117_SLICE_X48Y117_C2 = CLBLL_L_X34Y118_SLICE_X50Y118_CO6;
  assign CLBLM_R_X33Y117_SLICE_X48Y117_C3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X33Y117_SLICE_X48Y117_C4 = CLBLM_R_X33Y117_SLICE_X49Y117_BO6;
  assign CLBLM_R_X33Y117_SLICE_X48Y117_C5 = CLBLM_R_X33Y117_SLICE_X48Y117_DO6;
  assign CLBLM_R_X33Y117_SLICE_X48Y117_C6 = CLBLM_L_X32Y117_SLICE_X47Y117_AO6;
  assign CLBLM_R_X35Y125_SLICE_X52Y125_CX = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X35Y125_SLICE_X52Y125_D1 = 1'b1;
  assign CLBLM_R_X35Y125_SLICE_X52Y125_D2 = 1'b1;
  assign CLBLM_R_X35Y125_SLICE_X52Y125_D3 = LIOB33_X0Y145_IOB_X0Y145_I;
  assign CLBLM_R_X35Y125_SLICE_X52Y125_D4 = 1'b1;
  assign CLBLM_R_X35Y125_SLICE_X52Y125_D5 = 1'b1;
  assign CLBLM_R_X35Y125_SLICE_X52Y125_D6 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X35Y125_SLICE_X52Y125_DX = 1'b0;
  assign CLBLM_R_X33Y117_SLICE_X48Y117_D1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X33Y117_SLICE_X48Y117_D2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X33Y117_SLICE_X48Y117_D3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X33Y117_SLICE_X48Y117_D4 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X33Y117_SLICE_X48Y117_D5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X33Y117_SLICE_X48Y117_D6 = CLBLL_L_X36Y121_SLICE_X54Y121_AO5;
  assign CLBLM_R_X35Y119_SLICE_X52Y119_A4 = 1'b1;
  assign CLBLM_R_X35Y119_SLICE_X52Y119_A5 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_C1 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X37Y124_SLICE_X56Y124_C4 = CLBLL_L_X36Y120_SLICE_X55Y120_BO6;
  assign CLBLM_R_X37Y124_SLICE_X56Y124_C5 = CLBLM_R_X37Y120_SLICE_X56Y120_BO6;
  assign CLBLM_R_X35Y119_SLICE_X52Y119_A6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_C4 = CLBLM_R_X37Y118_SLICE_X56Y118_CO6;
  assign CLBLM_R_X37Y124_SLICE_X56Y124_C6 = CLBLL_L_X38Y124_SLICE_X58Y124_AO6;
  assign CLBLM_R_X35Y114_SLICE_X53Y114_A4 = 1'b1;
  assign CLBLM_R_X35Y114_SLICE_X53Y114_A5 = 1'b1;
  assign CLBLM_R_X35Y114_SLICE_X53Y114_A6 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_C5 = 1'b1;
  assign RIOB33_X105Y147_IOB_X1Y148_O = CLBLL_L_X36Y129_SLICE_X55Y129_DO6;
  assign RIOB33_X105Y147_IOB_X1Y147_O = CLBLM_R_X37Y126_SLICE_X56Y126_BO6;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_C6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X37Y124_SLICE_X56Y124_D1 = CLBLL_L_X36Y122_SLICE_X54Y122_BO6;
  assign CLBLM_R_X37Y124_SLICE_X56Y124_D2 = CLBLM_R_X37Y121_SLICE_X56Y121_CO6;
  assign CLBLM_R_X37Y124_SLICE_X56Y124_D3 = CLBLM_R_X35Y119_SLICE_X53Y119_AO6;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_D1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X37Y124_SLICE_X56Y124_D4 = CLBLM_R_X37Y124_SLICE_X56Y124_CO6;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_D2 = 1'b1;
  assign RIOI3_X105Y121_OLOGIC_X1Y121_T1 = 1'b1;
  assign CLBLM_R_X37Y124_SLICE_X56Y124_D5 = CLBLM_R_X33Y123_SLICE_X49Y123_AO6;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_D3 = 1'b1;
  assign CLBLM_R_X37Y124_SLICE_X56Y124_D6 = CLBLM_R_X33Y121_SLICE_X48Y121_AO6;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_D5 = 1'b1;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_D = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_D6 = CLBLL_L_X38Y119_SLICE_X58Y119_AO6;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_D = LIOB33_X0Y103_IOB_X0Y103_I;
  assign RIOI3_X105Y125_OLOGIC_X1Y126_D1 = CLBLL_L_X34Y121_SLICE_X51Y121_AO6;
  assign RIOI3_X105Y125_OLOGIC_X1Y126_T1 = 1'b1;
  assign CLBLL_L_X36Y125_SLICE_X54Y125_A1 = CLBLM_R_X35Y126_SLICE_X52Y126_AO6;
  assign CLBLL_L_X36Y125_SLICE_X54Y125_A2 = CLBLM_R_X35Y126_SLICE_X53Y126_A_XOR;
  assign CLBLL_L_X36Y125_SLICE_X54Y125_A3 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLL_L_X36Y125_SLICE_X54Y125_A4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X36Y125_SLICE_X54Y125_A5 = CLBLL_L_X36Y122_SLICE_X55Y122_AO6;
  assign CLBLL_L_X36Y125_SLICE_X54Y125_A6 = CLBLM_R_X35Y124_SLICE_X52Y124_A_XOR;
  assign RIOI3_X105Y125_OLOGIC_X1Y125_D1 = CLBLM_R_X33Y121_SLICE_X48Y121_AO6;
  assign CLBLL_L_X36Y125_SLICE_X54Y125_B1 = CLBLL_L_X36Y125_SLICE_X54Y125_DO6;
  assign CLBLL_L_X36Y125_SLICE_X54Y125_B2 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLL_L_X36Y125_SLICE_X54Y125_B3 = CLBLL_L_X36Y124_SLICE_X54Y124_AO6;
  assign CLBLL_L_X36Y125_SLICE_X54Y125_B4 = CLBLL_L_X34Y128_SLICE_X50Y128_AO6;
  assign CLBLL_L_X36Y125_SLICE_X54Y125_B5 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X36Y125_SLICE_X54Y125_B6 = CLBLM_R_X35Y126_SLICE_X53Y126_A_XOR;
  assign CLBLL_L_X36Y125_SLICE_X54Y125_C1 = CLBLL_L_X34Y125_SLICE_X50Y125_AO6;
  assign CLBLL_L_X36Y125_SLICE_X54Y125_C2 = CLBLL_L_X36Y124_SLICE_X54Y124_CO6;
  assign CLBLL_L_X36Y125_SLICE_X54Y125_C3 = CLBLL_L_X36Y124_SLICE_X55Y124_BO6;
  assign CLBLL_L_X36Y125_SLICE_X54Y125_C4 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X36Y125_SLICE_X54Y125_C5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X36Y125_SLICE_X54Y125_C6 = CLBLL_L_X34Y126_SLICE_X50Y126_AO6;
  assign CLBLM_L_X32Y117_SLICE_X47Y117_A4 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign RIOI3_X105Y125_OLOGIC_X1Y125_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_D1 = CLBLM_R_X35Y115_SLICE_X53Y115_AO6;
  assign CLBLL_L_X36Y125_SLICE_X54Y125_D1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X36Y125_SLICE_X54Y125_D2 = CLBLM_R_X35Y126_SLICE_X53Y126_A_XOR;
  assign CLBLL_L_X36Y125_SLICE_X54Y125_D3 = CLBLL_L_X36Y125_SLICE_X55Y125_AO6;
  assign CLBLL_L_X36Y125_SLICE_X54Y125_D4 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X36Y125_SLICE_X54Y125_D5 = 1'b1;
  assign CLBLL_L_X36Y125_SLICE_X54Y125_D6 = CLBLL_L_X36Y123_SLICE_X54Y123_AO5;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_T1 = 1'b1;
  assign CLBLM_L_X32Y117_SLICE_X47Y117_B1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_D1 = CLBLM_R_X33Y116_SLICE_X49Y116_AO6;
  assign CLBLM_L_X32Y117_SLICE_X47Y117_B2 = 1'b1;
  assign CLBLM_R_X35Y126_SLICE_X53Y126_A1 = 1'b1;
  assign CLBLM_R_X35Y126_SLICE_X53Y126_A2 = 1'b1;
  assign CLBLL_L_X36Y125_SLICE_X55Y125_A1 = CLBLL_L_X36Y125_SLICE_X55Y125_BO5;
  assign CLBLL_L_X36Y125_SLICE_X55Y125_A2 = CLBLL_L_X36Y124_SLICE_X55Y124_DO6;
  assign CLBLL_L_X36Y125_SLICE_X55Y125_A3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X36Y125_SLICE_X55Y125_A4 = CLBLM_R_X37Y123_SLICE_X56Y123_CO6;
  assign CLBLL_L_X36Y125_SLICE_X55Y125_A5 = 1'b1;
  assign CLBLL_L_X36Y125_SLICE_X55Y125_A6 = 1'b1;
  assign CLBLM_R_X35Y126_SLICE_X53Y126_A3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X35Y126_SLICE_X53Y126_A4 = LIOB33_X0Y137_IOB_X0Y138_I;
  assign CLBLM_R_X35Y126_SLICE_X53Y126_A5 = 1'b1;
  assign CLBLL_L_X36Y125_SLICE_X55Y125_B1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X36Y125_SLICE_X55Y125_B2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X36Y125_SLICE_X55Y125_B3 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLL_L_X36Y125_SLICE_X55Y125_B4 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X36Y125_SLICE_X55Y125_B5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X36Y125_SLICE_X55Y125_B6 = 1'b1;
  assign CLBLM_R_X33Y118_SLICE_X49Y118_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X33Y118_SLICE_X49Y118_A2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X33Y118_SLICE_X49Y118_A3 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X33Y118_SLICE_X49Y118_A4 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X33Y118_SLICE_X49Y118_A5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X36Y125_SLICE_X55Y125_C3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X36Y125_SLICE_X55Y125_C4 = CLBLM_R_X37Y125_SLICE_X56Y125_BO6;
  assign CLBLM_R_X33Y118_SLICE_X49Y118_A6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X36Y125_SLICE_X55Y125_C6 = CLBLL_L_X34Y126_SLICE_X50Y126_BO6;
  assign CLBLM_R_X33Y118_SLICE_X49Y118_B1 = CLBLL_L_X34Y117_SLICE_X51Y117_DO6;
  assign CLBLM_R_X33Y118_SLICE_X49Y118_B2 = CLBLL_L_X36Y116_SLICE_X55Y116_BO6;
  assign CLBLM_R_X33Y118_SLICE_X49Y118_B3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X33Y118_SLICE_X49Y118_B4 = CLBLM_R_X37Y118_SLICE_X57Y118_AO6;
  assign CLBLM_R_X33Y118_SLICE_X49Y118_B5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X33Y118_SLICE_X49Y118_B6 = CLBLM_R_X33Y118_SLICE_X48Y118_DO6;
  assign CLBLM_R_X33Y118_SLICE_X49Y118_C1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X36Y125_SLICE_X55Y125_D1 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X36Y125_SLICE_X55Y125_D2 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X36Y125_SLICE_X55Y125_D3 = CLBLL_L_X34Y126_SLICE_X50Y126_CO6;
  assign CLBLL_L_X36Y125_SLICE_X55Y125_D4 = CLBLL_L_X36Y121_SLICE_X54Y121_AO5;
  assign CLBLL_L_X36Y125_SLICE_X55Y125_D5 = CLBLL_L_X36Y116_SLICE_X54Y116_BO5;
  assign CLBLL_L_X36Y125_SLICE_X55Y125_D6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X33Y118_SLICE_X49Y118_C2 = CLBLL_L_X34Y117_SLICE_X51Y117_BO6;
  assign CLBLM_R_X33Y118_SLICE_X49Y118_C3 = CLBLM_R_X33Y118_SLICE_X48Y118_DO6;
  assign CLBLM_R_X33Y118_SLICE_X49Y118_C4 = CLBLL_L_X34Y117_SLICE_X51Y117_DO6;
  assign CLBLM_R_X33Y118_SLICE_X49Y118_C5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X33Y118_SLICE_X49Y118_C6 = CLBLM_R_X33Y117_SLICE_X49Y117_DO6;
  assign CLBLM_L_X32Y117_SLICE_X47Y117_C2 = 1'b1;
  assign CLBLM_R_X33Y118_SLICE_X49Y118_D1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X33Y118_SLICE_X49Y118_D2 = CLBLL_L_X36Y116_SLICE_X55Y116_BO6;
  assign CLBLM_R_X33Y118_SLICE_X49Y118_D3 = CLBLM_R_X33Y118_SLICE_X48Y118_DO6;
  assign CLBLM_R_X33Y118_SLICE_X49Y118_D4 = CLBLL_L_X34Y117_SLICE_X51Y117_DO6;
  assign CLBLM_R_X33Y118_SLICE_X49Y118_D5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X33Y118_SLICE_X49Y118_D6 = CLBLM_R_X33Y117_SLICE_X49Y117_DO6;
  assign CLBLM_L_X32Y117_SLICE_X47Y117_C3 = 1'b1;
  assign CLBLL_L_X34Y114_SLICE_X50Y114_A1 = 1'b1;
  assign CLBLL_L_X34Y114_SLICE_X50Y114_A2 = 1'b1;
  assign CLBLL_L_X34Y114_SLICE_X50Y114_A3 = 1'b1;
  assign CLBLL_L_X34Y114_SLICE_X50Y114_A4 = 1'b1;
  assign CLBLL_L_X34Y114_SLICE_X50Y114_A5 = 1'b1;
  assign CLBLL_L_X34Y114_SLICE_X50Y114_A6 = 1'b1;
  assign CLBLM_R_X33Y118_SLICE_X48Y118_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X33Y118_SLICE_X48Y118_A2 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X33Y118_SLICE_X48Y118_A4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X34Y114_SLICE_X50Y114_B1 = 1'b1;
  assign CLBLL_L_X34Y114_SLICE_X50Y114_B2 = 1'b1;
  assign CLBLL_L_X34Y114_SLICE_X50Y114_B3 = 1'b1;
  assign CLBLL_L_X34Y114_SLICE_X50Y114_B4 = 1'b1;
  assign CLBLL_L_X34Y114_SLICE_X50Y114_B5 = 1'b1;
  assign CLBLL_L_X34Y114_SLICE_X50Y114_B6 = 1'b1;
  assign CLBLM_R_X33Y118_SLICE_X48Y118_A5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X33Y118_SLICE_X48Y118_B1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X33Y118_SLICE_X48Y118_B3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X33Y118_SLICE_X48Y118_B4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X33Y118_SLICE_X48Y118_B5 = CLBLM_R_X33Y118_SLICE_X48Y118_AO6;
  assign CLBLM_R_X33Y118_SLICE_X48Y118_B6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X34Y114_SLICE_X50Y114_C1 = 1'b1;
  assign CLBLL_L_X34Y114_SLICE_X50Y114_C2 = 1'b1;
  assign CLBLL_L_X34Y114_SLICE_X50Y114_C3 = 1'b1;
  assign CLBLL_L_X34Y114_SLICE_X50Y114_C4 = 1'b1;
  assign CLBLL_L_X34Y114_SLICE_X50Y114_C5 = 1'b1;
  assign CLBLL_L_X34Y114_SLICE_X50Y114_C6 = 1'b1;
  assign CLBLM_R_X33Y118_SLICE_X48Y118_C1 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X33Y118_SLICE_X48Y118_C2 = CLBLM_R_X35Y118_SLICE_X52Y118_C_XOR;
  assign CLBLM_R_X33Y118_SLICE_X48Y118_C3 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_R_X33Y118_SLICE_X48Y118_C4 = CLBLM_R_X33Y118_SLICE_X48Y118_AO5;
  assign CLBLL_L_X34Y114_SLICE_X50Y114_D1 = 1'b1;
  assign CLBLL_L_X34Y114_SLICE_X50Y114_D2 = 1'b1;
  assign CLBLL_L_X34Y114_SLICE_X50Y114_D3 = 1'b1;
  assign CLBLL_L_X34Y114_SLICE_X50Y114_D4 = 1'b1;
  assign CLBLL_L_X34Y114_SLICE_X50Y114_D5 = 1'b1;
  assign CLBLL_L_X34Y114_SLICE_X50Y114_D6 = 1'b1;
  assign CLBLM_R_X33Y118_SLICE_X48Y118_C5 = CLBLM_R_X35Y120_SLICE_X53Y120_C_XOR;
  assign CLBLM_R_X33Y118_SLICE_X48Y118_D1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X33Y118_SLICE_X48Y118_D2 = 1'b1;
  assign CLBLM_R_X33Y118_SLICE_X48Y118_D3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X33Y118_SLICE_X48Y118_D4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X33Y118_SLICE_X48Y118_D5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X33Y118_SLICE_X48Y118_D6 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X35Y114_SLICE_X52Y114_B3 = 1'b1;
  assign LIOI3_X0Y111_ILOGIC_X0Y111_D = LIOB33_X0Y111_IOB_X0Y111_I;
  assign LIOI3_X0Y133_ILOGIC_X0Y134_D = LIOB33_X0Y133_IOB_X0Y134_I;
  assign CLBLM_R_X35Y114_SLICE_X52Y114_B4 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_C6 = CLBLM_R_X37Y118_SLICE_X56Y118_BO6;
  assign LIOI3_X0Y133_ILOGIC_X0Y133_D = LIOB33_X0Y133_IOB_X0Y133_I;
  assign CLBLL_L_X34Y114_SLICE_X51Y114_A1 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X34Y114_SLICE_X51Y114_A2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X34Y114_SLICE_X51Y114_A3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X34Y114_SLICE_X51Y114_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X34Y114_SLICE_X51Y114_A5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X34Y114_SLICE_X51Y114_A6 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_D3 = CLBLM_R_X37Y119_SLICE_X57Y119_BO6;
  assign CLBLL_L_X34Y114_SLICE_X51Y114_B1 = CLBLM_R_X35Y120_SLICE_X53Y120_A_XOR;
  assign CLBLL_L_X34Y114_SLICE_X51Y114_B2 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X34Y114_SLICE_X51Y114_B3 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X34Y114_SLICE_X51Y114_B4 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLL_L_X34Y114_SLICE_X51Y114_B5 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X34Y114_SLICE_X51Y114_B6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_D4 = CLBLL_L_X38Y118_SLICE_X58Y118_AO5;
  assign CLBLL_L_X34Y114_SLICE_X51Y114_C1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X34Y114_SLICE_X51Y114_C2 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X34Y114_SLICE_X51Y114_C3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X34Y114_SLICE_X51Y114_C4 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X34Y114_SLICE_X51Y114_C5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X34Y114_SLICE_X51Y114_C6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X35Y114_SLICE_X52Y114_C1 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_D6 = CLBLL_L_X36Y118_SLICE_X55Y118_AO5;
  assign CLBLM_R_X35Y114_SLICE_X52Y114_C2 = 1'b1;
  assign CLBLL_L_X34Y114_SLICE_X51Y114_D1 = 1'b1;
  assign CLBLL_L_X34Y114_SLICE_X51Y114_D2 = 1'b1;
  assign CLBLL_L_X34Y114_SLICE_X51Y114_D3 = 1'b1;
  assign CLBLL_L_X34Y114_SLICE_X51Y114_D4 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X34Y114_SLICE_X51Y114_D5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X34Y114_SLICE_X51Y114_D6 = 1'b1;
  assign CLBLM_R_X35Y114_SLICE_X52Y114_C3 = 1'b1;
  assign CLBLL_L_X36Y126_SLICE_X54Y126_A1 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLL_L_X36Y126_SLICE_X54Y126_A2 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X36Y126_SLICE_X54Y126_A3 = CLBLL_L_X34Y128_SLICE_X50Y128_AO6;
  assign CLBLL_L_X36Y126_SLICE_X54Y126_A4 = CLBLL_L_X36Y124_SLICE_X54Y124_BO6;
  assign CLBLL_L_X36Y126_SLICE_X54Y126_A5 = CLBLL_L_X36Y126_SLICE_X54Y126_CO6;
  assign CLBLL_L_X36Y126_SLICE_X54Y126_A6 = CLBLM_R_X35Y126_SLICE_X53Y126_B_XOR;
  assign CLBLL_L_X36Y126_SLICE_X54Y126_B1 = CLBLL_L_X36Y126_SLICE_X54Y126_DO6;
  assign CLBLL_L_X36Y126_SLICE_X54Y126_B2 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X36Y126_SLICE_X54Y126_B3 = CLBLL_L_X34Y128_SLICE_X50Y128_AO6;
  assign CLBLL_L_X36Y126_SLICE_X54Y126_B4 = CLBLM_R_X35Y126_SLICE_X53Y126_C_XOR;
  assign CLBLL_L_X36Y126_SLICE_X54Y126_B5 = CLBLL_L_X36Y125_SLICE_X54Y125_CO6;
  assign CLBLL_L_X36Y126_SLICE_X54Y126_B6 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLL_L_X36Y126_SLICE_X54Y126_C1 = 1'b1;
  assign CLBLL_L_X36Y126_SLICE_X54Y126_C2 = CLBLM_R_X37Y126_SLICE_X56Y126_AO6;
  assign CLBLL_L_X36Y126_SLICE_X54Y126_C3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X36Y126_SLICE_X54Y126_C4 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X36Y126_SLICE_X54Y126_C5 = CLBLL_L_X36Y125_SLICE_X55Y125_AO6;
  assign CLBLL_L_X36Y126_SLICE_X54Y126_C6 = CLBLM_R_X35Y126_SLICE_X53Y126_B_XOR;
  assign CLBLL_L_X36Y126_SLICE_X54Y126_D1 = CLBLL_L_X36Y125_SLICE_X55Y125_AO5;
  assign CLBLL_L_X36Y126_SLICE_X54Y126_D2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X36Y126_SLICE_X54Y126_D3 = CLBLM_R_X37Y126_SLICE_X56Y126_AO6;
  assign CLBLL_L_X36Y126_SLICE_X54Y126_D4 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X36Y126_SLICE_X54Y126_D5 = 1'b1;
  assign CLBLL_L_X36Y126_SLICE_X54Y126_D6 = CLBLM_R_X35Y126_SLICE_X53Y126_C_XOR;
  assign CLBLM_R_X33Y123_SLICE_X49Y123_C3 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X36Y126_SLICE_X55Y126_A1 = CLBLL_L_X36Y126_SLICE_X55Y126_DO6;
  assign CLBLL_L_X36Y126_SLICE_X55Y126_A2 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X36Y126_SLICE_X55Y126_A3 = CLBLM_R_X35Y126_SLICE_X53Y126_D_XOR;
  assign CLBLL_L_X36Y126_SLICE_X55Y126_A4 = CLBLL_L_X34Y128_SLICE_X50Y128_AO6;
  assign CLBLL_L_X36Y126_SLICE_X55Y126_A5 = CLBLL_L_X36Y125_SLICE_X55Y125_CO6;
  assign CLBLL_L_X36Y126_SLICE_X55Y126_A6 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLM_R_X33Y123_SLICE_X49Y123_C4 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLM_R_X35Y127_SLICE_X53Y127_A1 = 1'b1;
  assign CLBLM_R_X35Y127_SLICE_X53Y127_A2 = 1'b1;
  assign CLBLL_L_X36Y126_SLICE_X55Y126_B1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X36Y126_SLICE_X55Y126_B2 = CLBLL_L_X34Y126_SLICE_X50Y126_BO6;
  assign CLBLL_L_X36Y126_SLICE_X55Y126_B3 = CLBLL_L_X34Y126_SLICE_X50Y126_CO6;
  assign CLBLL_L_X36Y126_SLICE_X55Y126_B4 = CLBLM_R_X37Y127_SLICE_X56Y127_AO6;
  assign CLBLL_L_X36Y126_SLICE_X55Y126_B5 = CLBLM_R_X37Y125_SLICE_X56Y125_BO6;
  assign CLBLL_L_X36Y126_SLICE_X55Y126_B6 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X35Y127_SLICE_X53Y127_B1 = 1'b1;
  assign CLBLM_R_X35Y127_SLICE_X53Y127_B2 = LIOB33_X0Y143_IOB_X0Y143_I;
  assign CLBLM_R_X33Y119_SLICE_X49Y119_A1 = CLBLM_R_X33Y119_SLICE_X49Y119_BO6;
  assign CLBLL_L_X36Y126_SLICE_X55Y126_C1 = CLBLL_L_X34Y127_SLICE_X50Y127_AO6;
  assign CLBLL_L_X36Y126_SLICE_X55Y126_C2 = CLBLL_L_X36Y125_SLICE_X55Y125_DO6;
  assign CLBLL_L_X36Y126_SLICE_X55Y126_C3 = CLBLL_L_X36Y122_SLICE_X55Y122_AO5;
  assign CLBLL_L_X36Y126_SLICE_X55Y126_C4 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X36Y126_SLICE_X55Y126_C5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X36Y126_SLICE_X55Y126_C6 = CLBLM_R_X37Y127_SLICE_X56Y127_AO6;
  assign CLBLM_R_X33Y119_SLICE_X49Y119_A2 = CLBLL_L_X34Y119_SLICE_X50Y119_CO6;
  assign CLBLM_R_X33Y119_SLICE_X49Y119_A3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X33Y119_SLICE_X49Y119_A4 = CLBLM_R_X33Y118_SLICE_X48Y118_BO6;
  assign CLBLM_R_X33Y119_SLICE_X49Y119_A5 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X33Y119_SLICE_X49Y119_A6 = CLBLM_R_X33Y118_SLICE_X49Y118_CO6;
  assign CLBLM_R_X33Y119_SLICE_X49Y119_B1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X33Y119_SLICE_X49Y119_B2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X36Y126_SLICE_X55Y126_D1 = CLBLL_L_X36Y125_SLICE_X55Y125_AO5;
  assign CLBLL_L_X36Y126_SLICE_X55Y126_D2 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X36Y126_SLICE_X55Y126_D3 = 1'b1;
  assign CLBLL_L_X36Y126_SLICE_X55Y126_D4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X36Y126_SLICE_X55Y126_D5 = CLBLM_R_X37Y126_SLICE_X56Y126_AO5;
  assign CLBLL_L_X36Y126_SLICE_X55Y126_D6 = CLBLM_R_X35Y126_SLICE_X53Y126_D_XOR;
  assign CLBLM_R_X33Y119_SLICE_X49Y119_B4 = CLBLL_L_X36Y121_SLICE_X54Y121_AO5;
  assign CLBLM_R_X33Y119_SLICE_X49Y119_B5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X33Y119_SLICE_X49Y119_C1 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X33Y119_SLICE_X49Y119_C2 = CLBLL_L_X34Y119_SLICE_X50Y119_CO6;
  assign CLBLM_R_X33Y119_SLICE_X49Y119_C3 = CLBLM_R_X33Y118_SLICE_X49Y118_DO6;
  assign CLBLM_R_X33Y119_SLICE_X49Y119_C4 = CLBLL_L_X34Y119_SLICE_X51Y119_DO6;
  assign CLBLM_R_X33Y119_SLICE_X49Y119_C5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X33Y119_SLICE_X49Y119_C6 = CLBLM_R_X33Y118_SLICE_X48Y118_BO6;
  assign CLBLM_R_X35Y127_SLICE_X52Y127_A1 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X35Y127_SLICE_X52Y127_A2 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X33Y119_SLICE_X49Y119_D1 = 1'b1;
  assign CLBLM_R_X33Y119_SLICE_X49Y119_D2 = 1'b1;
  assign CLBLL_L_X34Y115_SLICE_X50Y115_A1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X34Y115_SLICE_X50Y115_A2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X34Y115_SLICE_X50Y115_A3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X34Y115_SLICE_X50Y115_A4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X34Y115_SLICE_X50Y115_A5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X34Y115_SLICE_X50Y115_A6 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X33Y119_SLICE_X49Y119_D3 = 1'b1;
  assign CLBLM_R_X33Y119_SLICE_X49Y119_D4 = 1'b1;
  assign CLBLM_R_X33Y119_SLICE_X49Y119_D5 = 1'b1;
  assign CLBLL_L_X34Y115_SLICE_X50Y115_B1 = CLBLM_R_X33Y117_SLICE_X48Y117_CO6;
  assign CLBLL_L_X34Y115_SLICE_X50Y115_B2 = CLBLL_L_X34Y128_SLICE_X50Y128_AO6;
  assign CLBLL_L_X34Y115_SLICE_X50Y115_B3 = CLBLM_R_X35Y121_SLICE_X53Y121_A_XOR;
  assign CLBLL_L_X34Y115_SLICE_X50Y115_B4 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLL_L_X34Y115_SLICE_X50Y115_B5 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X34Y115_SLICE_X50Y115_B6 = CLBLL_L_X34Y116_SLICE_X50Y116_AO5;
  assign CLBLM_R_X33Y119_SLICE_X48Y119_A1 = 1'b1;
  assign CLBLM_R_X33Y119_SLICE_X48Y119_A2 = 1'b1;
  assign CLBLM_R_X33Y119_SLICE_X48Y119_A3 = 1'b1;
  assign CLBLL_L_X34Y115_SLICE_X50Y115_C1 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X34Y115_SLICE_X50Y115_C2 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X34Y115_SLICE_X50Y115_C3 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X34Y115_SLICE_X50Y115_C4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X34Y115_SLICE_X50Y115_C5 = CLBLM_R_X35Y121_SLICE_X53Y121_A_XOR;
  assign CLBLL_L_X34Y115_SLICE_X50Y115_C6 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLM_R_X33Y119_SLICE_X48Y119_B1 = 1'b1;
  assign CLBLM_R_X33Y119_SLICE_X48Y119_B2 = 1'b1;
  assign CLBLM_R_X33Y119_SLICE_X48Y119_B3 = 1'b1;
  assign CLBLM_R_X33Y119_SLICE_X48Y119_B4 = 1'b1;
  assign CLBLM_R_X33Y119_SLICE_X48Y119_B5 = 1'b1;
  assign CLBLM_R_X33Y119_SLICE_X48Y119_B6 = 1'b1;
  assign CLBLL_L_X34Y115_SLICE_X50Y115_D1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X34Y115_SLICE_X50Y115_D2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X34Y115_SLICE_X50Y115_D3 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X34Y115_SLICE_X50Y115_D4 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X34Y115_SLICE_X50Y115_D5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X34Y115_SLICE_X50Y115_D6 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X33Y119_SLICE_X48Y119_C1 = 1'b1;
  assign CLBLM_R_X33Y119_SLICE_X48Y119_C2 = 1'b1;
  assign CLBLM_R_X33Y119_SLICE_X48Y119_C3 = 1'b1;
  assign CLBLM_R_X33Y119_SLICE_X48Y119_C4 = 1'b1;
  assign CLBLM_R_X33Y119_SLICE_X48Y119_C5 = 1'b1;
  assign CLBLM_R_X33Y119_SLICE_X48Y119_C6 = 1'b1;
  assign CLBLM_R_X33Y119_SLICE_X48Y119_D1 = 1'b1;
  assign CLBLM_R_X33Y119_SLICE_X48Y119_D2 = 1'b1;
  assign CLBLM_R_X33Y119_SLICE_X48Y119_D3 = 1'b1;
  assign CLBLM_R_X33Y119_SLICE_X48Y119_D4 = 1'b1;
  assign CLBLM_R_X33Y119_SLICE_X48Y119_D5 = 1'b1;
  assign CLBLM_R_X33Y119_SLICE_X48Y119_D6 = 1'b1;
  assign CLBLL_L_X34Y115_SLICE_X51Y115_A1 = CLBLM_R_X35Y115_SLICE_X52Y115_AO5;
  assign CLBLL_L_X34Y115_SLICE_X51Y115_A2 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X34Y115_SLICE_X51Y115_A3 = CLBLL_L_X34Y114_SLICE_X51Y114_BO6;
  assign CLBLL_L_X34Y115_SLICE_X51Y115_A4 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLL_L_X34Y115_SLICE_X51Y115_A5 = CLBLL_L_X34Y118_SLICE_X51Y118_DO6;
  assign CLBLL_L_X34Y115_SLICE_X51Y115_A6 = CLBLL_L_X34Y116_SLICE_X50Y116_BO6;
  assign CLBLL_L_X34Y115_SLICE_X51Y115_B1 = CLBLL_L_X34Y115_SLICE_X50Y115_CO6;
  assign CLBLL_L_X34Y115_SLICE_X51Y115_B2 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X34Y115_SLICE_X51Y115_B3 = CLBLL_L_X36Y122_SLICE_X55Y122_AO6;
  assign CLBLL_L_X34Y115_SLICE_X51Y115_B4 = CLBLM_R_X35Y121_SLICE_X53Y121_A_XOR;
  assign CLBLL_L_X34Y115_SLICE_X51Y115_B5 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLL_L_X34Y115_SLICE_X51Y115_B6 = CLBLM_R_X35Y119_SLICE_X52Y119_A_XOR;
  assign CLBLL_L_X34Y115_SLICE_X51Y115_C1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X34Y115_SLICE_X51Y115_C2 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLL_L_X34Y115_SLICE_X51Y115_C3 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLL_L_X34Y115_SLICE_X51Y115_C4 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X34Y115_SLICE_X51Y115_C5 = CLBLL_L_X34Y115_SLICE_X51Y115_DO6;
  assign CLBLL_L_X34Y115_SLICE_X51Y115_C6 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X34Y115_SLICE_X51Y115_D1 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X34Y115_SLICE_X51Y115_D2 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X34Y115_SLICE_X51Y115_D3 = CLBLM_R_X35Y121_SLICE_X53Y121_A_XOR;
  assign CLBLL_L_X34Y115_SLICE_X51Y115_D4 = CLBLM_R_X35Y119_SLICE_X52Y119_A_XOR;
  assign CLBLL_L_X34Y115_SLICE_X51Y115_D5 = CLBLL_L_X34Y114_SLICE_X51Y114_DO6;
  assign CLBLL_L_X34Y115_SLICE_X51Y115_D6 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign RIOB33_X105Y139_IOB_X1Y140_O = CLBLL_L_X38Y126_SLICE_X58Y126_AO6;
  assign RIOB33_X105Y139_IOB_X1Y139_O = CLBLM_R_X37Y125_SLICE_X57Y125_AO6;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_A1 = CLBLL_L_X36Y116_SLICE_X55Y116_AO5;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_A2 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_A3 = CLBLL_L_X36Y125_SLICE_X54Y125_BO6;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_A4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_A5 = CLBLL_L_X36Y125_SLICE_X54Y125_AO6;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_A6 = LIOB33_X0Y137_IOB_X0Y138_I;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_B1 = LIOB33_X0Y139_IOB_X0Y139_I;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_B2 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_B3 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_B4 = CLBLL_L_X36Y116_SLICE_X55Y116_AO5;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_B5 = CLBLL_L_X36Y126_SLICE_X54Y126_AO6;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_B6 = CLBLL_L_X36Y127_SLICE_X54Y127_CO6;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_C1 = CLBLL_L_X36Y122_SLICE_X55Y122_AO6;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_C2 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_C3 = CLBLM_R_X35Y124_SLICE_X52Y124_B_XOR;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_C4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_C5 = CLBLL_L_X36Y127_SLICE_X54Y127_DO6;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_C6 = CLBLM_R_X35Y126_SLICE_X53Y126_B_XOR;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_D1 = CLBLM_R_X35Y126_SLICE_X53Y126_B_XOR;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_D2 = LIOB33_X0Y139_IOB_X0Y139_I;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_D3 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_D4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_D5 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_D6 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_A2 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_A3 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_A4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_A5 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_A6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X35Y128_SLICE_X53Y128_A1 = CLBLM_R_X35Y127_SLICE_X53Y127_C_XOR;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_B1 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_B2 = CLBLM_R_X35Y127_SLICE_X53Y127_A_XOR;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_B3 = CLBLL_L_X36Y126_SLICE_X55Y126_BO6;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_B4 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_B5 = CLBLL_L_X36Y128_SLICE_X55Y128_DO6;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_B6 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X35Y128_SLICE_X53Y128_A2 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X35Y128_SLICE_X53Y128_A3 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_R_X35Y128_SLICE_X53Y128_A4 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_C1 = CLBLL_L_X34Y127_SLICE_X50Y127_AO6;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_C2 = CLBLL_L_X34Y126_SLICE_X50Y126_CO6;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_C3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_C4 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_C5 = CLBLL_L_X36Y127_SLICE_X55Y127_DO6;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_C6 = CLBLM_R_X37Y127_SLICE_X56Y127_AO6;
  assign CLBLM_R_X35Y128_SLICE_X53Y128_B1 = CLBLM_R_X35Y128_SLICE_X53Y128_DO6;
  assign CLBLM_R_X35Y128_SLICE_X53Y128_B2 = CLBLM_R_X35Y125_SLICE_X52Y125_A_XOR;
  assign CLBLM_R_X35Y128_SLICE_X53Y128_B3 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_R_X35Y128_SLICE_X53Y128_B4 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X33Y123_SLICE_X48Y123_D5 = CLBLM_R_X33Y124_SLICE_X48Y124_AO5;
  assign CLBLM_R_X35Y128_SLICE_X53Y128_B5 = CLBLM_R_X35Y127_SLICE_X53Y127_A_XOR;
  assign CLBLM_R_X35Y128_SLICE_X53Y128_B6 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_D1 = 1'b1;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_D2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_D3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_D4 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_D5 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_D6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X38Y118_SLICE_X59Y118_D6 = 1'b1;
  assign CLBLM_R_X33Y123_SLICE_X48Y123_D6 = CLBLL_L_X34Y123_SLICE_X50Y123_AO5;
  assign CLBLM_R_X35Y128_SLICE_X53Y128_D1 = 1'b1;
  assign CLBLM_R_X35Y128_SLICE_X53Y128_D2 = LIOB33_X0Y141_IOB_X0Y142_I;
  assign CLBLM_R_X35Y128_SLICE_X53Y128_D3 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X35Y128_SLICE_X53Y128_D4 = 1'b1;
  assign CLBLM_R_X35Y128_SLICE_X53Y128_D5 = 1'b1;
  assign CLBLM_R_X35Y128_SLICE_X53Y128_D6 = 1'b1;
  assign RIOI3_X105Y127_OLOGIC_X1Y128_T1 = 1'b1;
  assign CLBLL_L_X34Y116_SLICE_X50Y116_A1 = CLBLL_L_X34Y117_SLICE_X51Y117_CO6;
  assign CLBLL_L_X34Y116_SLICE_X50Y116_A2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X34Y116_SLICE_X50Y116_A3 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X34Y116_SLICE_X50Y116_A4 = CLBLL_L_X34Y116_SLICE_X51Y116_DO6;
  assign CLBLL_L_X34Y116_SLICE_X50Y116_A5 = CLBLM_R_X35Y121_SLICE_X53Y121_A_XOR;
  assign CLBLL_L_X34Y116_SLICE_X50Y116_A6 = 1'b1;
  assign CLBLM_R_X35Y128_SLICE_X52Y128_A1 = LIOB33_X0Y143_IOB_X0Y144_I;
  assign CLBLM_R_X35Y128_SLICE_X52Y128_A2 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X34Y116_SLICE_X50Y116_B1 = CLBLL_L_X34Y117_SLICE_X50Y117_AO6;
  assign CLBLL_L_X34Y116_SLICE_X50Y116_B2 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLL_L_X34Y116_SLICE_X50Y116_B3 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLL_L_X34Y116_SLICE_X50Y116_B4 = CLBLL_L_X34Y117_SLICE_X51Y117_AO6;
  assign CLBLL_L_X34Y116_SLICE_X50Y116_B5 = CLBLL_L_X34Y116_SLICE_X50Y116_AO6;
  assign CLBLL_L_X34Y116_SLICE_X50Y116_B6 = CLBLL_L_X34Y116_SLICE_X50Y116_CO6;
  assign CLBLM_R_X35Y128_SLICE_X52Y128_B1 = CLBLM_R_X35Y127_SLICE_X53Y127_D_XOR;
  assign CLBLM_R_X35Y128_SLICE_X52Y128_B2 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X34Y116_SLICE_X50Y116_C1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X34Y116_SLICE_X50Y116_C2 = CLBLL_L_X34Y116_SLICE_X51Y116_AO5;
  assign CLBLL_L_X34Y116_SLICE_X50Y116_C3 = CLBLL_L_X34Y117_SLICE_X50Y117_DO6;
  assign CLBLL_L_X34Y116_SLICE_X50Y116_C4 = CLBLL_L_X34Y115_SLICE_X50Y115_AO6;
  assign CLBLL_L_X34Y116_SLICE_X50Y116_C5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X34Y116_SLICE_X50Y116_C6 = CLBLL_L_X34Y114_SLICE_X51Y114_CO6;
  assign CLBLM_R_X35Y128_SLICE_X52Y128_C1 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X35Y128_SLICE_X52Y128_C2 = LIOB33_X0Y141_IOB_X0Y142_I;
  assign CLBLM_R_X35Y128_SLICE_X52Y128_C3 = CLBLM_R_X35Y128_SLICE_X53Y128_BO6;
  assign CLBLM_R_X35Y128_SLICE_X52Y128_C4 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLM_R_X35Y128_SLICE_X52Y128_C5 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X35Y128_SLICE_X52Y128_C6 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_D1 = CLBLL_L_X36Y122_SLICE_X55Y122_BO6;
  assign CLBLL_L_X34Y116_SLICE_X50Y116_D1 = 1'b1;
  assign CLBLL_L_X34Y116_SLICE_X50Y116_D2 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X34Y116_SLICE_X50Y116_D3 = 1'b1;
  assign CLBLL_L_X34Y116_SLICE_X50Y116_D4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X34Y116_SLICE_X50Y116_D5 = 1'b1;
  assign CLBLL_L_X34Y116_SLICE_X50Y116_D6 = CLBLL_L_X34Y117_SLICE_X50Y117_AO6;
  assign CLBLM_R_X33Y118_SLICE_X48Y118_A3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X35Y128_SLICE_X52Y128_D1 = 1'b1;
  assign CLBLM_R_X35Y128_SLICE_X52Y128_D2 = 1'b1;
  assign CLBLM_R_X35Y128_SLICE_X52Y128_D3 = 1'b1;
  assign CLBLM_R_X35Y128_SLICE_X52Y128_D4 = 1'b1;
  assign CLBLM_R_X35Y128_SLICE_X52Y128_D5 = 1'b1;
  assign CLBLM_R_X35Y128_SLICE_X52Y128_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_D1 = CLBLL_L_X36Y121_SLICE_X55Y121_BO6;
  assign CLBLM_R_X33Y118_SLICE_X48Y118_A6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_T1 = 1'b1;
  assign CLBLL_L_X34Y116_SLICE_X51Y116_A1 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X34Y116_SLICE_X51Y116_A2 = CLBLL_L_X34Y118_SLICE_X51Y118_CO6;
  assign CLBLL_L_X34Y116_SLICE_X51Y116_A3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X34Y116_SLICE_X51Y116_A4 = CLBLM_R_X35Y121_SLICE_X53Y121_B_XOR;
  assign CLBLL_L_X34Y116_SLICE_X51Y116_A5 = CLBLL_L_X34Y116_SLICE_X51Y116_DO6;
  assign CLBLL_L_X34Y116_SLICE_X51Y116_A6 = 1'b1;
  assign CLBLL_L_X34Y116_SLICE_X51Y116_B1 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X34Y116_SLICE_X51Y116_B2 = CLBLL_L_X36Y116_SLICE_X54Y116_BO5;
  assign CLBLL_L_X34Y116_SLICE_X51Y116_B3 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X34Y116_SLICE_X51Y116_B4 = CLBLL_L_X36Y121_SLICE_X54Y121_AO5;
  assign CLBLL_L_X34Y116_SLICE_X51Y116_B5 = CLBLM_R_X33Y117_SLICE_X49Y117_AO6;
  assign CLBLL_L_X34Y116_SLICE_X51Y116_B6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X34Y116_SLICE_X51Y116_C1 = CLBLL_L_X34Y116_SLICE_X51Y116_AO6;
  assign CLBLL_L_X34Y116_SLICE_X51Y116_C2 = CLBLL_L_X34Y128_SLICE_X50Y128_AO6;
  assign CLBLL_L_X34Y116_SLICE_X51Y116_C3 = CLBLM_R_X33Y117_SLICE_X49Y117_CO6;
  assign CLBLL_L_X34Y116_SLICE_X51Y116_C4 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X34Y116_SLICE_X51Y116_C5 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLL_L_X34Y116_SLICE_X51Y116_C6 = CLBLM_R_X35Y121_SLICE_X53Y121_B_XOR;
  assign CLBLM_R_X33Y118_SLICE_X48Y118_B2 = CLBLL_L_X36Y121_SLICE_X54Y121_AO5;
  assign CLBLL_L_X34Y116_SLICE_X51Y116_D1 = CLBLM_R_X35Y116_SLICE_X53Y116_AO6;
  assign CLBLL_L_X34Y116_SLICE_X51Y116_D2 = CLBLL_L_X34Y115_SLICE_X50Y115_DO6;
  assign CLBLL_L_X34Y116_SLICE_X51Y116_D3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X34Y116_SLICE_X51Y116_D4 = CLBLL_L_X34Y114_SLICE_X51Y114_AO6;
  assign CLBLL_L_X34Y116_SLICE_X51Y116_D5 = CLBLM_R_X35Y117_SLICE_X52Y117_AO6;
  assign CLBLL_L_X34Y116_SLICE_X51Y116_D6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_C3 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign LIOI3_X0Y145_ILOGIC_X0Y146_D = LIOB33_X0Y145_IOB_X0Y146_I;
  assign LIOI3_X0Y145_ILOGIC_X0Y145_D = LIOB33_X0Y145_IOB_X0Y145_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y116_D = LIOB33_X0Y115_IOB_X0Y116_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_D = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X33Y118_SLICE_X48Y118_C6 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y115_D = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X36Y128_SLICE_X54Y128_A1 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLL_L_X36Y128_SLICE_X54Y128_A2 = CLBLM_R_X35Y127_SLICE_X53Y127_B_XOR;
  assign CLBLL_L_X36Y128_SLICE_X54Y128_A3 = CLBLM_R_X35Y127_SLICE_X52Y127_AO6;
  assign CLBLL_L_X36Y128_SLICE_X54Y128_A4 = CLBLL_L_X36Y128_SLICE_X54Y128_BO6;
  assign CLBLL_L_X36Y128_SLICE_X54Y128_A5 = CLBLL_L_X34Y128_SLICE_X50Y128_AO6;
  assign CLBLL_L_X36Y128_SLICE_X54Y128_A6 = CLBLL_L_X36Y126_SLICE_X55Y126_CO6;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_D = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X36Y128_SLICE_X54Y128_B1 = CLBLL_L_X36Y116_SLICE_X55Y116_AO6;
  assign CLBLL_L_X36Y128_SLICE_X54Y128_B2 = CLBLM_R_X35Y127_SLICE_X53Y127_B_XOR;
  assign CLBLL_L_X36Y128_SLICE_X54Y128_B3 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X36Y128_SLICE_X54Y128_B4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X36Y128_SLICE_X54Y128_B5 = CLBLL_L_X36Y127_SLICE_X55Y127_AO6;
  assign CLBLL_L_X36Y128_SLICE_X54Y128_B6 = CLBLM_R_X37Y127_SLICE_X56Y127_BO6;
  assign CLBLL_L_X36Y128_SLICE_X54Y128_C1 = CLBLM_R_X35Y127_SLICE_X53Y127_B_XOR;
  assign CLBLL_L_X36Y128_SLICE_X54Y128_C2 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X36Y128_SLICE_X54Y128_C3 = CLBLL_L_X34Y128_SLICE_X50Y128_AO6;
  assign CLBLL_L_X36Y128_SLICE_X54Y128_C4 = CLBLL_L_X36Y127_SLICE_X55Y127_CO6;
  assign CLBLL_L_X36Y128_SLICE_X54Y128_C5 = CLBLL_L_X36Y128_SLICE_X54Y128_DO6;
  assign CLBLL_L_X36Y128_SLICE_X54Y128_C6 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLL_L_X36Y128_SLICE_X54Y128_D1 = CLBLL_L_X36Y127_SLICE_X55Y127_AO6;
  assign CLBLL_L_X36Y128_SLICE_X54Y128_D2 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X36Y128_SLICE_X54Y128_D3 = CLBLM_R_X37Y127_SLICE_X56Y127_BO6;
  assign CLBLL_L_X36Y128_SLICE_X54Y128_D4 = CLBLM_R_X35Y127_SLICE_X53Y127_B_XOR;
  assign CLBLL_L_X36Y128_SLICE_X54Y128_D5 = 1'b1;
  assign CLBLL_L_X36Y128_SLICE_X54Y128_D6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X35Y125_SLICE_X53Y125_B2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X35Y125_SLICE_X53Y125_B3 = 1'b1;
  assign CLBLM_R_X35Y125_SLICE_X53Y125_B4 = 1'b1;
  assign CLBLM_R_X35Y125_SLICE_X53Y125_B5 = 1'b1;
  assign CLBLM_R_X35Y125_SLICE_X53Y125_B6 = LIOB33_X0Y135_IOB_X0Y135_I;
  assign CLBLL_L_X36Y128_SLICE_X55Y128_A1 = CLBLL_L_X36Y128_SLICE_X55Y128_DO6;
  assign CLBLL_L_X36Y128_SLICE_X55Y128_A2 = CLBLL_L_X36Y126_SLICE_X55Y126_BO6;
  assign CLBLL_L_X36Y128_SLICE_X55Y128_A3 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X36Y128_SLICE_X55Y128_A4 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLL_L_X36Y128_SLICE_X55Y128_A5 = CLBLL_L_X34Y128_SLICE_X50Y128_AO6;
  assign CLBLL_L_X36Y128_SLICE_X55Y128_A6 = CLBLM_R_X35Y127_SLICE_X53Y127_A_XOR;
  assign CLBLM_R_X35Y125_SLICE_X53Y125_BX = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X36Y128_SLICE_X55Y128_B1 = CLBLM_R_X35Y129_SLICE_X52Y129_AO6;
  assign CLBLL_L_X36Y128_SLICE_X55Y128_B2 = CLBLM_R_X35Y128_SLICE_X52Y128_CO6;
  assign CLBLL_L_X36Y128_SLICE_X55Y128_B3 = CLBLL_L_X36Y126_SLICE_X55Y126_AO6;
  assign CLBLL_L_X36Y128_SLICE_X55Y128_B4 = CLBLL_L_X36Y128_SLICE_X54Y128_CO6;
  assign CLBLL_L_X36Y128_SLICE_X55Y128_B5 = CLBLL_L_X36Y128_SLICE_X55Y128_AO6;
  assign CLBLL_L_X36Y128_SLICE_X55Y128_B6 = CLBLM_R_X35Y127_SLICE_X52Y127_AO6;
  assign CLBLM_R_X35Y129_SLICE_X53Y129_A1 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLM_R_X35Y129_SLICE_X53Y129_A2 = CLBLM_R_X35Y125_SLICE_X52Y125_D_XOR;
  assign CLBLM_R_X35Y125_SLICE_X53Y125_C1 = 1'b1;
  assign CLBLL_L_X36Y128_SLICE_X55Y128_C1 = CLBLM_R_X35Y129_SLICE_X53Y129_AO6;
  assign CLBLL_L_X36Y128_SLICE_X55Y128_C2 = CLBLL_L_X36Y128_SLICE_X54Y128_CO6;
  assign CLBLL_L_X36Y128_SLICE_X55Y128_C3 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X36Y128_SLICE_X55Y128_C4 = CLBLM_R_X35Y128_SLICE_X52Y128_BO6;
  assign CLBLL_L_X36Y128_SLICE_X55Y128_C5 = CLBLM_R_X35Y127_SLICE_X52Y127_AO6;
  assign CLBLL_L_X36Y128_SLICE_X55Y128_C6 = CLBLM_R_X35Y129_SLICE_X53Y129_BO6;
  assign CLBLM_R_X35Y125_SLICE_X53Y125_C2 = 1'b1;
  assign CLBLM_R_X35Y129_SLICE_X53Y129_A6 = CLBLM_R_X35Y129_SLICE_X53Y129_CO6;
  assign CLBLM_R_X35Y125_SLICE_X53Y125_C3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X33Y121_SLICE_X49Y121_A1 = CLBLM_R_X33Y118_SLICE_X49Y118_DO6;
  assign CLBLM_R_X33Y121_SLICE_X49Y121_A2 = CLBLL_L_X34Y120_SLICE_X50Y120_CO6;
  assign CLBLM_R_X33Y121_SLICE_X49Y121_A3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X33Y121_SLICE_X49Y121_A4 = CLBLM_R_X33Y121_SLICE_X49Y121_BO6;
  assign CLBLM_R_X33Y121_SLICE_X49Y121_A5 = CLBLL_L_X34Y119_SLICE_X51Y119_DO6;
  assign CLBLL_L_X36Y128_SLICE_X55Y128_D1 = CLBLL_L_X36Y127_SLICE_X55Y127_AO6;
  assign CLBLL_L_X36Y128_SLICE_X55Y128_D2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X36Y128_SLICE_X55Y128_D3 = 1'b1;
  assign CLBLL_L_X36Y128_SLICE_X55Y128_D4 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X36Y128_SLICE_X55Y128_D5 = CLBLM_R_X37Y126_SLICE_X56Y126_AO5;
  assign CLBLL_L_X36Y128_SLICE_X55Y128_D6 = CLBLM_R_X35Y127_SLICE_X53Y127_A_XOR;
  assign CLBLM_R_X33Y121_SLICE_X49Y121_A6 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X33Y121_SLICE_X49Y121_B1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X33Y121_SLICE_X49Y121_B2 = CLBLL_L_X36Y121_SLICE_X54Y121_AO5;
  assign CLBLM_R_X33Y121_SLICE_X49Y121_B3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X33Y121_SLICE_X49Y121_B4 = CLBLM_R_X33Y122_SLICE_X49Y122_CO6;
  assign CLBLM_R_X33Y121_SLICE_X49Y121_B5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X33Y121_SLICE_X49Y121_B6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X33Y121_SLICE_X49Y121_C1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X33Y121_SLICE_X49Y121_C2 = 1'b1;
  assign CLBLM_R_X33Y121_SLICE_X49Y121_C3 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X33Y121_SLICE_X49Y121_C4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X33Y121_SLICE_X49Y121_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X34Y117_SLICE_X50Y117_A1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X34Y117_SLICE_X50Y117_A2 = CLBLM_R_X35Y117_SLICE_X52Y117_AO6;
  assign CLBLL_L_X34Y117_SLICE_X50Y117_A3 = CLBLL_L_X34Y119_SLICE_X50Y119_AO6;
  assign CLBLL_L_X34Y117_SLICE_X50Y117_A4 = CLBLL_L_X34Y119_SLICE_X50Y119_BO6;
  assign CLBLL_L_X34Y117_SLICE_X50Y117_A5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X34Y117_SLICE_X50Y117_A6 = CLBLL_L_X34Y114_SLICE_X51Y114_AO6;
  assign CLBLM_R_X33Y121_SLICE_X49Y121_C6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X33Y121_SLICE_X49Y121_D1 = 1'b1;
  assign CLBLL_L_X34Y117_SLICE_X50Y117_B1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X34Y117_SLICE_X50Y117_B2 = CLBLL_L_X34Y117_SLICE_X51Y117_BO6;
  assign CLBLL_L_X34Y117_SLICE_X50Y117_B3 = CLBLL_L_X34Y119_SLICE_X51Y119_CO6;
  assign CLBLL_L_X34Y117_SLICE_X50Y117_B4 = CLBLM_R_X33Y117_SLICE_X48Y117_AO6;
  assign CLBLL_L_X34Y117_SLICE_X50Y117_B5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X34Y117_SLICE_X50Y117_B6 = CLBLL_L_X34Y114_SLICE_X51Y114_CO6;
  assign CLBLM_R_X33Y121_SLICE_X49Y121_D2 = 1'b1;
  assign CLBLM_R_X33Y121_SLICE_X49Y121_D3 = 1'b1;
  assign CLBLM_R_X33Y121_SLICE_X49Y121_D4 = 1'b1;
  assign CLBLL_L_X34Y117_SLICE_X50Y117_C1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X34Y117_SLICE_X50Y117_C2 = CLBLM_R_X35Y117_SLICE_X52Y117_AO6;
  assign CLBLL_L_X34Y117_SLICE_X50Y117_C3 = CLBLL_L_X34Y115_SLICE_X50Y115_DO6;
  assign CLBLL_L_X34Y117_SLICE_X50Y117_C4 = CLBLL_L_X34Y114_SLICE_X51Y114_AO6;
  assign CLBLL_L_X34Y117_SLICE_X50Y117_C5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X34Y117_SLICE_X50Y117_C6 = CLBLL_L_X34Y119_SLICE_X50Y119_BO6;
  assign CLBLM_R_X33Y121_SLICE_X48Y121_A1 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLM_R_X33Y121_SLICE_X48Y121_A2 = CLBLL_L_X36Y116_SLICE_X55Y116_AO5;
  assign CLBLM_R_X33Y121_SLICE_X48Y121_A3 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLM_R_X33Y121_SLICE_X48Y121_A4 = CLBLM_R_X33Y121_SLICE_X48Y121_BO6;
  assign CLBLM_R_X33Y121_SLICE_X48Y121_A5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X33Y121_SLICE_X48Y121_A6 = CLBLM_R_X33Y121_SLICE_X48Y121_CO6;
  assign CLBLM_R_X33Y121_SLICE_X48Y121_B1 = CLBLL_L_X36Y122_SLICE_X55Y122_AO6;
  assign CLBLL_L_X34Y117_SLICE_X50Y117_D1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X34Y117_SLICE_X50Y117_D2 = 1'b1;
  assign CLBLL_L_X34Y117_SLICE_X50Y117_D3 = CLBLL_L_X34Y117_SLICE_X51Y117_BO6;
  assign CLBLL_L_X34Y117_SLICE_X50Y117_D4 = 1'b1;
  assign CLBLL_L_X34Y117_SLICE_X50Y117_D5 = 1'b1;
  assign CLBLL_L_X34Y117_SLICE_X50Y117_D6 = CLBLM_R_X33Y117_SLICE_X48Y117_AO6;
  assign CLBLM_R_X33Y121_SLICE_X48Y121_B2 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X33Y121_SLICE_X48Y121_B3 = CLBLM_R_X35Y120_SLICE_X52Y120_A_XOR;
  assign CLBLM_R_X33Y121_SLICE_X48Y121_B4 = CLBLM_R_X33Y121_SLICE_X48Y121_DO6;
  assign CLBLM_R_X33Y121_SLICE_X48Y121_B5 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLM_R_X33Y121_SLICE_X48Y121_B6 = CLBLM_R_X35Y122_SLICE_X53Y122_A_XOR;
  assign CLBLM_R_X33Y121_SLICE_X48Y121_C1 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLM_R_X33Y121_SLICE_X48Y121_C2 = CLBLM_R_X35Y122_SLICE_X53Y122_A_XOR;
  assign CLBLM_R_X33Y121_SLICE_X48Y121_C3 = CLBLL_L_X34Y128_SLICE_X50Y128_AO6;
  assign CLBLM_R_X33Y121_SLICE_X48Y121_C4 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_R_X33Y121_SLICE_X48Y121_C5 = CLBLM_R_X33Y121_SLICE_X49Y121_AO6;
  assign CLBLM_R_X33Y121_SLICE_X48Y121_C6 = CLBLL_L_X34Y121_SLICE_X50Y121_CO6;
  assign CLBLM_R_X35Y125_SLICE_X53Y125_D3 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X35Y125_SLICE_X53Y125_D4 = 1'b1;
  assign CLBLM_R_X35Y129_SLICE_X52Y129_D5 = 1'b1;
  assign CLBLM_R_X35Y125_SLICE_X53Y125_D5 = 1'b1;
  assign CLBLM_R_X33Y121_SLICE_X48Y121_D1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X33Y121_SLICE_X48Y121_D2 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLM_R_X33Y121_SLICE_X48Y121_D3 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLM_R_X33Y121_SLICE_X48Y121_D4 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_R_X33Y121_SLICE_X48Y121_D5 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X33Y121_SLICE_X48Y121_D6 = CLBLM_R_X35Y122_SLICE_X53Y122_A_XOR;
  assign CLBLM_R_X35Y125_SLICE_X53Y125_D6 = LIOB33_X0Y137_IOB_X0Y137_I;
  assign CLBLL_L_X34Y117_SLICE_X51Y117_A1 = CLBLM_R_X35Y120_SLICE_X53Y120_A_XOR;
  assign CLBLL_L_X34Y117_SLICE_X51Y117_A2 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X34Y117_SLICE_X51Y117_A3 = CLBLL_L_X36Y116_SLICE_X54Y116_BO5;
  assign CLBLL_L_X34Y117_SLICE_X51Y117_A4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X34Y117_SLICE_X51Y117_A5 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X34Y117_SLICE_X51Y117_A6 = CLBLL_L_X34Y119_SLICE_X51Y119_AO5;
  assign CLBLM_R_X37Y125_SLICE_X57Y125_B1 = CLBLM_R_X35Y125_SLICE_X53Y125_C_XOR;
  assign CLBLM_R_X37Y125_SLICE_X57Y125_B2 = CLBLL_L_X36Y122_SLICE_X55Y122_AO6;
  assign CLBLM_R_X35Y125_SLICE_X53Y125_DX = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X34Y117_SLICE_X51Y117_B1 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X34Y117_SLICE_X51Y117_B2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X34Y117_SLICE_X51Y117_B3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X34Y117_SLICE_X51Y117_B4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X34Y117_SLICE_X51Y117_B5 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X34Y117_SLICE_X51Y117_B6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X37Y125_SLICE_X57Y125_B3 = CLBLM_R_X35Y123_SLICE_X52Y123_C_XOR;
  assign CLBLM_R_X37Y125_SLICE_X57Y125_B4 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLL_L_X34Y117_SLICE_X51Y117_C1 = CLBLL_L_X34Y119_SLICE_X51Y119_CO6;
  assign CLBLL_L_X34Y117_SLICE_X51Y117_C2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X34Y117_SLICE_X51Y117_C3 = CLBLM_R_X33Y118_SLICE_X49Y118_AO6;
  assign CLBLL_L_X34Y117_SLICE_X51Y117_C4 = CLBLL_L_X34Y114_SLICE_X51Y114_CO6;
  assign CLBLL_L_X34Y117_SLICE_X51Y117_C5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X34Y117_SLICE_X51Y117_C6 = CLBLL_L_X34Y117_SLICE_X51Y117_BO6;
  assign CLBLM_R_X37Y125_SLICE_X57Y125_B5 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X37Y125_SLICE_X57Y125_B6 = CLBLM_R_X37Y125_SLICE_X57Y125_CO6;
  assign CLBLM_R_X35Y125_SLICE_X52Y125_A1 = LIOB33_X0Y141_IOB_X0Y142_I;
  assign CLBLL_L_X34Y117_SLICE_X51Y117_D1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X34Y117_SLICE_X51Y117_D2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X34Y117_SLICE_X51Y117_D3 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X34Y117_SLICE_X51Y117_D4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X34Y117_SLICE_X51Y117_D5 = 1'b1;
  assign CLBLL_L_X34Y117_SLICE_X51Y117_D6 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_C1 = CLBLM_R_X35Y124_SLICE_X53Y124_C_XOR;
  assign CLBLM_R_X35Y125_SLICE_X52Y125_A3 = 1'b1;
  assign CLBLM_R_X37Y125_SLICE_X57Y125_C1 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_R_X37Y125_SLICE_X57Y125_C2 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X37Y125_SLICE_X57Y125_C3 = LIOB33_X0Y135_IOB_X0Y136_I;
  assign CLBLM_R_X37Y125_SLICE_X57Y125_C4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X37Y125_SLICE_X57Y125_C5 = CLBLM_R_X35Y125_SLICE_X53Y125_C_XOR;
  assign CLBLM_R_X37Y125_SLICE_X57Y125_C6 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLM_R_X35Y125_SLICE_X52Y125_B1 = 1'b1;
  assign CLBLM_R_X35Y125_SLICE_X52Y125_B2 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X35Y125_SLICE_X52Y125_B3 = 1'b1;
  assign CLBLL_L_X36Y129_SLICE_X54Y129_A1 = CLBLL_L_X36Y116_SLICE_X55Y116_AO5;
  assign CLBLL_L_X36Y129_SLICE_X54Y129_A2 = CLBLL_L_X36Y128_SLICE_X55Y128_AO6;
  assign CLBLL_L_X36Y129_SLICE_X54Y129_A3 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X36Y129_SLICE_X54Y129_A4 = CLBLL_L_X36Y129_SLICE_X54Y129_BO6;
  assign CLBLL_L_X36Y129_SLICE_X54Y129_A5 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLL_L_X36Y129_SLICE_X54Y129_A6 = LIOB33_X0Y141_IOB_X0Y142_I;
  assign CLBLM_R_X35Y125_SLICE_X52Y125_B6 = LIOB33_X0Y143_IOB_X0Y143_I;
  assign CLBLL_L_X36Y129_SLICE_X54Y129_B1 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X36Y129_SLICE_X54Y129_B2 = CLBLM_R_X35Y125_SLICE_X52Y125_A_XOR;
  assign CLBLL_L_X36Y129_SLICE_X54Y129_B3 = CLBLL_L_X36Y122_SLICE_X55Y122_AO6;
  assign CLBLL_L_X36Y129_SLICE_X54Y129_B4 = CLBLM_R_X35Y127_SLICE_X53Y127_A_XOR;
  assign CLBLL_L_X36Y129_SLICE_X54Y129_B5 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLL_L_X36Y129_SLICE_X54Y129_B6 = CLBLL_L_X36Y129_SLICE_X54Y129_CO6;
  assign CLBLL_L_X36Y129_SLICE_X54Y129_C1 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X36Y129_SLICE_X54Y129_C2 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X36Y129_SLICE_X54Y129_C3 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X36Y129_SLICE_X54Y129_C4 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLL_L_X36Y129_SLICE_X54Y129_C5 = LIOB33_X0Y141_IOB_X0Y142_I;
  assign CLBLL_L_X36Y129_SLICE_X54Y129_C6 = CLBLM_R_X35Y127_SLICE_X53Y127_A_XOR;
  assign CLBLM_R_X35Y125_SLICE_X52Y125_C1 = LIOB33_X0Y143_IOB_X0Y144_I;
  assign CLBLM_R_X37Y125_SLICE_X57Y125_D5 = CLBLL_L_X36Y124_SLICE_X54Y124_DO6;
  assign CLBLL_L_X36Y129_SLICE_X54Y129_D1 = 1'b1;
  assign CLBLL_L_X36Y129_SLICE_X54Y129_D2 = 1'b1;
  assign CLBLL_L_X36Y129_SLICE_X54Y129_D3 = 1'b1;
  assign CLBLL_L_X36Y129_SLICE_X54Y129_D4 = 1'b1;
  assign CLBLL_L_X36Y129_SLICE_X54Y129_D5 = 1'b1;
  assign CLBLL_L_X36Y129_SLICE_X54Y129_D6 = 1'b1;
  assign CLBLM_R_X35Y125_SLICE_X52Y125_C2 = 1'b1;
  assign CLBLM_R_X37Y125_SLICE_X57Y125_D6 = CLBLM_R_X35Y125_SLICE_X53Y125_D_XOR;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_C2 = CLBLM_R_X37Y118_SLICE_X57Y118_CO6;
  assign CLBLM_R_X37Y125_SLICE_X56Y125_B1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X35Y125_SLICE_X52Y125_C6 = 1'b1;
  assign CLBLL_L_X36Y129_SLICE_X55Y129_A1 = CLBLL_L_X36Y116_SLICE_X55Y116_AO5;
  assign CLBLL_L_X36Y129_SLICE_X55Y129_A2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X36Y129_SLICE_X55Y129_A3 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLL_L_X36Y129_SLICE_X55Y129_A4 = CLBLL_L_X36Y129_SLICE_X55Y129_BO6;
  assign CLBLL_L_X36Y129_SLICE_X55Y129_A5 = CLBLL_L_X36Y126_SLICE_X55Y126_AO6;
  assign CLBLL_L_X36Y129_SLICE_X55Y129_A6 = LIOB33_X0Y141_IOB_X0Y141_I;
  assign CLBLM_R_X37Y125_SLICE_X56Y125_A1 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLL_L_X36Y129_SLICE_X55Y129_B1 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X36Y129_SLICE_X55Y129_B2 = CLBLM_R_X35Y126_SLICE_X53Y126_D_XOR;
  assign CLBLL_L_X36Y129_SLICE_X55Y129_B3 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLL_L_X36Y129_SLICE_X55Y129_B4 = CLBLL_L_X36Y122_SLICE_X55Y122_AO6;
  assign CLBLL_L_X36Y129_SLICE_X55Y129_B5 = CLBLM_R_X35Y124_SLICE_X52Y124_D_XOR;
  assign CLBLL_L_X36Y129_SLICE_X55Y129_B6 = CLBLL_L_X36Y129_SLICE_X55Y129_CO6;
  assign CLBLM_R_X37Y125_SLICE_X56Y125_A2 = CLBLM_R_X37Y124_SLICE_X56Y124_AO6;
  assign CLBLM_R_X37Y125_SLICE_X56Y125_A3 = CLBLL_L_X36Y120_SLICE_X55Y120_BO6;
  assign CLBLL_L_X36Y129_SLICE_X55Y129_C1 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X36Y129_SLICE_X55Y129_C2 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X36Y129_SLICE_X55Y129_C3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X36Y129_SLICE_X55Y129_C4 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLL_L_X36Y129_SLICE_X55Y129_C5 = LIOB33_X0Y141_IOB_X0Y141_I;
  assign CLBLL_L_X36Y129_SLICE_X55Y129_C6 = CLBLM_R_X35Y126_SLICE_X53Y126_D_XOR;
  assign CLBLM_R_X37Y125_SLICE_X56Y125_A4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X37Y125_SLICE_X56Y125_A5 = LIOB33_X0Y133_IOB_X0Y134_I;
  assign CLBLM_R_X33Y122_SLICE_X49Y122_A1 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X36Y129_SLICE_X55Y129_D1 = CLBLM_R_X35Y128_SLICE_X52Y128_BO6;
  assign CLBLL_L_X36Y129_SLICE_X55Y129_D2 = 1'b1;
  assign CLBLL_L_X36Y129_SLICE_X55Y129_D3 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X36Y129_SLICE_X55Y129_D4 = CLBLM_R_X35Y129_SLICE_X53Y129_BO6;
  assign CLBLL_L_X36Y129_SLICE_X55Y129_D5 = 1'b1;
  assign CLBLL_L_X36Y129_SLICE_X55Y129_D6 = CLBLM_R_X35Y129_SLICE_X53Y129_AO6;
  assign CLBLM_R_X33Y122_SLICE_X49Y122_A2 = CLBLL_L_X34Y128_SLICE_X50Y128_AO6;
  assign CLBLM_R_X33Y122_SLICE_X49Y122_A3 = CLBLL_L_X34Y122_SLICE_X50Y122_AO6;
  assign CLBLM_R_X33Y122_SLICE_X49Y122_A4 = CLBLM_R_X33Y122_SLICE_X49Y122_DO6;
  assign CLBLM_R_X33Y122_SLICE_X49Y122_A5 = CLBLM_R_X35Y122_SLICE_X53Y122_C_XOR;
  assign CLBLM_R_X33Y122_SLICE_X49Y122_A6 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLM_R_X33Y122_SLICE_X49Y122_B1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X33Y122_SLICE_X49Y122_B2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X33Y122_SLICE_X49Y122_B3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X33Y122_SLICE_X49Y122_B4 = CLBLL_L_X36Y121_SLICE_X54Y121_AO5;
  assign CLBLM_R_X33Y122_SLICE_X49Y122_B5 = CLBLM_R_X33Y123_SLICE_X48Y123_AO6;
  assign CLBLM_R_X33Y122_SLICE_X49Y122_B6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X33Y122_SLICE_X49Y122_C1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X34Y118_SLICE_X50Y118_A1 = CLBLM_R_X35Y118_SLICE_X53Y118_CO6;
  assign CLBLL_L_X34Y118_SLICE_X50Y118_A2 = CLBLM_R_X33Y118_SLICE_X49Y118_AO6;
  assign CLBLL_L_X34Y118_SLICE_X50Y118_A3 = CLBLL_L_X34Y118_SLICE_X51Y118_AO6;
  assign CLBLL_L_X34Y118_SLICE_X50Y118_A4 = CLBLM_R_X37Y118_SLICE_X57Y118_AO5;
  assign CLBLL_L_X34Y118_SLICE_X50Y118_A5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X34Y118_SLICE_X50Y118_A6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X33Y122_SLICE_X49Y122_C2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X33Y122_SLICE_X49Y122_C3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X33Y122_SLICE_X49Y122_C4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X34Y118_SLICE_X50Y118_B1 = CLBLL_L_X34Y114_SLICE_X51Y114_AO6;
  assign CLBLL_L_X34Y118_SLICE_X50Y118_B2 = CLBLL_L_X34Y119_SLICE_X50Y119_BO6;
  assign CLBLL_L_X34Y118_SLICE_X50Y118_B3 = CLBLL_L_X34Y119_SLICE_X50Y119_DO6;
  assign CLBLL_L_X34Y118_SLICE_X50Y118_B4 = CLBLM_R_X35Y117_SLICE_X52Y117_AO6;
  assign CLBLL_L_X34Y118_SLICE_X50Y118_B5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X34Y118_SLICE_X50Y118_B6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X33Y122_SLICE_X49Y122_D1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_L_X32Y123_SLICE_X47Y123_B3 = CLBLM_R_X33Y122_SLICE_X48Y122_AO6;
  assign CLBLL_L_X34Y118_SLICE_X50Y118_C1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X34Y118_SLICE_X50Y118_C2 = CLBLL_L_X34Y114_SLICE_X51Y114_AO6;
  assign CLBLL_L_X34Y118_SLICE_X50Y118_C3 = CLBLL_L_X34Y119_SLICE_X50Y119_DO6;
  assign CLBLL_L_X34Y118_SLICE_X50Y118_C4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X34Y118_SLICE_X50Y118_C5 = CLBLM_R_X33Y121_SLICE_X49Y121_CO6;
  assign CLBLL_L_X34Y118_SLICE_X50Y118_C6 = CLBLM_R_X35Y117_SLICE_X52Y117_AO6;
  assign CLBLM_R_X33Y122_SLICE_X48Y122_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X33Y122_SLICE_X48Y122_A2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_L_X32Y123_SLICE_X47Y123_B5 = CLBLM_L_X32Y123_SLICE_X47Y123_AO6;
  assign CLBLM_R_X33Y122_SLICE_X48Y122_A3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X33Y122_SLICE_X48Y122_A4 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X33Y122_SLICE_X48Y122_A5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X33Y122_SLICE_X48Y122_A6 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_B1 = 1'b1;
  assign CLBLL_L_X34Y118_SLICE_X50Y118_D1 = CLBLM_R_X33Y118_SLICE_X49Y118_AO6;
  assign CLBLL_L_X34Y118_SLICE_X50Y118_D2 = CLBLM_R_X35Y118_SLICE_X53Y118_CO6;
  assign CLBLL_L_X34Y118_SLICE_X50Y118_D3 = CLBLL_L_X34Y118_SLICE_X51Y118_AO6;
  assign CLBLL_L_X34Y118_SLICE_X50Y118_D4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X34Y118_SLICE_X50Y118_D5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X34Y118_SLICE_X50Y118_D6 = CLBLL_L_X34Y119_SLICE_X51Y119_CO6;
  assign CLBLM_R_X33Y122_SLICE_X48Y122_B1 = CLBLM_R_X33Y125_SLICE_X49Y125_BO5;
  assign CLBLM_R_X33Y122_SLICE_X48Y122_B2 = CLBLM_R_X33Y122_SLICE_X48Y122_AO5;
  assign CLBLM_R_X33Y122_SLICE_X48Y122_B3 = CLBLM_L_X32Y123_SLICE_X47Y123_AO5;
  assign CLBLM_R_X33Y122_SLICE_X48Y122_B4 = CLBLL_L_X34Y123_SLICE_X50Y123_BO6;
  assign CLBLM_R_X33Y122_SLICE_X48Y122_B5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X33Y122_SLICE_X48Y122_B6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X33Y122_SLICE_X48Y122_C3 = 1'b1;
  assign CLBLM_R_X33Y122_SLICE_X48Y122_C4 = 1'b1;
  assign CLBLM_R_X33Y122_SLICE_X48Y122_C5 = 1'b1;
  assign CLBLM_R_X33Y122_SLICE_X48Y122_C6 = 1'b1;
  assign CLBLM_R_X33Y122_SLICE_X48Y122_C1 = 1'b1;
  assign CLBLM_R_X33Y122_SLICE_X48Y122_C2 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_B5 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_B6 = 1'b1;
  assign CLBLM_R_X37Y125_SLICE_X56Y125_C1 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X33Y122_SLICE_X48Y122_D1 = 1'b1;
  assign CLBLM_R_X33Y122_SLICE_X48Y122_D2 = 1'b1;
  assign CLBLM_R_X33Y122_SLICE_X48Y122_D3 = 1'b1;
  assign CLBLM_R_X33Y122_SLICE_X48Y122_D4 = 1'b1;
  assign CLBLM_R_X33Y122_SLICE_X48Y122_D5 = 1'b1;
  assign CLBLM_R_X33Y122_SLICE_X48Y122_D6 = 1'b1;
  assign CLBLL_L_X34Y118_SLICE_X51Y118_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X34Y118_SLICE_X51Y118_A2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X34Y118_SLICE_X51Y118_A3 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X34Y118_SLICE_X51Y118_A4 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLL_L_X34Y118_SLICE_X51Y118_A5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X34Y118_SLICE_X51Y118_A6 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_C1 = 1'b1;
  assign CLBLL_L_X34Y118_SLICE_X51Y118_B1 = CLBLM_R_X35Y118_SLICE_X53Y118_CO6;
  assign CLBLL_L_X34Y118_SLICE_X51Y118_B2 = CLBLL_L_X36Y115_SLICE_X54Y115_AO6;
  assign CLBLL_L_X34Y118_SLICE_X51Y118_B3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X34Y118_SLICE_X51Y118_B4 = CLBLM_R_X37Y118_SLICE_X57Y118_AO5;
  assign CLBLL_L_X34Y118_SLICE_X51Y118_B5 = CLBLL_L_X34Y118_SLICE_X51Y118_AO6;
  assign CLBLL_L_X34Y118_SLICE_X51Y118_B6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_C2 = 1'b1;
  assign CLBLM_R_X37Y125_SLICE_X56Y125_C5 = CLBLL_L_X36Y116_SLICE_X54Y116_BO5;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_C3 = 1'b1;
  assign CLBLL_L_X34Y118_SLICE_X51Y118_C1 = CLBLL_L_X34Y118_SLICE_X51Y118_AO6;
  assign CLBLL_L_X34Y118_SLICE_X51Y118_C2 = CLBLL_L_X34Y119_SLICE_X51Y119_CO6;
  assign CLBLL_L_X34Y118_SLICE_X51Y118_C3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X34Y118_SLICE_X51Y118_C4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X34Y118_SLICE_X51Y118_C5 = CLBLM_R_X33Y118_SLICE_X49Y118_AO6;
  assign CLBLL_L_X34Y118_SLICE_X51Y118_C6 = CLBLL_L_X34Y117_SLICE_X51Y117_BO6;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_C4 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_C5 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_C6 = 1'b1;
  assign CLBLL_L_X34Y118_SLICE_X51Y118_D1 = CLBLM_R_X35Y118_SLICE_X52Y118_A_XOR;
  assign CLBLL_L_X34Y118_SLICE_X51Y118_D2 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X34Y118_SLICE_X51Y118_D3 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X34Y118_SLICE_X51Y118_D4 = 1'b1;
  assign CLBLL_L_X34Y118_SLICE_X51Y118_D5 = CLBLM_R_X35Y120_SLICE_X53Y120_A_XOR;
  assign CLBLL_L_X34Y118_SLICE_X51Y118_D6 = CLBLL_L_X34Y126_SLICE_X51Y126_D_CY;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_D1 = CLBLM_R_X35Y119_SLICE_X53Y119_AO6;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_T1 = 1'b1;
  assign CLBLM_R_X35Y120_SLICE_X52Y120_B4 = 1'b1;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_D1 = CLBLL_L_X34Y124_SLICE_X50Y124_AO6;
  assign CLBLM_R_X35Y120_SLICE_X52Y120_B5 = 1'b1;
  assign CLBLM_R_X37Y125_SLICE_X56Y125_D1 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign RIOI3_X105Y121_OLOGIC_X1Y122_D1 = CLBLM_R_X35Y116_SLICE_X53Y116_BO6;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_T1 = 1'b1;
  assign CLBLM_R_X35Y115_SLICE_X53Y115_B3 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLM_R_X37Y125_SLICE_X56Y125_D2 = CLBLL_L_X36Y124_SLICE_X54Y124_DO6;
  assign CLBLM_R_X37Y125_SLICE_X56Y125_D3 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_D1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_D1 = CLBLL_L_X36Y129_SLICE_X55Y129_AO6;
  assign CLBLM_R_X37Y125_SLICE_X56Y125_D4 = CLBLL_L_X36Y123_SLICE_X54Y123_DO6;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_D2 = 1'b1;
  assign CLBLM_R_X35Y115_SLICE_X53Y115_B6 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_D3 = 1'b1;
  assign CLBLM_R_X37Y125_SLICE_X56Y125_D5 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_T1 = 1'b1;
  assign CLBLM_R_X37Y125_SLICE_X56Y125_D6 = CLBLM_R_X35Y125_SLICE_X53Y125_D_XOR;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_D4 = 1'b1;
  assign CLBLM_R_X37Y125_SLICE_X56Y125_B3 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_D5 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_D1 = CLBLM_R_X35Y126_SLICE_X52Y126_BO6;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_T1 = 1'b1;
  assign RIOI3_X105Y121_OLOGIC_X1Y122_T1 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_A5 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_A6 = CLBLM_R_X37Y120_SLICE_X56Y120_CO6;
  assign RIOI3_X105Y121_OLOGIC_X1Y121_D1 = CLBLM_R_X35Y115_SLICE_X52Y115_BO6;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_B1 = CLBLM_R_X37Y120_SLICE_X56Y120_DO6;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_B2 = CLBLL_L_X34Y128_SLICE_X50Y128_AO6;
  assign LIOI3_X0Y147_ILOGIC_X0Y148_D = LIOB33_X0Y147_IOB_X0Y148_I;
  assign LIOI3_X0Y147_ILOGIC_X0Y147_D = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_B3 = CLBLM_R_X35Y124_SLICE_X53Y124_D_XOR;
  assign LIOI3_X0Y117_ILOGIC_X0Y118_D = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_B4 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign LIOI3_X0Y117_ILOGIC_X0Y117_D = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X33Y123_SLICE_X49Y123_A1 = CLBLL_L_X36Y116_SLICE_X55Y116_AO5;
  assign CLBLM_R_X33Y123_SLICE_X49Y123_A2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X33Y123_SLICE_X49Y123_A3 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLM_R_X33Y123_SLICE_X49Y123_A4 = CLBLM_R_X33Y123_SLICE_X49Y123_BO6;
  assign CLBLM_R_X33Y123_SLICE_X49Y123_A5 = CLBLM_R_X33Y122_SLICE_X49Y122_AO6;
  assign CLBLM_R_X33Y123_SLICE_X49Y123_A6 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_B5 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_B6 = CLBLL_L_X36Y120_SLICE_X55Y120_AO6;
  assign CLBLM_R_X37Y123_SLICE_X57Y123_A2 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLM_R_X33Y123_SLICE_X49Y123_B1 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLM_R_X33Y123_SLICE_X49Y123_B2 = CLBLL_L_X36Y122_SLICE_X55Y122_AO6;
  assign CLBLM_R_X33Y123_SLICE_X49Y123_B3 = CLBLM_R_X35Y122_SLICE_X53Y122_C_XOR;
  assign CLBLM_R_X33Y123_SLICE_X49Y123_B4 = CLBLM_R_X35Y120_SLICE_X52Y120_C_XOR;
  assign CLBLM_R_X33Y123_SLICE_X49Y123_B5 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X33Y123_SLICE_X49Y123_B6 = CLBLM_R_X33Y123_SLICE_X49Y123_CO6;
  assign CLBLL_L_X34Y119_SLICE_X50Y119_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X34Y119_SLICE_X50Y119_A2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X34Y119_SLICE_X50Y119_A3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X34Y119_SLICE_X50Y119_A4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X34Y119_SLICE_X50Y119_A5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X34Y119_SLICE_X50Y119_A6 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X33Y123_SLICE_X49Y123_C1 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLM_R_X33Y123_SLICE_X49Y123_C2 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X34Y119_SLICE_X50Y119_B1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X34Y119_SLICE_X50Y119_B2 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X34Y119_SLICE_X50Y119_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X34Y119_SLICE_X50Y119_B4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X34Y119_SLICE_X50Y119_B5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X34Y119_SLICE_X50Y119_B6 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X33Y123_SLICE_X49Y123_C5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X33Y123_SLICE_X49Y123_C6 = CLBLM_R_X35Y122_SLICE_X53Y122_C_XOR;
  assign CLBLL_L_X34Y119_SLICE_X50Y119_C1 = CLBLM_R_X35Y117_SLICE_X52Y117_AO6;
  assign CLBLL_L_X34Y119_SLICE_X50Y119_C2 = CLBLM_R_X33Y121_SLICE_X49Y121_CO6;
  assign CLBLL_L_X34Y119_SLICE_X50Y119_C3 = CLBLL_L_X34Y121_SLICE_X51Y121_DO6;
  assign CLBLL_L_X34Y119_SLICE_X50Y119_C4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X34Y119_SLICE_X50Y119_C5 = CLBLL_L_X34Y119_SLICE_X50Y119_DO6;
  assign CLBLL_L_X34Y119_SLICE_X50Y119_C6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X33Y123_SLICE_X49Y123_D1 = CLBLM_R_X33Y125_SLICE_X49Y125_AO6;
  assign CLBLM_R_X33Y123_SLICE_X49Y123_D2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X33Y123_SLICE_X49Y123_D3 = CLBLM_R_X33Y124_SLICE_X49Y124_AO5;
  assign CLBLM_R_X33Y123_SLICE_X49Y123_D4 = 1'b1;
  assign CLBLM_R_X33Y123_SLICE_X49Y123_D5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X33Y123_SLICE_X48Y123_A1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X33Y123_SLICE_X48Y123_A2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X33Y123_SLICE_X48Y123_A3 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X34Y119_SLICE_X50Y119_D1 = 1'b1;
  assign CLBLL_L_X34Y119_SLICE_X50Y119_D2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X34Y119_SLICE_X50Y119_D3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X34Y119_SLICE_X50Y119_D4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X34Y119_SLICE_X50Y119_D5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X34Y119_SLICE_X50Y119_D6 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X33Y123_SLICE_X48Y123_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X33Y123_SLICE_X48Y123_A5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X33Y123_SLICE_X48Y123_A6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X33Y123_SLICE_X48Y123_B1 = CLBLL_L_X34Y123_SLICE_X50Y123_AO6;
  assign CLBLM_R_X33Y123_SLICE_X48Y123_B2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X33Y123_SLICE_X48Y123_B3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X33Y123_SLICE_X48Y123_B4 = CLBLM_R_X33Y124_SLICE_X49Y124_AO6;
  assign CLBLM_R_X33Y123_SLICE_X48Y123_B5 = CLBLM_R_X33Y125_SLICE_X49Y125_AO6;
  assign CLBLM_R_X33Y123_SLICE_X48Y123_B6 = CLBLM_R_X33Y124_SLICE_X48Y124_AO5;
  assign CLBLM_R_X33Y123_SLICE_X48Y123_C1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X33Y123_SLICE_X48Y123_C2 = CLBLM_R_X33Y124_SLICE_X48Y124_AO5;
  assign CLBLM_R_X33Y123_SLICE_X48Y123_C3 = CLBLM_R_X33Y125_SLICE_X49Y125_AO5;
  assign CLBLM_R_X33Y123_SLICE_X48Y123_C4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X33Y123_SLICE_X48Y123_C5 = CLBLL_L_X34Y123_SLICE_X50Y123_AO6;
  assign CLBLM_R_X33Y123_SLICE_X48Y123_C6 = CLBLM_R_X33Y124_SLICE_X49Y124_AO6;
  assign CLBLM_R_X33Y123_SLICE_X49Y123_D6 = CLBLM_L_X32Y123_SLICE_X46Y123_AO6;
  assign CLBLM_R_X33Y123_SLICE_X48Y123_D1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X34Y119_SLICE_X51Y119_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X34Y119_SLICE_X51Y119_A2 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X34Y119_SLICE_X51Y119_A3 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLL_L_X34Y119_SLICE_X51Y119_A4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X34Y119_SLICE_X51Y119_A5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X34Y119_SLICE_X51Y119_A6 = 1'b1;
  assign CLBLM_R_X33Y123_SLICE_X48Y123_D2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X33Y123_SLICE_X48Y123_D3 = CLBLM_R_X33Y125_SLICE_X49Y125_AO5;
  assign CLBLM_R_X33Y123_SLICE_X48Y123_D4 = CLBLM_R_X33Y124_SLICE_X49Y124_AO6;
  assign CLBLL_L_X34Y119_SLICE_X51Y119_B1 = CLBLL_L_X34Y121_SLICE_X51Y121_DO6;
  assign CLBLL_L_X34Y119_SLICE_X51Y119_B2 = CLBLM_R_X35Y118_SLICE_X53Y118_AO5;
  assign CLBLL_L_X34Y119_SLICE_X51Y119_B3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X34Y119_SLICE_X51Y119_B4 = CLBLM_R_X37Y117_SLICE_X56Y117_AO5;
  assign CLBLL_L_X34Y119_SLICE_X51Y119_B5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X34Y119_SLICE_X51Y119_B6 = CLBLL_L_X36Y121_SLICE_X55Y121_AO6;
  assign CLBLM_R_X35Y115_SLICE_X52Y115_B4 = CLBLL_L_X34Y115_SLICE_X50Y115_BO6;
  assign CLBLL_L_X34Y119_SLICE_X51Y119_C1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X34Y119_SLICE_X51Y119_C2 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X34Y119_SLICE_X51Y119_C3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X34Y119_SLICE_X51Y119_C4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X34Y119_SLICE_X51Y119_C5 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLL_L_X34Y119_SLICE_X51Y119_C6 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X32Y123_SLICE_X46Y123_D3 = 1'b1;
  assign CLBLM_L_X32Y123_SLICE_X46Y123_D4 = 1'b1;
  assign CLBLM_R_X35Y115_SLICE_X52Y115_B5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X35Y115_SLICE_X52Y115_B6 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLM_L_X32Y123_SLICE_X46Y123_D5 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_D1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X34Y119_SLICE_X51Y119_D1 = CLBLM_R_X35Y118_SLICE_X53Y118_BO6;
  assign CLBLL_L_X34Y119_SLICE_X51Y119_D2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X34Y119_SLICE_X51Y119_D3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X34Y119_SLICE_X51Y119_D4 = CLBLL_L_X36Y121_SLICE_X54Y121_AO5;
  assign CLBLL_L_X34Y119_SLICE_X51Y119_D5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X34Y119_SLICE_X51Y119_D6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_D2 = CLBLM_R_X37Y118_SLICE_X57Y118_DO6;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_D3 = CLBLM_R_X35Y124_SLICE_X53Y124_D_XOR;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_D4 = CLBLM_R_X37Y118_SLICE_X56Y118_CO6;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_D5 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign LIOB33_X0Y65_IOB_X0Y65_O = CLBLL_L_X34Y115_SLICE_X51Y115_AO6;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_D6 = 1'b1;
  assign RIOI3_X105Y141_OLOGIC_X1Y141_D1 = CLBLL_L_X36Y127_SLICE_X54Y127_AO6;
  assign CLBLM_R_X33Y124_SLICE_X49Y124_B6 = CLBLM_R_X33Y124_SLICE_X49Y124_AO5;
  assign CLBLM_R_X33Y124_SLICE_X49Y124_C4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X33Y124_SLICE_X49Y124_C5 = CLBLM_R_X33Y124_SLICE_X48Y124_AO6;
  assign CLBLM_R_X33Y124_SLICE_X49Y124_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X33Y124_SLICE_X49Y124_A2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X33Y124_SLICE_X49Y124_A3 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X33Y124_SLICE_X49Y124_A4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X33Y124_SLICE_X49Y124_A5 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X33Y124_SLICE_X49Y124_A6 = 1'b1;
  assign CLBLM_R_X33Y124_SLICE_X49Y124_C6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X33Y124_SLICE_X49Y124_B1 = CLBLL_L_X34Y123_SLICE_X50Y123_AO6;
  assign CLBLM_R_X33Y124_SLICE_X49Y124_B2 = CLBLM_R_X33Y124_SLICE_X48Y124_AO6;
  assign CLBLL_L_X34Y120_SLICE_X50Y120_A1 = CLBLL_L_X34Y121_SLICE_X51Y121_DO6;
  assign CLBLL_L_X34Y120_SLICE_X50Y120_A2 = CLBLM_R_X33Y121_SLICE_X49Y121_CO6;
  assign CLBLL_L_X34Y120_SLICE_X50Y120_A3 = CLBLM_R_X35Y118_SLICE_X53Y118_AO5;
  assign CLBLL_L_X34Y120_SLICE_X50Y120_A4 = CLBLL_L_X36Y121_SLICE_X55Y121_AO6;
  assign CLBLL_L_X34Y120_SLICE_X50Y120_A5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X34Y120_SLICE_X50Y120_A6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X33Y124_SLICE_X49Y124_B3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X33Y124_SLICE_X49Y124_B4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X33Y124_SLICE_X49Y124_B5 = CLBLM_R_X33Y125_SLICE_X49Y125_AO6;
  assign CLBLL_L_X34Y120_SLICE_X50Y120_B1 = CLBLL_L_X34Y120_SLICE_X50Y120_DO6;
  assign CLBLL_L_X34Y120_SLICE_X50Y120_B2 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLL_L_X34Y120_SLICE_X50Y120_B3 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X34Y120_SLICE_X50Y120_B4 = CLBLM_R_X35Y121_SLICE_X53Y121_D_XOR;
  assign CLBLL_L_X34Y120_SLICE_X50Y120_B5 = CLBLL_L_X34Y128_SLICE_X50Y128_AO6;
  assign CLBLL_L_X34Y120_SLICE_X50Y120_B6 = CLBLM_R_X33Y119_SLICE_X49Y119_CO6;
  assign CLBLM_R_X33Y124_SLICE_X49Y124_C1 = CLBLM_R_X33Y124_SLICE_X49Y124_AO6;
  assign CLBLM_R_X33Y124_SLICE_X49Y124_C2 = CLBLM_R_X33Y125_SLICE_X49Y125_AO6;
  assign CLBLM_R_X33Y124_SLICE_X49Y124_C3 = CLBLL_L_X34Y123_SLICE_X50Y123_AO6;
  assign CLBLL_L_X34Y120_SLICE_X50Y120_C1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X34Y120_SLICE_X50Y120_C2 = CLBLM_R_X33Y121_SLICE_X49Y121_CO6;
  assign CLBLL_L_X34Y120_SLICE_X50Y120_C3 = CLBLL_L_X36Y121_SLICE_X55Y121_AO6;
  assign CLBLL_L_X34Y120_SLICE_X50Y120_C4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X34Y120_SLICE_X50Y120_C5 = CLBLL_L_X34Y121_SLICE_X51Y121_DO6;
  assign CLBLL_L_X34Y120_SLICE_X50Y120_C6 = CLBLL_L_X34Y119_SLICE_X50Y119_DO6;
  assign CLBLM_R_X33Y124_SLICE_X49Y124_D1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X33Y124_SLICE_X49Y124_D2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X33Y124_SLICE_X49Y124_D3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X33Y124_SLICE_X49Y124_D4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X33Y124_SLICE_X49Y124_D5 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X33Y124_SLICE_X49Y124_D6 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X34Y120_SLICE_X50Y120_D1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X34Y120_SLICE_X50Y120_D2 = CLBLL_L_X34Y118_SLICE_X50Y118_DO6;
  assign CLBLL_L_X34Y120_SLICE_X50Y120_D3 = CLBLM_R_X35Y117_SLICE_X52Y117_CO6;
  assign CLBLL_L_X34Y120_SLICE_X50Y120_D4 = 1'b1;
  assign CLBLL_L_X34Y120_SLICE_X50Y120_D5 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X34Y120_SLICE_X50Y120_D6 = CLBLM_R_X35Y121_SLICE_X53Y121_D_XOR;
  assign CLBLM_R_X33Y124_SLICE_X48Y124_A1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X33Y124_SLICE_X48Y124_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X33Y124_SLICE_X48Y124_A3 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X33Y124_SLICE_X48Y124_A4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X33Y124_SLICE_X48Y124_A5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X33Y124_SLICE_X48Y124_A6 = 1'b1;
  assign CLBLM_R_X33Y124_SLICE_X48Y124_B1 = CLBLM_R_X33Y125_SLICE_X49Y125_BO5;
  assign CLBLM_R_X33Y124_SLICE_X48Y124_B2 = CLBLL_L_X34Y123_SLICE_X50Y123_BO5;
  assign CLBLM_R_X33Y124_SLICE_X48Y124_B3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X33Y124_SLICE_X48Y124_B4 = CLBLM_L_X32Y123_SLICE_X47Y123_AO5;
  assign CLBLM_R_X33Y124_SLICE_X48Y124_B5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X33Y124_SLICE_X48Y124_B6 = CLBLM_R_X33Y122_SLICE_X48Y122_AO5;
  assign CLBLM_R_X33Y124_SLICE_X48Y124_C1 = 1'b1;
  assign CLBLM_R_X33Y124_SLICE_X48Y124_C2 = 1'b1;
  assign CLBLM_R_X33Y124_SLICE_X48Y124_C3 = 1'b1;
  assign CLBLM_R_X33Y124_SLICE_X48Y124_C4 = 1'b1;
  assign CLBLM_R_X33Y124_SLICE_X48Y124_C5 = 1'b1;
  assign CLBLM_R_X33Y124_SLICE_X48Y124_C6 = 1'b1;
  assign CLBLL_L_X34Y120_SLICE_X51Y120_A1 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLL_L_X34Y120_SLICE_X51Y120_A2 = CLBLL_L_X34Y120_SLICE_X50Y120_BO6;
  assign CLBLL_L_X34Y120_SLICE_X51Y120_A3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X34Y120_SLICE_X51Y120_A4 = CLBLL_L_X34Y120_SLICE_X51Y120_BO6;
  assign CLBLL_L_X34Y120_SLICE_X51Y120_A5 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLL_L_X34Y120_SLICE_X51Y120_A6 = CLBLL_L_X36Y116_SLICE_X55Y116_AO5;
  assign CLBLM_R_X33Y124_SLICE_X48Y124_D1 = 1'b1;
  assign CLBLM_R_X33Y124_SLICE_X48Y124_D2 = 1'b1;
  assign CLBLL_L_X34Y120_SLICE_X51Y120_B1 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X34Y120_SLICE_X51Y120_B2 = CLBLM_R_X35Y121_SLICE_X53Y121_D_XOR;
  assign CLBLL_L_X34Y120_SLICE_X51Y120_B3 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLL_L_X34Y120_SLICE_X51Y120_B4 = CLBLM_R_X35Y119_SLICE_X52Y119_D_XOR;
  assign CLBLL_L_X34Y120_SLICE_X51Y120_B5 = CLBLL_L_X36Y122_SLICE_X55Y122_AO6;
  assign CLBLL_L_X34Y120_SLICE_X51Y120_B6 = CLBLL_L_X34Y120_SLICE_X51Y120_CO6;
  assign CLBLM_R_X33Y124_SLICE_X48Y124_D4 = 1'b1;
  assign CLBLM_R_X33Y124_SLICE_X48Y124_D5 = 1'b1;
  assign CLBLL_L_X34Y120_SLICE_X51Y120_C1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X34Y120_SLICE_X51Y120_C2 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X34Y120_SLICE_X51Y120_C3 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X34Y120_SLICE_X51Y120_C4 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLL_L_X34Y120_SLICE_X51Y120_C5 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLL_L_X34Y120_SLICE_X51Y120_C6 = CLBLM_R_X35Y121_SLICE_X53Y121_D_XOR;
  assign CLBLL_L_X34Y120_SLICE_X51Y120_D1 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X34Y120_SLICE_X51Y120_D2 = CLBLL_L_X34Y118_SLICE_X51Y118_CO6;
  assign CLBLL_L_X34Y120_SLICE_X51Y120_D3 = CLBLM_R_X35Y121_SLICE_X53Y121_C_XOR;
  assign CLBLL_L_X34Y120_SLICE_X51Y120_D4 = 1'b1;
  assign CLBLL_L_X34Y120_SLICE_X51Y120_D5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X34Y120_SLICE_X51Y120_D6 = CLBLM_R_X35Y117_SLICE_X52Y117_CO6;
  assign CLBLM_R_X37Y125_SLICE_X56Y125_B4 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X33Y119_SLICE_X49Y119_B3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X36Y122_SLICE_X55Y122_A1 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X36Y122_SLICE_X55Y122_A2 = 1'b1;
  assign CLBLL_L_X36Y122_SLICE_X55Y122_A3 = 1'b1;
  assign CLBLM_R_X33Y119_SLICE_X49Y119_B6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_D1 = CLBLM_R_X37Y122_SLICE_X57Y122_AO6;
  assign RIOI3_X105Y141_OLOGIC_X1Y141_T1 = 1'b1;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_T1 = 1'b1;
  assign CLBLL_L_X36Y122_SLICE_X55Y122_B2 = CLBLL_L_X36Y119_SLICE_X54Y119_BO6;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_D1 = CLBLM_R_X37Y121_SLICE_X57Y121_AO6;
  assign CLBLL_L_X36Y122_SLICE_X55Y122_B3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X36Y122_SLICE_X55Y122_B4 = CLBLL_L_X36Y122_SLICE_X54Y122_CO6;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_T1 = 1'b1;
  assign CLBLL_L_X36Y122_SLICE_X55Y122_B5 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLL_L_X36Y122_SLICE_X55Y122_B6 = LIOB33_X0Y129_IOB_X0Y129_I;
  assign CLBLM_R_X33Y125_SLICE_X49Y125_A1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X33Y125_SLICE_X49Y125_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X33Y125_SLICE_X49Y125_A3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X33Y125_SLICE_X49Y125_A4 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X33Y125_SLICE_X49Y125_A5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X33Y125_SLICE_X49Y125_A6 = 1'b1;
  assign CLBLM_R_X33Y124_SLICE_X48Y124_D3 = 1'b1;
  assign CLBLL_L_X34Y121_SLICE_X50Y121_A1 = CLBLL_L_X34Y121_SLICE_X50Y121_DO6;
  assign CLBLL_L_X34Y121_SLICE_X50Y121_A2 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X34Y121_SLICE_X50Y121_A3 = CLBLL_L_X34Y128_SLICE_X50Y128_AO6;
  assign CLBLL_L_X34Y121_SLICE_X50Y121_A4 = CLBLL_L_X34Y121_SLICE_X50Y121_BO6;
  assign CLBLL_L_X34Y121_SLICE_X50Y121_A5 = CLBLM_R_X35Y122_SLICE_X53Y122_B_XOR;
  assign CLBLL_L_X34Y121_SLICE_X50Y121_A6 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLM_R_X33Y125_SLICE_X49Y125_B1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X33Y125_SLICE_X49Y125_B2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X34Y121_SLICE_X50Y121_B1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X34Y121_SLICE_X50Y121_B2 = CLBLM_R_X33Y118_SLICE_X49Y118_BO6;
  assign CLBLL_L_X34Y121_SLICE_X50Y121_B3 = CLBLM_R_X33Y121_SLICE_X49Y121_BO6;
  assign CLBLL_L_X34Y121_SLICE_X50Y121_B4 = CLBLM_R_X33Y122_SLICE_X49Y122_BO6;
  assign CLBLL_L_X34Y121_SLICE_X50Y121_B5 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X34Y121_SLICE_X50Y121_B6 = CLBLL_L_X34Y120_SLICE_X50Y120_CO6;
  assign CLBLM_R_X33Y124_SLICE_X48Y124_D6 = 1'b1;
  assign CLBLM_R_X33Y125_SLICE_X49Y125_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X33Y125_SLICE_X49Y125_C5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X34Y121_SLICE_X50Y121_C1 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X34Y121_SLICE_X50Y121_C2 = CLBLM_R_X35Y122_SLICE_X53Y122_A_XOR;
  assign CLBLL_L_X34Y121_SLICE_X50Y121_C3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X34Y121_SLICE_X50Y121_C4 = CLBLM_R_X35Y117_SLICE_X52Y117_DO6;
  assign CLBLL_L_X34Y121_SLICE_X50Y121_C5 = 1'b1;
  assign CLBLL_L_X34Y121_SLICE_X50Y121_C6 = CLBLL_L_X34Y118_SLICE_X50Y118_DO6;
  assign CLBLM_R_X33Y119_SLICE_X49Y119_D6 = 1'b1;
  assign CLBLM_R_X33Y125_SLICE_X49Y125_C6 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X33Y125_SLICE_X49Y125_D1 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X33Y125_SLICE_X49Y125_D2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X33Y125_SLICE_X49Y125_D3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X33Y125_SLICE_X49Y125_D4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X33Y125_SLICE_X49Y125_D5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X34Y121_SLICE_X50Y121_D1 = CLBLL_L_X34Y118_SLICE_X50Y118_AO6;
  assign CLBLL_L_X34Y121_SLICE_X50Y121_D2 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X34Y121_SLICE_X50Y121_D3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X34Y121_SLICE_X50Y121_D4 = CLBLM_R_X35Y117_SLICE_X52Y117_DO6;
  assign CLBLL_L_X34Y121_SLICE_X50Y121_D5 = CLBLM_R_X35Y122_SLICE_X53Y122_B_XOR;
  assign CLBLL_L_X34Y121_SLICE_X50Y121_D6 = 1'b1;
  assign CLBLM_R_X33Y125_SLICE_X48Y125_A1 = 1'b1;
  assign CLBLM_R_X33Y125_SLICE_X48Y125_A2 = 1'b1;
  assign CLBLM_R_X33Y125_SLICE_X48Y125_A3 = 1'b1;
  assign CLBLM_R_X33Y125_SLICE_X48Y125_A4 = 1'b1;
  assign CLBLM_R_X33Y125_SLICE_X48Y125_A5 = 1'b1;
  assign CLBLM_R_X33Y125_SLICE_X48Y125_A6 = 1'b1;
  assign CLBLM_R_X33Y125_SLICE_X48Y125_B1 = 1'b1;
  assign CLBLM_R_X33Y125_SLICE_X48Y125_B2 = 1'b1;
  assign CLBLM_R_X33Y125_SLICE_X48Y125_B3 = 1'b1;
  assign CLBLM_R_X33Y125_SLICE_X48Y125_B4 = 1'b1;
  assign CLBLM_R_X33Y125_SLICE_X48Y125_B5 = 1'b1;
  assign CLBLM_R_X33Y125_SLICE_X48Y125_B6 = 1'b1;
  assign CLBLM_R_X33Y125_SLICE_X48Y125_C1 = 1'b1;
  assign CLBLM_R_X33Y125_SLICE_X48Y125_C2 = 1'b1;
  assign CLBLM_R_X33Y125_SLICE_X48Y125_C3 = 1'b1;
  assign CLBLM_R_X33Y125_SLICE_X48Y125_C4 = 1'b1;
  assign CLBLM_R_X33Y125_SLICE_X48Y125_C5 = 1'b1;
  assign CLBLM_R_X33Y125_SLICE_X48Y125_C6 = 1'b1;
  assign CLBLL_L_X34Y121_SLICE_X51Y121_A1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X34Y121_SLICE_X51Y121_A2 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLL_L_X34Y121_SLICE_X51Y121_A3 = CLBLL_L_X34Y121_SLICE_X50Y121_AO6;
  assign CLBLL_L_X34Y121_SLICE_X51Y121_A4 = CLBLL_L_X34Y121_SLICE_X51Y121_BO6;
  assign CLBLL_L_X34Y121_SLICE_X51Y121_A5 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_L_X34Y121_SLICE_X51Y121_A6 = CLBLL_L_X36Y116_SLICE_X55Y116_AO5;
  assign CLBLM_R_X33Y125_SLICE_X48Y125_D1 = 1'b1;
  assign CLBLL_L_X34Y121_SLICE_X51Y121_B1 = CLBLL_L_X36Y122_SLICE_X55Y122_AO6;
  assign CLBLL_L_X34Y121_SLICE_X51Y121_B2 = CLBLM_R_X35Y122_SLICE_X53Y122_B_XOR;
  assign CLBLL_L_X34Y121_SLICE_X51Y121_B3 = CLBLM_R_X35Y120_SLICE_X52Y120_B_XOR;
  assign CLBLL_L_X34Y121_SLICE_X51Y121_B4 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLL_L_X34Y121_SLICE_X51Y121_B5 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X34Y121_SLICE_X51Y121_B6 = CLBLL_L_X34Y121_SLICE_X51Y121_CO6;
  assign CLBLM_R_X33Y119_SLICE_X48Y119_A4 = 1'b1;
  assign CLBLM_R_X33Y119_SLICE_X48Y119_A5 = 1'b1;
  assign CLBLM_R_X33Y125_SLICE_X48Y125_D2 = 1'b1;
  assign CLBLL_L_X34Y121_SLICE_X51Y121_C1 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_L_X34Y121_SLICE_X51Y121_C2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X34Y121_SLICE_X51Y121_C3 = CLBLM_R_X35Y122_SLICE_X53Y122_B_XOR;
  assign CLBLL_L_X34Y121_SLICE_X51Y121_C4 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X34Y121_SLICE_X51Y121_C5 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X34Y121_SLICE_X51Y121_C6 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLM_R_X33Y119_SLICE_X48Y119_A6 = 1'b1;
  assign LIOI3_X0Y121_ILOGIC_X0Y122_D = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X34Y121_SLICE_X51Y121_D1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X34Y121_SLICE_X51Y121_D2 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X34Y121_SLICE_X51Y121_D3 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X34Y121_SLICE_X51Y121_D4 = 1'b1;
  assign CLBLL_L_X34Y121_SLICE_X51Y121_D5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X34Y121_SLICE_X51Y121_D6 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign LIOI3_X0Y121_ILOGIC_X0Y121_D = LIOB33_X0Y121_IOB_X0Y121_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_D = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y145_OLOGIC_X1Y146_D1 = CLBLL_L_X36Y128_SLICE_X54Y128_AO6;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_D = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X35Y126_SLICE_X53Y126_A6 = 1'b1;
  assign CLBLM_R_X35Y126_SLICE_X53Y126_AX = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X35Y126_SLICE_X53Y126_B1 = LIOB33_X0Y139_IOB_X0Y139_I;
  assign CLBLM_R_X35Y126_SLICE_X53Y126_B2 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X35Y126_SLICE_X53Y126_B3 = 1'b1;
  assign CLBLM_R_X35Y126_SLICE_X53Y126_B4 = 1'b1;
  assign CLBLM_R_X35Y126_SLICE_X53Y126_B5 = 1'b1;
  assign CLBLM_R_X35Y126_SLICE_X53Y126_B6 = 1'b1;
  assign CLBLM_R_X35Y126_SLICE_X53Y126_BX = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X35Y126_SLICE_X53Y126_C1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X34Y122_SLICE_X50Y122_A1 = CLBLL_L_X36Y122_SLICE_X54Y122_AO5;
  assign CLBLL_L_X34Y122_SLICE_X50Y122_A2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X34Y122_SLICE_X50Y122_A3 = CLBLL_L_X34Y120_SLICE_X50Y120_AO6;
  assign CLBLL_L_X34Y122_SLICE_X50Y122_A4 = CLBLM_R_X33Y118_SLICE_X49Y118_BO6;
  assign CLBLL_L_X34Y122_SLICE_X50Y122_A5 = CLBLM_R_X33Y122_SLICE_X49Y122_BO6;
  assign CLBLL_L_X34Y122_SLICE_X50Y122_A6 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X35Y126_SLICE_X53Y126_C2 = 1'b1;
  assign CLBLM_R_X35Y126_SLICE_X53Y126_C3 = 1'b1;
  assign CLBLL_L_X34Y122_SLICE_X50Y122_B1 = CLBLL_L_X34Y122_SLICE_X50Y122_DO6;
  assign CLBLL_L_X34Y122_SLICE_X50Y122_B2 = CLBLL_L_X34Y128_SLICE_X50Y128_AO6;
  assign CLBLL_L_X34Y122_SLICE_X50Y122_B3 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLL_L_X34Y122_SLICE_X50Y122_B4 = CLBLM_R_X35Y122_SLICE_X53Y122_D_XOR;
  assign CLBLL_L_X34Y122_SLICE_X50Y122_B5 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X34Y122_SLICE_X50Y122_B6 = CLBLL_L_X34Y122_SLICE_X50Y122_CO6;
  assign CLBLM_R_X35Y126_SLICE_X53Y126_C4 = 1'b1;
  assign CLBLM_R_X35Y126_SLICE_X53Y126_C5 = 1'b1;
  assign CLBLL_L_X34Y122_SLICE_X50Y122_C1 = CLBLM_R_X35Y117_SLICE_X53Y117_AO6;
  assign CLBLL_L_X34Y122_SLICE_X50Y122_C2 = CLBLL_L_X36Y122_SLICE_X54Y122_AO5;
  assign CLBLL_L_X34Y122_SLICE_X50Y122_C3 = CLBLL_L_X34Y120_SLICE_X50Y120_AO6;
  assign CLBLL_L_X34Y122_SLICE_X50Y122_C4 = CLBLL_L_X36Y123_SLICE_X54Y123_AO6;
  assign CLBLL_L_X34Y122_SLICE_X50Y122_C5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X34Y122_SLICE_X50Y122_C6 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X35Y126_SLICE_X53Y126_C6 = LIOB33_X0Y139_IOB_X0Y140_I;
  assign CLBLM_R_X35Y126_SLICE_X53Y126_CIN = CLBLM_R_X35Y125_SLICE_X53Y125_D_CY;
  assign CLBLL_L_X34Y122_SLICE_X50Y122_D1 = CLBLM_R_X35Y117_SLICE_X52Y117_BO6;
  assign CLBLL_L_X34Y122_SLICE_X50Y122_D2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X34Y122_SLICE_X50Y122_D3 = CLBLL_L_X34Y118_SLICE_X51Y118_BO6;
  assign CLBLL_L_X34Y122_SLICE_X50Y122_D4 = CLBLM_R_X35Y122_SLICE_X53Y122_D_XOR;
  assign CLBLL_L_X34Y122_SLICE_X50Y122_D5 = 1'b1;
  assign CLBLL_L_X34Y122_SLICE_X50Y122_D6 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X35Y126_SLICE_X53Y126_CX = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X34Y122_SLICE_X51Y122_A1 = CLBLL_L_X34Y122_SLICE_X51Y122_DO6;
  assign CLBLL_L_X34Y122_SLICE_X51Y122_A2 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X34Y122_SLICE_X51Y122_A3 = CLBLL_L_X34Y122_SLICE_X51Y122_BO6;
  assign CLBLL_L_X34Y122_SLICE_X51Y122_A4 = CLBLL_L_X34Y128_SLICE_X50Y128_AO6;
  assign CLBLL_L_X34Y122_SLICE_X51Y122_A5 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLL_L_X34Y122_SLICE_X51Y122_A6 = CLBLM_R_X35Y123_SLICE_X53Y123_A_XOR;
  assign CLBLM_R_X35Y126_SLICE_X53Y126_D1 = 1'b1;
  assign CLBLM_R_X35Y126_SLICE_X53Y126_D2 = 1'b1;
  assign CLBLL_L_X34Y122_SLICE_X51Y122_B1 = CLBLM_R_X33Y123_SLICE_X49Y123_DO6;
  assign CLBLL_L_X34Y122_SLICE_X51Y122_B2 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X34Y122_SLICE_X51Y122_B3 = CLBLM_R_X35Y117_SLICE_X53Y117_AO6;
  assign CLBLL_L_X34Y122_SLICE_X51Y122_B4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X34Y122_SLICE_X51Y122_B5 = CLBLL_L_X34Y119_SLICE_X51Y119_BO6;
  assign CLBLL_L_X34Y122_SLICE_X51Y122_B6 = CLBLL_L_X36Y123_SLICE_X54Y123_AO6;
  assign CLBLM_R_X35Y126_SLICE_X53Y126_D3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X35Y126_SLICE_X53Y126_D4 = 1'b1;
  assign CLBLL_L_X34Y122_SLICE_X51Y122_C1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X34Y122_SLICE_X51Y122_C2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X34Y122_SLICE_X51Y122_C3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X34Y122_SLICE_X51Y122_C4 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X34Y122_SLICE_X51Y122_C5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X34Y122_SLICE_X51Y122_C6 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X35Y126_SLICE_X53Y126_D5 = 1'b1;
  assign CLBLM_R_X35Y126_SLICE_X53Y126_D6 = LIOB33_X0Y141_IOB_X0Y141_I;
  assign CLBLL_L_X34Y122_SLICE_X51Y122_D1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X34Y122_SLICE_X51Y122_D2 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X34Y122_SLICE_X51Y122_D3 = 1'b1;
  assign CLBLL_L_X34Y122_SLICE_X51Y122_D4 = CLBLM_R_X35Y123_SLICE_X53Y123_A_XOR;
  assign CLBLL_L_X34Y122_SLICE_X51Y122_D5 = CLBLL_L_X36Y117_SLICE_X55Y117_CO6;
  assign CLBLL_L_X34Y122_SLICE_X51Y122_D6 = CLBLL_L_X34Y118_SLICE_X51Y118_BO6;
  assign CLBLM_R_X37Y126_SLICE_X57Y126_B1 = CLBLM_R_X37Y126_SLICE_X57Y126_DO6;
  assign CLBLM_R_X37Y126_SLICE_X57Y126_B2 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLM_R_X35Y126_SLICE_X53Y126_DX = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X37Y126_SLICE_X57Y126_B3 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X37Y126_SLICE_X57Y126_B4 = CLBLM_R_X35Y125_SLICE_X53Y125_D_XOR;
  assign CLBLM_R_X37Y126_SLICE_X57Y126_B5 = CLBLM_R_X35Y123_SLICE_X52Y123_D_XOR;
  assign CLBLM_R_X37Y126_SLICE_X57Y126_B6 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_R_X35Y126_SLICE_X52Y126_A1 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLM_R_X35Y126_SLICE_X52Y126_A2 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_R_X35Y126_SLICE_X52Y126_A3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X35Y126_SLICE_X52Y126_A4 = LIOB33_X0Y137_IOB_X0Y138_I;
  assign CLBLM_R_X37Y126_SLICE_X57Y126_C1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X35Y126_SLICE_X52Y126_A5 = CLBLM_R_X35Y126_SLICE_X53Y126_A_XOR;
  assign CLBLM_R_X37Y126_SLICE_X57Y126_C2 = 1'b1;
  assign CLBLM_R_X35Y126_SLICE_X52Y126_A6 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X37Y126_SLICE_X57Y126_C4 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X37Y126_SLICE_X57Y126_C5 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X37Y126_SLICE_X57Y126_C6 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X35Y126_SLICE_X52Y126_B1 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLM_R_X35Y126_SLICE_X52Y126_B2 = LIOB33_X0Y139_IOB_X0Y140_I;
  assign CLBLM_R_X35Y126_SLICE_X52Y126_B3 = CLBLL_L_X36Y126_SLICE_X54Y126_BO6;
  assign CLBLM_R_X35Y126_SLICE_X52Y126_B4 = CLBLL_L_X36Y116_SLICE_X55Y116_AO5;
  assign CLBLM_R_X35Y126_SLICE_X52Y126_B5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X35Y126_SLICE_X52Y126_B6 = CLBLM_R_X35Y126_SLICE_X52Y126_CO6;
  assign CLBLM_R_X37Y126_SLICE_X57Y126_D3 = 1'b1;
  assign CLBLM_R_X37Y126_SLICE_X57Y126_D4 = 1'b1;
  assign CLBLM_R_X35Y126_SLICE_X52Y126_C1 = CLBLM_R_X35Y124_SLICE_X52Y124_C_XOR;
  assign CLBLM_R_X37Y126_SLICE_X57Y126_D5 = 1'b1;
  assign CLBLM_R_X35Y126_SLICE_X52Y126_C2 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLM_R_X37Y126_SLICE_X57Y126_D6 = LIOB33_X0Y137_IOB_X0Y137_I;
  assign CLBLM_R_X35Y126_SLICE_X52Y126_C3 = CLBLM_R_X35Y126_SLICE_X53Y126_C_XOR;
  assign CLBLM_R_X35Y126_SLICE_X52Y126_C4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X35Y126_SLICE_X52Y126_C5 = CLBLM_R_X35Y126_SLICE_X52Y126_DO6;
  assign CLBLM_R_X35Y126_SLICE_X52Y126_C6 = CLBLL_L_X36Y122_SLICE_X55Y122_AO6;
  assign CLBLM_R_X37Y126_SLICE_X56Y126_A1 = CLBLM_R_X37Y126_SLICE_X56Y126_DO6;
  assign LIOI3_SING_X0Y100_ILOGIC_X0Y100_D = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X37Y126_SLICE_X56Y126_A2 = 1'b1;
  assign CLBLM_R_X37Y126_SLICE_X56Y126_A3 = CLBLM_R_X37Y126_SLICE_X57Y126_CO6;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_A2 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_A3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_A4 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_A5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_A6 = 1'b1;
  assign CLBLM_R_X37Y126_SLICE_X56Y126_A4 = CLBLM_R_X37Y123_SLICE_X56Y123_DO6;
  assign CLBLM_R_X37Y126_SLICE_X56Y126_A5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_B1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_B2 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_B3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_B4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_B5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_B6 = 1'b1;
  assign CLBLM_R_X37Y126_SLICE_X56Y126_A6 = 1'b1;
  assign CLBLM_R_X35Y126_SLICE_X52Y126_D1 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_C1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_C2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_C3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_C4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_C5 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_C6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X35Y126_SLICE_X52Y126_D2 = CLBLM_R_X35Y126_SLICE_X53Y126_C_XOR;
  assign CLBLM_R_X35Y126_SLICE_X52Y126_D3 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLM_R_X35Y129_SLICE_X52Y129_D2 = 1'b1;
  assign CLBLM_R_X35Y126_SLICE_X52Y126_D4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_D1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_D2 = CLBLM_R_X33Y125_SLICE_X49Y125_BO6;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_D3 = CLBLM_L_X32Y123_SLICE_X47Y123_AO6;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_D4 = CLBLL_L_X34Y123_SLICE_X50Y123_CO6;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_D5 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X50Y123_D6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X35Y126_SLICE_X52Y126_D5 = LIOB33_X0Y139_IOB_X0Y140_I;
  assign CLBLM_R_X37Y121_SLICE_X57Y121_A5 = LIOB33_X0Y129_IOB_X0Y130_I;
  assign CLBLM_R_X35Y126_SLICE_X52Y126_D6 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X37Y121_SLICE_X57Y121_A6 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X37Y126_SLICE_X56Y126_B1 = CLBLM_R_X37Y127_SLICE_X56Y127_CO6;
  assign CLBLM_R_X37Y126_SLICE_X56Y126_B2 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign RIOI3_X105Y135_OLOGIC_X1Y136_D1 = CLBLM_R_X37Y123_SLICE_X57Y123_AO6;
  assign CLBLM_R_X35Y121_SLICE_X53Y121_D5 = 1'b1;
  assign CLBLM_R_X37Y126_SLICE_X56Y126_B3 = CLBLM_R_X35Y127_SLICE_X53Y127_C_XOR;
  assign CLBLM_R_X35Y121_SLICE_X53Y121_D6 = 1'b1;
  assign CLBLM_R_X37Y126_SLICE_X56Y126_B4 = CLBLL_L_X34Y128_SLICE_X50Y128_AO6;
  assign RIOI3_X105Y135_OLOGIC_X1Y136_T1 = 1'b1;
  assign CLBLM_R_X37Y126_SLICE_X56Y126_B5 = CLBLM_R_X35Y128_SLICE_X52Y128_AO6;
  assign CLBLM_R_X37Y121_SLICE_X57Y121_B1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X37Y126_SLICE_X56Y126_B6 = CLBLM_R_X37Y126_SLICE_X56Y126_CO6;
  assign CLBLM_R_X37Y121_SLICE_X57Y121_B2 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_D1 = CLBLM_R_X37Y123_SLICE_X56Y123_AO6;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_A1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_A2 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_A3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_A4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_A5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_A6 = 1'b1;
  assign CLBLM_R_X35Y121_SLICE_X53Y121_DX = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X37Y121_SLICE_X57Y121_B3 = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLM_R_X37Y121_SLICE_X57Y121_B4 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_D = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_B1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_B2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_B3 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_B4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_B5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_B6 = 1'b1;
  assign CLBLM_R_X37Y121_SLICE_X57Y121_B5 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X37Y124_SLICE_X56Y124_B4 = CLBLM_R_X35Y125_SLICE_X53Y125_A_XOR;
  assign CLBLM_R_X37Y121_SLICE_X57Y121_B6 = CLBLM_R_X37Y121_SLICE_X57Y121_CO6;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_C1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_C2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_C3 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_C4 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_C5 = LIOB33_X0Y119_IOB_X0Y119_I;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_C6 = 1'b1;
  assign CLBLM_R_X37Y126_SLICE_X56Y126_C1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X37Y126_SLICE_X56Y126_C2 = CLBLM_R_X37Y125_SLICE_X56Y125_CO6;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_D1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_D2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_D3 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_D4 = 1'b1;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_D5 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLL_L_X34Y123_SLICE_X51Y123_D6 = 1'b1;
  assign CLBLM_R_X37Y126_SLICE_X56Y126_C3 = CLBLL_L_X34Y127_SLICE_X50Y127_AO6;
  assign CLBLM_R_X37Y126_SLICE_X56Y126_C4 = CLBLL_L_X34Y126_SLICE_X50Y126_DO6;
  assign CLBLM_R_X37Y121_SLICE_X57Y121_C1 = CLBLM_R_X35Y124_SLICE_X53Y124_B_XOR;
  assign CLBLM_R_X37Y126_SLICE_X56Y126_C5 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X37Y121_SLICE_X57Y121_C2 = CLBLM_R_X35Y122_SLICE_X52Y122_B_XOR;
  assign CLBLM_R_X37Y123_SLICE_X57Y123_A4 = CLBLL_L_X36Y116_SLICE_X55Y116_AO5;
  assign CLBLM_R_X37Y125_SLICE_X56Y125_C4 = CLBLL_L_X36Y121_SLICE_X54Y121_AO5;
  assign CLBLM_R_X37Y126_SLICE_X56Y126_C6 = CLBLL_L_X36Y122_SLICE_X55Y122_AO5;
  assign CLBLM_R_X37Y121_SLICE_X57Y121_C3 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X37Y121_SLICE_X57Y121_C4 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_R_X37Y121_SLICE_X57Y121_C5 = CLBLM_R_X37Y121_SLICE_X57Y121_DO6;
  assign CLBLM_R_X37Y121_SLICE_X57Y121_C6 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLM_R_X37Y126_SLICE_X56Y126_D1 = 1'b1;
  assign CLBLM_R_X35Y116_SLICE_X53Y116_B3 = LIOB33_X0Y119_IOB_X0Y119_I;
  assign CLBLM_R_X37Y126_SLICE_X56Y126_D2 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X35Y116_SLICE_X53Y116_B4 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLM_R_X37Y126_SLICE_X56Y126_D3 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X37Y121_SLICE_X57Y121_D1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X35Y116_SLICE_X53Y116_B5 = CLBLL_L_X34Y116_SLICE_X51Y116_CO6;
  assign CLBLM_R_X37Y126_SLICE_X56Y126_D4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X37Y121_SLICE_X57Y121_D2 = 1'b1;
  assign CLBLM_R_X35Y116_SLICE_X53Y116_B6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X37Y126_SLICE_X56Y126_D5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X37Y126_SLICE_X56Y126_D6 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X37Y121_SLICE_X57Y121_D4 = LIOB33_X0Y127_IOB_X0Y128_I;
  assign CLBLM_R_X37Y124_SLICE_X56Y124_B5 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_L_X32Y116_SLICE_X47Y116_A1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X32Y116_SLICE_X47Y116_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X32Y116_SLICE_X47Y116_A3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_L_X32Y116_SLICE_X47Y116_A4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X32Y116_SLICE_X47Y116_A5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X32Y116_SLICE_X47Y116_A6 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X37Y121_SLICE_X57Y121_D5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X37Y121_SLICE_X57Y121_D6 = 1'b1;
  assign CLBLM_L_X32Y116_SLICE_X47Y116_B1 = 1'b1;
  assign CLBLM_L_X32Y116_SLICE_X47Y116_B2 = 1'b1;
  assign CLBLM_L_X32Y116_SLICE_X47Y116_B3 = 1'b1;
  assign CLBLM_L_X32Y116_SLICE_X47Y116_B4 = 1'b1;
  assign CLBLM_L_X32Y116_SLICE_X47Y116_B5 = 1'b1;
  assign CLBLM_L_X32Y116_SLICE_X47Y116_B6 = 1'b1;
  assign LIOI3_X0Y123_ILOGIC_X0Y124_D = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLM_L_X32Y116_SLICE_X47Y116_C1 = 1'b1;
  assign CLBLM_L_X32Y116_SLICE_X47Y116_C2 = 1'b1;
  assign CLBLM_L_X32Y116_SLICE_X47Y116_C3 = 1'b1;
  assign CLBLM_L_X32Y116_SLICE_X47Y116_C4 = 1'b1;
  assign CLBLM_L_X32Y116_SLICE_X47Y116_C5 = 1'b1;
  assign CLBLM_L_X32Y116_SLICE_X47Y116_C6 = 1'b1;
  assign LIOI3_X0Y123_ILOGIC_X0Y123_D = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLM_L_X32Y116_SLICE_X47Y116_D1 = 1'b1;
  assign CLBLM_L_X32Y116_SLICE_X47Y116_D2 = 1'b1;
  assign CLBLM_L_X32Y116_SLICE_X47Y116_D3 = 1'b1;
  assign CLBLM_L_X32Y116_SLICE_X47Y116_D4 = 1'b1;
  assign CLBLM_L_X32Y116_SLICE_X47Y116_D5 = 1'b1;
  assign CLBLM_L_X32Y116_SLICE_X47Y116_D6 = 1'b1;
  assign CLBLM_L_X32Y116_SLICE_X46Y116_A1 = 1'b1;
  assign CLBLM_L_X32Y116_SLICE_X46Y116_A2 = 1'b1;
  assign CLBLM_L_X32Y116_SLICE_X46Y116_A3 = 1'b1;
  assign CLBLM_L_X32Y116_SLICE_X46Y116_A4 = 1'b1;
  assign CLBLM_L_X32Y116_SLICE_X46Y116_A5 = 1'b1;
  assign CLBLM_L_X32Y116_SLICE_X46Y116_A6 = 1'b1;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_D = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_D = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X32Y116_SLICE_X46Y116_B1 = 1'b1;
  assign CLBLM_L_X32Y116_SLICE_X46Y116_B2 = 1'b1;
  assign CLBLM_L_X32Y116_SLICE_X46Y116_B3 = 1'b1;
  assign CLBLM_L_X32Y116_SLICE_X46Y116_B4 = 1'b1;
  assign CLBLM_L_X32Y116_SLICE_X46Y116_B5 = 1'b1;
  assign CLBLM_L_X32Y116_SLICE_X46Y116_B6 = 1'b1;
  assign CLBLM_R_X37Y121_SLICE_X56Y121_A4 = CLBLM_R_X37Y121_SLICE_X56Y121_BO6;
  assign CLBLM_R_X37Y121_SLICE_X56Y121_A5 = CLBLM_R_X35Y124_SLICE_X53Y124_A_XOR;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X32Y116_SLICE_X46Y116_C1 = 1'b1;
  assign CLBLM_L_X32Y116_SLICE_X46Y116_C2 = 1'b1;
  assign CLBLM_L_X32Y116_SLICE_X46Y116_C3 = 1'b1;
  assign CLBLM_L_X32Y116_SLICE_X46Y116_C4 = 1'b1;
  assign CLBLM_L_X32Y116_SLICE_X46Y116_C5 = 1'b1;
  assign CLBLM_L_X32Y116_SLICE_X46Y116_C6 = 1'b1;
  assign CLBLM_R_X37Y121_SLICE_X56Y121_A6 = CLBLM_R_X35Y122_SLICE_X52Y122_A_XOR;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D = LIOB33_X0Y107_IOB_X0Y107_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D = RIOB33_X105Y113_IOB_X1Y114_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X32Y116_SLICE_X46Y116_D1 = 1'b1;
  assign CLBLM_L_X32Y116_SLICE_X46Y116_D2 = 1'b1;
  assign CLBLM_L_X32Y116_SLICE_X46Y116_D3 = 1'b1;
  assign CLBLM_L_X32Y116_SLICE_X46Y116_D4 = 1'b1;
  assign CLBLM_L_X32Y116_SLICE_X46Y116_D5 = 1'b1;
  assign CLBLM_L_X32Y116_SLICE_X46Y116_D6 = 1'b1;
  assign LIOI3_X0Y141_ILOGIC_X0Y142_D = LIOB33_X0Y141_IOB_X0Y142_I;
  assign CLBLL_L_X34Y124_SLICE_X50Y124_A1 = CLBLL_L_X36Y116_SLICE_X55Y116_AO5;
  assign CLBLL_L_X34Y124_SLICE_X50Y124_A2 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X34Y124_SLICE_X50Y124_A3 = CLBLL_L_X34Y122_SLICE_X51Y122_AO6;
  assign CLBLL_L_X34Y124_SLICE_X50Y124_A4 = CLBLL_L_X34Y124_SLICE_X50Y124_BO6;
  assign CLBLL_L_X34Y124_SLICE_X50Y124_A5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X34Y124_SLICE_X50Y124_A6 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLM_R_X37Y121_SLICE_X56Y121_B1 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X37Y121_SLICE_X56Y121_B2 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign LIOI3_X0Y141_ILOGIC_X0Y141_D = LIOB33_X0Y141_IOB_X0Y141_I;
  assign CLBLL_L_X34Y124_SLICE_X50Y124_B1 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLL_L_X34Y124_SLICE_X50Y124_B2 = CLBLL_L_X36Y122_SLICE_X55Y122_AO6;
  assign CLBLL_L_X34Y124_SLICE_X50Y124_B3 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLL_L_X34Y124_SLICE_X50Y124_B4 = CLBLM_R_X35Y121_SLICE_X52Y121_A_XOR;
  assign CLBLL_L_X34Y124_SLICE_X50Y124_B5 = CLBLL_L_X34Y124_SLICE_X50Y124_CO6;
  assign CLBLL_L_X34Y124_SLICE_X50Y124_B6 = CLBLM_R_X35Y123_SLICE_X53Y123_A_XOR;
  assign CLBLM_R_X37Y121_SLICE_X56Y121_B3 = LIOB33_X0Y129_IOB_X0Y130_I;
  assign CLBLM_R_X37Y121_SLICE_X56Y121_B4 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_D = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X34Y124_SLICE_X50Y124_C1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X34Y124_SLICE_X50Y124_C2 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X34Y124_SLICE_X50Y124_C3 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLL_L_X34Y124_SLICE_X50Y124_C4 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X34Y124_SLICE_X50Y124_C5 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X34Y124_SLICE_X50Y124_C6 = CLBLM_R_X35Y123_SLICE_X53Y123_A_XOR;
  assign CLBLM_R_X37Y121_SLICE_X56Y121_B5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X37Y121_SLICE_X56Y121_B6 = CLBLM_R_X35Y124_SLICE_X53Y124_A_XOR;
  assign CLBLL_L_X34Y124_SLICE_X50Y124_D1 = CLBLM_R_X33Y124_SLICE_X49Y124_DO6;
  assign CLBLL_L_X34Y124_SLICE_X50Y124_D2 = CLBLL_L_X34Y123_SLICE_X50Y123_AO5;
  assign CLBLL_L_X34Y124_SLICE_X50Y124_D3 = CLBLM_R_X33Y124_SLICE_X48Y124_AO5;
  assign CLBLL_L_X34Y124_SLICE_X50Y124_D4 = CLBLM_R_X33Y125_SLICE_X49Y125_AO5;
  assign CLBLL_L_X34Y124_SLICE_X50Y124_D5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X34Y124_SLICE_X50Y124_D6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign LIOI3_SING_X0Y149_ILOGIC_X0Y149_D = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_D = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X37Y121_SLICE_X56Y121_C1 = CLBLM_R_X37Y119_SLICE_X56Y119_AO6;
  assign CLBLM_R_X37Y121_SLICE_X56Y121_C2 = CLBLM_R_X37Y118_SLICE_X56Y118_AO6;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_D = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X37Y121_SLICE_X56Y121_C3 = CLBLM_R_X37Y121_SLICE_X57Y121_BO6;
  assign CLBLL_L_X34Y124_SLICE_X51Y124_A1 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X34Y124_SLICE_X51Y124_A2 = 1'b1;
  assign CLBLL_L_X34Y124_SLICE_X51Y124_A3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X34Y124_SLICE_X51Y124_A4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X34Y124_SLICE_X51Y124_A5 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_L_X34Y124_SLICE_X51Y124_A6 = 1'b1;
  assign CLBLM_R_X37Y121_SLICE_X56Y121_C4 = CLBLL_L_X38Y121_SLICE_X58Y121_BO6;
  assign CLBLM_R_X37Y121_SLICE_X56Y121_C5 = CLBLM_R_X37Y121_SLICE_X56Y121_DO6;
  assign CLBLL_L_X34Y124_SLICE_X51Y124_B1 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_L_X34Y124_SLICE_X51Y124_B2 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X34Y124_SLICE_X51Y124_B3 = 1'b1;
  assign CLBLL_L_X34Y124_SLICE_X51Y124_B4 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLL_L_X34Y124_SLICE_X51Y124_B5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X34Y124_SLICE_X51Y124_B6 = 1'b1;
  assign CLBLM_R_X37Y121_SLICE_X56Y121_C6 = CLBLL_L_X36Y119_SLICE_X55Y119_AO6;
  assign CLBLL_L_X34Y124_SLICE_X51Y124_C1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X34Y124_SLICE_X51Y124_C2 = 1'b1;
  assign CLBLL_L_X34Y124_SLICE_X51Y124_C3 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLL_L_X34Y124_SLICE_X51Y124_C4 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X34Y124_SLICE_X51Y124_C5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X34Y124_SLICE_X51Y124_C6 = 1'b1;
  assign CLBLL_L_X34Y124_SLICE_X51Y124_CIN = CLBLL_L_X34Y123_SLICE_X51Y123_D_CY;
  assign LIOI3_TBYTESRC_X0Y143_ILOGIC_X0Y144_D = LIOB33_X0Y143_IOB_X0Y144_I;
  assign CLBLM_R_X35Y129_SLICE_X53Y129_B5 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X34Y124_SLICE_X51Y124_D1 = LIOB33_X0Y127_IOB_X0Y128_I;
  assign CLBLL_L_X34Y124_SLICE_X51Y124_D2 = LIOB33_X0Y129_IOB_X0Y129_I;
  assign CLBLL_L_X34Y124_SLICE_X51Y124_D3 = 1'b1;
  assign CLBLL_L_X34Y124_SLICE_X51Y124_D4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X34Y124_SLICE_X51Y124_D5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X34Y124_SLICE_X51Y124_D6 = 1'b1;
  assign CLBLM_R_X35Y116_SLICE_X52Y116_B3 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign LIOI3_TBYTESRC_X0Y143_ILOGIC_X0Y143_D = LIOB33_X0Y143_IOB_X0Y143_I;
  assign CLBLM_R_X35Y129_SLICE_X53Y129_B6 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X35Y116_SLICE_X52Y116_B5 = CLBLL_L_X36Y122_SLICE_X55Y122_AO6;
  assign CLBLM_R_X35Y116_SLICE_X52Y116_B6 = CLBLM_R_X35Y116_SLICE_X52Y116_CO6;
  assign CLBLM_R_X37Y121_SLICE_X56Y121_D1 = LIOB33_X0Y129_IOB_X0Y130_I;
  assign CLBLM_R_X37Y121_SLICE_X56Y121_D2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X38Y118_SLICE_X58Y118_A1 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLL_L_X38Y118_SLICE_X58Y118_A2 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X38Y118_SLICE_X58Y118_A3 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X38Y118_SLICE_X58Y118_A4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X38Y118_SLICE_X58Y118_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X38Y118_SLICE_X58Y118_A6 = 1'b1;
  assign CLBLM_R_X37Y121_SLICE_X56Y121_D3 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X37Y121_SLICE_X56Y121_D4 = CLBLL_L_X34Y127_SLICE_X50Y127_DO6;
  assign CLBLL_L_X38Y118_SLICE_X58Y118_B1 = 1'b1;
  assign CLBLL_L_X38Y118_SLICE_X58Y118_B2 = 1'b1;
  assign CLBLL_L_X38Y118_SLICE_X58Y118_B3 = 1'b1;
  assign CLBLL_L_X38Y118_SLICE_X58Y118_B4 = 1'b1;
  assign CLBLL_L_X38Y118_SLICE_X58Y118_B5 = 1'b1;
  assign CLBLL_L_X38Y118_SLICE_X58Y118_B6 = 1'b1;
  assign CLBLM_R_X37Y121_SLICE_X56Y121_D5 = CLBLM_R_X37Y122_SLICE_X56Y122_CO6;
  assign CLBLM_R_X37Y121_SLICE_X56Y121_D6 = CLBLL_L_X34Y129_SLICE_X50Y129_AO6;
  assign CLBLL_L_X38Y118_SLICE_X58Y118_C1 = 1'b1;
  assign CLBLL_L_X38Y118_SLICE_X58Y118_C2 = 1'b1;
  assign CLBLL_L_X38Y118_SLICE_X58Y118_C3 = 1'b1;
  assign CLBLL_L_X38Y118_SLICE_X58Y118_C4 = 1'b1;
  assign CLBLL_L_X38Y118_SLICE_X58Y118_C5 = 1'b1;
  assign CLBLL_L_X38Y118_SLICE_X58Y118_C6 = 1'b1;
  assign CLBLL_L_X38Y118_SLICE_X58Y118_D1 = 1'b1;
  assign CLBLL_L_X38Y118_SLICE_X58Y118_D2 = 1'b1;
  assign CLBLL_L_X38Y118_SLICE_X58Y118_D3 = 1'b1;
  assign CLBLL_L_X38Y118_SLICE_X58Y118_D4 = 1'b1;
  assign CLBLL_L_X38Y118_SLICE_X58Y118_D5 = 1'b1;
  assign CLBLL_L_X38Y118_SLICE_X58Y118_D6 = 1'b1;
  assign CLBLM_R_X35Y123_SLICE_X53Y123_C4 = 1'b1;
  assign CLBLM_L_X32Y117_SLICE_X47Y117_A1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X38Y118_SLICE_X59Y118_A1 = 1'b1;
  assign CLBLL_L_X38Y118_SLICE_X59Y118_A2 = 1'b1;
  assign CLBLL_L_X38Y118_SLICE_X59Y118_A3 = 1'b1;
  assign CLBLM_L_X32Y117_SLICE_X47Y117_A5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_L_X32Y117_SLICE_X47Y117_A6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X38Y118_SLICE_X59Y118_A4 = 1'b1;
  assign CLBLL_L_X38Y118_SLICE_X59Y118_A5 = 1'b1;
  assign CLBLL_L_X38Y118_SLICE_X59Y118_A6 = 1'b1;
  assign CLBLM_L_X32Y117_SLICE_X47Y117_A2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_L_X32Y117_SLICE_X47Y117_A3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X32Y117_SLICE_X47Y117_B3 = 1'b1;
  assign CLBLM_L_X32Y117_SLICE_X47Y117_B4 = 1'b1;
  assign CLBLM_L_X32Y117_SLICE_X47Y117_B5 = 1'b1;
  assign CLBLM_L_X32Y117_SLICE_X47Y117_B6 = 1'b1;
  assign CLBLL_L_X38Y118_SLICE_X59Y118_B1 = 1'b1;
  assign CLBLL_L_X38Y118_SLICE_X59Y118_B2 = 1'b1;
  assign CLBLL_L_X38Y118_SLICE_X59Y118_B3 = 1'b1;
  assign CLBLL_L_X38Y118_SLICE_X59Y118_B4 = 1'b1;
  assign CLBLL_L_X38Y118_SLICE_X59Y118_B5 = 1'b1;
  assign CLBLL_L_X38Y118_SLICE_X59Y118_B6 = 1'b1;
  assign CLBLM_L_X32Y117_SLICE_X47Y117_C4 = 1'b1;
  assign CLBLM_L_X32Y117_SLICE_X47Y117_C5 = 1'b1;
  assign CLBLL_L_X38Y118_SLICE_X59Y118_C1 = 1'b1;
  assign CLBLL_L_X38Y118_SLICE_X59Y118_C2 = 1'b1;
  assign CLBLL_L_X38Y118_SLICE_X59Y118_C3 = 1'b1;
  assign CLBLL_L_X38Y118_SLICE_X59Y118_C4 = 1'b1;
  assign CLBLL_L_X38Y118_SLICE_X59Y118_C5 = 1'b1;
  assign CLBLL_L_X38Y118_SLICE_X59Y118_C6 = 1'b1;
  assign CLBLM_L_X32Y117_SLICE_X47Y117_C6 = 1'b1;
  assign CLBLM_L_X32Y117_SLICE_X47Y117_D1 = 1'b1;
  assign CLBLM_L_X32Y117_SLICE_X47Y117_D2 = 1'b1;
  assign CLBLM_L_X32Y117_SLICE_X47Y117_D3 = 1'b1;
  assign CLBLM_L_X32Y117_SLICE_X47Y117_D4 = 1'b1;
  assign CLBLM_L_X32Y117_SLICE_X47Y117_D5 = 1'b1;
  assign CLBLM_L_X32Y117_SLICE_X47Y117_D6 = 1'b1;
  assign CLBLL_L_X38Y118_SLICE_X59Y118_D4 = 1'b1;
  assign CLBLL_L_X38Y118_SLICE_X59Y118_D1 = 1'b1;
  assign CLBLL_L_X38Y118_SLICE_X59Y118_D2 = 1'b1;
  assign CLBLL_L_X38Y118_SLICE_X59Y118_D3 = 1'b1;
  assign CLBLL_L_X38Y118_SLICE_X59Y118_D5 = 1'b1;
  assign CLBLM_L_X32Y117_SLICE_X46Y117_A1 = 1'b1;
  assign CLBLM_L_X32Y117_SLICE_X46Y117_A2 = 1'b1;
  assign CLBLM_L_X32Y117_SLICE_X46Y117_A3 = 1'b1;
  assign CLBLM_L_X32Y117_SLICE_X46Y117_A4 = 1'b1;
  assign CLBLM_L_X32Y117_SLICE_X46Y117_A5 = 1'b1;
  assign CLBLM_L_X32Y117_SLICE_X46Y117_A6 = 1'b1;
  assign CLBLM_R_X35Y129_SLICE_X53Y129_C1 = 1'b1;
  assign CLBLM_R_X33Y125_SLICE_X49Y125_B3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X32Y117_SLICE_X46Y117_B1 = 1'b1;
  assign CLBLM_L_X32Y117_SLICE_X46Y117_B2 = 1'b1;
  assign CLBLM_L_X32Y117_SLICE_X46Y117_B3 = 1'b1;
  assign CLBLM_L_X32Y117_SLICE_X46Y117_B4 = 1'b1;
  assign CLBLM_L_X32Y117_SLICE_X46Y117_B5 = 1'b1;
  assign CLBLM_L_X32Y117_SLICE_X46Y117_B6 = 1'b1;
  assign CLBLM_R_X33Y125_SLICE_X49Y125_B4 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X33Y125_SLICE_X49Y125_B5 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_L_X32Y117_SLICE_X46Y117_C1 = 1'b1;
  assign CLBLM_L_X32Y117_SLICE_X46Y117_C2 = 1'b1;
  assign CLBLM_L_X32Y117_SLICE_X46Y117_C3 = 1'b1;
  assign CLBLM_L_X32Y117_SLICE_X46Y117_C4 = 1'b1;
  assign CLBLM_L_X32Y117_SLICE_X46Y117_C5 = 1'b1;
  assign CLBLM_L_X32Y117_SLICE_X46Y117_C6 = 1'b1;
  assign CLBLM_R_X33Y125_SLICE_X49Y125_B6 = 1'b1;
  assign CLBLM_R_X35Y129_SLICE_X53Y129_C2 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_A1 = 1'b1;
  assign CLBLM_L_X32Y117_SLICE_X46Y117_D1 = 1'b1;
  assign CLBLM_L_X32Y117_SLICE_X46Y117_D2 = 1'b1;
  assign CLBLM_L_X32Y117_SLICE_X46Y117_D3 = 1'b1;
  assign CLBLM_L_X32Y117_SLICE_X46Y117_D4 = 1'b1;
  assign CLBLM_L_X32Y117_SLICE_X46Y117_D5 = 1'b1;
  assign CLBLM_L_X32Y117_SLICE_X46Y117_D6 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_A2 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_A3 = 1'b1;
  assign CLBLM_R_X35Y129_SLICE_X53Y129_C3 = 1'b1;
  assign CLBLL_L_X34Y125_SLICE_X50Y125_A1 = CLBLM_R_X33Y125_SLICE_X49Y125_AO5;
  assign CLBLL_L_X34Y125_SLICE_X50Y125_A2 = CLBLM_R_X33Y124_SLICE_X49Y124_DO6;
  assign CLBLL_L_X34Y125_SLICE_X50Y125_A3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X34Y125_SLICE_X50Y125_A4 = CLBLL_L_X34Y123_SLICE_X50Y123_AO5;
  assign CLBLL_L_X34Y125_SLICE_X50Y125_A5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X34Y125_SLICE_X50Y125_A6 = CLBLM_R_X33Y125_SLICE_X49Y125_DO6;
  assign CLBLM_R_X33Y125_SLICE_X49Y125_C1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X33Y125_SLICE_X49Y125_C2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_B4 = 1'b1;
  assign CLBLL_L_X34Y125_SLICE_X50Y125_B1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X34Y125_SLICE_X50Y125_B2 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X34Y125_SLICE_X50Y125_B3 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X34Y125_SLICE_X50Y125_B4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X34Y125_SLICE_X50Y125_B5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X34Y125_SLICE_X50Y125_B6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X33Y125_SLICE_X49Y125_C3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_C2 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_C4 = 1'b1;
  assign CLBLL_L_X34Y125_SLICE_X50Y125_C1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X34Y125_SLICE_X50Y125_C2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X34Y125_SLICE_X50Y125_C3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X34Y125_SLICE_X50Y125_C4 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X34Y125_SLICE_X50Y125_C5 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X34Y125_SLICE_X50Y125_C6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X35Y123_SLICE_X53Y123_C5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X35Y129_SLICE_X53Y129_C4 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_D1 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_D2 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_D3 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_D4 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_D5 = 1'b1;
  assign CLBLL_L_X34Y125_SLICE_X50Y125_D1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X34Y125_SLICE_X50Y125_D2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X34Y125_SLICE_X50Y125_D3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X34Y125_SLICE_X50Y125_D4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X34Y125_SLICE_X50Y125_D5 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X34Y125_SLICE_X50Y125_D6 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_A2 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_A3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_A4 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_A5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_A6 = 1'b1;
  assign CLBLM_R_X35Y129_SLICE_X53Y129_C5 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_B1 = 1'b1;
  assign CLBLM_R_X35Y129_SLICE_X52Y129_D3 = 1'b1;
endmodule
