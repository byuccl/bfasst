
module chip (input \sum_o[14] , input io_0_3_0, input io_0_3_1, input io_0_4_0, input io_0_4_1, input \a_i[15] , output \b_i[14] , output io_0_6_0, output io_0_6_1, output io_0_7_1, output \b_i[15] , output \sum_o[11] , output \sum_o[12] , output \sum_o[13] , output \b_i[13] , output \sum_o[9] , output \a_i[14] , input \sum_o[10] , input io_0_14_0, input \sum_o[3] , input \b_i[2] , input \a_i[5] , input \b_i[0] , output \a_i[0] , input \sum_o[4] , output \sum_o[7] , output \sum_o[8] , input \a_i[6] , input \a_i[8] , input \sum_o[2] , input \sum_o[0] , input \b_i[7] , input \a_i[7] , output \sum_o[6] , output \a_i[1] , output \a_i[9] , input \sum_o[5] , input \b_i[10] , input clk_i, input \b_i[8] , input \a_i[4] , input \b_i[11] , input \b_i[4] , input \b_i[6] , input \a_i[10] , input \a_i[12] , input \a_i[11] , input \b_i[9] , input io_3_33_0, input \b_i[1] , input io_4_33_0, input \sum_o[1] , input \b_i[5] , input \sum_o[15] , input \b_i[12] , input \a_i[13] , input \b_i[3] , input cin_i, input \a_i[2] , input cout_o, input \a_i[3] );

wire \sum_o[14] , io_0_3_0, io_0_3_1, io_0_4_0, io_0_4_1, \a_i[15] , \sum_o[10] , io_0_14_0, \sum_o[3] , n30;
wire n31, n32, \b_i[2] , \a_i[5] , \b_i[0] , n37, n38, n41, \sum_o[4] , n49;
wire \a_i[6] , \a_i[8] , \sum_o[2] , n57, \sum_o[0] , \b_i[7] , \a_i[7] , \sum_o[5] , \b_i[10] , clk_i;
wire \b_i[8] , \a_i[4] , \b_i[11] , \b_i[4] , \b_i[6] , \a_i[10] , n75, n77, n78, n79;
wire n80, n81, n82, \a_i[12] , n84, n85, n86, n87, n88, n89;
wire n90, n91, n92, n97, n99, n100, n101, n102, \a_i[11] , \b_i[9] ;
wire n108, n109, n110, n111, n112, n113, n114, n115, n116, n117;
wire n118, n119, n121, n122, n123, n124, n125, n126, n127, n128;
wire io_3_33_0, n132, n133, n134, \b_i[1] , io_4_33_0, n137, n138, n139, n140;
wire n141, n142, n143, n144, n145, n146, n147, n148, n149, n150;
wire n151, n152, n153, n154, n155, n156, n157, n158, n159, n160;
wire n161, n162, n163, n164, n165, n166, n167, n168, n169, n170;
wire n171, n172, n173, n174, n175, n176, n177, n178, n179, n180;
wire n181, n182, n183, n184, n185, n186, n187, n188, n189, n190;
wire n191, n192, n193, n194, n195, n196, n197, n198, n199, n200;
wire n201, n202, n203, n204, n205, n206, n207, n208, n209, n210;
wire n211, n212, n213, n214, n215, n216, n217, n218;
reg \b_i[14]  = 0, io_0_6_0 = 0, io_0_6_1 = 0, io_0_7_1 = 0, \b_i[15]  = 0, \sum_o[11]  = 0, \sum_o[12]  = 0, \sum_o[13]  = 0, \b_i[13]  = 0, \sum_o[9]  = 0;
reg \a_i[14]  = 0, n19 = 0, n22 = 0, n23 = 0, n24 = 0, n25 = 0, n26 = 0, n27 = 0, n28 = 0, n29 = 0;
reg n36 = 0, \a_i[0]  = 0, n40 = 0, n43 = 0, \sum_o[7]  = 0, \sum_o[8]  = 0, n46 = 0, n47 = 0, n48 = 0, n53 = 0;
reg n54 = 0, n55 = 0, n56 = 0, n58 = 0, \sum_o[6]  = 0, \a_i[1]  = 0, \a_i[9]  = 0, n74 = 0, n76 = 0, n93 = 0;
reg n94 = 0, n95 = 0, n96 = 0, n98 = 0, n103 = 0, n104 = 0, n105 = 0, n120 = 0, n129 = 0, n130 = 0;
assign n160 = 0;

assign n159 = /* LUT    2 16  0 */ 1'b0;
assign n137 = /* LUT    3 16  0 */ !n120;
assign n138 = /* LUT    1 19  0 */ \b_i[4] ;
assign n139 = /* LUT    1 15  6 */ \sum_o[3] ;
assign n140 = /* LUT    1 16  6 */ !n26;
assign n141 = /* LUT    2 19  0 */ \b_i[6] ;
assign n142 = /* LUT    2 16  5 */ (n115 ? (n22 ? n103 : !n103) : (n22 ? !n103 : n103));
assign n143 = /* LUT    1 15  5 */ io_0_4_0;
assign n144 = /* LUT    1 16  7 */ (n24 ? n26 : !n26);
assign n145 = /* LUT    2 16  4 */ (n114 ? (n38 ? n96 : !n96) : (n38 ? !n96 : n96));
assign n146 = /* LUT    1 15  4 */ io_0_14_0;
assign n88  = /* LUT    1 16  4 */ (n86 ? (n55 ? n54 : !n54) : (n55 ? !n54 : n54));
assign n148 = /* LUT    2 19  2 */ \b_i[7] ;
assign n149 = /* LUT    1 14  7 */ io_0_3_1;
assign n150 = /* LUT    2 16  7 */ (n117 ? (n110 ? n40 : !n40) : (n110 ? !n40 : n40));
assign n151 = /* LUT    1 16  5 */ (n85 ? (n88 ? 1'b1 : (n87 ? n84 : 1'b0)) : 1'b0);
assign n152 = /* LUT    2 19  7 */ \a_i[10] ;
assign n153 = /* LUT    2 16  6 */ (n116 ? (n109 ? n29 : !n29) : (n109 ? !n29 : n29));
assign n154 = /* LUT    2 16  1 */ (n111 ? (n76 ? n25 : !n25) : (n76 ? !n25 : n25));
assign n155 = /* LUT    2 17  6 */ (n126 ? (n94 ? n31 : !n31) : (n94 ? !n31 : n31));
assign n156 = /* LUT    1 18  0 */ \a_i[8] ;
assign n157 = /* LUT    2 18  4 */ (n82 ? (n134 ? 1'b1 : !n81) : (n134 ? 1'b0 : n81));
assign n161 = /* LUT    3 17  7 */ \b_i[1] ;
assign n162 = /* LUT    2 17  7 */ (n127 ? (n32 ? n23 : !n23) : (n32 ? !n23 : n23));
assign n163 = /* LUT    1 18  1 */ (n91 ? (n92 ? n97 : !n97) : n92);
assign n164 = /* LUT    3 17  6 */ \b_i[10] ;
assign n165 = /* LUT    2 16  3 */ (n113 ? (n37 ? n95 : !n95) : (n37 ? !n95 : n95));
assign n166 = /* LUT    1 18  2 */ n90;
assign n167 = /* LUT    2 17  4 */ (n124 ? (n49 ? n53 : !n53) : (n49 ? !n53 : n53));
assign n168 = /* LUT    3 17  5 */ (n100 ? n89 : (n81 ? (n89 ? n82 : 1'b0) : 1'b0));
assign n169 = /* LUT    2 16  2 */ (n112 ? (n41 ? n36 : !n36) : (n41 ? !n36 : n36));
assign n170 = /* LUT    3 17  4 */ (n130 ? n120 : !n120);
assign n171 = /* LUT    1 18  3 */ \b_i[9] ;
assign n172 = /* LUT    2 17  5 */ (n125 ? (n55 ? n54 : !n54) : (n55 ? !n54 : n54));
assign n173 = /* LUT    2 15  0 */ \a_i[12] ;
assign n174 = /* LUT    1 18  4 */ n97;
assign n175 = /* LUT    2 17  2 */ (n122 ? (n102 ? n27 : !n27) : (n102 ? !n27 : n27));
assign n176 = /* LUT    3 17  3 */ (n129 ? 1'b1 : (n130 ? 1'b1 : n120));
assign n177 = /* LUT    2 15  1 */ (n75 ? n79 : (n77 ? (n79 ? n78 : 1'b0) : 1'b0));
assign n178 = /* LUT    1 17  1 */ (n91 ? n97 : !n97);
assign n134 = /* LUT    2 18  3 */ (n90 ? (n47 ? n43 : !n43) : (n47 ? !n43 : n43));
assign n179 = /* LUT    3 18  3 */ \sum_o[0] ;
assign n180 = /* LUT    1 18  5 */ \sum_o[2] ;
assign n181 = /* LUT    2 17  3 */ (n123 ? (n101 ? n104 : !n104) : (n101 ? !n104 : n104));
assign n182 = /* LUT    2 15  2 */ (n22 ? (n77 ? (n103 ? n80 : !n80) : (n103 ? !n80 : n80)) : (n77 ? (n103 ? !n80 : n80) : (n103 ? n80 : !n80)));
assign n183 = /* LUT    2 18  2 */ (n99 ? (n133 ? 1'b1 : (n92 ? n91 : 1'b0)) : 1'b0);
assign n184 = /* LUT    1 17  0 */ (n86 ? (n57 ? (n87 ? !n84 : n84) : n87) : (n57 ? n87 : (n87 ? !n84 : n84)));
assign n185 = /* LUT    1 19  7 */ \b_i[11] ;
assign n186 = /* LUT    1 18  6 */ \a_i[11] ;
assign n187 = /* LUT    2 17  0 */ (n118 ? (n119 ? n93 : !n93) : (n119 ? !n93 : n93));
assign n188 = /* LUT    2 15  3 */ n80;
assign n189 = /* LUT    1 17  3 */ (n48 ? n98 : !n98);
assign n133 = /* LUT    2 18  1 */ n132;
assign n190 = /* LUT    2 17  1 */ (n121 ? (n43 ? n47 : !n47) : (n43 ? !n47 : n47));
assign n191 = /* LUT    1 18  7 */ (n56 ? 1'b1 : (n58 ? 1'b1 : n105));
assign n192 = /* LUT    3 17  0 */ io_4_33_0;
assign n193 = /* LUT    2 18  0 */ (n128 ? (n30 ? n19 : !n19) : (n30 ? !n19 : n19));
assign n194 = /* LUT    1 17  2 */ \sum_o[4] ;
assign n108 = /* LUT    2 15  5 */ (n80 ? (n22 ? n103 : !n103) : (n22 ? !n103 : n103));
assign n195 = /* LUT    1 17  5 */ (n90 ? (n43 ? (n81 ? n47 : !n47) : (n81 ? !n47 : n47)) : (n43 ? (n81 ? !n47 : n47) : (n81 ? n47 : !n47)));
assign n196 = /* LUT    1 19  4 */ (n55 ? !n54 : n54);
assign n197 = /* LUT    2 18  7 */ !n105;
assign n198 = /* LUT    1 15  2 */ io_0_4_1;
assign n199 = /* LUT    1 16  2 */ \a_i[5] ;
assign n200 = /* LUT    2 19  4 */ clk_i;
assign n201 = /* LUT    2 15  6 */ (n78 ? (n108 ? 1'b1 : !n77) : (n108 ? 1'b0 : n77));
assign n202 = /* LUT    1 17  4 */ (n46 ? 1'b1 : (n48 ? 1'b1 : n98));
assign n203 = /* LUT    1 19  3 */ \a_i[4] ;
assign n204 = /* LUT    2 18  6 */ io_3_33_0;
assign n205 = /* LUT    1 15  1 */ io_0_3_0;
assign n206 = /* LUT    1 16  3 */ (n24 ? 1'b1 : (n28 ? 1'b1 : n26));
assign n207 = /* LUT    2 19  5 */ \b_i[0] ;
assign n208 = /* LUT    2 15  7 */ \sum_o[10] ;
assign n209 = /* LUT    1 17  7 */ !n98;
assign n210 = /* LUT    1 19  2 */ \b_i[8] ;
assign n211 = /* LUT    2 18  5 */ (n58 ? n105 : !n105);
assign n212 = /* LUT    1 15  0 */ \b_i[2] ;
assign n213 = /* LUT    1 16  0 */ n86;
assign n214 = /* LUT    3 18  5 */ \sum_o[5] ;
assign n215 = /* LUT    1 17  6 */ \a_i[6] ;
assign n216 = /* LUT    1 19  1 */ \a_i[7] ;
assign n217 = /* LUT    1 15  7 */ \a_i[15] ;
assign n218 = /* LUT    1 16  1 */ (n84 ? (n55 ? (n54 ? n86 : !n86) : (n54 ? !n86 : n86)) : (n55 ? (n54 ? !n86 : n86) : (n54 ? n86 : !n86)));
assign n116 = /* CARRY  2 16  5 */ (n103 & n22) | ((n103 | n22) & n115);
assign n115 = /* CARRY  2 16  4 */ (n96 & n38) | ((n96 | n38) & n114);
assign n118 = /* CARRY  2 16  7 */ (n40 & n110) | ((n40 | n110) & n117);
assign n117 = /* CARRY  2 16  6 */ (n29 & n109) | ((n29 | n109) & n116);
assign n112 = /* CARRY  2 16  1 */ (n25 & n76) | ((n25 | n76) & n111);
assign n127 = /* CARRY  2 17  6 */ (n31 & n94) | ((n31 | n94) & n126);
assign n111 = /* CARRY  2 16  0 */ (n74 & n74) | ((n74 | n74) & n160);
assign n128 = /* CARRY  2 17  7 */ (n23 & n32) | ((n23 | n32) & n127);
assign n114 = /* CARRY  2 16  3 */ (n95 & n37) | ((n95 | n37) & n113);
assign n125 = /* CARRY  2 17  4 */ (n53 & n49) | ((n53 | n49) & n124);
assign n113 = /* CARRY  2 16  2 */ (n36 & n41) | ((n36 | n41) & n112);
assign n126 = /* CARRY  2 17  5 */ (n54 & n55) | ((n54 | n55) & n125);
assign n123 = /* CARRY  2 17  2 */ (n27 & n102) | ((n27 | n102) & n122);
assign n124 = /* CARRY  2 17  3 */ (n104 & n101) | ((n104 | n101) & n123);
assign n121 = /* CARRY  2 17  0 */ (n93 & n119) | ((n93 | n119) & n118);
assign n122 = /* CARRY  2 17  1 */ (n47 & n43) | ((n47 | n43) & n121);
assign n132 = /* CARRY  2 18  0 */ (n19 & n30) | ((n19 | n30) & n128);
/* FF  3 16  0 */ assign n109 = n137;
/* FF  1 19  0 */ always @(posedge \sum_o[14] ) if (1'b1) n53 <= 1'b0 ? 1'b0 : n138;
/* FF  1 15  6 */ always @(posedge \sum_o[14] ) if (1'b1) n27 <= 1'b0 ? 1'b0 : n139;
/* FF  1 16  6 */ assign n31 = n140;
/* FF  2 19  0 */ always @(posedge \sum_o[14] ) if (1'b1) n104 <= 1'b0 ? 1'b0 : n141;
/* FF  2 16  5 */ assign n80 = n142;
/* FF  1 15  5 */ always @(posedge \sum_o[14] ) if (1'b1) n26 <= 1'b0 ? 1'b0 : n143;
/* FF  1 16  7 */ assign n32 = n144;
/* FF  2 16  4 */ assign n79 = n145;
/* FF  1 15  4 */ always @(posedge \sum_o[14] ) if (1'b1) n25 <= 1'b0 ? 1'b0 : n146;
/* FF  1 16  4 */ assign n147 = n88;
/* FF  2 19  2 */ always @(posedge \sum_o[14] ) if (1'b1) n105 <= 1'b0 ? 1'b0 : n148;
/* FF  1 14  7 */ always @(posedge \sum_o[14] ) if (1'b1) n19 <= 1'b0 ? 1'b0 : n149;
/* FF  2 16  7 */ assign n82 = n150;
/* FF  1 16  5 */ always @(posedge \sum_o[14] ) if (1'b1) io_0_6_0 <= 1'b0 ? 1'b0 : n151;
/* FF  2 19  7 */ always @(posedge \sum_o[14] ) if (1'b1) n103 <= 1'b0 ? 1'b0 : n152;
/* FF  2 16  6 */ assign n81 = n153;
/* FF  2 16  1 */ always @(posedge \sum_o[14] ) if (1'b1) \a_i[9]  <= 1'b0 ? 1'b0 : n154;
/* FF  2 17  6 */ assign n91 = n155;
/* FF  1 18  0 */ always @(posedge \sum_o[14] ) if (1'b1) n43 <= 1'b0 ? 1'b0 : n156;
/* FF  2 18  4 */ always @(posedge \sum_o[14] ) if (1'b1) \sum_o[6]  <= 1'b0 ? 1'b0 : n157;
/* FF  2 16  0 */ assign n158 = n159;
/* FF  3 17  7 */ always @(posedge \sum_o[14] ) if (1'b1) n96 <= 1'b0 ? 1'b0 : n161;
/* FF  2 17  7 */ assign n92 = n162;
/* FF  1 18  1 */ always @(posedge \sum_o[14] ) if (1'b1) \sum_o[7]  <= 1'b0 ? 1'b0 : n163;
/* FF  3 17  6 */ always @(posedge \sum_o[14] ) if (1'b1) n120 <= 1'b0 ? 1'b0 : n164;
/* FF  2 16  3 */ assign n78 = n165;
/* FF  1 18  2 */ always @(posedge \sum_o[14] ) if (1'b1) \sum_o[8]  <= 1'b0 ? 1'b0 : n166;
/* FF  2 17  4 */ assign n85 = n167;
/* FF  3 17  5 */ always @(posedge \sum_o[14] ) if (1'b1) \a_i[1]  <= 1'b0 ? 1'b0 : n168;
/* FF  2 16  2 */ assign n77 = n169;
/* FF  3 17  4 */ assign n110 = n170;
/* FF  1 18  3 */ always @(posedge \sum_o[14] ) if (1'b1) n46 <= 1'b0 ? 1'b0 : n171;
/* FF  2 17  5 */ assign n86 = n172;
/* FF  2 15  0 */ always @(posedge \sum_o[14] ) if (1'b1) n74 <= 1'b0 ? 1'b0 : n173;
/* FF  1 18  4 */ always @(posedge \sum_o[14] ) if (1'b1) \b_i[14]  <= 1'b0 ? 1'b0 : n174;
/* FF  2 17  2 */ assign n84 = n175;
/* FF  3 17  3 */ assign n119 = n176;
/* FF  2 15  1 */ always @(posedge \sum_o[14] ) if (1'b1) \sum_o[9]  <= 1'b0 ? 1'b0 : n177;
/* FF  1 17  1 */ always @(posedge \sum_o[14] ) if (1'b1) \b_i[15]  <= 1'b0 ? 1'b0 : n178;
/* FF  2 18  3 */ assign n100 = n134;
/* FF  3 18  3 */ always @(posedge \sum_o[14] ) if (1'b1) n129 <= 1'b0 ? 1'b0 : n179;
/* FF  1 18  5 */ always @(posedge \sum_o[14] ) if (1'b1) n47 <= 1'b0 ? 1'b0 : n180;
/* FF  2 17  3 */ assign n87 = n181;
/* FF  2 15  2 */ always @(posedge \sum_o[14] ) if (1'b1) \sum_o[12]  <= 1'b0 ? 1'b0 : n182;
/* FF  2 18  2 */ always @(posedge \sum_o[14] ) if (1'b1) io_0_7_1 <= 1'b0 ? 1'b0 : n183;
/* FF  1 17  0 */ always @(posedge \sum_o[14] ) if (1'b1) \sum_o[13]  <= 1'b0 ? 1'b0 : n184;
/* FF  1 19  7 */ always @(posedge \sum_o[14] ) if (1'b1) n58 <= 1'b0 ? 1'b0 : n185;
/* FF  1 18  6 */ always @(posedge \sum_o[14] ) if (1'b1) n48 <= 1'b0 ? 1'b0 : n186;
/* FF  2 17  0 */ assign n89 = n187;
/* FF  2 15  3 */ always @(posedge \sum_o[14] ) if (1'b1) \a_i[14]  <= 1'b0 ? 1'b0 : n188;
/* FF  1 17  3 */ assign n37 = n189;
/* FF  2 18  1 */ assign n97 = n133;
/* FF  2 17  1 */ assign n90 = n190;
/* FF  1 18  7 */ assign n49 = n191;
/* FF  3 17  0 */ always @(posedge \sum_o[14] ) if (1'b1) n95 <= 1'b0 ? 1'b0 : n192;
/* FF  2 18  0 */ assign n99 = n193;
/* FF  1 17  2 */ always @(posedge \sum_o[14] ) if (1'b1) n36 <= 1'b0 ? 1'b0 : n194;
/* FF  2 15  5 */ assign n75 = n108;
/* FF  1 17  5 */ always @(posedge \sum_o[14] ) if (1'b1) \a_i[0]  <= 1'b0 ? 1'b0 : n195;
/* FF  1 19  4 */ assign n57 = n196;
/* FF  2 18  7 */ assign n102 = n197;
/* FF  1 15  2 */ always @(posedge \sum_o[14] ) if (1'b1) n24 <= 1'b0 ? 1'b0 : n198;
/* FF  1 16  2 */ always @(posedge \sum_o[14] ) if (1'b1) n29 <= 1'b0 ? 1'b0 : n199;
/* FF  2 19  4 */ always @(posedge \sum_o[14] ) if (1'b1) n93 <= 1'b0 ? 1'b0 : n200;
/* FF  2 15  6 */ always @(posedge \sum_o[14] ) if (1'b1) \b_i[13]  <= 1'b0 ? 1'b0 : n201;
/* FF  1 17  4 */ assign n38 = n202;
/* FF  1 19  3 */ always @(posedge \sum_o[14] ) if (1'b1) n56 <= 1'b0 ? 1'b0 : n203;
/* FF  2 18  6 */ always @(posedge \sum_o[14] ) if (1'b1) n98 <= 1'b0 ? 1'b0 : n204;
/* FF  1 15  1 */ always @(posedge \sum_o[14] ) if (1'b1) n23 <= 1'b0 ? 1'b0 : n205;
/* FF  1 16  3 */ assign n30 = n206;
/* FF  2 19  5 */ always @(posedge \sum_o[14] ) if (1'b1) n94 <= 1'b0 ? 1'b0 : n207;
/* FF  2 15  7 */ always @(posedge \sum_o[14] ) if (1'b1) n76 <= 1'b0 ? 1'b0 : n208;
/* FF  1 17  7 */ assign n41 = n209;
/* FF  1 19  2 */ always @(posedge \sum_o[14] ) if (1'b1) n55 <= 1'b0 ? 1'b0 : n210;
/* FF  2 18  5 */ assign n101 = n211;
/* FF  1 15  0 */ always @(posedge \sum_o[14] ) if (1'b1) n22 <= 1'b0 ? 1'b0 : n212;
/* FF  1 16  0 */ always @(posedge \sum_o[14] ) if (1'b1) io_0_6_1 <= 1'b0 ? 1'b0 : n213;
/* FF  3 18  5 */ always @(posedge \sum_o[14] ) if (1'b1) n130 <= 1'b0 ? 1'b0 : n214;
/* FF  1 17  6 */ always @(posedge \sum_o[14] ) if (1'b1) n40 <= 1'b0 ? 1'b0 : n215;
/* FF  1 19  1 */ always @(posedge \sum_o[14] ) if (1'b1) n54 <= 1'b0 ? 1'b0 : n216;
/* FF  1 15  7 */ always @(posedge \sum_o[14] ) if (1'b1) n28 <= 1'b0 ? 1'b0 : n217;
/* FF  1 16  1 */ always @(posedge \sum_o[14] ) if (1'b1) \sum_o[11]  <= 1'b0 ? 1'b0 : n218;

// Warning: unmatched port '\sum_o[1] '
// Warning: unmatched port '\b_i[5] '
// Warning: unmatched port '\sum_o[15] '
// Warning: unmatched port '\b_i[12] '
// Warning: unmatched port '\a_i[13] '
// Warning: unmatched port '\b_i[3] '
// Warning: unmatched port 'cin_i'
// Warning: unmatched port '\a_i[2] '
// Warning: unmatched port 'cout_o'
// Warning: unmatched port '\a_i[3] '

endmodule

