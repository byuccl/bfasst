
module chip (input clk, output \cypher[31] , output \cypher[5] , output \cypher[6] , output \cypher[26] , output \cypher[27] , output \cypher[24] , output \cypher[25] , output \cypher[20] , output \cypher[21] , output \cypher[12] , output \cypher[13] , output \cypher[3] , output \cypher[4] , output \cypher[16] , output \cypher[17] , output \cypher[22] , output \cypher[23] , output \cypher[18] , output ready, output \cypher[19] , output \cypher[14] , output \cypher[15] , output \cypher[7] , output \cypher[8] , output \cypher[2] , output \cypher[28] , input reset, output \cypher[9] , input \inMod[5] , input ds, output \cypher[0] , output \cypher[30] , output \cypher[29] , output \cypher[11] , input \inMod[6] , input \inExp[0] , output \cypher[10] , output \cypher[1] , input \inMod[8] , input \inMod[7] , input \inMod[4] , input \inMod[31] , input \indata[15] , input \inMod[30] , input \inMod[3] , input \indata[18] , input \inMod[14] , input \inMod[13] , input \indata[21] , input \inMod[12] , input \inMod[11] , input \inMod[10] , input \inMod[1] , input \inMod[0] , input \indata[22] , input \inMod[21] , input \inMod[20] , input \inMod[2] , input \indata[24] , input \inMod[18] , input \inMod[19] , input \indata[5] , input \inMod[17] , input \inMod[16] , input \indata[1] , input \indata[29] , input \inMod[15] , input \inMod[22] , input \indata[31] , input \inMod[28] , input \inMod[29] , input \inMod[23] , input \indata[2] , input \indata[10] , input \indata[0] , input \indata[30] , input \indata[28] , input \indata[11] , input \indata[14] , input \inMod[25] , input \inMod[24] , input \indata[4] , input \inMod[26] , input \inMod[27] , input \indata[6] , input \indata[27] , input \indata[9] , input \indata[8] , input \indata[12] , input \indata[3] , input \indata[23] , input \indata[13] , input \indata[19] , input \inMod[9] , input \inExp[11] , input \indata[26] , input \indata[7] , input \indata[25] , input \inExp[12] , input \inExp[13] , input \inExp[14] , input \indata[20] , input \indata[16] , input \indata[17] , input \inExp[15] , input \inExp[29] , input \inExp[5] , input \inExp[30] , input \inExp[31] , input \inExp[7] , input \inExp[20] , input \inExp[19] , input \inExp[16] , input \inExp[1] , input \inExp[21] , input \inExp[28] , input \inExp[26] , input \inExp[10] , input \inExp[8] , input \inExp[23] , input \inExp[22] , input \inExp[9] , input \inExp[18] , input \inExp[6] , input \inExp[25] , input \inExp[24] , input \inExp[17] , input \inExp[3] , input \inExp[2] , input \inExp[27] , input \inExp[4] );

wire clk, n2, n3, \cypher[31] , \cypher[5] , n6, n7, n8, \cypher[6] , \cypher[26] ;
wire n11, \cypher[27] , n13, \cypher[24] , n15, \cypher[25] , n17, \cypher[20] , n19, \cypher[21] ;
wire n21, \cypher[12] , n23, \cypher[13] , n25, \cypher[3] , n27, \cypher[4] , n29, \cypher[16] ;
wire n31, \cypher[17] , n33, \cypher[22] , n35, n36, \cypher[23] , n38, \cypher[18] , n40;
wire \cypher[19] , \cypher[14] , n44, \cypher[15] , n46, \cypher[7] , n48, n51, n53, n54;
wire \cypher[8] , \cypher[2] , n57, n58, n59, n60, n61, n62, n63, n64;
wire n67, \cypher[28] , n69, n70, n71, n72, n73, n74, n75, n76;
wire n79, n80, n81, n82, n83, reset, n85, \cypher[9] , n87, n88;
wire n89, n90, n91, n92, n93, n94, n97, n100, n102, n103;
wire n104, \inMod[5] , n106, n107, ds, n109, \cypher[0] , n111, \cypher[30] , n113;
wire n114, n115, n116, n117, n118, n119, n120, n121, n122, n123;
wire n124, n125, n128, n129, \cypher[29] , \cypher[11] , n132, n133, n135, n136;
wire n137, n138, n141, \inMod[6] , n144, n145, n146, \inExp[0] , n148, n149;
wire n150, n151, n152, n153, n154, n155, n156, n157, n159, n160;
wire n161, n162, \cypher[10] , n164, \cypher[1] , n166, n167, n168, n169, n170;
wire n171, n172, n173, n177, n178, n181, n182, n185, n186, n187;
wire n189, \inMod[8] , \inMod[7] , n193, n194, n195, n196, n197, n198, n199;
wire n201, n203, n204, n206, n207, n208, n210, n211, n212, n213;
wire n214, n215, n216, n217, n218, n219, n224, n226, \inMod[4] , \inMod[31] ;
wire n230, n231, n232, n233, n234, n235, \indata[15] , n242, n245, n246;
wire n247, n248, n253, \inMod[30] , \inMod[3] , \indata[18] , \inMod[14] , \inMod[13] , \indata[21] , \inMod[12] ;
wire \inMod[11] , \inMod[10] , \inMod[1] , \inMod[0] , n272, \indata[22] , n274, n276, n277, n278;
wire n279, n280, n281, n282, n283, n284, n285, n286, n287, n288;
wire n290, n291, n292, n293, n294, n295, n296, n297, n298, n299;
wire n300, n301, n302, n303, n307, n308, n309, n310, n311, n312;
wire n313, n314, n315, n316, n317, n318, n319, n321, n322, n324;
wire n326, n327, n328, n329, n330, n331, n332, n333, n334, n335;
wire n336, n337, n338, n339, n340, n342, n343, n344, n345, n346;
wire n347, n348, n349, n350, n351, n352, n353, n354, n355, n356;
wire n357, n358, n361, n362, n363, n364, n365, n366, n367, n368;
wire n369, n370, n371, n372, n373, n374, n375, n376, n377, n379;
wire n380, n382, n383, n384, n385, n386, n387, n388, n389, n390;
wire n391, n392, n393, n394, n395, n401, n402, n403, n404, n405;
wire n406, n407, n408, n409, n410, n411, n412, n418, n419, n420;
wire n421, n422, n423, n424, n425, n426, n427, n428, n429, n430;
wire n433, n434, n436, n437, \inMod[21] , \inMod[20] , \inMod[2] , n443, n450, n451;
wire n452, n453, n457, n458, n459, n460, n461, n462, n464, n466;
wire n469, n472, n473, n474, n475, n476, n477, n478, n479, n483;
wire n484, n485, n486, n487, n488, n489, n490, n491, n495, n496;
wire n497, n498, n499, n500, n501, n502, n504, n505, n506, n507;
wire n508, n509, n510, n511, n512, n513, n514, n515, n516, n519;
wire n525, \indata[24] , n529, \inMod[18] , \inMod[19] , n545, n561, n562, n563, n564;
wire \indata[5] , n570, n571, n572, n573, n574, n575, n576, n577, n579;
wire n580, n581, n582, n583, n585, n593, n599, n601, n602, n604;
wire n607, n608, n609, n610, n613, n614, n615, n616, n617, n619;
wire n620, n622, \inMod[17] , \inMod[16] , n627, n628, n643, n644, n646, n648;
wire n650, n651, n652, n653, n657, n658, \indata[1] , n669, \indata[29] , n679;
wire n680, n681, n682, n683, n684, n685, n688, n689, n690, n691;
wire n692, n693, n694, n695, n697, n698, n699, n700, n701, n702;
wire n703, n704, n705, n706, n708, n709, n710, n711, n712, n713;
wire n714, n715, n716, n717, n720, n721, n722, n723, \inMod[15] , \inMod[22] ;
wire \indata[31] , n727, n731, n734, n735, n737, n745, n746, n747, n748;
wire n750, n752, n753, n754, n755, n756, n757, n759, n760, n761;
wire n763, n767, n769, n770, n771, n776, n777, n779, n780, n781;
wire n785, n786, n792, n793, n794, n795, n796, n797, n798, n799;
wire n800, n801, n802, n803, n804, n805, n806, n807, n808, n809;
wire n810, n811, n812, n813, n814, n815, n816, n817, n818, n819;
wire n820, n821, n822, n823, n824, n825, n826, n827, n828, n829;
wire \inMod[28] , \inMod[29] , \inMod[23] , \indata[2] , n834, n835, \indata[10] , n838, n839, \indata[0] ;
wire n845, n849, n850, \indata[30] , n852, n853, n854, n855, n858, n859;
wire n860, n861, n862, n863, n869, n870, n871, n872, n873, n874;
wire n875, n876, n878, \indata[28] , n880, n886, n887, \indata[11] , n889, n890;
wire n892, n893, n894, \indata[14] , n896, n900, n901, n905, n906, \inMod[25] ;
wire \inMod[24] , n910, n911, n912, n913, n915, n918, n919, n920, n921;
wire n922, n923, n924, n925, n926, n927, n928, n929, n930, n931;
wire n932, n933, n934, n935, n936, n937, n938, n939, \indata[4] , n941;
wire \inMod[26] , \inMod[27] , n947, n948, n949, \indata[6] , \indata[27] , n954, n955, n956;
wire n958, n959, \indata[9] , n962, \indata[8] , n970, n971, n972, \indata[12] , n978;
wire n979, n981, n982, n983, n984, n985, \indata[3] , n989, n990, \indata[23] ;
wire n994, n995, n996, n999, n1000, n1002, n1003, n1004, n1005, n1008;
wire n1010, n1012, n1013, n1014, n1015, n1016, n1017, n1019, n1021, n1022;
wire n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032;
wire \indata[13] , n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042;
wire n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052;
wire n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1061, n1062, n1063;
wire n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073;
wire n1074, n1075, n1076, n1077, n1078, \indata[19] , n1081, n1082, n1083, n1084;
wire n1085, \inMod[9] , \inExp[11] , \indata[26] , n1090, n1091, n1092, n1093, n1094, n1095;
wire n1096, n1097, n1098, n1099, n1100, n1101, n1106, n1107, n1109, n1111;
wire n1112, n1113, n1116, n1117, n1121, n1123, \indata[7] , n1125, n1126, n1127;
wire \indata[25] , n1129, n1130, n1131, n1132, n1133, n1134, n1137, n1138, n1139;
wire n1140, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150;
wire n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160;
wire n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170;
wire n1171, n1172, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181;
wire n1182, n1183, n1184, n1185, \inExp[12] , \inExp[13] , \inExp[14] , n1190, n1191, n1194;
wire n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1206, n1207;
wire n1208, n1209, n1210, n1213, n1215, n1216, n1217, n1218, n1219, n1220;
wire n1221, n1222, n1223, n1224, n1225, n1228, n1229, n1230, n1231, n1232;
wire n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242;
wire n1243, n1244, n1245, n1246, n1247, n1249, n1251, n1253, n1255, n1256;
wire n1257, n1258, n1259, n1260, n1261, n1262, n1267, n1268, n1269, n1270;
wire n1271, n1272, n1273, n1274, \indata[20] , n1278, n1280, n1281, n1282, n1286;
wire n1289, n1290, n1291, n1292, n1294, n1296, n1297, n1298, n1299, n1300;
wire n1301, n1302, n1303, n1311, n1312, n1313, n1314, n1315, n1316, n1317;
wire n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1328;
wire n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338;
wire \indata[16] , \indata[17] , n1342, n1343, n1344, \inExp[15] , n1346, n1347, n1348, n1349;
wire n1350, n1351, n1352, n1354, n1355, n1356, \inExp[29] , n1358, n1359, n1360;
wire n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375;
wire n1376, n1377, n1378, n1380, n1381, n1382, n1383, n1384, n1385, n1386;
wire n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396;
wire n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406;
wire n1407, n1408, n1409, n1410, n1411, \inExp[5] , n1415, n1426, n1427, n1429;
wire n1430, n1431, n1437, n1438, n1439, n1441, n1444, n1445, \inExp[30] , \inExp[31] ;
wire \inExp[7] , \inExp[20] , n1459, \inExp[19] , n1472, n1473, n1474, \inExp[16] , \inExp[1] , \inExp[21] ;
wire \inExp[28] , \inExp[26] , \inExp[10] , \inExp[8] , \inExp[23] , \inExp[22] , n1484, \inExp[9] , \inExp[18] , \inExp[6] ;
wire \inExp[25] , \inExp[24] , n1495, n1496, n1498, \inExp[17] , \inExp[3] , \inExp[2] , \inExp[27] , n1507;
wire n1508, \inExp[4] , n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549;
wire n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559;
wire n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569;
wire n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579;
wire n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589;
wire n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599;
wire n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609;
wire n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619;
wire n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629;
wire n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639;
wire n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649;
wire n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659;
wire n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669;
wire n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679;
wire n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689;
wire n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699;
wire n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709;
wire n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719;
wire n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729;
wire n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739;
wire n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749;
wire n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759;
wire n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769;
wire n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779;
wire n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789;
wire n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799;
wire n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809;
wire n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819;
wire n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829;
wire n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839;
wire n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849;
wire n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859;
wire n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869;
wire n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879;
wire n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889;
wire n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899;
wire n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909;
wire n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919;
wire n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929;
wire n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939;
wire n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949;
wire n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959;
wire n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969;
wire n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979;
wire n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989;
wire n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999;
wire n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009;
wire n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019;
wire n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029;
wire n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039;
wire n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049;
wire n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059;
wire n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069;
wire n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079;
wire n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089;
wire n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099;
wire n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109;
wire n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119;
wire n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129;
wire n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139;
wire n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149;
wire n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159;
wire n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169;
wire n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179;
wire n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189;
wire n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199;
wire n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209;
wire n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219;
wire n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229;
wire n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239;
wire n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249;
wire n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259;
wire n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269;
wire n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279;
wire n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289;
wire n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299;
wire n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309;
wire n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319;
wire n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329;
wire n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339;
wire n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349;
wire n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359;
wire n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369;
wire n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379;
wire n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389;
wire n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399;
wire n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409;
wire n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419;
wire n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429;
wire n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439;
wire n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449;
wire n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459;
wire n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469;
wire n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479;
wire n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489;
wire n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499;
wire n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509;
wire n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519;
wire n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529;
wire n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539;
wire n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549;
wire n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559;
wire n2560, n2561, n2562, n2563;
reg ready = 0, n49 = 0, n50 = 0, n52 = 0, n65 = 0, n66 = 0, n77 = 0, n78 = 0, n95 = 0, n96 = 0;
reg n98 = 0, n99 = 0, n101 = 0, n126 = 0, n127 = 0, n134 = 0, n139 = 0, n140 = 0, n142 = 0, n158 = 0;
reg n174 = 0, n175 = 0, n176 = 0, n179 = 0, n180 = 0, n183 = 0, n184 = 0, n188 = 0, n190 = 0, n200 = 0;
reg n202 = 0, n205 = 0, n209 = 0, n220 = 0, n221 = 0, n222 = 0, n223 = 0, n225 = 0, n227 = 0, n236 = 0;
reg n237 = 0, n238 = 0, n239 = 0, n240 = 0, n243 = 0, n244 = 0, n249 = 0, n250 = 0, n251 = 0, n252 = 0;
reg n254 = 0, n255 = 0, n256 = 0, n257 = 0, n261 = 0, n262 = 0, n265 = 0, n275 = 0, n289 = 0, n304 = 0;
reg n305 = 0, n306 = 0, n320 = 0, n323 = 0, n325 = 0, n341 = 0, n359 = 0, n360 = 0, n378 = 0, n381 = 0;
reg n396 = 0, n397 = 0, n398 = 0, n399 = 0, n400 = 0, n413 = 0, n414 = 0, n415 = 0, n416 = 0, n417 = 0;
reg n431 = 0, n432 = 0, n435 = 0, n438 = 0, n439 = 0, n444 = 0, n445 = 0, n446 = 0, n447 = 0, n448 = 0;
reg n449 = 0, n454 = 0, n455 = 0, n456 = 0, n463 = 0, n465 = 0, n467 = 0, n468 = 0, n470 = 0, n471 = 0;
reg n480 = 0, n481 = 0, n482 = 0, n492 = 0, n493 = 0, n494 = 0, n503 = 0, n517 = 0, n518 = 0, n520 = 0;
reg n521 = 0, n522 = 0, n523 = 0, n524 = 0, n526 = 0, n527 = 0, n530 = 0, n531 = 0, n532 = 0, n533 = 0;
reg n534 = 0, n535 = 0, n536 = 0, n537 = 0, n538 = 0, n541 = 0, n542 = 0, n543 = 0, n544 = 0, n546 = 0;
reg n547 = 0, n548 = 0, n549 = 0, n550 = 0, n551 = 0, n552 = 0, n553 = 0, n554 = 0, n555 = 0, n556 = 0;
reg n557 = 0, n558 = 0, n559 = 0, n560 = 0, n565 = 0, n566 = 0, n568 = 0, n569 = 0, n578 = 0, n584 = 0;
reg n586 = 0, n587 = 0, n588 = 0, n589 = 0, n590 = 0, n591 = 0, n592 = 0, n594 = 0, n595 = 0, n596 = 0;
reg n597 = 0, n598 = 0, n600 = 0, n603 = 0, n605 = 0, n606 = 0, n611 = 0, n612 = 0, n618 = 0, n621 = 0;
reg n623 = 0, n624 = 0, n629 = 0, n630 = 0, n631 = 0, n632 = 0, n633 = 0, n634 = 0, n635 = 0, n636 = 0;
reg n637 = 0, n638 = 0, n639 = 0, n640 = 0, n641 = 0, n642 = 0, n645 = 0, n647 = 0, n649 = 0, n654 = 0;
reg n655 = 0, n656 = 0, n659 = 0, n660 = 0, n661 = 0, n662 = 0, n663 = 0, n665 = 0, n666 = 0, n667 = 0;
reg n668 = 0, n670 = 0, n671 = 0, n672 = 0, n673 = 0, n674 = 0, n675 = 0, n676 = 0, n678 = 0, n686 = 0;
reg n687 = 0, n696 = 0, n707 = 0, n718 = 0, n719 = 0, n728 = 0, n729 = 0, n730 = 0, n732 = 0, n733 = 0;
reg n736 = 0, n738 = 0, n739 = 0, n740 = 0, n741 = 0, n742 = 0, n743 = 0, n744 = 0, n749 = 0, n751 = 0;
reg n758 = 0, n762 = 0, n764 = 0, n765 = 0, n766 = 0, n768 = 0, n772 = 0, n773 = 0, n774 = 0, n775 = 0;
reg n778 = 0, n782 = 0, n783 = 0, n784 = 0, n787 = 0, n788 = 0, n789 = 0, n790 = 0, n791 = 0, n837 = 0;
reg n841 = 0, n842 = 0, n843 = 0, n844 = 0, n846 = 0, n847 = 0, n848 = 0, n856 = 0, n857 = 0, n864 = 0;
reg n865 = 0, n866 = 0, n867 = 0, n868 = 0, n877 = 0, n881 = 0, n882 = 0, n883 = 0, n884 = 0, n885 = 0;
reg n891 = 0, n897 = 0, n898 = 0, n899 = 0, n902 = 0, n903 = 0, n904 = 0, n907 = 0, n914 = 0, n916 = 0;
reg n917 = 0, n942 = 0, n945 = 0, n946 = 0, n952 = 0, n953 = 0, n957 = 0, n960 = 0, n963 = 0, n965 = 0;
reg n966 = 0, n967 = 0, n968 = 0, n969 = 0, n973 = 0, n974 = 0, n975 = 0, n976 = 0, n980 = 0, n987 = 0;
reg n988 = 0, n992 = 0, n993 = 0, n997 = 0, n998 = 0, n1001 = 0, n1006 = 0, n1007 = 0, n1009 = 0, n1011 = 0;
reg n1018 = 0, n1020 = 0, n1060 = 0, n1079 = 0, n1086 = 0, n1102 = 0, n1103 = 0, n1104 = 0, n1105 = 0, n1108 = 0;
reg n1110 = 0, n1114 = 0, n1115 = 0, n1118 = 0, n1119 = 0, n1120 = 0, n1122 = 0, n1135 = 0, n1136 = 0, n1141 = 0;
reg n1173 = 0, n1189 = 0, n1192 = 0, n1193 = 0, n1195 = 0, n1196 = 0, n1205 = 0, n1211 = 0, n1212 = 0, n1214 = 0;
reg n1226 = 0, n1227 = 0, n1248 = 0, n1250 = 0, n1252 = 0, n1254 = 0, n1263 = 0, n1264 = 0, n1265 = 0, n1266 = 0;
reg n1275 = 0, n1276 = 0, n1279 = 0, n1283 = 0, n1284 = 0, n1285 = 0, n1287 = 0, n1288 = 0, n1293 = 0, n1295 = 0;
reg n1304 = 0, n1305 = 0, n1306 = 0, n1307 = 0, n1308 = 0, n1309 = 0, n1310 = 0, n1327 = 0, n1340 = 0, n1353 = 0;
reg n1361 = 0, n1362 = 0, n1363 = 0, n1364 = 0, n1365 = 0, n1379 = 0, n1412 = 0, n1413 = 0, n1416 = 0, n1417 = 0;
reg n1418 = 0, n1419 = 0, n1420 = 0, n1421 = 0, n1422 = 0, n1423 = 0, n1424 = 0, n1425 = 0, n1428 = 0, n1432 = 0;
reg n1433 = 0, n1434 = 0, n1435 = 0, n1436 = 0, n1440 = 0, n1442 = 0, n1443 = 0, n1446 = 0, n1450 = 0, n1451 = 0;
reg n1452 = 0, n1453 = 0, n1454 = 0, n1455 = 0, n1456 = 0, n1457 = 0, n1461 = 0, n1462 = 0, n1463 = 0, n1464 = 0;
reg n1465 = 0, n1466 = 0, n1467 = 0, n1468 = 0, n1469 = 0, n1470 = 0, n1471 = 0, n1485 = 0, n1486 = 0, n1487 = 0;
reg n1488 = 0, n1489 = 0, n1497 = 0, n1499 = 0, n1500 = 0, n1501 = 0, n1502 = 0;
assign n1608 = 1;
assign n792 = 1;
assign n276 = 1;
assign n2011 = 1;
assign n2188 = 0;
assign n2216 = 0;
assign n2414 = 1;
assign n1143 = 1;

// IO Cell (0, 5, 1)
reg n1510;
always @(posedge clk) if (n6) n1510 <= n13;
assign \cypher[24]  = n1510;

// IO Cell (0, 22, 0)
reg n1511;
always @(posedge clk) if (n6) n1511 <= n162;
assign \cypher[10]  = n1511;

// IO Cell (0, 12, 1)
reg n1512;
always @(posedge clk) if (n6) n1512 <= n35;
assign \cypher[14]  = n1512;

// IO Cell (0, 19, 0)
reg n1513;
always @(posedge clk) if (n6) n1513 <= n109;
assign \cypher[0]  = n1513;

// IO Cell (0, 16, 0)
reg n1514;
always @(posedge clk) if (n6) n1514 <= n54;
assign \cypher[8]  = n1514;

// IO Cell (0, 9, 1)
reg n1515;
always @(posedge clk) if (n6) n1515 <= n29;
assign \cypher[16]  = n1515;

// IO Cell (0, 7, 0)
reg n1516;
always @(posedge clk) if (n6) n1516 <= n19;
assign \cypher[21]  = n1516;

// IO Cell (0, 4, 0)
reg n1517;
always @(posedge clk) if (n6) n1517 <= n8;
assign \cypher[6]  = n1517;

// IO Cell (0, 11, 0)
reg n1518;
always @(posedge clk) if (n6) n1518 <= n36;
assign \cypher[23]  = n1518;

// IO Cell (0, 8, 0)
reg n1519;
always @(posedge clk) if (n6) n1519 <= n23;
assign \cypher[13]  = n1519;

// IO Cell (0, 6, 1)
reg n1520;
always @(posedge clk) if (n6) n1520 <= n17;
assign \cypher[20]  = n1520;

// IO Cell (0, 3, 1)
reg n1521;
always @(posedge clk) if (n6) n1521 <= n2;
assign \cypher[5]  = n1521;

// IO Cell (0, 20, 0)
reg n1522;
always @(posedge clk) if (n6) n1522 <= n123;
assign \cypher[29]  = n1522;

// IO Cell (0, 10, 1)
reg n1523;
always @(posedge clk) if (n6) n1523 <= n33;
assign \cypher[22]  = n1523;

// IO Cell (0, 5, 0)
reg n1524;
always @(posedge clk) if (n6) n1524 <= n11;
assign \cypher[27]  = n1524;

// IO Cell (0, 22, 1)
reg n1525;
always @(posedge clk) if (n6) n1525 <= n164;
assign \cypher[1]  = n1525;

// IO Cell (0, 12, 0)
reg n1526;
always @(posedge clk) if (n6) n1526 <= n40;
assign \cypher[19]  = n1526;

// IO Cell (0, 16, 1)
reg n1527;
always @(posedge clk) if (n6) n1527 <= n48;
assign \cypher[2]  = n1527;

// IO Cell (0, 19, 1)
reg n1528;
always @(posedge clk) if (n6) n1528 <= n111;
assign \cypher[30]  = n1528;

// IO Cell (0, 9, 0)
reg n1529;
always @(posedge clk) if (n6) n1529 <= n27;
assign \cypher[4]  = n1529;

// IO Cell (0, 4, 1)
reg n1530;
always @(posedge clk) if (n6) n1530 <= n7;
assign \cypher[26]  = n1530;

// IO Cell (0, 7, 1)
reg n1531;
always @(posedge clk) if (n6) n1531 <= n21;
assign \cypher[12]  = n1531;

// IO Cell (0, 14, 1)
reg n1532;
always @(posedge clk) if (n6) n1532 <= n46;
assign \cypher[7]  = n1532;

// IO Cell (0, 18, 0)
reg n1533;
always @(posedge clk) if (n6) n1533 <= n85;
assign \cypher[9]  = n1533;

// IO Cell (0, 8, 1)
reg n1534;
always @(posedge clk) if (n6) n1534 <= n25;
assign \cypher[3]  = n1534;

// IO Cell (0, 11, 1)
reg n1535;
always @(posedge clk) if (n6) n1535 <= n38;
assign \cypher[18]  = n1535;

// IO Cell (0, 6, 0)
reg n1536;
always @(posedge clk) if (n6) n1536 <= n15;
assign \cypher[25]  = n1536;

// IO Cell (0, 3, 0)
reg n1537;
always @(posedge clk) if (n6) n1537 <= n3;
assign \cypher[31]  = n1537;

// IO Cell (0, 20, 1)
reg n1538;
always @(posedge clk) if (n6) n1538 <= n129;
assign \cypher[11]  = n1538;

// IO Cell (0, 13, 0)
reg n1539;
always @(posedge clk) if (n6) n1539 <= n44;
assign \cypher[15]  = n1539;

// IO Cell (0, 10, 0)
reg n1540;
always @(posedge clk) if (n6) n1540 <= n31;
assign \cypher[17]  = n1540;

// IO Cell (0, 17, 1)
reg n1541;
always @(posedge clk) if (n6) n1541 <= n67;
assign \cypher[28]  = n1541;

assign n1797 = /* LUT   10 22  5 */ 1'b1;
assign n2010 = /* LUT    2 21  0 */ 1'b0;
assign n2413 = /* LUT   11 21  0 */ 1'b0;
assign n1542 = /* LUT    6 19  1 */ (n643 ? (ready ? \indata[30]  : 1'b1) : (ready ? \indata[30]  : 1'b0));
assign n938  = /* LUT    7 24  4 */ (n934 ? (n786 ? 1'b1 : !n811) : (n786 ? n811 : 1'b0));
assign n1544 = /* LUT   18 20  7 */ (n1465 ? 1'b1 : (n1461 ? 1'b1 : (n1471 ? 1'b1 : n1451)));
assign n1545 = /* LUT    4 25  6 */ (ds ? (n691 ? (ready ? 1'b0 : n77) : 1'b0) : (n691 ? (ready ? 1'b1 : n77) : 1'b0));
assign n1546 = /* LUT    9 23  2 */ (\indata[12]  ? (n1036 ? (\inExp[0]  ? 1'b1 : !ready) : (\inExp[0]  ? ready : 1'b0)) : (n1036 ? !ready : 1'b0));
assign n922  = /* LUT    7 22  0 */ (n878 ? 1'b0 : (reset ? 1'b0 : (n142 ? n49 : 1'b0)));
assign n1547 = /* LUT   10 22  7 */ !n1018;
assign n1548 = /* LUT    4 22  7 */ !n494;
assign n1426 = /* LUT   14 21  2 */ (n918 ? n1122 : n1201);
assign n1550 = /* LUT    5 24  5 */ (n529 ? (n253 ? n568 : 1'b1) : (n253 ? n568 : 1'b0));
assign n1551 = /* LUT   10 16  7 */ (n288 ? (ready ? \indata[6]  : 1'b1) : (ready ? \indata[6]  : 1'b0));
assign n1552 = /* LUT    5 19  4 */ (n643 ? (ds ? (ready ? 1'b0 : n77) : (ready ? 1'b1 : n77)) : 1'b0);
assign n1553 = /* LUT    2 25  3 */ (n523 ? n524 : 1'b0);
assign n1554 = /* LUT   10 26  7 */ (n1182 ? (n1078 ? n781 : !n781) : (n1078 ? !n781 : n781));
assign n1555 = /* LUT   11 17  4 */ \inMod[11] ;
assign n1556 = /* LUT   13 21  5 */ (n1373 ? (n955 ? n1307 : !n1307) : (n955 ? !n1307 : n1307));
assign n460  = /* LUT    2 19  3 */ (n88 ? (n133 ? n182 : 1'b1) : (n133 ? n182 : 1'b0));
assign n1558 = /* LUT   11 23  0 */ (n1247 ? (n177 ? n1065 : !n1065) : (n177 ? !n1065 : n1065));
assign n1559 = /* LUT    4 30  0 */ \inMod[15] ;
assign n1560 = /* LUT    5 17  5 */ !n636;
assign n1561 = /* LUT    1 25  2 */ (n423 ? (n421 ? n237 : !n237) : (n421 ? !n237 : n237));
assign n1562 = /* LUT   15 21  5 */ (n1423 ? (n568 ? 1'b1 : (n49 ? !n142 : 1'b1)) : (n568 ? (n49 ? n142 : 1'b0) : 1'b0));
assign n1133 = /* LUT   10 21  3 */ (n861 ? n1132 : n1130);
assign n1563 = /* LUT    6 18  6 */ (n741 ? (reset ? 1'b1 : (n99 ? 1'b1 : !n290)) : (reset ? 1'b0 : (n99 ? n290 : 1'b0)));
assign n1564 = /* LUT    5 27  1 */ (n801 ? (n178 ? n597 : !n597) : (n178 ? !n597 : n597));
assign n771  = /* LUT    5 22  6 */ (n708 ? (n507 ? n667 : 1'b1) : (n507 ? n667 : 1'b0));
assign n1566 = /* LUT   14 22  0 */ (n1135 ? n732 : 1'b0);
assign n1567 = /* LUT    2 26  7 */ (n530 ? n524 : 1'b0);
assign n1568 = /* LUT    6 20  6 */ (ready ? (\indata[1]  ? \inExp[0]  : 1'b0) : n872);
assign n572  = /* LUT    3 20  3 */ (n74 ? (n171 ? 1'b1 : !n133) : (n171 ? n133 : 1'b0));
assign n1570 = /* LUT    2 20  7 */ (n113 ? (n210 ? 1'b1 : !n133) : (n210 ? n133 : 1'b0));
assign n1571 = /* LUT    6 25  5 */ (n784 ? n524 : 1'b0);
assign n1572 = /* LUT   11 18  6 */ (n1192 ? n732 : 1'b0);
assign n1344 = /* LUT   12 27  5 */ (n861 ? n1343 : n1138);
assign n1573 = /* LUT   14 19  2 */ (n918 ? n1227 : 1'b0);
assign n1574 = /* LUT    5 30  1 */ (n624 ? (n717 ? 1'b1 : n507) : (n717 ? !n507 : 1'b0));
assign n1575 = /* LUT    3 22  6 */ (n253 ? (n190 ? (reset ? n481 : 1'b1) : (reset ? n481 : 1'b0)) : n481);
assign n1576 = /* LUT   13 16  0 */ (n44 ? (n1283 ? (n839 ? !n53 : 1'b1) : (n839 ? 1'b0 : n53)) : (n1283 ? !n53 : 1'b0));
assign n1577 = /* LUT   11 27  0 */ (n1142 ? (n1024 ? 1'b1 : (n861 ? n811 : 1'b1)) : (n1024 ? (n861 ? !n811 : 1'b0) : 1'b0));
assign n1578 = /* LUT    9 19  7 */ (n290 ? n945 : n1005);
assign n1579 = /* LUT    7 26  7 */ !n877;
assign n1580 = /* LUT    4 27  5 */ (n242 ? (ds ? (n77 ? !ready : 1'b0) : (n77 ? 1'b1 : ready)) : 1'b0);
assign n1581 = /* LUT    9 21  7 */ (n646 ? (ready ? \indata[9]  : 1'b1) : (ready ? \indata[9]  : 1'b0));
assign n1582 = /* LUT    7 16  7 */ (n835 ? 1'b0 : !reset);
assign n1583 = /* LUT    4 16  4 */ (n275 ? (n65 ? 1'b1 : (n49 ? n50 : 1'b0)) : (n65 ? (n49 ? !n50 : 1'b1) : 1'b0));
assign n1584 = /* LUT    5 23  1 */ (n598 ? (n751 ? 1'b1 : (n49 ? !n142 : 1'b1)) : (n751 ? (n49 ? n142 : 1'b0) : 1'b0));
assign n1585 = /* LUT   12 22  5 */ (n1332 ? (n585 ? n1310 : !n1310) : (n585 ? !n1310 : n1310));
assign n1586 = /* LUT    1 22  3 */ (n366 ? (n362 ? n360 : !n360) : (n362 ? !n360 : n360));
assign n1587 = /* LUT   13 19  6 */ (n1293 ? n732 : 1'b0);
assign n1588 = /* LUT   10 24  0 */ (n1151 ? (n1057 ? n850 : !n850) : (n1057 ? !n850 : n850));
assign n1589 = /* LUT    3 27  0 */ !n265;
assign n1590 = /* LUT    7 25  3 */ (n237 ? (n650 ? !n106 : (n106 ? 1'b0 : !n157)) : (n650 ? (n106 ? 1'b0 : n157) : 1'b0));
assign n1591 = /* LUT    4 18  5 */ \inMod[6] ;
assign n1592 = /* LUT    7 23  3 */ (n469 ? (ready ? \indata[29]  : 1'b1) : (ready ? \indata[29]  : 1'b0));
assign n1593 = /* LUT   14 18  5 */ (n1279 ? (n1410 ? 1'b1 : n290) : (n1410 ? !n290 : 1'b0));
assign n1594 = /* LUT    1 20  6 */ (n332 ? (n208 ? n217 : !n217) : (n208 ? !n217 : n217));
assign n680  = /* LUT    4 24  1 */ (n507 ? n673 : n599);
assign n1596 = /* LUT    4 21  6 */ (n116 ? (n213 ? 1'b1 : !n133) : (n213 ? n133 : 1'b0));
assign n1597 = /* LUT   14 20  1 */ (n1417 ? (n142 ? (n49 ? n174 : 1'b1) : 1'b1) : (n142 ? (n49 ? n174 : 1'b0) : 1'b0));
assign n1598 = /* LUT    5 25  6 */ (n676 ? (n693 ? 1'b1 : n507) : (n693 ? !n507 : 1'b0));
assign n1599 = /* LUT    5 20  5 */ (ready ? (n754 ? !ds : 1'b0) : (n754 ? n77 : 1'b0));
assign n1600 = /* LUT    1 17  7 */ (n284 ? (n155 ? n181 : !n181) : (n155 ? !n181 : n181));
assign n1601 = /* LUT    2 24  0 */ (n502 ? (n233 ? n210 : !n210) : (n233 ? !n210 : n210));
assign n1602 = /* LUT   13 22  4 */ (n1383 ? (n1117 ? n974 : !n974) : (n1117 ? !n974 : n974));
assign n1603 = /* LUT   16 23  6 */ (n1413 ? (n719 ? 1'b1 : (n49 ? !n142 : 1'b1)) : (n719 ? (n49 ? n142 : 1'b0) : 1'b0));
assign n1604 = /* LUT    2 18  4 */ (n339 ? (n451 ? 1'b1 : !n324) : (n451 ? n324 : 1'b0));
assign n1218 = /* LUT   11 20  1 */ (n649 ? (n918 ? 1'b1 : n1210) : (n918 ? 1'b0 : n1210));
assign n1606 = /* LUT    5 18  4 */ !n739;
assign n1607 = /* LUT   12 19  0 */ (n732 ? n1195 : 1'b0);
assign n1609 = /* LUT    5 28  0 */ (n808 ? (n234 ? n667 : !n667) : (n234 ? !n667 : n667));
assign n1610 = /* LUT   10 20  0 */ (n46 ? (\indata[7]  ? (ready ? \inExp[0]  : 1'b1) : !ready) : (\indata[7]  ? (ready ? \inExp[0]  : 1'b0) : 1'b0));
assign n1611 = /* LUT    6 23  7 */ (n820 ? (n885 ? 1'b1 : !n253) : (n885 ? n253 : 1'b0));
assign n582  = /* LUT    3 21  4 */ (n117 ? (n214 ? 1'b1 : !n133) : (n214 ? n133 : 1'b0));
assign n1613 = /* LUT    4 20  1 */ (reset ? n140 : (n140 ? (n253 ? n456 : 1'b1) : (n253 ? n456 : 1'b0)));
assign n1614 = /* LUT    2 23  6 */ (n500 ? (n128 ? n198 : !n198) : (n128 ? !n198 : n198));
assign n889  = /* LUT    6 24  6 */ (n507 ? n778 : n698);
assign n1616 = /* LUT   16 25  3 */ (n242 ? (ready ? \indata[16]  : 1'b1) : (ready ? \indata[16]  : 1'b0));
assign n1083 = /* LUT    9 27  4 */ (n811 ? n906 : n1052);
assign n1209 = /* LUT   11 19  5 */ (n1207 ? (n918 ? n1115 : 1'b1) : (n918 ? n1115 : 1'b0));
assign n1619 = /* LUT   17 21  5 */ (ready ? (ds ? \inExp[31]  : 1'b0) : 1'b0);
assign n1620 = /* LUT   13 23  3 */ (n1392 ? (n1286 ? n1060 : !n1060) : (n1286 ? !n1060 : n1060));
assign n1621 = /* LUT    3 23  5 */ (n256 ? (n506 ? 1'b1 : n507) : (n506 ? !n507 : 1'b0));
assign n1622 = /* LUT   15 23  2 */ (n1433 ? (n678 ? 1'b1 : (n142 ? !n49 : 1'b1)) : (n678 ? (n142 ? n49 : 1'b0) : 1'b0));
assign n1623 = /* LUT    6 16  3 */ (n546 ? (n50 ? (n49 ? n537 : 1'b1) : 1'b1) : (n50 ? (n49 ? n537 : 1'b0) : 1'b0));
assign n1624 = /* LUT    4 28  6 */ (n439 ? (n617 ? 1'b1 : n507) : (n617 ? !n507 : 1'b0));
assign n1625 = /* LUT   11 24  1 */ (n1267 ? (n1076 ? n981 : !n981) : (n1076 ? !n981 : n981));
assign n1626 = /* LUT    9 22  6 */ (n157 ? (n175 ? n253 : 1'b0) : n969);
assign n1627 = /* LUT    4 23  5 */ (reset ? n591 : (n591 ? (n290 ? n238 : 1'b1) : (n290 ? n238 : 1'b0)));
assign n1628 = /* LUT    7 15  4 */ (n838 ? (n49 ? 1'b0 : n50) : (n913 ? (n49 ? 1'b0 : n50) : (n49 ? !n50 : 1'b1)));
assign n1629 = /* LUT    9 24  6 */ (\indata[4]  ? (n1048 ? (\inExp[0]  ? 1'b1 : !ready) : (\inExp[0]  ? ready : 1'b0)) : (n1048 ? !ready : 1'b0));
assign n1630 = /* LUT   10 17  5 */ (n650 ? (ready ? \indata[26]  : 1'b1) : (ready ? \indata[26]  : 1'b0));
assign n1631 = /* LUT   12 21  4 */ (n1322 ? (n1288 ? n849 : !n849) : (n1288 ? !n849 : n849));
assign n1632 = /* LUT   18 19  4 */ (n1488 ? (\inExp[9]  ? 1'b1 : (ready ? !ds : 1'b1)) : (\inExp[9]  ? (ready ? ds : 1'b0) : 1'b0));
assign n1633 = /* LUT    1 23  4 */ (n385 ? (n380 ? n126 : !n126) : (n380 ? !n126 : n126));
assign n1634 = /* LUT    2 22  1 */ (n483 ? (n292 ? n167 : !n167) : (n292 ? !n167 : n167));
assign n1635 = /* LUT   13 20  7 */ (n25 ? (n839 ? 1'b0 : (n53 ? 1'b1 : n1309)) : (n839 ? 1'b0 : (n53 ? 1'b0 : n1309)));
assign n1185 = /* LUT   10 27  1 */ (n1184 ? (n1085 ? n344 : !n344) : (n1085 ? !n344 : n344));
assign n1507 = /* LUT   19 20  2 */ (n1467 ? 1'b1 : (n1469 ? 1'b1 : (n1466 ? 1'b1 : n1468)));
assign n1637 = /* LUT    3 24  1 */ (n434 ? (n220 ? !n106 : (n157 ? !n106 : 1'b0)) : (n220 ? (n157 ? 1'b0 : !n106) : 1'b0));
assign n1638 = /* LUT    7 30  2 */ \inMod[24] ;
assign n1639 = /* LUT   11 22  0 */ (n1237 ? (n932 ? n1057 : !n1057) : (n932 ? !n1057 : n1057));
assign n1640 = /* LUT    7 20  2 */ (n123 ? (n53 ? !n839 : n663) : (n53 ? 1'b0 : n663));
assign n1641 = /* LUT    9 17  0 */ (n8 ? (\indata[6]  ? (\inExp[0]  ? 1'b1 : !ready) : !ready) : (\indata[6]  ? (\inExp[0]  ? ready : 1'b0) : 1'b0));
assign n1642 = /* LUT    5 16  7 */ (n729 ? (n50 ? (n49 ? n647 : 1'b1) : 1'b1) : (n50 ? (n49 ? n647 : 1'b0) : 1'b0));
assign n1643 = /* LUT    1 21  5 */ (n70 ? (n167 ? 1'b1 : !n133) : (n167 ? n133 : 1'b0));
assign n1644 = /* LUT    1 24  6 */ (n407 ? (n224 ? n225 : !n225) : (n224 ? !n225 : n225));
assign n1645 = /* LUT    5 26  7 */ (n799 ? (n181 ? n673 : !n673) : (n181 ? !n673 : n673));
assign n1111 = /* LUT   10 18  1 */ (n1110 ? (n956 ? 1'b1 : n918) : (n956 ? !n918 : 1'b0));
assign n1647 = /* LUT   14 23  0 */ (n1141 ? (n918 ? 1'b1 : n1229) : (n918 ? 1'b0 : n1229));
assign n1648 = /* LUT    5 21  6 */ (n77 ? (n761 ? (ready ? !ds : 1'b1) : 1'b0) : (n761 ? (ready ? !ds : 1'b0) : 1'b0));
assign n1649 = /* LUT    1 18  6 */ (n298 ? (n172 ? n104 : !n104) : (n172 ? !n104 : n104));
assign n1650 = /* LUT   19 19  4 */ (n1489 ? (\inExp[26]  ? 1'b1 : (ds ? !ready : 1'b1)) : (\inExp[26]  ? (ds ? ready : 1'b0) : 1'b0));
assign n1651 = /* LUT    6 21  2 */ (n337 ? (n874 ? 1'b1 : !n324) : (n874 ? n324 : 1'b0));
assign n1459 = /* LUT   16 22  5 */ (n1432 ? 1'b1 : (n1365 ? 1'b1 : (n1436 ? 1'b1 : n1419)));
assign n1653 = /* LUT    2 21  5 */ (n476 ? (n80 ? n153 : !n153) : (n80 ? !n153 : n153));
assign n1654 = /* LUT   11 21  6 */ (n1235 ? (n121 ? n1042 : !n1042) : (n121 ? !n1042 : n1042));
assign n1655 = /* LUT   12 20  3 */ (n1313 ? (n1095 ? n1115 : !n1115) : (n1095 ? !n1115 : n1115));
assign n1656 = /* LUT    5 19  3 */ (n77 ? (n747 ? (ds ? !ready : 1'b1) : 1'b0) : (n747 ? (ds ? 1'b0 : ready) : 1'b0));
assign n1291 = /* LUT   12 18  3 */ (n1195 ? (n1290 ? n344 : !n344) : (n1290 ? !n344 : n344));
assign n1658 = /* LUT    5 29  3 */ (n824 ? (n145 ? n623 : !n623) : (n145 ? !n623 : n623));
assign n1659 = /* LUT    3 25  6 */ (ready ? (n609 ? !ds : 1'b0) : (n609 ? n77 : 1'b0));
assign n1660 = /* LUT    2 19  4 */ (n342 ? (n460 ? 1'b1 : !n324) : (n460 ? n324 : 1'b0));
assign n1661 = /* LUT    6 28  4 */ (n707 ? (n712 ? 1'b1 : n507) : (n712 ? !n507 : 1'b0));
assign n1662 = /* LUT   10 23  1 */ (n1144 ? (n1041 ? n1094 : !n1094) : (n1041 ? !n1094 : n1094));
assign n1663 = /* LUT    6 22  0 */ (n524 ? n774 : 1'b0);
assign n1664 = /* LUT    7 21  5 */ (n60 ? (n151 ? 1'b1 : !n133) : (n151 ? n133 : 1'b0));
assign n1665 = /* LUT    3 18  5 */ !n559;
assign n1666 = /* LUT    7 19  1 */ !n738;
assign n1667 = /* LUT    9 20  5 */ (n605 ? n524 : 1'b0);
assign n1668 = /* LUT    1 19  1 */ (n308 ? (n182 ? n185 : !n185) : (n182 ? !n185 : n185));
assign n1669 = /* LUT   12 23  7 */ (n1108 ? n732 : 1'b0);
assign n1670 = /* LUT   13 24  2 */ (n1400 ? (n1249 ? n1103 : !n1103) : (n1249 ? !n1103 : n1103));
assign n1671 = /* LUT    3 20  4 */ (n349 ? (n572 ? 1'b1 : !n324) : (n572 ? n324 : 1'b0));
assign n1672 = /* LUT   19 22  1 */ (n1500 ? (\inExp[17]  ? 1'b1 : (ds ? !ready : 1'b1)) : (\inExp[17]  ? (ds ? ready : 1'b0) : 1'b0));
assign n1673 = /* LUT    6 25  2 */ (n707 ? n524 : 1'b0);
assign n1674 = /* LUT   13 18  2 */ (n290 ? n988 : n1349);
assign n1675 = /* LUT   10 25  0 */ (n1162 ? (n1065 ? n767 : !n767) : (n1065 ? !n767 : n767));
assign n1676 = /* LUT    6 19  2 */ (ready ? (\inExp[0]  ? \indata[31]  : 1'b0) : n3);
assign n1677 = /* LUT    3 26  0 */ (n602 ? (ready ? \indata[21]  : 1'b1) : (ready ? \indata[21]  : 1'b0));
assign n939  = /* LUT    7 24  5 */ (n861 ? n938 : n933);
assign n1678 = /* LUT   18 20  6 */ (n1467 ? (\inExp[24]  ? 1'b1 : (ds ? !ready : 1'b1)) : (\inExp[24]  ? (ds ? ready : 1'b0) : 1'b0));
assign n1679 = /* LUT    4 19  7 */ (n146 ? (n157 ? !n106 : (n320 ? !n106 : 1'b0)) : (n157 ? 1'b0 : (n320 ? !n106 : 1'b0)));
assign n1680 = /* LUT    4 25  7 */ (n601 ? (ready ? !ds : n77) : 1'b0);
assign n1036 = /* LUT    9 23  1 */ (n982 ? (n1035 ? 1'b1 : !n861) : (n1035 ? n861 : 1'b0));
assign n1681 = /* LUT   10 22  6 */ (n21 ? (n53 ? !n839 : n974) : (n53 ? 1'b0 : n974));
assign n1682 = /* LUT    7 22  1 */ (n756 ? (n922 ? 1'b0 : (n360 ? 1'b1 : n157)) : (n922 ? 1'b0 : (n360 ? !n157 : 1'b0)));
assign n1683 = /* LUT    4 22  6 */ (n586 ? (n253 ? (reset ? 1'b1 : n671) : 1'b1) : (n253 ? (reset ? 1'b0 : n671) : 1'b0));
assign n1684 = /* LUT   14 21  3 */ (n743 ? (n1426 ? 1'b1 : n290) : (n1426 ? !n290 : 1'b0));
assign n1685 = /* LUT    5 24  2 */ (n439 ? n524 : 1'b0);
assign n1686 = /* LUT    2 25  0 */ (n515 ? (n291 ? n230 : !n230) : (n291 ? !n230 : n230));
assign n1687 = /* LUT   10 26  6 */ (n1181 ? (n1077 ? n737 : !n737) : (n1077 ? !n737 : n737));
assign n1688 = /* LUT   11 17  3 */ \inMod[10] ;
assign n1689 = /* LUT   13 21  4 */ (n1372 ? (n954 ? n1308 : !n1308) : (n954 ? !n1308 : n1308));
assign n1690 = /* LUT   19 21  5 */ (n1443 ? 1'b1 : (n1450 ? 1'b1 : (n1463 ? 1'b1 : n1457)));
assign n1691 = /* LUT    4 16  3 */ (n633 ? (n446 ? 1'b1 : (n50 ? !n49 : 1'b1)) : (n446 ? (n50 ? n49 : 1'b0) : 1'b0));
assign n1692 = /* LUT   11 23  3 */ (n1257 ? (n734 ? n906 : !n906) : (n734 ? !n906 : n906));
assign n1693 = /* LUT    4 30  3 */ \inMod[18] ;
assign n1694 = /* LUT    1 22  4 */ (n367 ? (n179 ? n363 : !n363) : (n179 ? !n363 : n363));
assign n1695 = /* LUT    1 25  5 */ (n426 ? (n419 ? n415 : !n415) : (n419 ? !n415 : n415));
assign n1696 = /* LUT   15 21  4 */ (n142 ? (n49 ? n535 : n1442) : n1442);
assign n1697 = /* LUT   14 22  7 */ (n1009 ? (n1431 ? 1'b1 : n290) : (n1431 ? !n290 : 1'b0));
assign n1698 = /* LUT    5 27  0 */ (n800 ? (n292 ? n596 : !n596) : (n292 ? !n596 : n596));
assign n1131 = /* LUT   10 21  0 */ (n1061 ? (n811 ? n1075 : 1'b1) : (n811 ? n1075 : 1'b0));
assign n1700 = /* LUT    5 22  7 */ (n174 ? (n771 ? 1'b1 : n253) : (n771 ? !n253 : 1'b0));
assign n871  = /* LUT    6 20  1 */ (n616 ? (n861 ? 1'b1 : n858) : (n861 ? 1'b0 : n858));
assign n1701 = /* LUT   11 18  7 */ !n1193;
assign n1702 = /* LUT   12 27  2 */ (\indata[16]  ? (n1342 ? (\inExp[0]  ? 1'b1 : !ready) : (\inExp[0]  ? ready : 1'b0)) : (n1342 ? !ready : 1'b0));
assign n753  = /* LUT    5 20  2 */ (n133 ? n148 : (n57 ? (n148 ? 1'b1 : n324) : (n148 ? !n324 : 1'b0)));
assign n1703 = /* LUT   14 19  3 */ (n1214 ? n732 : 1'b0);
assign n1704 = /* LUT    3 22  7 */ (n482 ? (reset ? 1'b1 : (n176 ? 1'b1 : !n253)) : (reset ? 1'b0 : (n176 ? n253 : 1'b0)));
assign n451  = /* LUT    2 18  3 */ (n64 ? (n155 ? 1'b1 : !n133) : (n155 ? n133 : 1'b0));
assign n1706 = /* LUT   13 16  1 */ (n8 ? (n1284 ? !n839 : (n53 ? !n839 : 1'b0)) : (n1284 ? (n53 ? 1'b0 : !n839) : 1'b0));
assign n1707 = /* LUT    3 28  7 */ (n614 ? (n535 ? 1'b1 : !n253) : (n535 ? n253 : 1'b0));
assign n1708 = /* LUT   11 27  3 */ (n1153 ? (n1280 ? 1'b1 : !n861) : (n1280 ? n861 : 1'b0));
assign n1709 = /* LUT    6 17  1 */ !n765;
assign n1710 = /* LUT    7 26  4 */ !n902;
assign n1711 = /* LUT    3 19  6 */ (ready ? ds : 1'b1);
assign n1005 = /* LUT    9 19  6 */ (n918 ? n952 : n1002);
assign n1713 = /* LUT    7 16  0 */ (n736 ? (n569 ? 1'b1 : (n50 ? !n49 : 1'b1)) : (n569 ? (n50 ? n49 : 1'b0) : 1'b0));
assign n1714 = /* LUT   12 24  0 */ (n29 ? (n53 ? !n839 : n1263) : (n53 ? 1'b0 : n1263));
assign n1715 = /* LUT    9 21  6 */ (n67 ? (\inExp[0]  ? (\indata[28]  ? 1'b1 : !ready) : !ready) : (\inExp[0]  ? (\indata[28]  ? ready : 1'b0) : 1'b0));
assign n1716 = /* LUT    5 23  0 */ (n200 ? (n202 ? 1'b1 : (n142 ? !n49 : 1'b1)) : (n202 ? (n142 ? n49 : 1'b0) : 1'b0));
assign n1717 = /* LUT   12 22  4 */ (n1331 ? (n684 ? n1001 : !n1001) : (n684 ? !n1001 : n1001));
assign n1718 = /* LUT   13 25  1 */ (n1407 ? (n1398 ? n1340 : !n1340) : (n1398 ? !n1340 : n1340));
assign n1719 = /* LUT    3 21  3 */ (ready ? (n581 ? !ds : 1'b0) : (n581 ? n77 : 1'b0));
assign n1720 = /* LUT   13 19  5 */ (n290 ? n1006 : n1359);
assign n1721 = /* LUT   10 24  3 */ (n1157 ? (n433 ? n1095 : !n1095) : (n433 ? !n1095 : n1095));
assign n1722 = /* LUT    3 27  3 */ !n533;
assign n1723 = /* LUT    4 18  4 */ \inMod[5] ;
assign n1724 = /* LUT    7 23  2 */ (\indata[29]  ? (n929 ? (\inExp[0]  ? 1'b1 : !ready) : (\inExp[0]  ? ready : 1'b0)) : (n929 ? !ready : 1'b0));
assign n1725 = /* LUT    4 24  0 */ (n673 ? n524 : 1'b0);
assign n1726 = /* LUT    1 20  7 */ (n333 ? (n215 ? n291 : !n291) : (n215 ? !n291 : n291));
assign n1410 = /* LUT   14 18  4 */ (n1310 ? (n918 ? 1'b1 : n1239) : (n918 ? 1'b0 : n1239));
assign n1728 = /* LUT    4 21  7 */ (n469 ? (n415 ? !n106 : (n157 ? !n106 : 1'b0)) : (n415 ? (n157 ? 1'b0 : !n106) : 1'b0));
assign n1729 = /* LUT   14 20  0 */ (n1361 ? 1'b1 : (n1363 ? 1'b1 : (n783 ? 1'b1 : n1362)));
assign n1730 = /* LUT    5 25  1 */ (n589 ? (n507 ? 1'b1 : n692) : (n507 ? 1'b0 : n692));
assign n1731 = /* LUT   10 19  7 */ (n78 ? (n654 ? 1'b1 : (n49 ? !n50 : 1'b1)) : (n654 ? (n49 ? n50 : 1'b0) : 1'b0));
assign n1073 = /* LUT    9 26  4 */ (n1056 ? (n1069 ? 1'b1 : !n811) : (n1069 ? n811 : 1'b0));
assign n1733 = /* LUT    1 17  6 */ (n283 ? (n154 ? n274 : !n274) : (n154 ? !n274 : n274));
assign n1734 = /* LUT    2 24  3 */ (n510 ? (n160 ? n213 : !n213) : (n160 ? !n213 : n213));
assign n1735 = /* LUT   13 22  5 */ (n1384 ? (n996 ? n967 : !n967) : (n996 ? !n967 : n967));
assign n1736 = /* LUT    4 23  2 */ (n666 ? n524 : 1'b0);
assign n1737 = /* LUT   11 20  2 */ (n290 ? n1211 : n1218);
assign n1738 = /* LUT    5 18  5 */ (reset ? n640 : (n640 ? (n253 ? n554 : 1'b1) : (n253 ? n554 : 1'b0)));
assign n1739 = /* LUT    1 23  3 */ (n384 ? (n340 ? n378 : !n378) : (n340 ? !n378 : n378));
assign n1740 = /* LUT   12 19  1 */ (n1296 ? (n1094 ? n1122 : !n1122) : (n1094 ? !n1122 : n1122));
assign n1741 = /* LUT    1 26  4 */ !n236;
assign n1742 = /* LUT    5 28  1 */ (n812 ? (n185 ? n668 : !n668) : (n185 ? !n668 : n668));
assign n1127 = /* LUT   10 20  3 */ (n861 ? n1126 : n1123);
assign n1743 = /* LUT    6 23  0 */ (n780 ? (n253 ? n503 : 1'b1) : (n253 ? n503 : 1'b0));
assign n1744 = /* LUT    4 20  0 */ (n565 ? (reset ? 1'b1 : (n553 ? 1'b1 : !n253)) : (reset ? 1'b0 : (n553 ? n253 : 1'b0)));
assign n1745 = /* LUT    2 23  7 */ (n501 ? (n235 ? n199 : !n199) : (n235 ? !n199 : n199));
assign n1746 = /* LUT    7 18  3 */ !n741;
assign n1747 = /* LUT    9 27  3 */ (n303 ? (ready ? \indata[18]  : 1'b1) : (ready ? \indata[18]  : 1'b0));
assign n1748 = /* LUT   11 19  4 */ (n1115 ? n732 : 1'b0);
assign n1749 = /* LUT   17 21  4 */ (n1443 ? (ds ? (\inExp[15]  ? 1'b1 : !ready) : 1'b1) : (ds ? (\inExp[15]  ? ready : 1'b0) : 1'b0));
assign n759  = /* LUT    5 21  1 */ (n115 ? (n212 ? 1'b1 : !n133) : (n212 ? n133 : 1'b0));
assign n1751 = /* LUT   13 23  2 */ (n1391 ? (n947 ? n1248 : !n1248) : (n947 ? !n1248 : n1248));
assign n1752 = /* LUT    2 21  2 */ (n473 ? (n277 ? n150 : !n150) : (n277 ? !n150 : n150));
assign n1753 = /* LUT   15 23  5 */ (n1436 ? (n885 ? 1'b1 : (n49 ? !n142 : 1'b1)) : (n885 ? (n49 ? n142 : 1'b0) : 1'b0));
assign n1754 = /* LUT    4 28  5 */ (n523 ? (n507 ? 1'b1 : n714) : (n507 ? 1'b0 : n714));
assign n1755 = /* LUT   11 24  2 */ (n1268 ? (n893 ? n900 : !n900) : (n893 ? !n900 : n900));
assign n700  = /* LUT    4 26  1 */ (n699 ? (n507 ? n257 : 1'b1) : (n507 ? n257 : 1'b0));
assign n1757 = /* LUT    9 24  7 */ (n755 ? (ready ? \indata[4]  : 1'b1) : (ready ? \indata[4]  : 1'b0));
assign n1099 = /* LUT   10 17  2 */ (n995 ? (n894 ? 1'b1 : !n811) : (n894 ? n811 : 1'b0));
assign n1759 = /* LUT   12 21  5 */ (n1323 ? (n890 ? n957 : !n957) : (n890 ? !n957 : n957));
assign n1760 = /* LUT    3 18  2 */ (n325 ? (n453 ? !n106 : (n157 ? 1'b0 : !n106)) : (n453 ? (n157 ? !n106 : 1'b0) : 1'b0));
assign n1761 = /* LUT    2 22  0 */ (n479 ? (n181 ? n166 : !n166) : (n181 ? !n166 : n166));
assign n1762 = /* LUT   13 20  4 */ (n1306 ? (n164 ? !n839 : (n839 ? 1'b0 : !n53)) : (n164 ? (n839 ? 1'b0 : n53) : 1'b0));
assign n1763 = /* LUT   10 27  2 */ (n1041 ? (n1185 ? 1'b1 : n1025) : (n1185 ? 1'b0 : n1025));
assign n1508 = /* LUT   19 20  3 */ (n1496 ? 1'b1 : (n1507 ? 1'b1 : (n1472 ? 1'b1 : n1473)));
assign n1765 = /* LUT    3 24  2 */ (n221 ? (n242 ? !n106 : (n106 ? 1'b0 : !n157)) : (n242 ? (n106 ? 1'b0 : n157) : 1'b0));
assign n1766 = /* LUT    4 17  5 */ (n50 ? (n240 ? (n547 ? 1'b1 : n49) : (n547 ? !n49 : 1'b0)) : n547);
assign n1767 = /* LUT    7 30  3 */ \inMod[25] ;
assign n1768 = /* LUT   11 22  1 */ (n1240 ? (n850 ? n970 : !n970) : (n850 ? !n970 : n970));
assign n1769 = /* LUT    5 16  4 */ (n548 ? (n50 ? (n656 ? 1'b1 : !n49) : 1'b1) : (n50 ? (n656 ? n49 : 1'b0) : 1'b0));
assign n1770 = /* LUT   19 22  6 */ (n1499 ? (\inExp[16]  ? 1'b1 : (ready ? !ds : 1'b1)) : (\inExp[16]  ? (ready ? ds : 1'b0) : 1'b0));
assign n1771 = /* LUT    1 24  7 */ (n408 ? (n355 ? n220 : !n220) : (n355 ? !n220 : n220));
assign n1772 = /* LUT    5 26  0 */ (n792 ? (n83 ? n589 : !n589) : (n83 ? !n589 : n589));
assign n1773 = /* LUT   10 18  0 */ (n997 ? n732 : 1'b0);
assign n1437 = /* LUT   14 23  1 */ (n1327 ? (n1228 ? 1'b1 : n918) : (n1228 ? !n918 : 1'b0));
assign n1775 = /* LUT   18 20  1 */ (n1470 ? (\inExp[19]  ? 1'b1 : (ready ? !ds : 1'b1)) : (\inExp[19]  ? (ready ? ds : 1'b0) : 1'b0));
assign n1776 = /* LUT    1 18  7 */ (n299 ? (n173 ? n107 : !n107) : (n173 ? !n107 : n107));
assign n875  = /* LUT    6 21  3 */ (n873 ? (n324 ? 1'b1 : n156) : (n324 ? 1'b0 : n156));
assign n1777 = /* LUT    4 22  1 */ (ds ? 1'b1 : !ready);
assign n1778 = /* LUT   11 21  5 */ (n1234 ? (n669 ? n1040 : !n1040) : (n669 ? !n1040 : n1040));
assign n1779 = /* LUT   12 20  2 */ (n1312 ? (n1106 ? n1114 : !n1114) : (n1106 ? !n1114 : n1114));
assign n747  = /* LUT    5 19  2 */ (n648 ? (n124 ? 1'b1 : n324) : (n124 ? !n324 : 1'b0));
assign n1780 = /* LUT    6 26  7 */ !n789;
assign n1290 = /* LUT   12 18  2 */ !n1196;
assign n1781 = /* LUT    5 29  2 */ (n823 ? (n160 ? n530 : !n530) : (n160 ? !n530 : n530));
assign n609  = /* LUT    3 25  5 */ (n319 ? (n324 ? 1'b1 : n390) : (n324 ? 1'b0 : n390));
assign n461  = /* LUT    2 19  5 */ (n318 ? (n324 ? 1'b1 : n343) : (n324 ? 1'b0 : n343));
assign n1782 = /* LUT   10 23  2 */ (n1145 ? (n745 ? n853 : !n853) : (n745 ? !n853 : n853));
assign n1783 = /* LUT    6 22  7 */ !n762;
assign n1784 = /* LUT    7 19  0 */ !n846;
assign n1785 = /* LUT    9 20  2 */ (n520 ? n524 : 1'b0);
assign n1786 = /* LUT    1 19  0 */ (n300 ? (n193 ? n234 : !n234) : (n193 ? !n234 : n234));
assign n1787 = /* LUT   12 23  4 */ (n1119 ? n732 : 1'b0);
assign n1788 = /* LUT   13 24  3 */ (n1401 ? (n1253 ? n1104 : !n1104) : (n1253 ? !n1104 : n1104));
assign n573  = /* LUT    3 20  5 */ (n317 ? (n324 ? 1'b1 : n350) : (n324 ? 1'b0 : n350));
assign n1350 = /* LUT   13 18  3 */ (n918 ? n1287 : n1222);
assign n1790 = /* LUT   10 25  1 */ (n1163 ? (n1066 ? n1019 : !n1019) : (n1066 ? !n1019 : n1019));
assign n1791 = /* LUT   15 20  4 */ (n1422 ? (n538 ? 1'b1 : (n49 ? !n142 : 1'b1)) : (n538 ? (n49 ? n142 : 1'b0) : 1'b0));
assign n1792 = /* LUT    6 19  3 */ (n652 ? (ready ? \indata[31]  : 1'b1) : (ready ? \indata[31]  : 1'b0));
assign n1793 = /* LUT    7 24  6 */ (\indata[15]  ? (n939 ? (\inExp[0]  ? 1'b1 : !ready) : (\inExp[0]  ? ready : 1'b0)) : (n939 ? !ready : 1'b0));
assign n1794 = /* LUT    4 19  4 */ !n560;
assign n688  = /* LUT    4 25  0 */ (n90 ? (n195 ? 1'b1 : !n133) : (n195 ? n133 : 1'b0));
assign n1796 = /* LUT    7 22  6 */ (n755 ? (n924 ? !n106 : (n179 ? !n106 : 1'b0)) : (n924 ? 1'b0 : (n179 ? !n106 : 1'b0)));
assign n1035 = /* LUT    9 23  0 */ (n1034 ? (n1030 ? 1'b1 : !n811) : (n1030 ? n811 : 1'b0));
assign n1799 = /* LUT   14 21  0 */ (n1194 ? (n290 ? n744 : 1'b1) : (n290 ? n744 : 1'b0));
assign n1800 = /* LUT    5 24  3 */ (n682 ? (n253 ? n670 : 1'b1) : (n253 ? n670 : 1'b0));
assign n1801 = /* LUT   10 16  1 */ (n861 ? n1092 : n1091);
assign n1802 = /* LUT    9 25  4 */ !n527;
assign n562  = /* LUT    3 19  1 */ (n336 ? (n561 ? 1'b1 : !n324) : (n561 ? n324 : 1'b0));
assign n1803 = /* LUT    2 25  1 */ (n525 ? (n344 ? n231 : !n231) : (n344 ? !n231 : n231));
assign n1804 = /* LUT   10 26  5 */ (n1180 ? (n779 ? n585 : !n585) : (n779 ? !n585 : n585));
assign n1805 = /* LUT   11 17  2 */ \inMod[1] ;
assign n1806 = /* LUT   13 21  7 */ (n1375 ? (n1294 ? n1305 : !n1305) : (n1294 ? !n1305 : n1305));
assign n1807 = /* LUT    4 16  2 */ (n634 ? (n603 ? 1'b1 : (n49 ? !n50 : 1'b1)) : (n603 ? (n49 ? n50 : 1'b0) : 1'b0));
assign n1808 = /* LUT    5 23  7 */ (n253 ? n751 : n777);
assign n1809 = /* LUT   11 23  2 */ (n1256 ? (n1019 ? n1059 : !n1059) : (n1019 ? !n1059 : n1059));
assign n1810 = /* LUT    4 30  2 */ \inMod[17] ;
assign n1811 = /* LUT    5 17  7 */ !n641;
assign n1812 = /* LUT    1 22  5 */ (n368 ? (n187 ? n183 : !n183) : (n187 ? !n183 : n183));
assign n1813 = /* LUT    1 25  4 */ (n425 ? (n245 ? n243 : !n243) : (n245 ? !n243 : n243));
assign n1814 = /* LUT   15 21  3 */ (n49 ? (n541 ? (n142 ? 1'b1 : n1365) : (n142 ? 1'b0 : n1365)) : n1365);
assign n1815 = /* LUT   10 21  1 */ (n861 ? n1131 : n1129);
assign n1816 = /* LUT    6 18  4 */ (n740 ? (reset ? 1'b1 : (n554 ? 1'b1 : !n290)) : (reset ? 1'b0 : (n554 ? n290 : 1'b0)));
assign n1817 = /* LUT    5 27  7 */ (n807 ? (n107 ? n666 : !n666) : (n107 ? !n666 : n666));
assign n1431 = /* LUT   14 22  6 */ (n918 ? n1136 : n1225);
assign n1819 = /* LUT    2 26  5 */ (n524 ? n256 : 1'b0);
assign n1820 = /* LUT   11 28  0 */ \inMod[9] ;
assign n1821 = /* LUT    4 21  0 */ !n565;
assign n1822 = /* LUT   11 18  4 */ (n190 ? (n290 ? (reset ? n1105 : 1'b1) : n1105) : (n290 ? (reset ? n1105 : 1'b0) : n1105));
assign n1823 = /* LUT    5 20  3 */ (ready ? (n753 ? 1'b1 : ds) : (n753 ? 1'b1 : !n77));
assign n1824 = /* LUT    1 17  1 */ (n278 ? (n149 ? n277 : !n277) : (n149 ? !n277 : n277));
assign n1825 = /* LUT   14 19  4 */ (n1212 ? n732 : 1'b0);
assign n1826 = /* LUT    5 30  3 */ (n530 ? (n715 ? 1'b1 : n507) : (n715 ? !n507 : 1'b0));
assign n1827 = /* LUT    3 22  4 */ (n480 ? (n290 ? (reset ? 1'b1 : n262) : 1'b1) : (n290 ? (reset ? 1'b0 : n262) : 1'b0));
assign n1280 = /* LUT   11 27  2 */ (n1064 ? (n1078 ? 1'b1 : !n811) : (n1078 ? n811 : 1'b0));
assign n1829 = /* LUT    3 15  7 */ (n52 ? (n468 ? 1'b1 : (n49 ? !n50 : 1'b1)) : (n468 ? (n49 ? n50 : 1'b0) : 1'b0));
assign n1830 = /* LUT    9 19  5 */ (n952 ? n732 : 1'b0);
assign n1831 = /* LUT   12 19  6 */ (n1301 ? (n855 ? n866 : !n866) : (n855 ? !n866 : n866));
assign n1832 = /* LUT    7 26  5 */ !n904;
assign n1833 = /* LUT    7 16  1 */ (n543 ? (n445 ? 1'b1 : (n49 ? !n50 : 1'b1)) : (n445 ? (n49 ? n50 : 1'b0) : 1'b0));
assign n1834 = /* LUT   12 24  7 */ (n31 ? (n1266 ? (n839 ? !n53 : 1'b1) : (n839 ? 1'b0 : n53)) : (n1266 ? !n53 : 1'b0));
assign n1835 = /* LUT    9 21  1 */ (n861 ? n1015 : n971);
assign n1836 = /* LUT   12 22  7 */ (n1334 ? (n781 ? n1214 : !n1214) : (n781 ? !n1214 : n1214));
assign n1837 = /* LUT   13 25  0 */ (n1406 ? (n766 ? n1352 : !n1352) : (n766 ? !n1352 : n1352));
assign n1838 = /* LUT    6 24  0 */ (n604 ? (n782 ? 1'b1 : !n253) : (n782 ? n253 : 1'b0));
assign n1839 = /* LUT    4 20  7 */ (n643 ? (n106 ? 1'b0 : (n250 ? 1'b1 : n157)) : (n106 ? 1'b0 : (n250 ? !n157 : 1'b0)));
assign n1840 = /* LUT    2 23  0 */ (n490 ? (n107 ? n193 : !n193) : (n107 ? !n193 : n193));
assign n581  = /* LUT    3 21  2 */ (n324 ? n580 : n394);
assign n1359 = /* LUT   13 19  4 */ (n866 ? (n918 ? 1'b1 : n1203) : (n918 ? 1'b0 : n1203));
assign n1842 = /* LUT   10 24  2 */ (n1156 ? (n1045 ? n1106 : !n1106) : (n1045 ? !n1106 : n1106));
assign n1843 = /* LUT    4 18  7 */ \inMod[8] ;
assign n931  = /* LUT    7 23  5 */ (n861 ? n930 : n925);
assign n1844 = /* LUT    4 24  7 */ (n491 ? (n678 ? 1'b1 : !n253) : (n678 ? n253 : 1'b0));
assign n1845 = /* LUT    1 20  4 */ (n330 ? (n214 ? n326 : !n326) : (n214 ? !n326 : n326));
assign n1846 = /* LUT   14 18  3 */ (n1347 ? (n881 ? 1'b1 : !n290) : (n881 ? n290 : 1'b0));
assign n1847 = /* LUT   14 20  3 */ (n1412 ? (n142 ? (n49 ? n251 : 1'b1) : 1'b1) : (n142 ? (n49 ? n251 : 1'b0) : 1'b0));
assign n1074 = /* LUT    9 26  5 */ (n861 ? n1073 : n990);
assign n1848 = /* LUT   10 19  0 */ (n843 ? (n463 ? 1'b1 : (n50 ? !n49 : 1'b1)) : (n463 ? (n50 ? n49 : 1'b0) : 1'b0));
assign n1849 = /* LUT    5 25  0 */ !n788;
assign n1850 = /* LUT    2 24  2 */ (n509 ? (n232 ? n212 : !n212) : (n232 ? !n212 : n212));
assign n1851 = /* LUT   13 22  6 */ (n1385 ? (n999 ? n758 : !n758) : (n999 ? !n758 : n758));
assign n1852 = /* LUT   16 23  4 */ (n49 ? (n142 ? n665 : n969) : n969);
assign n1219 = /* LUT   11 20  3 */ (n1119 ? (n918 ? 1'b1 : n1217) : (n918 ? 1'b0 : n1217));
assign n1854 = /* LUT    4 29  3 */ (n722 ? (n718 ? 1'b1 : !n253) : (n718 ? n253 : 1'b0));
assign n1855 = /* LUT    5 18  6 */ (n641 ? (reset ? 1'b1 : (n555 ? 1'b1 : !n253)) : (reset ? 1'b0 : (n555 ? n253 : 1'b0)));
assign n1856 = /* LUT    1 23  2 */ (n383 ? (n204 ? n209 : !n209) : (n204 ? !n209 : n209));
assign n1857 = /* LUT    2 22  7 */ (n489 ? (n104 ? n173 : !n173) : (n104 ? !n173 : n173));
assign n1858 = /* LUT   19 20  4 */ (n1474 ? 1'b1 : (n1508 ? 1'b1 : (n1484 ? 1'b1 : n1495)));
assign n1859 = /* LUT    1 26  5 */ !n432;
assign n1860 = /* LUT    5 28  6 */ (n817 ? (n784 ? n235 : !n235) : (n784 ? !n235 : n235));
assign n1861 = /* LUT    6 29  5 */ (n605 ? (n711 ? 1'b1 : n507) : (n711 ? !n507 : 1'b0));
assign n1126 = /* LUT   10 20  2 */ (n1022 ? (n1057 ? 1'b1 : !n811) : (n1057 ? n811 : 1'b0));
assign n1863 = /* LUT   11 22  6 */ (n1245 ? (n785 ? n593 : !n593) : (n785 ? !n593 : n593));
assign n1864 = /* LUT    6 23  1 */ (n772 ? n524 : 1'b0);
assign n1865 = /* LUT    7 18  0 */ (n844 ? (reset ? 1'b1 : (n290 ? n98 : 1'b1)) : (reset ? 1'b0 : (n290 ? n98 : 1'b0)));
assign n1866 = /* LUT    9 27  2 */ (\indata[18]  ? (n1082 ? (\inExp[0]  ? 1'b1 : !ready) : (\inExp[0]  ? ready : 1'b0)) : (n1082 ? !ready : 1'b0));
assign n1867 = /* LUT   11 19  7 */ (n1110 ? n732 : 1'b0);
assign n1868 = /* LUT   17 21  7 */ (ready ? (n1456 ? (ds ? \inExp[29]  : 1'b1) : (ds ? \inExp[29]  : 1'b0)) : n1456);
assign n1869 = /* LUT    3 17  7 */ (ready ? (n286 ? !ds : 1'b0) : (n286 ? n77 : 1'b0));
assign n1870 = /* LUT    1 18  0 */ (n285 ? (n166 ? n292 : !n292) : (n166 ? !n292 : n292));
assign n1871 = /* LUT   12 16  4 */ (n918 ? n1285 : n1198);
assign n1872 = /* LUT   13 23  1 */ (n1390 ? (n1121 ? n1266 : !n1266) : (n1121 ? !n1266 : n1266));
assign n1873 = /* LUT    3 23  7 */ (n595 ? n524 : 1'b0);
assign n1874 = /* LUT    2 21  3 */ (n474 ? (n272 ? n151 : !n151) : (n272 ? !n151 : n151));
assign n1875 = /* LUT   15 23  4 */ (n1435 ? (n884 ? 1'b1 : (n142 ? !n49 : 1'b1)) : (n884 ? (n142 ? n49 : 1'b0) : 1'b0));
assign n1876 = /* LUT    6 16  5 */ (n50 ? (n645 ? (n49 ? 1'b1 : n444) : (n49 ? 1'b0 : n444)) : n444);
assign n1877 = /* LUT    4 28  4 */ (n534 ? (n619 ? 1'b1 : n507) : (n619 ? !n507 : 1'b0));
assign n1878 = /* LUT    7 27  6 */ !n532;
assign n1879 = /* LUT   11 24  3 */ (n1269 ? (n894 ? n1171 : !n1171) : (n894 ? !n1171 : n1171));
assign n1880 = /* LUT   12 18  5 */ (n290 ? (n1195 ? (n53 ? n662 : 1'b1) : (n53 ? n662 : 1'b0)) : (n1195 ? !n53 : 1'b0));
assign n1881 = /* LUT    4 26  0 */ (n611 ? (n437 ? 1'b1 : n507) : (n437 ? !n507 : 1'b0));
assign n1882 = /* LUT    9 22  0 */ (n53 ? (n23 ? !n839 : 1'b0) : n967);
assign n1047 = /* LUT    9 24  4 */ (n1027 ? (n1043 ? 1'b1 : !n811) : (n1043 ? n811 : 1'b0));
assign n1100 = /* LUT   10 17  3 */ (n861 ? n1099 : n1097);
assign n1884 = /* LUT   12 21  6 */ (n1324 ? (n892 ? n1135 : !n1135) : (n892 ? !n1135 : n1135));
assign n1885 = /* LUT   18 19  6 */ (n910 ? (n50 ? n142 : 1'b0) : 1'b0);
assign n1886 = /* LUT   13 20  5 */ (n2 ? (n1307 ? !n839 : (n53 ? !n839 : 1'b0)) : (n1307 ? (n53 ? 1'b0 : !n839) : 1'b0));
assign n1887 = /* LUT   10 27  3 */ (n40 ? (n53 ? !n839 : n1060) : (n53 ? 1'b0 : n1060));
assign n1888 = /* LUT    3 24  3 */ (n302 ? (n222 ? !n106 : (n157 ? !n106 : 1'b0)) : (n222 ? (n157 ? 1'b0 : !n106) : 1'b0));
assign n1889 = /* LUT    4 17  6 */ (n49 ? (n50 ? n558 : n542) : n542);
assign n1890 = /* LUT    7 30  0 */ \inMod[22] ;
assign n1891 = /* LUT    1 19  7 */ (n314 ? (n199 ? n233 : !n233) : (n199 ? !n233 : n233));
assign n1892 = /* LUT    5 16  5 */ (n49 ? (n304 ? (n50 ? 1'b1 : n544) : (n50 ? 1'b0 : n544)) : n544);
assign n1893 = /* LUT    1 21  7 */ (n92 ? (n133 ? n197 : 1'b1) : (n133 ? n197 : 1'b0));
assign n1894 = /* LUT   19 22  7 */ (n1501 ? (\inExp[1]  ? 1'b1 : (ds ? !ready : 1'b1)) : (\inExp[1]  ? (ds ? ready : 1'b0) : 1'b0));
assign n1895 = /* LUT   13 18  4 */ (n290 ? n1276 : n1350);
assign n1896 = /* LUT   10 25  6 */ (n1168 ? (n1067 ? n892 : !n892) : (n1067 ? !n892 : n892));
assign n1897 = /* LUT    1 24  4 */ (n405 ? (n356 ? n400 : !n400) : (n356 ? !n400 : n400));
assign n1898 = /* LUT    5 26  1 */ (n793 ? (n277 ? n439 : !n439) : (n277 ? !n439 : n439));
assign n1899 = /* LUT   10 18  7 */ (n883 ? (n1113 ? 1'b1 : n290) : (n1113 ? !n290 : 1'b0));
assign n1900 = /* LUT   14 23  2 */ (n290 ? n1011 : n1437);
assign n1901 = /* LUT   19 19  6 */ (n1486 ? (\inExp[27]  ? 1'b1 : (ds ? !ready : 1'b1)) : (\inExp[27]  ? (ds ? ready : 1'b0) : 1'b0));
assign n1902 = /* LUT    6 21  0 */ (n77 ? (n757 ? (ds ? !ready : 1'b1) : 1'b0) : (n757 ? (ds ? 1'b0 : ready) : 1'b0));
assign n1903 = /* LUT    2 27  3 */ (n536 ? n524 : 1'b0);
assign n1904 = /* LUT    4 22  0 */ (reset ? n584 : (n253 ? n101 : n584));
assign n1905 = /* LUT   11 21  4 */ (n1233 ? (n854 ? n1043 : !n1043) : (n854 ? !n1043 : n1043));
assign n1906 = /* LUT   12 20  1 */ (n1311 ? (n577 ? n1192 : !n1192) : (n577 ? !n1192 : n1192));
assign n1907 = /* LUT    5 19  1 */ (n324 ? n746 : n186);
assign n1908 = /* LUT    6 26  6 */ (n588 ? (n253 ? (reset ? n790 : 1'b1) : n790) : (n253 ? (reset ? n790 : 1'b0) : n790));
assign n1909 = /* LUT    2 25  6 */ (n414 ? (reset ? 1'b1 : (n253 ? n238 : 1'b1)) : (reset ? 1'b0 : (n253 ? n238 : 1'b0)));
assign n1910 = /* LUT   19 21  3 */ (n1499 ? 1'b1 : (n1502 ? 1'b1 : (n1501 ? 1'b1 : n1500)));
assign n1911 = /* LUT    5 29  5 */ (n826 ? (n322 ? n257 : !n257) : (n322 ? !n257 : n257));
assign n1912 = /* LUT    3 25  4 */ (n375 ? (n608 ? 1'b1 : !n324) : (n608 ? n324 : 1'b0));
assign n1913 = /* LUT    2 19  6 */ (ready ? (n461 ? !ds : 1'b0) : (n461 ? n77 : 1'b0));
assign n1914 = /* LUT    6 28  6 */ (n612 ? (n694 ? 1'b1 : n507) : (n694 ? !n507 : 1'b0));
assign n1915 = /* LUT   11 23  5 */ (n1259 ? (n1070 ? n849 : !n849) : (n1070 ? !n849 : n849));
assign n1916 = /* LUT   10 23  3 */ (n1146 ? (n1031 ? n854 : !n854) : (n1031 ? !n854 : n854));
assign n1917 = /* LUT    6 22  6 */ (reset ? n765 : (n765 ? (n600 ? 1'b1 : !n290) : (n600 ? n290 : 1'b0)));
assign n1918 = /* LUT   11 26  6 */ (n1053 ? (n1068 ? 1'b1 : !n811) : (n1068 ? n811 : 1'b0));
assign n1919 = /* LUT    7 19  3 */ !n864;
assign n1920 = /* LUT   12 25  1 */ (ready ? \indata[20]  : n601);
assign n1921 = /* LUT    9 20  3 */ (n687 ? n524 : 1'b0);
assign n769  = /* LUT    5 22  1 */ (n704 ? (n507 ? n687 : 1'b1) : (n507 ? n687 : 1'b0));
assign n1923 = /* LUT   12 23  5 */ (n33 ? (n839 ? (n53 ? 1'b0 : n1252) : (n53 ? 1'b1 : n1252)) : (n53 ? 1'b0 : n1252));
assign n1924 = /* LUT   13 24  0 */ (n1397 ? (n1336 ? n1020 : !n1020) : (n1336 ? !n1020 : n1020));
assign n1925 = /* LUT    3 20  6 */ (n77 ? (n573 ? (ready ? !ds : 1'b1) : 1'b0) : (n573 ? (ready ? !ds : 1'b0) : 1'b0));
assign n1926 = /* LUT    6 25  0 */ (n821 ? (n253 ? n526 : 1'b1) : (n253 ? n526 : 1'b0));
assign n1927 = /* LUT   15 20  5 */ (n1424 ? (n587 ? 1'b1 : (n142 ? !n49 : 1'b1)) : (n587 ? (n142 ? n49 : 1'b0) : 1'b0));
assign n862  = /* LUT    6 19  4 */ (n859 ? (n745 ? 1'b1 : !n811) : (n745 ? n811 : 1'b0));
assign n1929 = /* LUT    7 24  7 */ (n301 ? (ready ? \indata[15]  : 1'b1) : (ready ? \indata[15]  : 1'b0));
assign n1930 = /* LUT    4 19  5 */ (n644 ? (n157 ? !n106 : (n209 ? !n106 : 1'b0)) : (n157 ? 1'b0 : (n209 ? !n106 : 1'b0)));
assign n1931 = /* LUT   12 17  4 */ (n1190 ? (n290 ? n963 : 1'b1) : (n290 ? n963 : 1'b0));
assign n1932 = /* LUT    7 22  7 */ (n757 ? (n183 ? !n106 : (n106 ? 1'b0 : n157)) : (n183 ? (n106 ? 1'b0 : !n157) : 1'b0));
assign n1933 = /* LUT    9 23  7 */ (n146 ? (ready ? \indata[13]  : 1'b1) : (ready ? \indata[13]  : 1'b0));
assign n689  = /* LUT    4 25  1 */ (n324 ? n688 : n373);
assign n1934 = /* LUT   14 21  1 */ (n1122 ? n732 : 1'b0);
assign n1935 = /* LUT    5 24  0 */ (n783 ? (n341 ? 1'b1 : (n49 ? !n142 : 1'b1)) : (n341 ? (n49 ? n142 : 1'b0) : 1'b0));
assign n1092 = /* LUT   10 16  0 */ (n994 ? (n1040 ? 1'b1 : !n811) : (n1040 ? n811 : 1'b0));
assign n561  = /* LUT    3 19  0 */ (n59 ? (n150 ? 1'b1 : !n133) : (n150 ? n133 : 1'b0));
assign n1938 = /* LUT   10 26  4 */ (n1179 ? (n1014 ? n684 : !n684) : (n1014 ? !n684 : n684));
assign n1939 = /* LUT   11 17  1 */ \inMod[0] ;
assign n1940 = /* LUT   13 21  6 */ (n1374 ? (n959 ? n1284 : !n1284) : (n959 ? !n1284 : n1284));
assign n1941 = /* LUT    4 16  1 */ (n551 ? (n470 ? 1'b1 : (n50 ? !n49 : 1'b1)) : (n470 ? (n50 ? n49 : 1'b0) : 1'b0));
assign n777  = /* LUT    5 23  6 */ (n672 ? (n507 ? 1'b1 : n504) : (n507 ? 1'b0 : n504));
assign n1943 = /* LUT    4 30  5 */ \inMod[2] ;
assign n1944 = /* LUT    5 17  6 */ (n253 ? (reset ? n636 : n642) : n636);
assign n1945 = /* LUT    1 22  6 */ (n369 ? (n361 ? n359 : !n359) : (n361 ? !n359 : n359));
assign n1946 = /* LUT   10 24  5 */ (n1159 ? (n972 ? n593 : !n593) : (n972 ? !n593 : n593));
assign n1947 = /* LUT   13 19  3 */ (n1285 ? n732 : 1'b0);
assign n1948 = /* LUT    1 25  7 */ (n428 ? (n418 ? n244 : !n244) : (n418 ? !n244 : n244));
assign n1949 = /* LUT   15 21  2 */ (n1421 ? (n526 ? 1'b1 : (n142 ? !n49 : 1'b1)) : (n526 ? (n142 ? n49 : 1'b0) : 1'b0));
assign n1950 = /* LUT   10 21  6 */ (n13 ? (\indata[24]  ? (\inExp[0]  ? 1'b1 : !ready) : !ready) : (\indata[24]  ? (\inExp[0]  ? ready : 1'b0) : 1'b0));
assign n1951 = /* LUT    6 18  3 */ (reset ? n739 : (n739 ? (n253 ? n837 : 1'b1) : (n253 ? n837 : 1'b0)));
assign n1952 = /* LUT    5 27  6 */ (n806 ? (n104 ? n687 : !n687) : (n104 ? !n687 : n687));
assign n1953 = /* LUT   14 22  5 */ (n1136 ? n732 : 1'b0);
assign n1954 = /* LUT    2 26  4 */ (n432 ? (n438 ? 1'b1 : (reset ? 1'b1 : !n253)) : (n438 ? (reset ? 1'b0 : n253) : 1'b0));
assign n1955 = /* LUT    6 20  3 */ (n644 ? (\indata[10]  ? 1'b1 : !ready) : (\indata[10]  ? ready : 1'b0));
assign n1956 = /* LUT    4 21  1 */ (n462 ? (n126 ? !n106 : (n157 ? !n106 : 1'b0)) : (n126 ? (n157 ? 1'b0 : !n106) : 1'b0));
assign n1957 = /* LUT   11 18  5 */ !n1105;
assign n752  = /* LUT    5 20  0 */ (n93 ? (n198 ? 1'b1 : !n133) : (n198 ? n133 : 1'b0));
assign n1959 = /* LUT    1 17  0 */ (n276 ? (n83 ? n148 : !n148) : (n83 ? !n148 : n148));
assign n1960 = /* LUT    2 24  5 */ (n512 ? (n326 ? n161 : !n161) : (n326 ? !n161 : n161));
assign n1961 = /* LUT   14 19  5 */ (n1310 ? n732 : 1'b0);
assign n1962 = /* LUT    5 30  4 */ (n710 ? (n507 ? n696 : 1'b1) : (n507 ? n696 : 1'b0));
assign n1963 = /* LUT    3 22  5 */ !n481;
assign n1964 = /* LUT    2 18  1 */ (n307 ? (n450 ? 1'b1 : !n324) : (n450 ? n324 : 1'b0));
assign n1965 = /* LUT   11 20  4 */ (n290 ? n1205 : n1219);
assign n1966 = /* LUT   15 22  4 */ (n1412 ? 1'b1 : (n1433 ? 1'b1 : (n1422 ? 1'b1 : n1424)));
assign n1967 = /* LUT    6 17  7 */ (n53 ? (n655 ? n290 : 1'b0) : n736);
assign n1968 = /* LUT    7 26  2 */ (reset ? n898 : (n898 ? (n290 ? n252 : 1'b1) : (n290 ? n252 : 1'b0)));
assign n622  = /* LUT    3 28  1 */ (n621 ? (n620 ? 1'b1 : n507) : (n620 ? !n507 : 1'b0));
assign n1970 = /* LUT    9 19  4 */ (n953 ? n732 : 1'b0);
assign n1281 = /* LUT   11 27  5 */ (n1063 ? (n1077 ? 1'b1 : !n811) : (n1077 ? n811 : 1'b0));
assign n1972 = /* LUT   12 19  7 */ (n1302 ? (n932 ? n1293 : !n1293) : (n932 ? !n1293 : n1293));
assign n1015 = /* LUT    9 21  0 */ (n1012 ? (n1014 ? 1'b1 : !n811) : (n1014 ? n811 : 1'b0));
assign n1974 = /* LUT   12 22  6 */ (n1333 ? (n737 ? n1212 : !n1212) : (n737 ? !n1212 : n1212));
assign n580  = /* LUT    3 21  1 */ (n118 ? (n133 ? n161 : 1'b1) : (n133 ? n161 : 1'b0));
assign n1976 = /* LUT    4 20  6 */ !n566;
assign n1977 = /* LUT    2 23  1 */ (n495 ? (n234 ? n182 : !n182) : (n234 ? !n182 : n182));
assign n1349 = /* LUT   13 18  1 */ (n917 ? (n918 ? 1'b1 : n1221) : (n918 ? 1'b0 : n1221));
assign n1979 = /* LUT    4 18  6 */ \inMod[7] ;
assign n1980 = /* LUT    7 25  0 */ !n897;
assign n1981 = /* LUT    4 24  6 */ (n679 ? (n253 ? n578 : 1'b1) : (n253 ? n578 : 1'b0));
assign n1982 = /* LUT   14 18  2 */ (n1409 ? (n960 ? 1'b1 : !n290) : (n960 ? n290 : 1'b0));
assign n1983 = /* LUT    1 20  5 */ (n331 ? (n161 ? n322 : !n322) : (n161 ? !n322 : n322));
assign n930  = /* LUT    7 23  4 */ (n887 ? (n433 ? 1'b1 : !n811) : (n433 ? n811 : 1'b0));
assign n1985 = /* LUT   14 20  2 */ (n1416 ? (n142 ? (n670 ? 1'b1 : !n49) : 1'b1) : (n142 ? (n670 ? n49 : 1'b0) : 1'b0));
assign n1986 = /* LUT    9 26  6 */ (\indata[23]  ? (n1074 ? (\inExp[0]  ? 1'b1 : !ready) : (\inExp[0]  ? ready : 1'b0)) : (n1074 ? !ready : 1'b0));
assign n1987 = /* LUT   10 19  1 */ (n914 ? (n465 ? 1'b1 : (n49 ? !n50 : 1'b1)) : (n465 ? (n49 ? n50 : 1'b0) : 1'b0));
assign n1988 = /* LUT    5 25  3 */ (n507 ? n597 : n697);
assign n1989 = /* LUT   13 22  7 */ (n1386 ? (n949 ? n1283 : !n1283) : (n949 ? !n1283 : n1283));
assign n1990 = /* LUT   16 23  5 */ (n1446 ? (n606 ? 1'b1 : (n142 ? !n49 : 1'b1)) : (n606 ? (n142 ? n49 : 1'b0) : 1'b0));
assign n1991 = /* LUT    4 23  0 */ (n589 ? (n341 ? (n157 ? n253 : 1'b1) : !n157) : (n341 ? (n157 ? n253 : 1'b0) : 1'b0));
assign n1992 = /* LUT    4 29  4 */ (n623 ? n524 : 1'b0);
assign n1993 = /* LUT    5 18  7 */ !n638;
assign n1994 = /* LUT    1 23  1 */ (n382 ? (n207 ? n127 : !n127) : (n207 ? !n127 : n127));
assign n1995 = /* LUT    2 22  6 */ (n488 ? (n97 ? n172 : !n172) : (n97 ? !n172 : n172));
assign n1996 = /* LUT   13 20  2 */ (n54 ? (n1304 ? !n839 : (n839 ? 1'b0 : n53)) : (n1304 ? (n839 ? 1'b0 : !n53) : 1'b0));
assign n1997 = /* LUT    1 26  6 */ !n431;
assign n1998 = /* LUT    5 28  7 */ (n818 ? (n233 ? n621 : !n621) : (n233 ? !n621 : n621));
assign n1999 = /* LUT   10 20  5 */ (n287 ? (\indata[7]  ? 1'b1 : !ready) : (\indata[7]  ? ready : 1'b0));
assign n2000 = /* LUT   11 22  7 */ (n1246 ? (n763 ? n786 : !n786) : (n763 ? !n786 : n786));
assign n2001 = /* LUT   16 20  1 */ (n524 ? 1'b1 : (n1416 ? 1'b1 : (n1413 ? 1'b1 : n1417)));
assign n2002 = /* LUT    7 18  1 */ (n637 ? 1'b1 : (n52 ? 1'b1 : (n633 ? 1'b1 : n916)));
assign n1082 = /* LUT    9 27  1 */ (n978 ? (n1081 ? 1'b1 : !n861) : (n1081 ? n861 : 1'b0));
assign n2003 = /* LUT   11 19  6 */ (n290 ? n965 : n1209);
assign n2004 = /* LUT   17 21  6 */ (n1455 ? (ds ? (\inExp[30]  ? 1'b1 : !ready) : 1'b1) : (ds ? (\inExp[30]  ? ready : 1'b0) : 1'b0));
assign n760  = /* LUT    5 21  3 */ (n575 ? (n324 ? 1'b1 : n376) : (n324 ? 1'b0 : n376));
assign n2005 = /* LUT    3 17  6 */ (n287 ? (ds ? (n77 ? !ready : 1'b0) : (n77 ? 1'b1 : ready)) : 1'b0);
assign n2006 = /* LUT   19 19  1 */ (ready ? (\inExp[22]  ? (n1461 ? 1'b1 : ds) : (n1461 ? !ds : 1'b0)) : n1461);
assign n2007 = /* LUT    1 18  1 */ (n293 ? (n167 ? n178 : !n178) : (n167 ? !n178 : n178));
assign n2008 = /* LUT   13 23  0 */ (n1387 ? (n1251 ? n1263 : !n1263) : (n1251 ? !n1263 : n1263));
assign n2012 = /* LUT   11 21  3 */ (n1232 ? (n1031 ? n853 : !n853) : (n1031 ? !n853 : n853));
assign n2013 = /* LUT   15 23  7 */ (n396 ? (n521 ? 1'b1 : (n49 ? !n142 : 1'b1)) : (n521 ? (n49 ? n142 : 1'b0) : 1'b0));
assign n2014 = /* LUT    6 16  4 */ (n631 ? (n50 ? (n239 ? 1'b1 : !n49) : 1'b1) : (n50 ? (n239 ? n49 : 1'b0) : 1'b0));
assign n2015 = /* LUT    4 28  3 */ (n253 ? (n265 ? (reset ? 1'b1 : n618) : (reset ? 1'b0 : n618)) : n265);
assign n2016 = /* LUT    7 27  1 */ (reset ? n903 : (n253 ? n907 : n903));
assign n2017 = /* LUT   11 24  4 */ (n1270 ? (n905 ? n1014 : !n1014) : (n905 ? !n1014 : n1014));
assign n2018 = /* LUT   12 18  4 */ (n918 ? n1195 : n1291);
assign n2019 = /* LUT    4 26  3 */ (n253 ? n175 : n610);
assign n1048 = /* LUT    9 24  5 */ (n941 ? (n1047 ? 1'b1 : !n861) : (n1047 ? n861 : 1'b0));
assign n1098 = /* LUT   10 17  0 */ (n1062 ? (n893 ? 1'b1 : !n811) : (n893 ? n811 : 1'b0));
assign n2021 = /* LUT   12 21  7 */ (n1325 ? (n901 ? n1136 : !n1136) : (n901 ? !n1136 : n1136));
assign n2022 = /* LUT    3 18  0 */ (n287 ? (n157 ? !n106 : (n323 ? !n106 : 1'b0)) : (n157 ? 1'b0 : (n323 ? !n106 : 1'b0)));
assign n2023 = /* LUT    3 24  4 */ (n303 ? (n157 ? !n106 : (n399 ? !n106 : 1'b0)) : (n157 ? 1'b0 : (n399 ? !n106 : 1'b0)));
assign n2024 = /* LUT    4 17  7 */ (n549 ? (n454 ? 1'b1 : (n50 ? !n49 : 1'b1)) : (n454 ? (n50 ? n49 : 1'b0) : 1'b0));
assign n2025 = /* LUT    7 30  1 */ \inMod[23] ;
assign n2026 = /* LUT    1 19  6 */ (n313 ? (n198 ? n235 : !n235) : (n198 ? !n235 : n235));
assign n2027 = /* LUT   12 23  2 */ (n1118 ? n732 : 1'b0);
assign n2028 = /* LUT    7 20  5 */ (n162 ? (n865 ? !n839 : (n839 ? 1'b0 : n53)) : (n865 ? (n839 ? 1'b0 : !n53) : 1'b0));
assign n2029 = /* LUT    9 17  5 */ (n2 ? (\indata[5]  ? (ready ? \inExp[0]  : 1'b1) : !ready) : (\indata[5]  ? (ready ? \inExp[0]  : 1'b0) : 1'b0));
assign n2030 = /* LUT    1 21  6 */ (n120 ? (n133 ? n215 : 1'b1) : (n133 ? n215 : 1'b0));
assign n2031 = /* LUT   19 22  4 */ (n1462 ? (\inExp[4]  ? 1'b1 : (ready ? !ds : 1'b1)) : (\inExp[4]  ? (ready ? ds : 1'b0) : 1'b0));
assign n2032 = /* LUT   13 18  5 */ (n1288 ? n732 : 1'b0);
assign n2033 = /* LUT   10 25  7 */ (n1169 ? (n1069 ? n901 : !n901) : (n1069 ? !n901 : n901));
assign n2034 = /* LUT    1 24  5 */ (n406 ? (n218 ? n223 : !n223) : (n218 ? !n223 : n223));
assign n2035 = /* LUT    5 26  2 */ (n794 ? (n272 ? n676 : !n676) : (n272 ? !n676 : n676));
assign n2036 = /* LUT   14 23  3 */ (n1388 ? (n993 ? 1'b1 : !n290) : (n993 ? n290 : 1'b0));
assign n1113 = /* LUT   10 18  6 */ (n918 ? n998 : n958);
assign n2038 = /* LUT   18 20  3 */ (n1485 ? (\inExp[21]  ? 1'b1 : (ready ? !ds : 1'b1)) : (\inExp[21]  ? (ready ? ds : 1'b0) : 1'b0));
assign n874  = /* LUT    6 21  1 */ (n61 ? (n152 ? 1'b1 : !n133) : (n152 ? n133 : 1'b0));
assign n2040 = /* LUT   16 22  6 */ (n1444 ? 1'b1 : (n1459 ? 1'b1 : (n1429 ? 1'b1 : n1445)));
assign n2041 = /* LUT    4 22  3 */ !n584;
assign n2042 = /* LUT   14 21  6 */ (n290 ? n975 : n1427);
assign n2043 = /* LUT   12 20  0 */ (n1303 ? (n850 ? n1285 : !n1285) : (n850 ? !n1285 : n1285));
assign n746  = /* LUT    5 19  0 */ (n119 ? (n133 ? n208 : 1'b1) : (n133 ? n208 : 1'b0));
assign n2045 = /* LUT    6 26  5 */ !n790;
assign n2046 = /* LUT    2 25  7 */ !n413;
assign n2047 = /* LUT   10 26  3 */ (n1178 ? (n894 ? n905 : !n905) : (n894 ? !n905 : n905));
assign n2048 = /* LUT   13 21  1 */ (n1369 ? (n1366 ? n1306 : !n1306) : (n1366 ? !n1306 : n1306));
assign n2049 = /* LUT    5 29  4 */ (n825 ? (n326 ? n624 : !n624) : (n326 ? !n624 : n624));
assign n608  = /* LUT    3 25  3 */ (n94 ? (n199 ? 1'b1 : !n133) : (n199 ? n133 : 1'b0));
assign n2051 = /* LUT    2 19  7 */ (ready ? (n302 ? !ds : 1'b0) : (n302 ? n77 : 1'b0));
assign n2052 = /* LUT   10 23  4 */ (n1147 ? (n1043 ? n669 : !n669) : (n1043 ? !n669 : n669));
assign n2053 = /* LUT   11 23  4 */ (n1258 ? (n1068 ? n852 : !n852) : (n1068 ? !n852 : n852));
assign n2054 = /* LUT    6 22  5 */ (n764 ? (reset ? 1'b1 : (n290 ? n96 : 1'b1)) : (reset ? 1'b0 : (n290 ? n96 : 1'b0)));
assign n2055 = /* LUT   11 26  7 */ (n1054 ? (n1070 ? 1'b1 : !n811) : (n1070 ? n811 : 1'b0));
assign n2056 = /* LUT    7 19  2 */ !n740;
assign n2057 = /* LUT    9 20  0 */ (n321 ? (ready ? \indata[1]  : 1'b1) : (ready ? \indata[1]  : 1'b0));
assign n2058 = /* LUT    5 22  2 */ (n253 ? n768 : n769);
assign n2059 = /* LUT   14 24  0 */ (n85 ? (n53 ? !n839 : (n1379 ? !n839 : 1'b0)) : (n53 ? 1'b0 : (n1379 ? !n839 : 1'b0)));
assign n2060 = /* LUT    2 26  3 */ (n431 ? (reset ? 1'b1 : (n253 ? n252 : 1'b1)) : (reset ? 1'b0 : (n253 ? n252 : 1'b0)));
assign n2061 = /* LUT   13 24  1 */ (n1399 ? (n1389 ? n1102 : !n1102) : (n1389 ? !n1102 : n1102));
assign n2062 = /* LUT    3 20  7 */ (n146 ? (ready ? !ds : n77) : 1'b0);
assign n2063 = /* LUT    2 20  3 */ (n72 ? (n169 ? 1'b1 : !n133) : (n169 ? n133 : 1'b0));
assign n2064 = /* LUT   11 18  2 */ (n7 ? (n1103 ? (n839 ? !n53 : 1'b1) : (n839 ? 1'b0 : n53)) : (n1103 ? !n53 : 1'b0));
assign n2065 = /* LUT   15 20  6 */ (n49 ? (n142 ? n718 : n1440) : n1440);
assign n2066 = /* LUT    3 26  7 */ (n516 ? (\indata[24]  ? 1'b1 : !ready) : (\indata[24]  ? ready : 1'b0));
assign n863  = /* LUT    6 19  5 */ (n861 ? n862 : n860);
assign n2067 = /* LUT    4 19  2 */ (n559 ? (reset ? 1'b1 : (n99 ? 1'b1 : !n253)) : (reset ? 1'b0 : (n99 ? n253 : 1'b0)));
assign n936  = /* LUT    7 24  0 */ (n935 ? (n785 ? 1'b1 : !n811) : (n785 ? n811 : 1'b0));
assign n2069 = /* LUT   12 17  5 */ (n1197 ? (n992 ? 1'b1 : !n290) : (n992 ? n290 : 1'b0));
assign n2070 = /* LUT    4 25  2 */ (ds ? (n689 ? (ready ? 1'b0 : n77) : 1'b0) : (n689 ? (ready ? 1'b1 : n77) : 1'b0));
assign n2071 = /* LUT    9 23  6 */ (\indata[13]  ? (n1038 ? (\inExp[0]  ? 1'b1 : !ready) : (\inExp[0]  ? ready : 1'b0)) : (n1038 ? !ready : 1'b0));
assign n2072 = /* LUT   10 22  3 */ (n13 ? (n1020 ? (n53 ? !n839 : 1'b1) : (n53 ? !n839 : 1'b0)) : (n1020 ? !n53 : 1'b0));
assign n923  = /* LUT    7 22  4 */ (n141 ? (n142 ? !n49 : 1'b0) : (n142 ? !n49 : !n443));
assign n2073 = /* LUT    5 24  1 */ (n524 ? n589 : 1'b0);
assign n2074 = /* LUT   10 16  3 */ (n757 ? (ready ? \indata[5]  : 1'b1) : (ready ? \indata[5]  : 1'b0));
assign n563  = /* LUT    3 19  3 */ (n133 ? n149 : n58);
assign n2076 = /* LUT   11 17  0 */ !n1189;
assign n2077 = /* LUT    4 16  0 */ (n629 ? (n552 ? 1'b1 : (n49 ? !n50 : 1'b1)) : (n552 ? (n49 ? n50 : 1'b0) : 1'b0));
assign n2078 = /* LUT    5 23  5 */ (n49 ? n142 : 1'b0);
assign n2079 = /* LUT   12 22  1 */ (n1328 ? (n900 ? n1141 : !n1141) : (n900 ? !n1141 : n1141));
assign n2080 = /* LUT    4 30  4 */ \inMod[19] ;
assign n2081 = /* LUT    5 17  1 */ !n635;
assign n2082 = /* LUT    1 22  7 */ (n370 ? (n189 ? n323 : !n323) : (n189 ? !n323 : n323));
assign n2083 = /* LUT   13 19  2 */ (n1007 ? (n1358 ? 1'b1 : n290) : (n1358 ? !n290 : 1'b0));
assign n2084 = /* LUT   10 24  4 */ (n1158 ? (n1030 ? n1021 : !n1021) : (n1030 ? !n1021 : n1021));
assign n2085 = /* LUT    1 25  6 */ (n427 ? (n246 ? n250 : !n250) : (n246 ? !n250 : n250));
assign n2086 = /* LUT   15 21  1 */ (n1420 ? (n775 ? 1'b1 : (n49 ? !n142 : 1'b1)) : (n775 ? (n49 ? n142 : 1'b0) : 1'b0));
assign n2087 = /* LUT   10 21  7 */ (n658 ? (ready ? \indata[25]  : 1'b1) : (ready ? \indata[25]  : 1'b0));
assign n2088 = /* LUT    6 18  2 */ (n738 ? (reset ? 1'b1 : (n95 ? 1'b1 : !n290)) : (reset ? 1'b0 : (n95 ? n290 : 1'b0)));
assign n2089 = /* LUT    5 27  5 */ (n805 ? (n97 ? n773 : !n773) : (n97 ? !n773 : n773));
assign n2090 = /* LUT   14 22  4 */ (n1154 ? (n290 ? n942 : 1'b1) : (n290 ? n942 : 1'b0));
assign n2091 = /* LUT    6 20  2 */ (ready ? (\indata[10]  ? \inExp[0]  : 1'b0) : n871);
assign n2092 = /* LUT    4 21  2 */ (n579 ? (n227 ? !n106 : (n106 ? 1'b0 : n157)) : (n227 ? (n106 ? 1'b0 : !n157) : 1'b0));
assign n2093 = /* LUT   14 20  5 */ (n49 ? (n674 ? (n142 ? 1'b1 : n1361) : (n142 ? 1'b0 : n1361)) : n1361);
assign n1342 = /* LUT   12 27  1 */ (n1172 ? (n861 ? 1'b1 : n1137) : (n861 ? 1'b0 : n1137));
assign n2094 = /* LUT    5 20  1 */ (n324 ? n752 : n352);
assign n2095 = /* LUT    1 17  3 */ (n280 ? (n151 ? n79 : !n79) : (n151 ? !n79 : n79));
assign n2096 = /* LUT    2 24  4 */ (n511 ? (n145 ? n214 : !n214) : (n145 ? !n214 : n214));
assign n2097 = /* LUT   13 22  0 */ (n1376 ? (n1292 ? n1304 : !n1304) : (n1292 ? !n1304 : n1304));
assign n2098 = /* LUT   14 19  6 */ (n1001 ? n732 : 1'b0);
assign n2099 = /* LUT    5 30  5 */ (n623 ? (n716 ? 1'b1 : n507) : (n716 ? !n507 : 1'b0));
assign n2100 = /* LUT    3 22  2 */ (n180 ? (n290 ? (reset ? 1'b1 : n588) : 1'b1) : (n290 ? (reset ? 1'b0 : n588) : 1'b0));
assign n450  = /* LUT    2 18  0 */ (n69 ? (n166 ? 1'b1 : !n133) : (n166 ? n133 : 1'b0));
assign n2102 = /* LUT   11 20  5 */ (n1120 ? n732 : 1'b0);
assign n2103 = /* LUT   15 22  5 */ (n1418 ? 1'b1 : (n396 ? 1'b1 : (n1226 ? 1'b1 : n1421)));
assign n2104 = /* LUT    3 28  2 */ (n253 ? n251 : n622);
assign n2105 = /* LUT    7 26  3 */ (reset ? n899 : (n899 ? (n642 ? 1'b1 : !n290) : (n642 ? n290 : 1'b0)));
assign n2106 = /* LUT    9 19  3 */ (n290 ? n976 : n1004);
assign n2107 = /* LUT   12 19  4 */ (n1299 ? (n669 ? n953 : !n953) : (n669 ? !n953 : n953));
assign n915  = /* LUT    7 16  3 */ (n842 ? 1'b1 : (n914 ? 1'b1 : (n447 ? 1'b1 : n551)));
assign n2109 = /* LUT   12 24  5 */ (n19 ? (n1265 ? (n839 ? !n53 : 1'b1) : (n839 ? 1'b0 : n53)) : (n1265 ? !n53 : 1'b0));
assign n1017 = /* LUT    9 21  3 */ (n861 ? n1016 : n962);
assign n2110 = /* LUT    3 21  0 */ (n466 ? (ds ? (n77 ? !ready : 1'b0) : (n77 ? 1'b1 : ready)) : 1'b0);
assign n2111 = /* LUT    4 20  5 */ (n653 ? (n188 ? (n253 ? !n157 : 1'b1) : (n253 ? 1'b0 : n157)) : (n188 ? !n157 : 1'b0));
assign n2112 = /* LUT    2 23  2 */ (n496 ? (n185 ? n194 : !n194) : (n185 ? !n194 : n194));
assign n2113 = /* LUT    7 18  6 */ (n290 ? (reset ? n848 : n456) : n848);
assign n2114 = /* LUT    6 24  2 */ (n524 ? n696 : 1'b0);
assign n2115 = /* LUT   11 19  1 */ (n1114 ? n732 : 1'b0);
assign n2116 = /* LUT    3 27  4 */ (n532 ? (n290 ? (reset ? 1'b1 : n255) : 1'b1) : (n290 ? (reset ? 1'b0 : n255) : 1'b0));
assign n2117 = /* LUT    4 18  1 */ \inMod[30] ;
assign n2118 = /* LUT   12 16  2 */ (n1189 ? (reset ? 1'b1 : (n594 ? 1'b1 : !n290)) : (reset ? 1'b0 : (n594 ? n290 : 1'b0)));
assign n2119 = /* LUT   13 23  7 */ (n1396 ? (n1378 ? n966 : !n966) : (n1378 ? !n966 : n966));
assign n2120 = /* LUT    7 23  7 */ (n466 ? (ready ? \indata[11]  : 1'b1) : (ready ? \indata[11]  : 1'b0));
assign n2121 = /* LUT    4 24  5 */ (n416 ? (n681 ? 1'b1 : n253) : (n681 ? !n253 : 1'b0));
assign n2122 = /* LUT    1 20  2 */ (n328 ? (n212 ? n160 : !n160) : (n212 ? !n160 : n160));
assign n1409 = /* LUT   14 18  1 */ (n1108 ? (n1213 ? 1'b1 : n918) : (n1213 ? !n918 : 1'b0));
assign n2124 = /* LUT    9 26  7 */ (n434 ? (ready ? \indata[23]  : 1'b1) : (ready ? \indata[23]  : 1'b0));
assign n2125 = /* LUT   10 19  2 */ (n730 ? (n139 ? 1'b1 : (n50 ? !n49 : 1'b1)) : (n139 ? (n50 ? n49 : 1'b0) : 1'b0));
assign n2126 = /* LUT   16 23  2 */ (n1442 ? 1'b1 : (n1435 ? 1'b1 : (n200 ? 1'b1 : n1446)));
assign n2127 = /* LUT    4 23  1 */ (n596 ? n524 : 1'b0);
assign n2128 = /* LUT    7 15  0 */ (n910 ? 1'b0 : (reset ? 1'b0 : (n911 ? !ready : 1'b0)));
assign n2129 = /* LUT    9 24  2 */ (\indata[3]  ? (n1046 ? (\inExp[0]  ? 1'b1 : !ready) : (\inExp[0]  ? ready : 1'b0)) : (n1046 ? !ready : 1'b0));
assign n2130 = /* LUT   12 21  0 */ (n1318 ? (n767 ? n1119 : !n1119) : (n767 ? !n1119 : n1119));
assign n2131 = /* LUT    4 29  5 */ (n624 ? n524 : 1'b0);
assign n2132 = /* LUT    1 23  0 */ (n371 ? (n201 ? n205 : !n205) : (n201 ? !n205 : n205));
assign n2133 = /* LUT    2 22  5 */ (n487 ? (n102 ? n171 : !n171) : (n102 ? !n171 : n171));
assign n2134 = /* LUT   13 20  3 */ (n46 ? (n1305 ? !n839 : (n53 ? !n839 : 1'b0)) : (n1305 ? (n53 ? 1'b0 : !n839) : 1'b0));
assign n2135 = /* LUT    1 26  7 */ (n253 ? (reset ? n236 : n254) : n236);
assign n2136 = /* LUT    5 28  4 */ (n815 ? (n247 ? n605 : !n605) : (n247 ? !n605 : n605));
assign n2137 = /* LUT   10 20  4 */ (ready ? (\indata[8]  ? \inExp[0]  : 1'b0) : n1127);
assign n2138 = /* LUT   11 22  4 */ (n1243 ? (n1030 ? n1095 : !n1095) : (n1030 ? !n1095 : n1095));
assign n886  = /* LUT    6 23  3 */ (n772 ? (n507 ? 1'b1 : n702) : (n507 ? 1'b0 : n702));
assign n2140 = /* LUT    1 24  2 */ (n403 ? (n216 ? n399 : !n399) : (n216 ? !n399 : n399));
assign n2141 = /* LUT   14 23  4 */ (n1141 ? n732 : 1'b0);
assign n1081 = /* LUT    9 27  0 */ (n811 ? n1059 : n1051);
assign n2143 = /* LUT   17 21  1 */ (ready ? (n1452 ? (ds ? \inExp[12]  : 1'b1) : (ds ? \inExp[12]  : 1'b0)) : n1452);
assign n2144 = /* LUT    5 21  2 */ (n391 ? (n759 ? 1'b1 : !n324) : (n759 ? n324 : 1'b0));
assign n2145 = /* LUT    1 18  2 */ (n294 ? (n168 ? n103 : !n103) : (n168 ? !n103 : n103));
assign n2146 = /* LUT   19 19  0 */ (n1486 ? 1'b1 : (n1488 ? 1'b1 : (n1485 ? 1'b1 : n1487)));
assign n876  = /* LUT    6 21  6 */ (n62 ? (n153 ? 1'b1 : !n133) : (n153 ? n133 : 1'b0));
assign n2148 = /* LUT    3 23  1 */ (n324 ? n574 : n410);
assign n2149 = /* LUT    2 21  1 */ (n472 ? (n83 ? n149 : !n149) : (n83 ? !n149 : n149));
assign n2150 = /* LUT   11 21  2 */ (n1231 ? (n745 ? n1094 : !n1094) : (n745 ? !n1094 : n1094));
assign n2151 = /* LUT   12 20  7 */ (n1317 ? (n177 ? n649 : !n649) : (n177 ? !n649 : n649));
assign n2152 = /* LUT   15 23  6 */ (n1364 ? (n768 ? 1'b1 : (n142 ? !n49 : 1'b1)) : (n768 ? (n142 ? n49 : 1'b0) : 1'b0));
assign n2153 = /* LUT    6 16  7 */ (n729 ? 1'b1 : (n548 ? 1'b1 : (n730 ? 1'b1 : n65)));
assign n2154 = /* LUT    7 27  0 */ (n902 ? (reset ? 1'b1 : (n261 ? 1'b1 : !n290)) : (reset ? 1'b0 : (n261 ? n290 : 1'b0)));
assign n2155 = /* LUT   11 24  5 */ (n1271 ? (n684 ? n779 : !n779) : (n684 ? !n779 : n779));
assign n2156 = /* LUT   12 18  7 */ (n1118 ? (n1238 ? 1'b1 : n918) : (n1238 ? !n918 : 1'b0));
assign n2157 = /* LUT    4 26  2 */ (n253 ? n665 : n700);
assign n2158 = /* LUT    9 22  2 */ (n53 ? (n36 ? !n839 : 1'b0) : n966);
assign n2159 = /* LUT   13 15  4 */ (n910 ? (ds ? 1'b0 : ready) : (ds ? (n911 ? !ready : 1'b0) : (n911 ? 1'b1 : ready)));
assign n2160 = /* LUT   10 17  1 */ (n861 ? n1098 : n1096);
assign n2161 = /* LUT   18 19  0 */ (n1471 ? (\inExp[23]  ? 1'b1 : (ready ? !ds : 1'b1)) : (\inExp[23]  ? (ready ? ds : 1'b0) : 1'b0));
assign n2162 = /* LUT    3 18  1 */ !n449;
assign n2163 = /* LUT    7 19  5 */ !n847;
assign n2164 = /* LUT    3 24  5 */ (n516 ? (n106 ? 1'b0 : (n157 ? 1'b1 : n417)) : (n106 ? 1'b0 : (n157 ? 1'b0 : n417)));
assign n2165 = /* LUT    4 17  0 */ (n546 ? 1'b1 : (n542 ? 1'b1 : (n78 ? 1'b1 : n547)));
assign n2166 = /* LUT    7 30  6 */ \inMod[28] ;
assign n2167 = /* LUT    1 19  5 */ (n312 ? (n197 ? n128 : !n128) : (n197 ? !n128 : n128));
assign n2168 = /* LUT   12 23  3 */ (n129 ? (n1250 ? (n53 ? !n839 : 1'b1) : (n53 ? !n839 : 1'b0)) : (n1250 ? !n53 : 1'b0));
assign n2169 = /* LUT   13 24  6 */ (n1404 ? (n1354 ? n1086 : !n1086) : (n1354 ? !n1086 : n1086));
assign n2170 = /* LUT    5 16  3 */ (n447 ? (n50 ? (n49 ? n289 : 1'b1) : 1'b1) : (n50 ? (n49 ? n289 : 1'b0) : 1'b0));
assign n2171 = /* LUT    1 21  1 */ (n345 ? (n231 ? n344 : !n344) : (n231 ? !n344 : n344));
assign n2172 = /* LUT   19 22  5 */ (n1502 ? (\inExp[3]  ? 1'b1 : (ds ? !ready : 1'b1)) : (\inExp[3]  ? (ds ? ready : 1'b0) : 1'b0));
assign n2173 = /* LUT   10 25  4 */ (n1166 ? (n1068 ? n849 : !n849) : (n1068 ? !n849 : n849));
assign n1351 = /* LUT   13 18  6 */ (n1134 ? (n918 ? n1288 : 1'b1) : (n918 ? n1288 : 1'b0));
assign n2175 = /* LUT    5 26  3 */ (n795 ? (n534 ? n79 : !n79) : (n534 ? !n79 : n79));
assign n2176 = /* LUT   10 18  5 */ (n998 ? n732 : 1'b0);
assign n2177 = /* LUT   11 25  2 */ (ready ? ds : 1'b0);
assign n2178 = /* LUT   18 20  2 */ (n1487 ? (\inExp[25]  ? 1'b1 : (ds ? !ready : 1'b1)) : (\inExp[25]  ? (ds ? ready : 1'b0) : 1'b0));
assign n2179 = /* LUT    4 22  2 */ !n586;
assign n2180 = /* LUT   14 21  7 */ (n867 ? n732 : 1'b0);
assign n2181 = /* LUT    5 24  6 */ (n534 ? n524 : 1'b0);
assign n2182 = /* LUT    9 25  1 */ !n891;
assign n2183 = /* LUT    5 19  7 */ (n71 ? (n168 ? 1'b1 : !n133) : (n168 ? n133 : 1'b0));
assign n2184 = /* LUT    2 25  4 */ (n492 ? n524 : 1'b0);
assign n2185 = /* LUT   10 26  2 */ (n1177 ? (n893 ? n1171 : !n1171) : (n893 ? !n1171 : n1171));
assign n2186 = /* LUT   11 17  7 */ \inMod[14] ;
assign n2187 = /* LUT   13 21  0 */ (n1200 ? !n1254 : n1254);
assign n2189 = /* LUT    5 29  7 */ (n828 ? (n291 ? n256 : !n256) : (n291 ? !n256 : n256));
assign n2190 = /* LUT   10 23  5 */ (n1148 ? (n1040 ? n121 : !n121) : (n1040 ? !n121 : n121));
assign n458  = /* LUT    2 19  0 */ (n76 ? (n173 ? 1'b1 : !n133) : (n173 ? n133 : 1'b0));
assign n2192 = /* LUT   11 23  7 */ (n1261 ? (n1069 ? n892 : !n892) : (n1069 ? !n892 : n892));
assign n2193 = /* LUT    6 22  4 */ (n651 ? (n157 ? !n106 : (n249 ? !n106 : 1'b0)) : (n157 ? 1'b0 : (n249 ? !n106 : 1'b0)));
assign n2194 = /* LUT    7 21  1 */ (n861 ? n921 : n919);
assign n2195 = /* LUT    1 25  1 */ (n422 ? (n420 ? n158 : !n158) : (n420 ? !n158 : n158));
assign n1337 = /* LUT   12 25  3 */ (n1175 ? (n861 ? 1'b1 : n1140) : (n861 ? 1'b0 : n1140));
assign n2196 = /* LUT    9 20  1 */ (n866 ? n732 : 1'b0);
assign n770  = /* LUT    5 22  3 */ (n666 ? (n507 ? 1'b1 : n705) : (n507 ? 1'b0 : n705));
assign n872  = /* LUT    6 20  5 */ (n870 ? (n861 ? 1'b1 : n869) : (n861 ? 1'b0 : n869));
assign n570  = /* LUT    3 20  0 */ (n73 ? (n170 ? 1'b1 : !n133) : (n170 ? n133 : 1'b0));
assign n2199 = /* LUT    2 20  2 */ (n443 ? (n142 ? !n49 : 1'b0) : (n142 ? !n49 : !n141));
assign n896  = /* LUT    6 25  6 */ (n507 ? n784 : n706);
assign n2201 = /* LUT   11 18  3 */ (n53 ? (n11 ? !n839 : 1'b0) : n1104);
assign n2202 = /* LUT   12 27  6 */ (\indata[17]  ? (n1344 ? (\inExp[0]  ? 1'b1 : !ready) : (\inExp[0]  ? ready : 1'b0)) : (n1344 ? !ready : 1'b0));
assign n2203 = /* LUT    6 19  6 */ (ready ? (\inExp[0]  ? \indata[2]  : 1'b0) : n863);
assign n937  = /* LUT    7 24  1 */ (n861 ? n936 : n685);
assign n2204 = /* LUT    4 19  3 */ (n646 ? (n157 ? !n106 : (n127 ? !n106 : 1'b0)) : (n157 ? 1'b0 : (n127 ? !n106 : 1'b0)));
assign n924  = /* LUT    7 22  5 */ (reset ? 1'b0 : !n923);
assign n1038 = /* LUT    9 23  5 */ (n983 ? (n1037 ? 1'b1 : !n861) : (n1037 ? n861 : 1'b0));
assign n690  = /* LUT    4 25  3 */ (n91 ? (n196 ? 1'b1 : !n133) : (n196 ? n133 : 1'b0));
assign n2206 = /* LUT   10 22  2 */ !n844;
assign n2207 = /* LUT   15 22  2 */ !n1428;
assign n2208 = /* LUT    3 19  2 */ (ds ? (n562 ? (n77 ? !ready : 1'b0) : 1'b0) : (n562 ? (n77 ? 1'b1 : ready) : 1'b0));
assign n2209 = /* LUT    7 16  4 */ (n731 ? 1'b1 : (n915 ? 1'b1 : (n628 ? 1'b1 : n735)));
assign n2210 = /* LUT    5 23  4 */ (n672 ? n524 : 1'b0);
assign n2211 = /* LUT   12 22  0 */ (n1326 ? (n981 ? n1327 : !n1327) : (n981 ? !n1327 : n1327));
assign n2212 = /* LUT   13 25  5 */ (n732 ? n1327 : 1'b0);
assign n2213 = /* LUT    4 30  7 */ \inMod[21] ;
assign n2214 = /* LUT    5 17  0 */ (n253 ? (reset ? n635 : n557) : n635);
assign n2215 = /* LUT    1 22  0 */ (n357 ? !n188 : n188);
assign n2217 = /* LUT    9 18  5 */ (n957 ? n732 : 1'b0);
assign n2218 = /* LUT   10 24  7 */ (n1161 ? (n786 ? n177 : !n177) : (n786 ? !n177 : n177));
assign n1358 = /* LUT   13 19  1 */ (n1204 ? (n918 ? n1293 : 1'b1) : (n918 ? n1293 : 1'b0));
assign n2220 = /* LUT   15 21  0 */ (n1419 ? (n787 ? 1'b1 : (n142 ? !n49 : 1'b1)) : (n787 ? (n142 ? n49 : 1'b0) : 1'b0));
assign n2221 = /* LUT   10 21  4 */ (\indata[25]  ? (n1133 ? (\inExp[0]  ? 1'b1 : !ready) : (\inExp[0]  ? ready : 1'b0)) : (n1133 ? !ready : 1'b0));
assign n2222 = /* LUT    5 27  4 */ (n804 ? (n102 ? n772 : !n772) : (n102 ? !n772 : n772));
assign n2223 = /* LUT    6 18  1 */ !n639;
assign n2224 = /* LUT    4 21  3 */ (n658 ? (n158 ? !n106 : (n157 ? !n106 : 1'b0)) : (n158 ? (n157 ? 1'b0 : !n106) : 1'b0));
assign n2225 = /* LUT   14 20  4 */ (n1226 ? (n142 ? (n686 ? 1'b1 : !n49) : 1'b1) : (n142 ? (n686 ? n49 : 1'b0) : 1'b0));
assign n2226 = /* LUT    5 25  5 */ (n612 ? n524 : 1'b0);
assign n1071 = /* LUT    9 26  0 */ (n1055 ? (n1067 ? 1'b1 : !n811) : (n1067 ? n811 : 1'b0));
assign n2228 = /* LUT    5 20  6 */ (n627 ? (ds ? (n77 ? !ready : 1'b0) : (n77 ? 1'b1 : ready)) : 1'b0);
assign n2229 = /* LUT    1 17  2 */ (n279 ? (n150 ? n272 : !n272) : (n150 ? !n272 : n272));
assign n2230 = /* LUT    2 24  7 */ (n514 ? (n217 ? n215 : !n215) : (n217 ? !n215 : n215));
assign n2231 = /* LUT   13 22  1 */ (n1380 ? (n1107 ? n1379 : !n1379) : (n1107 ? !n1379 : n1379));
assign n2232 = /* LUT    3 22  3 */ (n464 ? (n157 ? !n106 : (n381 ? !n106 : 1'b0)) : (n157 ? 1'b0 : (n381 ? !n106 : 1'b0)));
assign n1220 = /* LUT   11 20  6 */ (n1216 ? (n918 ? n1120 : 1'b1) : (n918 ? n1120 : 1'b0));
assign n2234 = /* LUT    3 28  3 */ (n615 ? (n538 ? 1'b1 : !n253) : (n538 ? n253 : 1'b0));
assign n2235 = /* LUT   11 27  7 */ (n1086 ? (n1282 ? !n839 : (n839 ? 1'b0 : !n53)) : (n1282 ? (n839 ? 1'b0 : n53) : 1'b0));
assign n2236 = /* LUT    7 26  0 */ (reset ? n897 : (n897 ? (n290 ? n618 : 1'b1) : (n290 ? n618 : 1'b0)));
assign n1004 = /* LUT    9 19  2 */ (n867 ? (n918 ? 1'b1 : n750) : (n918 ? 1'b0 : n750));
assign n2238 = /* LUT   12 19  5 */ (n1300 ? (n121 ? n952 : !n952) : (n121 ? !n952 : n952));
assign n2239 = /* LUT    1 26  0 */ (n429 ? (n397 ? n430 : !n430) : (n397 ? !n430 : n430));
assign n2240 = /* LUT   12 24  4 */ (n17 ? (n53 ? !n839 : n1264) : (n53 ? 1'b0 : n1264));
assign n1016 = /* LUT    9 21  2 */ (n1013 ? (n970 ? 1'b1 : !n811) : (n970 ? n811 : 1'b0));
assign n2242 = /* LUT    6 23  4 */ (n253 ? n884 : n886);
assign n2243 = /* LUT    6 24  5 */ (n778 ? n524 : 1'b0);
assign n2244 = /* LUT    2 23  3 */ (n497 ? (n125 ? n195 : !n195) : (n125 ? !n195 : n195));
assign n2245 = /* LUT    3 21  7 */ (n316 ? (n347 ? 1'b1 : n324) : (n347 ? !n324 : 1'b0));
assign n2246 = /* LUT   11 19  0 */ (n1101 ? (n290 ? n749 : 1'b1) : (n290 ? n749 : 1'b0));
assign n2247 = /* LUT    9 27  7 */ (n579 ? (ready ? \indata[19]  : 1'b1) : (ready ? \indata[19]  : 1'b0));
assign n2248 = /* LUT   12 26  5 */ (n111 ? (\indata[30]  ? (ready ? \inExp[0]  : 1'b1) : !ready) : (\indata[30]  ? (ready ? \inExp[0]  : 1'b0) : 1'b0));
assign n2249 = /* LUT    7 18  7 */ !n848;
assign n2250 = /* LUT    4 18  0 */ \inMod[3] ;
assign n2251 = /* LUT    7 25  6 */ !n898;
assign n2252 = /* LUT   13 23  6 */ (n1395 ? (n1377 ? n1252 : !n1252) : (n1377 ? !n1252 : n1252));
assign n2253 = /* LUT    7 23  6 */ (\indata[11]  ? (n931 ? (\inExp[0]  ? 1'b1 : !ready) : (\inExp[0]  ? ready : 1'b0)) : (n931 ? !ready : 1'b0));
assign n681  = /* LUT    4 24  4 */ (n596 ? (n519 ? 1'b1 : n507) : (n519 ? !n507 : 1'b0));
assign n2255 = /* LUT    1 20  3 */ (n329 ? (n213 ? n145 : !n145) : (n213 ? !n145 : n145));
assign n2256 = /* LUT   14 18  0 */ (n1001 ? (n918 ? 1'b1 : n1215) : (n918 ? 1'b0 : n1215));
assign n2257 = /* LUT   15 23  1 */ (n578 ? (n1425 ? 1'b1 : (n49 ? n142 : 1'b0)) : (n1425 ? (n49 ? !n142 : 1'b1) : 1'b0));
assign n2258 = /* LUT   10 19  3 */ (n916 ? (n659 ? 1'b1 : (n49 ? !n50 : 1'b1)) : (n659 ? (n49 ? n50 : 1'b0) : 1'b0));
assign n1498 = /* LUT   18 21  6 */ (n1470 ? 1'b1 : (n1452 ? 1'b1 : (n77 ? 1'b1 : n1464)));
assign n2260 = /* LUT   16 23  3 */ (n1440 ? 1'b1 : (n1434 ? 1'b1 : (n969 ? 1'b1 : n1423)));
assign n2261 = /* LUT    4 23  6 */ (n253 ? (reset ? n592 : n594) : n592);
assign n913  = /* LUT    7 15  3 */ (n845 ? 1'b1 : (n912 ? 1'b1 : (n727 ? 1'b1 : n545)));
assign n2262 = /* LUT    9 24  3 */ (ready ? \indata[3]  : n756);
assign n2263 = /* LUT   10 17  6 */ (n7 ? (\indata[26]  ? (\inExp[0]  ? 1'b1 : !ready) : !ready) : (\indata[26]  ? (\inExp[0]  ? ready : 1'b0) : 1'b0));
assign n2264 = /* LUT   12 21  1 */ (n1319 ? (n1019 ? n1120 : !n1120) : (n1019 ? !n1120 : n1120));
assign n2265 = /* LUT    5 18  1 */ (reset ? n638 : (n638 ? (n253 ? n467 : 1'b1) : (n253 ? n467 : 1'b0)));
assign n2266 = /* LUT    1 23  7 */ (n388 ? (n377 ? n134 : !n134) : (n377 ? !n134 : n134));
assign n2267 = /* LUT    2 22  4 */ (n486 ? (n100 ? n170 : !n170) : (n100 ? !n170 : n170));
assign n2268 = /* LUT   10 27  6 */ (n1028 ? (n1044 ? 1'b1 : !n811) : (n1044 ? n811 : 1'b0));
assign n2269 = /* LUT    5 28  5 */ (n816 ? (n128 ? n707 : !n707) : (n128 ? !n707 : n707));
assign n2270 = /* LUT   10 20  7 */ (n286 ? (\indata[8]  ? 1'b1 : !ready) : (\indata[8]  ? ready : 1'b0));
assign n2271 = /* LUT   11 22  5 */ (n1244 ? (n972 ? n1021 : !n1021) : (n972 ? !n1021 : n1021));
assign n2272 = /* LUT    1 24  3 */ (n404 ? (n219 ? n227 : !n227) : (n219 ? !n227 : n227));
assign n2273 = /* LUT    5 26  4 */ (n796 ? (n80 ? n612 : !n612) : (n80 ? !n612 : n612));
assign n2274 = /* LUT   17 21  0 */ (\inExp[11]  ? (ds ? (n1451 ? 1'b1 : ready) : n1451) : (ds ? (n1451 ? !ready : 1'b0) : n1451));
assign n761  = /* LUT    5 21  5 */ (n576 ? (n324 ? 1'b1 : n392) : (n324 ? 1'b0 : n392));
assign n2275 = /* LUT    1 18  3 */ (n295 ? (n169 ? n100 : !n100) : (n169 ? !n100 : n100));
assign n2276 = /* LUT    6 21  7 */ (n324 ? n876 : n159);
assign n2277 = /* LUT    3 23  0 */ (n133 ? (n231 ? n324 : 1'b0) : 1'b0);
assign n2278 = /* LUT    2 21  6 */ (n477 ? (n81 ? n154 : !n154) : (n81 ? !n154 : n154));
assign n2279 = /* LUT   11 21  1 */ (n1230 ? (n1041 ? n979 : !n979) : (n1041 ? !n979 : n979));
assign n2280 = /* LUT   12 20  6 */ (n1316 ? (n763 ? n998 : !n998) : (n763 ? !n998 : n998));
assign n2281 = /* LUT    6 16  6 */ (n66 ? (n49 ? (n50 ? 1'b1 : n728) : n728) : (n49 ? (n50 ? 1'b0 : n728) : n728));
assign n2282 = /* LUT   11 24  6 */ (n1272 ? (n585 ? n1077 : !n1077) : (n585 ? !n1077 : n1077));
assign n2283 = /* LUT   12 18  6 */ (n1196 ? (n675 ? 1'b1 : (reset ? 1'b1 : !n290)) : (n675 ? (reset ? 1'b0 : n290) : 1'b0));
assign n2284 = /* LUT    9 22  3 */ (n67 ? (n968 ? (n839 ? !n53 : 1'b1) : (n839 ? 1'b0 : n53)) : (n968 ? !n53 : 1'b0));
assign n2285 = /* LUT    6 22  3 */ !n180;
assign n2286 = /* LUT   18 19  1 */ (ready ? (\inExp[5]  ? (ds ? 1'b1 : n1469) : (ds ? 1'b0 : n1469)) : n1469);
assign n2287 = /* LUT    3 18  6 */ (n253 ? (reset ? n449 : n95) : n449);
assign n2288 = /* LUT    6 27  4 */ (n810 ? (n253 ? n521 : 1'b1) : (n253 ? n521 : 1'b0));
assign n2289 = /* LUT   11 16  1 */ (n841 ? (n660 ? 1'b1 : (n49 ? !n50 : 1'b1)) : (n660 ? (n49 ? n50 : 1'b0) : 1'b0));
assign n2290 = /* LUT   12 25  4 */ (\indata[21]  ? (n1337 ? (\inExp[0]  ? 1'b1 : !ready) : (\inExp[0]  ? ready : 1'b0)) : (n1337 ? !ready : 1'b0));
assign n2291 = /* LUT    7 19  4 */ !n482;
assign n2292 = /* LUT    3 24  6 */ (n601 ? (n157 ? !n106 : (n400 ? !n106 : 1'b0)) : (n157 ? 1'b0 : (n400 ? !n106 : 1'b0)));
assign n2293 = /* LUT    4 17  1 */ (n632 ? (n305 ? 1'b1 : (n50 ? !n49 : 1'b1)) : (n305 ? (n50 ? n49 : 1'b0) : 1'b0));
assign n2294 = /* LUT    7 30  7 */ \inMod[29] ;
assign n2295 = /* LUT    1 19  4 */ (n311 ? (n196 ? n247 : !n247) : (n196 ? !n247 : n247));
assign n2296 = /* LUT   12 23  0 */ (n1335 ? (n344 ? n1227 : !n1227) : (n344 ? !n1227 : n1227));
assign n2297 = /* LUT    9 20  6 */ (n621 ? n524 : 1'b0);
assign n2298 = /* LUT   13 24  7 */ (n1405 ? (n1348 ? n1173 : !n1173) : (n1348 ? !n1173 : n1173));
assign n2299 = /* LUT    5 16  0 */ (n544 ? 1'b1 : (n630 ? 1'b1 : (n629 ? 1'b1 : n631)));
assign n2300 = /* LUT    1 21  0 */ (n334 ? (n230 ? n344 : !n344) : (n230 ? !n344 : n344));
assign n2301 = /* LUT   19 22  2 */ (n1466 ? (\inExp[18]  ? 1'b1 : (ready ? !ds : 1'b1)) : (\inExp[18]  ? (ready ? ds : 1'b0) : 1'b0));
assign n2302 = /* LUT   13 18  7 */ (n1275 ? (n1351 ? 1'b1 : n290) : (n1351 ? !n290 : 1'b0));
assign n2303 = /* LUT   10 25  5 */ (n1167 ? (n1070 ? n890 : !n890) : (n1070 ? !n890 : n890));
assign n1441 = /* LUT   15 20  0 */ (n598 ? 1'b1 : (n1420 ? 1'b1 : (n1425 ? 1'b1 : n1364)));
assign n2305 = /* LUT   10 18  4 */ (n290 ? n868 : n1112);
assign n2306 = /* LUT   11 25  1 */ (n1278 ? (n1085 ? n344 : !n344) : (n1085 ? !n344 : n344));
assign n2307 = /* LUT   18 20  5 */ (ready ? (n1468 ? (\inExp[20]  ? 1'b1 : !ds) : (\inExp[20]  ? ds : 1'b0)) : n1468);
assign n2308 = /* LUT    7 22  2 */ (n288 ? (n359 ? !n106 : (n157 ? !n106 : 1'b0)) : (n359 ? (n157 ? 1'b0 : !n106) : 1'b0));
assign n2309 = /* LUT    4 25  4 */ (n374 ? (n690 ? 1'b1 : !n324) : (n690 ? n324 : 1'b0));
assign n2310 = /* LUT    4 22  5 */ !n140;
assign n2311 = /* LUT   14 21  4 */ (n1295 ? n732 : 1'b0);
assign n2312 = /* LUT    9 25  0 */ (n788 ? (reset ? 1'b1 : (n253 ? n306 : 1'b1)) : (reset ? 1'b0 : (n253 ? n306 : 1'b0)));
assign n2313 = /* LUT   10 16  5 */ (n861 ? n1093 : n1090);
assign n2314 = /* LUT    5 24  7 */ (n683 ? (n253 ? n518 : 1'b1) : (n253 ? n518 : 1'b0));
assign n2315 = /* LUT    5 19  6 */ (ready ? (n748 ? !ds : 1'b0) : (n748 ? n77 : 1'b0));
assign n2316 = /* LUT    6 26  3 */ (n789 ? (reset ? 1'b1 : (n255 ? 1'b1 : !n253)) : (reset ? 1'b0 : (n255 ? n253 : 1'b0)));
assign n2317 = /* LUT    2 25  5 */ (reset ? n413 : (n522 ? (n413 ? 1'b1 : n253) : (n413 ? !n253 : 1'b0)));
assign n2318 = /* LUT   10 26  1 */ (n1176 ? (n1076 ? n900 : !n900) : (n1076 ? !n900 : n900));
assign n2319 = /* LUT   11 17  6 */ \inMod[13] ;
assign n2320 = /* LUT   13 21  3 */ (n1371 ? (n1368 ? n1309 : !n1309) : (n1368 ? !n1309 : n1309));
assign n2321 = /* LUT    5 29  6 */ (n827 ? (n611 ? n217 : !n217) : (n611 ? !n217 : n217));
assign n2322 = /* LUT    3 25  1 */ (n324 ? n607 : n372);
assign n459  = /* LUT    2 19  1 */ (n324 ? n458 : n351);
assign n2323 = /* LUT    6 28  3 */ (n668 ? (n507 ? 1'b1 : n709) : (n507 ? 1'b0 : n709));
assign n2324 = /* LUT   10 23  6 */ (n1149 ? (n1042 ? n855 : !n855) : (n1042 ? !n855 : n855));
assign n2325 = /* LUT   11 23  6 */ (n1260 ? (n1067 ? n890 : !n890) : (n1067 ? !n890 : n890));
assign n2326 = /* LUT   11 26  5 */ (n3 ? (n53 ? !n839 : (n839 ? 1'b0 : n1173)) : (n53 ? 1'b0 : (n839 ? 1'b0 : n1173)));
assign n921  = /* LUT    7 21  0 */ (n811 ? n920 : n880);
assign n2328 = /* LUT    1 25  0 */ (n409 ? (n411 ? n417 : !n417) : (n411 ? !n417 : n417));
assign n2329 = /* LUT   15 21  7 */ (n1418 ? (n782 ? 1'b1 : (n49 ? !n142 : 1'b1)) : (n782 ? (n49 ? n142 : 1'b0) : 1'b0));
assign n2330 = /* LUT    5 27  3 */ (n803 ? (n100 ? n520 : !n520) : (n100 ? !n520 : n520));
assign n2331 = /* LUT   14 22  2 */ (n290 ? n980 : n1430);
assign n2332 = /* LUT    5 22  4 */ (n253 ? n674 : n770);
assign n2333 = /* LUT   14 24  2 */ (n1353 ? n732 : 1'b0);
assign n2334 = /* LUT    2 26  1 */ (n524 ? n493 : 1'b0);
assign n2335 = /* LUT    6 20  4 */ (n109 ? (\inExp[0]  ? (ready ? \indata[0]  : 1'b1) : 1'b1) : (\inExp[0]  ? (ready ? \indata[0]  : 1'b0) : ready));
assign n2336 = /* LUT    6 25  7 */ (n791 ? (n896 ? 1'b1 : n253) : (n896 ? !n253 : 1'b0));
assign n2337 = /* LUT    2 20  5 */ (n89 ? (n194 ? 1'b1 : !n133) : (n194 ? n133 : 1'b0));
assign n571  = /* LUT    3 20  1 */ (n324 ? n570 : n348);
assign n2338 = /* LUT   11 18  0 */ (n1192 ? (n1199 ? 1'b1 : n918) : (n1199 ? !n918 : 1'b0));
assign n2339 = /* LUT   12 27  7 */ (n302 ? (ready ? \indata[17]  : 1'b1) : (ready ? \indata[17]  : 1'b0));
assign n2340 = /* LUT    6 19  7 */ (n453 ? (ready ? \indata[2]  : 1'b1) : (ready ? \indata[2]  : 1'b0));
assign n2341 = /* LUT    7 24  2 */ (\indata[14]  ? (n937 ? (\inExp[0]  ? 1'b1 : !ready) : (\inExp[0]  ? ready : 1'b0)) : (n937 ? !ready : 1'b0));
assign n2342 = /* LUT    4 19  0 */ (n560 ? (reset ? 1'b1 : (n96 ? 1'b1 : !n253)) : (reset ? 1'b0 : (n96 ? n253 : 1'b0)));
assign n2343 = /* LUT   14 19  0 */ (n918 ? n1214 : n1029);
assign n1037 = /* LUT    9 23  4 */ (n1032 ? (n972 ? 1'b1 : !n811) : (n972 ? n811 : 1'b0));
assign n2345 = /* LUT   10 22  1 */ (reset ? n1018 : (n1018 ? (n290 ? n176 : 1'b1) : (n290 ? n176 : 1'b0)));
assign n2346 = /* LUT   15 22  3 */ (reset ? n1428 : (n290 ? n671 : n1428));
assign n2347 = /* LUT    3 19  5 */ (ready ? (n564 ? !ds : 1'b0) : (n564 ? n77 : 1'b0));
assign n2348 = /* LUT    7 16  5 */ (n835 ? 1'b0 : (reset ? 1'b0 : (n49 ? n50 : 1'b0)));
assign n2349 = /* LUT    9 21  5 */ (n457 ? (ready ? \indata[28]  : 1'b1) : (ready ? \indata[28]  : 1'b0));
assign n2350 = /* LUT    5 23  3 */ (n253 ? n202 : n776);
assign n2351 = /* LUT   12 22  3 */ (n1330 ? (n905 ? n1108 : !n1108) : (n905 ? !n1108 : n1108));
assign n2352 = /* LUT   13 25  4 */ (n49 ? n50 : 1'b0);
assign n2353 = /* LUT    4 30  6 */ \inMod[20] ;
assign n2354 = /* LUT    5 17  3 */ !n640;
assign n2355 = /* LUT    1 22  1 */ (n364 ? (n354 ? n184 : !n184) : (n354 ? !n184 : n184));
assign n2356 = /* LUT    9 18  6 */ (n917 ? n732 : 1'b0);
assign n2357 = /* LUT   10 24  6 */ (n1160 ? (n785 ? n763 : !n763) : (n785 ? !n763 : n763));
assign n929  = /* LUT    7 23  1 */ (n861 ? n928 : n926);
assign n2358 = /* LUT   14 18  7 */ (n742 ? (n1411 ? 1'b1 : n290) : (n1411 ? !n290 : 1'b0));
assign n2359 = /* LUT    4 21  4 */ (n230 ? (n132 ? 1'b1 : n133) : (n132 ? !n133 : 1'b0));
assign n1072 = /* LUT    9 26  1 */ (n861 ? n1071 : n989);
assign n2360 = /* LUT   10 19  4 */ (n842 ? (n661 ? 1'b1 : (n50 ? !n49 : 1'b1)) : (n661 ? (n50 ? n49 : 1'b0) : 1'b0));
assign n2361 = /* LUT    5 25  4 */ (n597 ? n524 : 1'b0);
assign n2362 = /* LUT    1 17  5 */ (n282 ? (n153 ? n81 : !n81) : (n153 ? !n81 : n81));
assign n2363 = /* LUT    2 24  6 */ (n513 ? (n322 ? n208 : !n208) : (n322 ? !n208 : n208));
assign n2364 = /* LUT   13 22  2 */ (n1381 ? (n1008 ? n865 : !n865) : (n1008 ? !n865 : n865));
assign n2365 = /* LUT    3 22  0 */ !n480;
assign n2366 = /* LUT    2 18  6 */ (ready ? (n452 ? !ds : 1'b0) : (n452 ? n77 : 1'b0));
assign n2367 = /* LUT   11 20  7 */ (n987 ? (n1220 ? 1'b1 : n290) : (n1220 ? !n290 : 1'b0));
assign n1282 = /* LUT   11 27  6 */ (n861 ? n1281 : n1152);
assign n2368 = /* LUT    9 19  1 */ (n290 ? n946 : n1003);
assign n2369 = /* LUT   12 19  2 */ (n1297 ? (n853 ? n1295 : !n1295) : (n853 ? !n1295 : n1295));
assign n2370 = /* LUT    1 26  1 */ (n436 ? (n412 ? n398 : !n398) : (n412 ? !n398 : n398));
assign n2371 = /* LUT    5 28  2 */ (n813 ? (n125 ? n696 : !n696) : (n125 ? !n696 : n696));
assign n1438 = /* LUT   15 16  6 */ (n49 ? 1'b0 : (n50 ? n142 : 1'b0));
assign n2372 = /* LUT    6 23  5 */ (n773 ? n524 : 1'b0);
assign n2373 = /* LUT    3 21  6 */ (n77 ? (n583 ? (ready ? !ds : 1'b1) : 1'b0) : (n583 ? (ready ? !ds : 1'b0) : 1'b0));
assign n2374 = /* LUT    4 20  3 */ (n253 ? (n556 ? (reset ? n566 : 1'b1) : (reset ? n566 : 1'b0)) : n566);
assign n2375 = /* LUT    2 23  4 */ (n498 ? (n122 ? n196 : !n196) : (n122 ? !n196 : n196));
assign n2376 = /* LUT    7 18  4 */ (n846 ? (reset ? 1'b1 : (n290 ? n101 : 1'b1)) : (reset ? 1'b0 : (n290 ? n101 : 1'b0)));
assign n2377 = /* LUT    9 27  6 */ (\indata[19]  ? (n1084 ? (\inExp[0]  ? 1'b1 : !ready) : (\inExp[0]  ? ready : 1'b0)) : (n1084 ? !ready : 1'b0));
assign n2378 = /* LUT    6 24  4 */ (n723 ? (n787 ? 1'b1 : !n253) : (n787 ? n253 : 1'b0));
assign n2379 = /* LUT    3 27  6 */ (reset ? n533 : (n253 ? n262 : n533));
assign n2380 = /* LUT    7 25  5 */ (n891 ? (reset ? 1'b1 : (n290 ? n907 : 1'b1)) : (reset ? 1'b0 : (n290 ? n907 : 1'b0)));
assign n2381 = /* LUT    4 18  3 */ \inMod[4] ;
assign n2382 = /* LUT   11 19  3 */ (n882 ? (n1208 ? 1'b1 : n290) : (n1208 ? !n290 : 1'b0));
assign n2383 = /* LUT   13 23  5 */ (n1394 ? (n948 ? n1265 : !n1265) : (n948 ? !n1265 : n1265));
assign n2384 = /* LUT    1 20  0 */ (n315 ? (n210 ? n144 : !n144) : (n210 ? !n144 : n144));
assign n2385 = /* LUT   15 23  0 */ (n416 ? (n1432 ? 1'b1 : (n142 ? n49 : 1'b0)) : (n1432 ? (n142 ? !n49 : 1'b1) : 1'b0));
assign n2386 = /* LUT   18 21  7 */ (n1454 ? 1'b1 : (n1498 ? 1'b1 : (n1455 ? 1'b1 : n1497)));
assign n2387 = /* LUT    4 26  4 */ (n524 ? n611 : 1'b0);
assign n2388 = /* LUT    4 23  7 */ !n592;
assign n912  = /* LUT    7 15  2 */ (n732 ? 1'b1 : (n550 ? 1'b1 : (n841 ? 1'b1 : n632)));
assign n2390 = /* LUT   12 21  2 */ (n1320 ? (n734 ? n917 : !n917) : (n734 ? !n917 : n917));
assign n2391 = /* LUT   10 17  7 */ (n651 ? (ready ? \indata[27]  : 1'b1) : (ready ? \indata[27]  : 1'b0));
assign n2392 = /* LUT    4 29  7 */ (n721 ? (n606 ? 1'b1 : !n253) : (n606 ? n253 : 1'b0));
assign n2393 = /* LUT    5 18  2 */ (n639 ? (reset ? 1'b1 : (n555 ? 1'b1 : !n290)) : (reset ? 1'b0 : (n555 ? n290 : 1'b0)));
assign n2394 = /* LUT    1 23  6 */ (n387 ? (n379 ? n381 : !n381) : (n379 ? !n381 : n381));
assign n2395 = /* LUT    2 22  3 */ (n485 ? (n103 ? n169 : !n169) : (n103 ? !n169 : n169));
assign n2396 = /* LUT   10 27  7 */ (n1039 ? (n1045 ? 1'b1 : !n811) : (n1045 ? n811 : 1'b0));
assign n2397 = /* LUT    6 29  1 */ (n773 ? (n703 ? 1'b1 : n507) : (n703 ? !n507 : 1'b0));
assign n2398 = /* LUT   11 22  2 */ (n1241 ? (n577 ? n1045 : !n1045) : (n577 ? !n1045 : n1045));
assign n2399 = /* LUT    7 20  0 */ (n48 ? (n53 ? !n839 : (n857 ? !n839 : 1'b0)) : (n53 ? 1'b0 : (n857 ? !n839 : 1'b0)));
assign n2400 = /* LUT   10 15  7 */ (n838 ? (n50 ? !n49 : 1'b0) : (n50 ? !n49 : !n834));
assign n2401 = /* LUT    1 24  0 */ (n389 ? (n401 ? n221 : !n221) : (n401 ? !n221 : n221));
assign n2402 = /* LUT    5 26  5 */ (n797 ? (n81 ? n774 : !n774) : (n81 ? !n774 : n774));
assign n1112 = /* LUT   10 18  3 */ (n1109 ? (n918 ? n997 : 1'b1) : (n918 ? n997 : 1'b0));
assign n2404 = /* LUT   17 21  3 */ (ready ? (n1454 ? (ds ? \inExp[14]  : 1'b1) : (ds ? \inExp[14]  : 1'b0)) : n1454);
assign n2405 = /* LUT    5 21  4 */ (n77 ? (n760 ? (ready ? !ds : 1'b1) : 1'b0) : (n760 ? (ready ? !ds : 1'b0) : 1'b0));
assign n2406 = /* LUT    1 18  4 */ (n296 ? (n170 ? n102 : !n102) : (n170 ? !n102 : n102));
assign n2407 = /* LUT   19 19  2 */ (n1457 ? (\inExp[28]  ? 1'b1 : (ds ? !ready : 1'b1)) : (\inExp[28]  ? (ds ? ready : 1'b0) : 1'b0));
assign n2408 = /* LUT    6 21  4 */ (n77 ? (n875 ? (ds ? !ready : 1'b1) : 1'b0) : (n875 ? (ds ? 1'b0 : ready) : 1'b0));
assign n2409 = /* LUT    2 27  7 */ !n531;
assign n2410 = /* LUT    3 23  3 */ (n493 ? n507 : 1'b0);
assign n2411 = /* LUT    2 21  7 */ (n478 ? (n274 ? n155 : !n155) : (n274 ? !n155 : n155));
assign n2415 = /* LUT   12 20  5 */ (n1315 ? (n593 ? n997 : !n997) : (n593 ? !n997 : n997));
assign n2416 = /* LUT    7 27  2 */ !n903;
assign n2417 = /* LUT    4 28  0 */ (n713 ? (n507 ? n536 : 1'b1) : (n507 ? n536 : 1'b0));
assign n2418 = /* LUT   11 24  7 */ (n1273 ? (n737 ? n1078 : !n1078) : (n737 ? !n1078 : n1078));
assign n2419 = /* LUT    5 29  1 */ (n822 ? (n232 ? n536 : !n536) : (n232 ? !n536 : n536));
assign n2420 = /* LUT   13 15  2 */ (n1346 ? (ds ? !n49 : (n49 ? 1'b0 : !ready)) : (ds ? (n49 ? 1'b0 : ready) : 1'b0));
assign n2421 = /* LUT   11 26  2 */ !n1079;
assign n2422 = /* LUT   18 19  2 */ (n1464 ? (\inExp[7]  ? 1'b1 : (ready ? !ds : 1'b1)) : (\inExp[7]  ? (ready ? ds : 1'b0) : 1'b0));
assign n2423 = /* LUT    3 18  7 */ (n205 ? (n286 ? !n106 : (n106 ? 1'b0 : !n157)) : (n286 ? (n106 ? 1'b0 : n157) : 1'b0));
assign n2424 = /* LUT    7 19  7 */ !n856;
assign n1338 = /* LUT   12 25  5 */ (n1174 ? (n861 ? 1'b1 : n1139) : (n861 ? 1'b0 : n1139));
assign n2425 = /* LUT    3 24  7 */ (n602 ? (n223 ? !n106 : (n157 ? !n106 : 1'b0)) : (n223 ? (n157 ? 1'b0 : !n106) : 1'b0));
assign n2426 = /* LUT    4 17  2 */ (n550 ? (n455 ? 1'b1 : (n49 ? !n50 : 1'b1)) : (n455 ? (n49 ? n50 : 1'b0) : 1'b0));
assign n2427 = /* LUT    7 30  4 */ \inMod[26] ;
assign n2428 = /* LUT    1 19  3 */ (n310 ? (n195 ? n122 : !n122) : (n195 ? !n122 : n122));
assign n2429 = /* LUT   12 23  1 */ (n38 ? (n1248 ? (n53 ? !n839 : 1'b1) : (n53 ? !n839 : 1'b0)) : (n1248 ? !n53 : 1'b0));
assign n2430 = /* LUT   13 24  4 */ (n1402 ? (n1356 ? n968 : !n968) : (n1356 ? !n968 : n968));
assign n2431 = /* LUT    5 16  1 */ (n630 ? (n50 ? (n49 ? n733 : 1'b1) : 1'b1) : (n50 ? (n49 ? n733 : 1'b0) : 1'b0));
assign n2432 = /* LUT    1 21  3 */ (n63 ? (n154 ? 1'b1 : !n133) : (n154 ? n133 : 1'b0));
assign n2433 = /* LUT   19 22  3 */ (n1497 ? (\inExp[2]  ? 1'b1 : (ds ? !ready : 1'b1)) : (\inExp[2]  ? (ds ? ready : 1'b0) : 1'b0));
assign n2434 = /* LUT   13 18  0 */ (n1287 ? n732 : 1'b0);
assign n2435 = /* LUT   10 25  2 */ (n1164 ? (n1059 ? n734 : !n734) : (n1059 ? !n734 : n734));
assign n2436 = /* LUT   15 20  1 */ (n1439 ? 1'b1 : (n1441 ? 1'b1 : (n1415 ? 1'b1 : n1360)));
assign n2437 = /* LUT   11 25  0 */ (n1274 ? (n781 ? n920 : !n920) : (n781 ? !n920 : n920));
assign n2438 = /* LUT   18 20  4 */ (n1463 ? (\inExp[6]  ? 1'b1 : (ds ? !ready : 1'b1)) : (\inExp[6]  ? (ds ? ready : 1'b0) : 1'b0));
assign n2439 = /* LUT    7 22  3 */ (reset ? n877 : (n877 ? (n290 ? n306 : 1'b1) : (n290 ? n306 : 1'b0)));
assign n2440 = /* LUT    9 23  3 */ (n462 ? (ready ? \indata[12]  : 1'b1) : (ready ? \indata[12]  : 1'b0));
assign n691  = /* LUT    4 25  5 */ (n138 ? (n324 ? 1'b1 : n206) : (n324 ? 1'b0 : n206));
assign n2441 = /* LUT    4 22  4 */ !n591;
assign n1427 = /* LUT   14 21  5 */ (n1202 ? (n918 ? n1295 : 1'b1) : (n918 ? n1295 : 1'b0));
assign n2443 = /* LUT    5 24  4 */ (n676 ? n524 : 1'b0);
assign n2444 = /* LUT    9 25  3 */ (n1026 ? (n811 ? n1031 : 1'b1) : (n811 ? n1031 : 1'b0));
assign n1093 = /* LUT   10 16  4 */ (n1000 ? (n1042 ? 1'b1 : !n811) : (n1042 ? n811 : 1'b0));
assign n2446 = /* LUT   13 27  2 */ (n811 ? (n861 ? n1085 : 1'b0) : 1'b0);
assign n748  = /* LUT    5 19  5 */ (n136 ? (n324 ? 1'b1 : n346) : (n324 ? 1'b0 : n346));
assign n2447 = /* LUT    6 26  2 */ (reset ? n494 : (n494 ? (n253 ? n600 : 1'b1) : (n253 ? n600 : 1'b0)));
assign n2448 = /* LUT    2 25  2 */ !n414;
assign n2449 = /* LUT   13 21  2 */ (n1370 ? (n1367 ? n857 : !n857) : (n1367 ? !n857 : n857));
assign n2450 = /* LUT   11 17  5 */ \inMod[12] ;
assign n2451 = /* LUT   10 26  0 */ (n1170 ? (n1075 ? n981 : !n981) : (n1075 ? !n981 : n981));
assign n607  = /* LUT    3 25  0 */ (n87 ? (n193 ? 1'b1 : !n133) : (n193 ? n133 : 1'b0));
assign n2453 = /* LUT    2 19  2 */ (ready ? (n459 ? !ds : 1'b0) : (n459 ? n77 : 1'b0));
assign n2454 = /* LUT   10 23  7 */ (n1150 ? (n1044 ? n932 : !n932) : (n1044 ? !n932 : n932));
assign n2455 = /* LUT   11 23  1 */ (n1255 ? (n767 ? n1066 : !n1066) : (n767 ? !n1066 : n1066));
assign n2456 = /* LUT    4 30  1 */ \inMod[16] ;
assign n2457 = /* LUT    1 25  3 */ (n424 ? (n248 ? n249 : !n249) : (n248 ? !n249 : n249));
assign n2458 = /* LUT   15 21  6 */ (n1363 ? (n518 ? 1'b1 : (n142 ? !n49 : 1'b1)) : (n518 ? (n142 ? n49 : 1'b0) : 1'b0));
assign n2459 = /* LUT    5 27  2 */ (n802 ? (n595 ? n103 : !n103) : (n595 ? !n103 : n103));
assign n1132 = /* LUT   10 21  2 */ (n1023 ? (n811 ? n1076 : 1'b1) : (n811 ? n1076 : 1'b0));
assign n1430 = /* LUT   14 22  1 */ (n957 ? (n1223 ? 1'b1 : n918) : (n1223 ? !n918 : 1'b0));
assign n2462 = /* LUT    5 22  5 */ (n667 ? n524 : 1'b0);
assign n2463 = /* LUT    2 26  0 */ (n257 ? n524 : 1'b0);
assign n2464 = /* LUT    6 20  7 */ (n653 ? (\indata[0]  ? 1'b1 : !ready) : (\indata[0]  ? ready : 1'b0));
assign n2465 = /* LUT    3 20  2 */ (n77 ? (n571 ? (ready ? !ds : 1'b1) : 1'b0) : (n571 ? (ready ? !ds : 1'b0) : 1'b0));
assign n2466 = /* LUT    2 20  4 */ (n75 ? (n133 ? n172 : 1'b1) : (n133 ? n172 : 1'b0));
assign n2467 = /* LUT    6 25  4 */ (n809 ? (n253 ? n541 : 1'b1) : (n253 ? n541 : 1'b0));
assign n2468 = /* LUT   11 18  1 */ (n53 ? (n15 ? !n839 : 1'b0) : n1102);
assign n1343 = /* LUT   12 27  4 */ (n1050 ? (n1066 ? 1'b1 : !n811) : (n1066 ? n811 : 1'b0));
assign n2470 = /* LUT    7 24  3 */ (n464 ? (ready ? \indata[14]  : 1'b1) : (ready ? \indata[14]  : 1'b0));
assign n2471 = /* LUT    4 19  1 */ (n652 ? (n157 ? !n106 : (n244 ? !n106 : 1'b0)) : (n157 ? 1'b0 : (n244 ? !n106 : 1'b0)));
assign n2472 = /* LUT   14 19  1 */ (n1227 ? n732 : 1'b0);
assign n2473 = /* LUT    5 30  0 */ (n829 ? (n493 ? n344 : !n344) : (n493 ? !n344 : n344));
assign n2474 = /* LUT   10 22  0 */ !n764;
assign n2475 = /* LUT    6 17  3 */ (n448 ? 1'b1 : (n736 ? 1'b1 : (n549 ? 1'b1 : n843)));
assign n2476 = /* LUT    7 26  6 */ !n899;
assign n564  = /* LUT    3 19  4 */ (n324 ? n563 : n335);
assign n2477 = /* LUT    9 21  4 */ (\inExp[0]  ? (n1017 ? (\indata[9]  ? 1'b1 : !ready) : (\indata[9]  ? ready : 1'b0)) : (n1017 ? !ready : 1'b0));
assign n2478 = /* LUT   12 24  2 */ (n109 ? (n53 ? !n839 : (n1254 ? !n839 : 1'b0)) : (n53 ? 1'b0 : (n1254 ? !n839 : 1'b0)));
assign n776  = /* LUT    5 23  2 */ (n774 ? (n507 ? 1'b1 : n695) : (n507 ? 1'b0 : n695));
assign n2480 = /* LUT   12 22  2 */ (n1329 ? (n1171 ? n1118 : !n1118) : (n1171 ? !n1118 : n1118));
assign n2481 = /* LUT   13 25  7 */ (n1079 ? (reset ? 1'b1 : (n290 ? n557 : 1'b1)) : (reset ? 1'b0 : (n290 ? n557 : 1'b0)));
assign n2482 = /* LUT    9 18  7 */ (n649 ? n732 : 1'b0);
assign n2483 = /* LUT    1 22  2 */ (n365 ? (n358 ? n325 : !n325) : (n358 ? !n325 : n325));
assign n2484 = /* LUT   10 24  1 */ (n1155 ? (n970 ? n577 : !n577) : (n970 ? !n577 : n577));
assign n2485 = /* LUT    3 27  1 */ (n253 ? (n531 ? (n98 ? 1'b1 : reset) : (n98 ? !reset : 1'b0)) : n531);
assign n2486 = /* LUT    4 24  2 */ (n253 ? n587 : n680);
assign n928  = /* LUT    7 23  0 */ (n927 ? (n779 ? 1'b1 : !n811) : (n779 ? n811 : 1'b0));
assign n1411 = /* LUT   14 18  6 */ (n1212 ? (n918 ? 1'b1 : n1191) : (n918 ? 1'b0 : n1191));
assign n2489 = /* LUT    4 21  5 */ (n114 ? (n211 ? 1'b1 : !n133) : (n211 ? n133 : 1'b0));
assign n2490 = /* LUT   14 20  6 */ (n791 ? (n49 ? (n142 ? 1'b1 : n1362) : n1362) : (n49 ? (n142 ? 1'b0 : n1362) : n1362));
assign n2491 = /* LUT    9 26  2 */ (\indata[22]  ? (n1072 ? (\inExp[0]  ? 1'b1 : !ready) : (\inExp[0]  ? ready : 1'b0)) : (n1072 ? !ready : 1'b0));
assign n2492 = /* LUT   10 19  5 */ (n448 ? (n471 ? 1'b1 : (n49 ? !n50 : 1'b1)) : (n471 ? (n49 ? n50 : 1'b0) : 1'b0));
assign n2493 = /* LUT    5 25  7 */ (n527 ? (reset ? 1'b1 : (n290 ? n438 : 1'b1)) : (reset ? 1'b0 : (n290 ? n438 : 1'b0)));
assign n754  = /* LUT    5 20  4 */ (n137 ? (n395 ? 1'b1 : n324) : (n395 ? !n324 : 1'b0));
assign n2494 = /* LUT    1 17  4 */ (n281 ? (n152 ? n80 : !n80) : (n152 ? !n80 : n80));
assign n2495 = /* LUT    2 24  1 */ (n508 ? (n144 ? n211 : !n211) : (n144 ? !n211 : n211));
assign n2496 = /* LUT   13 22  3 */ (n1382 ? (n1116 ? n1250 : !n1250) : (n1116 ? !n1250 : n1250));
assign n2497 = /* LUT    3 22  1 */ (n321 ? (n157 ? !n106 : (n184 ? !n106 : 1'b0)) : (n157 ? 1'b0 : (n184 ? !n106 : 1'b0)));
assign n452  = /* LUT    2 18  5 */ (n135 ? (n324 ? 1'b1 : n338) : (n324 ? 1'b0 : n338));
assign n2498 = /* LUT    4 29  0 */ (n720 ? (n253 ? n719 : 1'b1) : (n253 ? n719 : 1'b0));
assign n1003 = /* LUT    9 19  0 */ (n953 ? (n918 ? 1'b1 : n657) : (n918 ? 1'b0 : n657));
assign n2500 = /* LUT   12 19  3 */ (n1298 ? (n854 ? n867 : !n867) : (n854 ? !n867 : n867));
assign n2501 = /* LUT    1 26  2 */ !n435;
assign n2502 = /* LUT    5 28  3 */ (n814 ? (n122 ? n778 : !n778) : (n122 ? !n778 : n778));
assign n2503 = /* LUT   10 20  1 */ (n1010 ? (n861 ? 1'b1 : n1125) : (n861 ? 1'b0 : n1125));
assign n2504 = /* LUT    6 29  6 */ (n520 ? (n507 ? 1'b1 : n701) : (n507 ? 1'b0 : n701));
assign n2505 = /* LUT   15 16  7 */ (n910 ? (n1438 ? (ready ? ds : 1'b1) : (ready ? ds : 1'b0)) : (ready ? ds : 1'b0));
assign n2506 = /* LUT    6 24  7 */ (n253 ? n775 : n889);
assign n2507 = /* LUT    4 20  2 */ (n627 ? (n225 ? !n106 : (n157 ? !n106 : 1'b0)) : (n225 ? (n157 ? 1'b0 : !n106) : 1'b0));
assign n2508 = /* LUT    2 23  5 */ (n499 ? (n247 ? n197 : !n197) : (n247 ? !n197 : n197));
assign n2509 = /* LUT    7 18  5 */ (n556 ? (n847 ? 1'b1 : (reset ? 1'b0 : n290)) : (n847 ? (reset ? 1'b1 : !n290) : 1'b0));
assign n1084 = /* LUT    9 27  5 */ (n1058 ? (n1083 ? 1'b1 : !n861) : (n1083 ? n861 : 1'b0));
assign n583  = /* LUT    3 21  5 */ (n393 ? (n582 ? 1'b1 : !n324) : (n582 ? n324 : 1'b0));
assign n1208 = /* LUT   11 19  2 */ (n918 ? n1114 : n1206);
assign n2511 = /* LUT    4 18  2 */ \inMod[31] ;
assign n2512 = /* LUT   13 23  4 */ (n1393 ? (n1289 ? n1264 : !n1264) : (n1289 ? !n1264 : n1264));
assign n2513 = /* LUT    1 20  1 */ (n327 ? (n211 ? n232 : !n232) : (n211 ? !n232 : n232));
assign n2514 = /* LUT   15 23  3 */ (n1434 ? (n503 ? 1'b1 : (n49 ? !n142 : 1'b1)) : (n503 ? (n49 ? n142 : 1'b0) : 1'b0));
assign n2515 = /* LUT    6 16  0 */ (n543 ? 1'b1 : (n634 ? 1'b1 : (n444 ? 1'b1 : n728)));
assign n2516 = /* LUT    7 27  5 */ (n290 ? (n904 ? (reset ? 1'b1 : n254) : (reset ? 1'b0 : n254)) : n904);
assign n2517 = /* LUT   11 24  0 */ (n1262 ? (n1075 ? n901 : !n901) : (n1075 ? !n901 : n901));
assign n2518 = /* LUT   18 21  4 */ (n1489 ? 1'b1 : (n1462 ? 1'b1 : (n1453 ? 1'b1 : n1456)));
assign n2519 = /* LUT    4 26  7 */ (n613 ? (n253 ? n686 : 1'b1) : (n253 ? n686 : 1'b0));
assign n2520 = /* LUT    9 22  5 */ (n35 ? (n758 ? (n839 ? !n53 : 1'b1) : (n839 ? 1'b0 : n53)) : (n758 ? !n53 : 1'b0));
assign n2521 = /* LUT    4 23  4 */ (n590 ? (reset ? 1'b1 : (n253 ? n675 : 1'b1)) : (reset ? 1'b0 : (n253 ? n675 : 1'b0)));
assign n1046 = /* LUT    9 24  1 */ (n984 ? (n985 ? 1'b1 : n861) : (n985 ? !n861 : 1'b0));
assign n2522 = /* LUT   10 17  4 */ (\indata[27]  ? (n1100 ? (\inExp[0]  ? 1'b1 : !ready) : (\inExp[0]  ? ready : 1'b0)) : (n1100 ? !ready : 1'b0));
assign n2523 = /* LUT   12 21  3 */ (n1321 ? (n852 ? n1287 : !n1287) : (n852 ? !n1287 : n1287));
assign n2524 = /* LUT    5 18  3 */ (n466 ? (n157 ? !n106 : (n378 ? !n106 : 1'b0)) : (n157 ? 1'b0 : (n378 ? !n106 : 1'b0)));
assign n2525 = /* LUT    1 23  5 */ (n386 ? (n203 ? n320 : !n320) : (n203 ? !n320 : n320));
assign n2526 = /* LUT    2 22  2 */ (n484 ? (n178 ? n168 : !n168) : (n178 ? !n168 : n168));
assign n2527 = /* LUT   13 20  6 */ (n27 ? (n1308 ? !n839 : (n839 ? 1'b0 : n53)) : (n1308 ? (n839 ? 1'b0 : !n53) : 1'b0));
assign n2528 = /* LUT   10 27  0 */ (n1183 ? (n920 ? n344 : !n344) : (n920 ? !n344 : n344));
assign n2529 = /* LUT    3 24  0 */ !n590;
assign n2530 = /* LUT   11 22  3 */ (n1242 ? (n433 ? n1106 : !n1106) : (n433 ? !n1106 : n1106));
assign n2531 = /* LUT    7 20  1 */ (n864 ? (reset ? 1'b1 : (n290 ? n522 : 1'b1)) : (reset ? 1'b0 : (n290 ? n522 : 1'b0)));
assign n2532 = /* LUT    1 24  1 */ (n402 ? (n353 ? n222 : !n222) : (n353 ? !n222 : n222));
assign n2533 = /* LUT    5 26  6 */ (n798 ? (n274 ? n672 : !n672) : (n274 ? !n672 : n672));
assign n2534 = /* LUT   10 18  2 */ (n290 ? n973 : n1111);
assign n2535 = /* LUT   17 21  2 */ (n1453 ? (ds ? (\inExp[13]  ? 1'b1 : !ready) : 1'b1) : (ds ? (\inExp[13]  ? ready : 1'b0) : 1'b0));
assign n2536 = /* LUT    5 21  7 */ (n650 ? (ready ? !ds : n77) : 1'b0);
assign n2537 = /* LUT    1 18  5 */ (n297 ? (n171 ? n97 : !n97) : (n171 ? !n97 : n97));
assign n2538 = /* LUT    2 27  0 */ (n435 ? (reset ? 1'b1 : (n261 ? 1'b1 : !n253)) : (reset ? 1'b0 : (n261 ? n253 : 1'b0)));
assign n2539 = /* LUT   19 19  5 */ (n1450 ? (\inExp[10]  ? 1'b1 : (ready ? !ds : 1'b1)) : (\inExp[10]  ? (ready ? ds : 1'b0) : 1'b0));
assign n2540 = /* LUT    6 21  5 */ (n755 ? (ds ? (ready ? 1'b0 : n77) : (ready ? 1'b1 : n77)) : 1'b0);
assign n2541 = /* LUT    3 23  2 */ (n507 ? n595 : n505);
assign n2542 = /* LUT    5 14  6 */ (n627 ? (ready ? \indata[22]  : 1'b1) : (ready ? \indata[22]  : 1'b0));
assign n2543 = /* LUT    2 21  4 */ (n475 ? (n79 ? n152 : !n152) : (n79 ? !n152 : n152));
assign n2544 = /* LUT   11 21  7 */ (n1236 ? (n855 ? n1044 : !n1044) : (n855 ? !n1044 : n1044));
assign n2545 = /* LUT   12 20  4 */ (n1314 ? (n1021 ? n1110 : !n1110) : (n1021 ? !n1110 : n1110));
assign n2546 = /* LUT   12 18  0 */ (n1193 ? (reset ? 1'b1 : (n837 ? 1'b1 : !n290)) : (reset ? 1'b0 : (n837 ? n290 : 1'b0)));
assign n2547 = /* LUT    5 29  0 */ (n819 ? (n144 ? n523 : !n523) : (n144 ? !n523 : n523));
assign n2548 = /* LUT    3 25  7 */ (n434 ? (n77 ? (ds ? !ready : 1'b1) : (ds ? 1'b0 : ready)) : 1'b0);
assign n2549 = /* LUT   10 23  0 */ (n1143 ? (n979 ? n1142 : !n1142) : (n979 ? !n1142 : n1142));
assign n2550 = /* LUT    6 22  1 */ (n762 ? (reset ? 1'b1 : (n290 ? n467 : 1'b1)) : (reset ? 1'b0 : (n290 ? n467 : 1'b0)));
assign n2551 = /* LUT   11 26  3 */ (n1049 ? (n1065 ? 1'b1 : !n811) : (n1065 ? n811 : 1'b0));
assign n2552 = /* LUT   18 19  3 */ (n1465 ? (ready ? (ds ? \inExp[8]  : 1'b1) : 1'b1) : (ready ? (ds ? \inExp[8]  : 1'b0) : 1'b0));
assign n2553 = /* LUT    3 18  4 */ (n457 ? (n157 ? !n106 : (n243 ? !n106 : 1'b0)) : (n157 ? 1'b0 : (n243 ? !n106 : 1'b0)));
assign n2554 = /* LUT    7 19  6 */ (n290 ? (n553 ? (n856 ? 1'b1 : !reset) : (n856 ? reset : 1'b0)) : n856);
assign n2555 = /* LUT   12 25  6 */ (\indata[20]  ? (n1338 ? (\inExp[0]  ? 1'b1 : !ready) : (\inExp[0]  ? ready : 1'b0)) : (n1338 ? !ready : 1'b0));
assign n2556 = /* LUT    9 20  4 */ (n524 ? n668 : 1'b0);
assign n2557 = /* LUT    4 17  3 */ (n637 ? (n517 ? 1'b1 : (n50 ? !n49 : 1'b1)) : (n517 ? (n50 ? n49 : 1'b0) : 1'b0));
assign n2558 = /* LUT    7 30  5 */ \inMod[27] ;
assign n2559 = /* LUT    1 19  2 */ (n309 ? (n194 ? n125 : !n125) : (n194 ? !n125 : n125));
assign n2560 = /* LUT   12 23  6 */ (n1135 ? (n918 ? 1'b1 : n1224) : (n918 ? 1'b0 : n1224));
assign n2561 = /* LUT   13 24  5 */ (n1403 ? (n1355 ? n663 : !n663) : (n1355 ? !n663 : n663));
assign n2562 = /* LUT    1 21  2 */ (n134 ? (n301 ? !n106 : (n106 ? 1'b0 : !n157)) : (n301 ? (n106 ? 1'b0 : n157) : 1'b0));
assign n2563 = /* LUT   10 25  3 */ (n1165 ? (n906 ? n852 : !n852) : (n906 ? !n852 : n852));
assign n1183 = /* CARRY 10 26  7 */ (n781 & n1078) | ((n781 | n1078) & n1182);
assign n1374 = /* CARRY 13 21  5 */ (n1307 & n955) | ((n1307 | n955) & n1373);
assign n1255 = /* CARRY 11 23  0 */ (n1065 & n177) | ((n1065 | n177) & n1247);
assign n424  = /* CARRY  1 25  2 */ (n237 & n421) | ((n237 | n421) & n423);
assign n802  = /* CARRY  5 27  1 */ (n597 & n178) | ((n597 | n178) & n801);
assign n1333 = /* CARRY 12 22  5 */ (n1310 & n585) | ((n1310 | n585) & n1332);
assign n367  = /* CARRY  1 22  3 */ (n360 & n362) | ((n360 | n362) & n366);
assign n1155 = /* CARRY 10 24  0 */ (n850 & n1057) | ((n850 | n1057) & n1151);
assign n333  = /* CARRY  1 20  6 */ (n217 & n208) | ((n217 | n208) & n332);
assign n285  = /* CARRY  1 17  7 */ (n181 & n155) | ((n181 | n155) & n284);
assign n508  = /* CARRY  2 24  0 */ (n210 & n233) | ((n210 | n233) & n502);
assign n1384 = /* CARRY 13 22  4 */ (n974 & n1117) | ((n974 | n1117) & n1383);
assign n1296 = /* CARRY 12 19  0 */ (n979 & n1195) | ((n979 | n1195) & n1608);
assign n812  = /* CARRY  5 28  0 */ (n667 & n234) | ((n667 | n234) & n808);
assign n501  = /* CARRY  2 23  6 */ (n198 & n128) | ((n198 | n128) & n500);
assign n1393 = /* CARRY 13 23  3 */ (n1060 & n1286) | ((n1060 | n1286) & n1392);
assign n1268 = /* CARRY 11 24  1 */ (n981 & n1076) | ((n981 | n1076) & n1267);
assign n1323 = /* CARRY 12 21  4 */ (n849 & n1288) | ((n849 | n1288) & n1322);
assign n386  = /* CARRY  1 23  4 */ (n126 & n380) | ((n126 | n380) & n385);
assign n484  = /* CARRY  2 22  1 */ (n167 & n292) | ((n167 | n292) & n483);
assign n1240 = /* CARRY 11 22  0 */ (n1057 & n932) | ((n1057 | n932) & n1237);
assign n408  = /* CARRY  1 24  6 */ (n225 & n224) | ((n225 | n224) & n407);
assign n800  = /* CARRY  5 26  7 */ (n673 & n181) | ((n673 | n181) & n799);
assign n299  = /* CARRY  1 18  6 */ (n104 & n172) | ((n104 | n172) & n298);
assign n477  = /* CARRY  2 21  5 */ (n153 & n80) | ((n153 | n80) & n476);
assign n1236 = /* CARRY 11 21  6 */ (n1042 & n121) | ((n1042 | n121) & n1235);
assign n1314 = /* CARRY 12 20  3 */ (n1115 & n1095) | ((n1115 | n1095) & n1313);
assign n825  = /* CARRY  5 29  3 */ (n623 & n145) | ((n623 | n145) & n824);
assign n1145 = /* CARRY 10 23  1 */ (n1094 & n1041) | ((n1094 | n1041) & n1144);
assign n309  = /* CARRY  1 19  1 */ (n185 & n182) | ((n185 | n182) & n308);
assign n1401 = /* CARRY 13 24  2 */ (n1103 & n1249) | ((n1103 | n1249) & n1400);
assign n1163 = /* CARRY 10 25  0 */ (n767 & n1065) | ((n767 | n1065) & n1162);
assign n525  = /* CARRY  2 25  0 */ (n230 & n291) | ((n230 | n291) & n515);
assign n1182 = /* CARRY 10 26  6 */ (n737 & n1077) | ((n737 | n1077) & n1181);
assign n1373 = /* CARRY 13 21  4 */ (n1308 & n954) | ((n1308 | n954) & n1372);
assign n1258 = /* CARRY 11 23  3 */ (n906 & n734) | ((n906 | n734) & n1257);
assign n368  = /* CARRY  1 22  4 */ (n363 & n179) | ((n363 | n179) & n367);
assign n427  = /* CARRY  1 25  5 */ (n415 & n419) | ((n415 | n419) & n426);
assign n801  = /* CARRY  5 27  0 */ (n596 & n292) | ((n596 | n292) & n800);
assign n1332 = /* CARRY 12 22  4 */ (n1001 & n684) | ((n1001 | n684) & n1331);
assign n1158 = /* CARRY 10 24  3 */ (n1095 & n433) | ((n1095 | n433) & n1157);
assign n334  = /* CARRY  1 20  7 */ (n291 & n215) | ((n291 | n215) & n333);
assign n284  = /* CARRY  1 17  6 */ (n274 & n154) | ((n274 | n154) & n283);
assign n511  = /* CARRY  2 24  3 */ (n213 & n160) | ((n213 | n160) & n510);
assign n1385 = /* CARRY 13 22  5 */ (n967 & n996) | ((n967 | n996) & n1384);
assign n385  = /* CARRY  1 23  3 */ (n378 & n340) | ((n378 | n340) & n384);
assign n1297 = /* CARRY 12 19  1 */ (n1122 & n1094) | ((n1122 | n1094) & n1296);
assign n813  = /* CARRY  5 28  1 */ (n668 & n185) | ((n668 | n185) & n812);
assign n502  = /* CARRY  2 23  7 */ (n199 & n235) | ((n199 | n235) & n501);
assign n1392 = /* CARRY 13 23  2 */ (n1248 & n947) | ((n1248 | n947) & n1391);
assign n474  = /* CARRY  2 21  2 */ (n150 & n277) | ((n150 | n277) & n473);
assign n1269 = /* CARRY 11 24  2 */ (n900 & n893) | ((n900 | n893) & n1268);
assign n1324 = /* CARRY 12 21  5 */ (n957 & n890) | ((n957 | n890) & n1323);
assign n483  = /* CARRY  2 22  0 */ (n166 & n181) | ((n166 | n181) & n479);
assign n1241 = /* CARRY 11 22  1 */ (n970 & n850) | ((n970 | n850) & n1240);
assign n409  = /* CARRY  1 24  7 */ (n220 & n355) | ((n220 | n355) & n408);
assign n793  = /* CARRY  5 26  0 */ (n589 & n83) | ((n589 | n83) & n792);
assign n300  = /* CARRY  1 18  7 */ (n107 & n173) | ((n107 | n173) & n299);
assign n1235 = /* CARRY 11 21  5 */ (n1040 & n669) | ((n1040 | n669) & n1234);
assign n1313 = /* CARRY 12 20  2 */ (n1114 & n1106) | ((n1114 | n1106) & n1312);
assign n824  = /* CARRY  5 29  2 */ (n530 & n160) | ((n530 | n160) & n823);
assign n1146 = /* CARRY 10 23  2 */ (n853 & n745) | ((n853 | n745) & n1145);
assign n308  = /* CARRY  1 19  0 */ (n234 & n193) | ((n234 | n193) & n300);
assign n1402 = /* CARRY 13 24  3 */ (n1104 & n1253) | ((n1104 | n1253) & n1401);
assign n1164 = /* CARRY 10 25  1 */ (n1019 & n1066) | ((n1019 | n1066) & n1163);
assign n1181 = /* CARRY 10 26  5 */ (n585 & n779) | ((n585 | n779) & n1180);
assign n1376 = /* CARRY 13 21  7 */ (n1305 & n1294) | ((n1305 | n1294) & n1375);
assign n1257 = /* CARRY 11 23  2 */ (n1059 & n1019) | ((n1059 | n1019) & n1256);
assign n369  = /* CARRY  1 22  5 */ (n183 & n187) | ((n183 | n187) & n368);
assign n426  = /* CARRY  1 25  4 */ (n243 & n245) | ((n243 | n245) & n425);
assign n808  = /* CARRY  5 27  7 */ (n666 & n107) | ((n666 | n107) & n807);
assign n279  = /* CARRY  1 17  1 */ (n277 & n149) | ((n277 | n149) & n278);
assign n1302 = /* CARRY 12 19  6 */ (n866 & n855) | ((n866 | n855) & n1301);
assign n1335 = /* CARRY 12 22  7 */ (n1214 & n781) | ((n1214 | n781) & n1334);
assign n1407 = /* CARRY 13 25  0 */ (n1352 & n766) | ((n1352 | n766) & n1406);
assign n495  = /* CARRY  2 23  0 */ (n193 & n107) | ((n193 | n107) & n490);
assign n1157 = /* CARRY 10 24  2 */ (n1106 & n1045) | ((n1106 | n1045) & n1156);
assign n331  = /* CARRY  1 20  4 */ (n326 & n214) | ((n326 | n214) & n330);
assign n510  = /* CARRY  2 24  2 */ (n212 & n232) | ((n212 | n232) & n509);
assign n1386 = /* CARRY 13 22  6 */ (n758 & n999) | ((n758 | n999) & n1385);
assign n384  = /* CARRY  1 23  2 */ (n209 & n204) | ((n209 | n204) & n383);
assign n490  = /* CARRY  2 22  7 */ (n173 & n104) | ((n173 | n104) & n489);
assign n818  = /* CARRY  5 28  6 */ (n235 & n784) | ((n235 | n784) & n817);
assign n1246 = /* CARRY 11 22  6 */ (n593 & n785) | ((n593 | n785) & n1245);
assign n293  = /* CARRY  1 18  0 */ (n292 & n166) | ((n292 | n166) & n285);
assign n1391 = /* CARRY 13 23  1 */ (n1266 & n1121) | ((n1266 | n1121) & n1390);
assign n475  = /* CARRY  2 21  3 */ (n151 & n272) | ((n151 | n272) & n474);
assign n1270 = /* CARRY 11 24  3 */ (n1171 & n894) | ((n1171 | n894) & n1269);
assign n1325 = /* CARRY 12 21  6 */ (n1135 & n892) | ((n1135 | n892) & n1324);
assign n315  = /* CARRY  1 19  7 */ (n233 & n199) | ((n233 | n199) & n314);
assign n1169 = /* CARRY 10 25  6 */ (n892 & n1067) | ((n892 | n1067) & n1168);
assign n406  = /* CARRY  1 24  4 */ (n400 & n356) | ((n400 | n356) & n405);
assign n794  = /* CARRY  5 26  1 */ (n439 & n277) | ((n439 | n277) & n793);
assign n1234 = /* CARRY 11 21  4 */ (n1043 & n854) | ((n1043 | n854) & n1233);
assign n1312 = /* CARRY 12 20  1 */ (n1192 & n577) | ((n1192 | n577) & n1311);
assign n827  = /* CARRY  5 29  5 */ (n257 & n322) | ((n257 | n322) & n826);
assign n1260 = /* CARRY 11 23  5 */ (n849 & n1070) | ((n849 | n1070) & n1259);
assign n1147 = /* CARRY 10 23  3 */ (n854 & n1031) | ((n854 | n1031) & n1146);
assign n1399 = /* CARRY 13 24  0 */ (n1020 & n1336) | ((n1020 | n1336) & n1397);
assign n1180 = /* CARRY 10 26  4 */ (n684 & n1014) | ((n684 | n1014) & n1179);
assign n1375 = /* CARRY 13 21  6 */ (n1284 & n959) | ((n1284 | n959) & n1374);
assign n370  = /* CARRY  1 22  6 */ (n359 & n361) | ((n359 | n361) & n369);
assign n1160 = /* CARRY 10 24  5 */ (n593 & n972) | ((n593 | n972) & n1159);
assign n429  = /* CARRY  1 25  7 */ (n244 & n418) | ((n244 | n418) & n428);
assign n807  = /* CARRY  5 27  6 */ (n687 & n104) | ((n687 | n104) & n806);
assign n278  = /* CARRY  1 17  0 */ (n148 & n83) | ((n148 | n83) & n276);
assign n513  = /* CARRY  2 24  5 */ (n161 & n326) | ((n161 | n326) & n512);
assign n1303 = /* CARRY 12 19  7 */ (n1293 & n932) | ((n1293 | n932) & n1302);
assign n1334 = /* CARRY 12 22  6 */ (n1212 & n737) | ((n1212 | n737) & n1333);
assign n496  = /* CARRY  2 23  1 */ (n182 & n234) | ((n182 | n234) & n495);
assign n332  = /* CARRY  1 20  5 */ (n322 & n161) | ((n322 | n161) & n331);
assign n1387 = /* CARRY 13 22  7 */ (n1283 & n949) | ((n1283 | n949) & n1386);
assign n383  = /* CARRY  1 23  1 */ (n127 & n207) | ((n127 | n207) & n382);
assign n489  = /* CARRY  2 22  6 */ (n172 & n97) | ((n172 | n97) & n488);
assign n819  = /* CARRY  5 28  7 */ (n621 & n233) | ((n621 | n233) & n818);
assign n1247 = /* CARRY 11 22  7 */ (n786 & n763) | ((n786 | n763) & n1246);
assign n294  = /* CARRY  1 18  1 */ (n178 & n167) | ((n178 | n167) & n293);
assign n1390 = /* CARRY 13 23  0 */ (n1263 & n1251) | ((n1263 | n1251) & n1387);
assign n472  = /* CARRY  2 21  0 */ (n148 & n344) | ((n148 | n344) & n2011);
assign n1233 = /* CARRY 11 21  3 */ (n853 & n1031) | ((n853 | n1031) & n1232);
assign n1271 = /* CARRY 11 24  4 */ (n1014 & n905) | ((n1014 | n905) & n1270);
assign n1326 = /* CARRY 12 21  7 */ (n1136 & n901) | ((n1136 | n901) & n1325);
assign n314  = /* CARRY  1 19  6 */ (n235 & n198) | ((n235 | n198) & n313);
assign n1170 = /* CARRY 10 25  7 */ (n901 & n1069) | ((n901 | n1069) & n1169);
assign n407  = /* CARRY  1 24  5 */ (n223 & n218) | ((n223 | n218) & n406);
assign n795  = /* CARRY  5 26  2 */ (n676 & n272) | ((n676 | n272) & n794);
assign n1311 = /* CARRY 12 20  0 */ (n1285 & n850) | ((n1285 | n850) & n1303);
assign n1179 = /* CARRY 10 26  3 */ (n905 & n894) | ((n905 | n894) & n1178);
assign n1370 = /* CARRY 13 21  1 */ (n1306 & n1366) | ((n1306 | n1366) & n1369);
assign n826  = /* CARRY  5 29  4 */ (n624 & n326) | ((n624 | n326) & n825);
assign n1148 = /* CARRY 10 23  4 */ (n669 & n1043) | ((n669 | n1043) & n1147);
assign n1259 = /* CARRY 11 23  4 */ (n852 & n1068) | ((n852 | n1068) & n1258);
assign n1400 = /* CARRY 13 24  1 */ (n1102 & n1389) | ((n1102 | n1389) & n1399);
assign n1329 = /* CARRY 12 22  1 */ (n1141 & n900) | ((n1141 | n900) & n1328);
assign n371  = /* CARRY  1 22  7 */ (n323 & n189) | ((n323 | n189) & n370);
assign n1159 = /* CARRY 10 24  4 */ (n1021 & n1030) | ((n1021 | n1030) & n1158);
assign n428  = /* CARRY  1 25  6 */ (n250 & n246) | ((n250 | n246) & n427);
assign n806  = /* CARRY  5 27  5 */ (n773 & n97) | ((n773 | n97) & n805);
assign n281  = /* CARRY  1 17  3 */ (n79 & n151) | ((n79 | n151) & n280);
assign n512  = /* CARRY  2 24  4 */ (n214 & n145) | ((n214 | n145) & n511);
assign n1380 = /* CARRY 13 22  0 */ (n1304 & n1292) | ((n1304 | n1292) & n1376);
assign n1300 = /* CARRY 12 19  4 */ (n953 & n669) | ((n953 | n669) & n1299);
assign n497  = /* CARRY  2 23  2 */ (n194 & n185) | ((n194 | n185) & n496);
assign n1397 = /* CARRY 13 23  7 */ (n966 & n1378) | ((n966 | n1378) & n1396);
assign n329  = /* CARRY  1 20  2 */ (n160 & n212) | ((n160 | n212) & n328);
assign n1319 = /* CARRY 12 21  0 */ (n1119 & n767) | ((n1119 | n767) & n1318);
assign n382  = /* CARRY  1 23  0 */ (n205 & n201) | ((n205 | n201) & n371);
assign n488  = /* CARRY  2 22  5 */ (n171 & n102) | ((n171 | n102) & n487);
assign n816  = /* CARRY  5 28  4 */ (n605 & n247) | ((n605 | n247) & n815);
assign n1244 = /* CARRY 11 22  4 */ (n1095 & n1030) | ((n1095 | n1030) & n1243);
assign n404  = /* CARRY  1 24  2 */ (n399 & n216) | ((n399 | n216) & n403);
assign n295  = /* CARRY  1 18  2 */ (n103 & n168) | ((n103 | n168) & n294);
assign n473  = /* CARRY  2 21  1 */ (n149 & n83) | ((n149 | n83) & n472);
assign n1232 = /* CARRY 11 21  2 */ (n1094 & n745) | ((n1094 | n745) & n1231);
assign n1318 = /* CARRY 12 20  7 */ (n649 & n177) | ((n649 | n177) & n1317);
assign n1272 = /* CARRY 11 24  5 */ (n779 & n684) | ((n779 | n684) & n1271);
assign n313  = /* CARRY  1 19  5 */ (n128 & n197) | ((n128 | n197) & n312);
assign n1405 = /* CARRY 13 24  6 */ (n1086 & n1354) | ((n1086 | n1354) & n1404);
assign n1167 = /* CARRY 10 25  4 */ (n849 & n1068) | ((n849 | n1068) & n1166);
assign n796  = /* CARRY  5 26  3 */ (n79 & n534) | ((n79 | n534) & n795);
assign n1178 = /* CARRY 10 26  2 */ (n1171 & n893) | ((n1171 | n893) & n1177);
assign n1369 = /* CARRY 13 21  0 */ (n1254 & n1200) | ((n1254 | n1200) & n2188);
assign n829  = /* CARRY  5 29  7 */ (n256 & n291) | ((n256 | n291) & n828);
assign n1149 = /* CARRY 10 23  5 */ (n121 & n1040) | ((n121 | n1040) & n1148);
assign n1262 = /* CARRY 11 23  7 */ (n892 & n1069) | ((n892 | n1069) & n1261);
assign n423  = /* CARRY  1 25  1 */ (n158 & n420) | ((n158 | n420) & n422);
assign n1328 = /* CARRY 12 22  0 */ (n1327 & n981) | ((n1327 | n981) & n1326);
assign n364  = /* CARRY  1 22  0 */ (n188 & n357) | ((n188 | n357) & n2216);
assign n1162 = /* CARRY 10 24  7 */ (n177 & n786) | ((n177 | n786) & n1161);
assign n805  = /* CARRY  5 27  4 */ (n772 & n102) | ((n772 | n102) & n804);
assign n280  = /* CARRY  1 17  2 */ (n272 & n150) | ((n272 | n150) & n279);
assign n515  = /* CARRY  2 24  7 */ (n215 & n217) | ((n215 | n217) & n514);
assign n1381 = /* CARRY 13 22  1 */ (n1379 & n1107) | ((n1379 | n1107) & n1380);
assign n1301 = /* CARRY 12 19  5 */ (n952 & n121) | ((n952 | n121) & n1300);
assign n436  = /* CARRY  1 26  0 */ (n430 & n397) | ((n430 | n397) & n429);
assign n498  = /* CARRY  2 23  3 */ (n195 & n125) | ((n195 | n125) & n497);
assign n1396 = /* CARRY 13 23  6 */ (n1252 & n1377) | ((n1252 | n1377) & n1395);
assign n330  = /* CARRY  1 20  3 */ (n145 & n213) | ((n145 | n213) & n329);
assign n1320 = /* CARRY 12 21  1 */ (n1120 & n1019) | ((n1120 | n1019) & n1319);
assign n389  = /* CARRY  1 23  7 */ (n134 & n377) | ((n134 | n377) & n388);
assign n487  = /* CARRY  2 22  4 */ (n170 & n100) | ((n170 | n100) & n486);
assign n817  = /* CARRY  5 28  5 */ (n707 & n128) | ((n707 | n128) & n816);
assign n1245 = /* CARRY 11 22  5 */ (n1021 & n972) | ((n1021 | n972) & n1244);
assign n405  = /* CARRY  1 24  3 */ (n227 & n219) | ((n227 | n219) & n404);
assign n797  = /* CARRY  5 26  4 */ (n612 & n80) | ((n612 | n80) & n796);
assign n296  = /* CARRY  1 18  3 */ (n100 & n169) | ((n100 | n169) & n295);
assign n478  = /* CARRY  2 21  6 */ (n154 & n81) | ((n154 | n81) & n477);
assign n1231 = /* CARRY 11 21  1 */ (n979 & n1041) | ((n979 | n1041) & n1230);
assign n1317 = /* CARRY 12 20  6 */ (n998 & n763) | ((n998 | n763) & n1316);
assign n1273 = /* CARRY 11 24  6 */ (n1077 & n585) | ((n1077 | n585) & n1272);
assign n312  = /* CARRY  1 19  4 */ (n247 & n196) | ((n247 | n196) & n311);
assign n1406 = /* CARRY 13 24  7 */ (n1173 & n1348) | ((n1173 | n1348) & n1405);
assign n345  = /* CARRY  1 21  0 */ (n344 & n230) | ((n344 | n230) & n334);
assign n1168 = /* CARRY 10 25  5 */ (n890 & n1070) | ((n890 | n1070) & n1167);
assign n1177 = /* CARRY 10 26  1 */ (n900 & n1076) | ((n900 | n1076) & n1176);
assign n1372 = /* CARRY 13 21  3 */ (n1309 & n1368) | ((n1309 | n1368) & n1371);
assign n828  = /* CARRY  5 29  6 */ (n217 & n611) | ((n217 | n611) & n827);
assign n1150 = /* CARRY 10 23  6 */ (n855 & n1042) | ((n855 | n1042) & n1149);
assign n1261 = /* CARRY 11 23  6 */ (n890 & n1067) | ((n890 | n1067) & n1260);
assign n422  = /* CARRY  1 25  0 */ (n417 & n411) | ((n417 | n411) & n409);
assign n804  = /* CARRY  5 27  3 */ (n520 & n100) | ((n520 | n100) & n803);
assign n1331 = /* CARRY 12 22  3 */ (n1108 & n905) | ((n1108 | n905) & n1330);
assign n365  = /* CARRY  1 22  1 */ (n184 & n354) | ((n184 | n354) & n364);
assign n1161 = /* CARRY 10 24  6 */ (n763 & n785) | ((n763 | n785) & n1160);
assign n283  = /* CARRY  1 17  5 */ (n81 & n153) | ((n81 | n153) & n282);
assign n514  = /* CARRY  2 24  6 */ (n208 & n322) | ((n208 | n322) & n513);
assign n1382 = /* CARRY 13 22  2 */ (n865 & n1008) | ((n865 | n1008) & n1381);
assign n1298 = /* CARRY 12 19  2 */ (n1295 & n853) | ((n1295 | n853) & n1297);
assign n814  = /* CARRY  5 28  2 */ (n696 & n125) | ((n696 | n125) & n813);
assign n499  = /* CARRY  2 23  4 */ (n196 & n122) | ((n196 | n122) & n498);
assign n1395 = /* CARRY 13 23  5 */ (n1265 & n948) | ((n1265 | n948) & n1394);
assign n327  = /* CARRY  1 20  0 */ (n144 & n210) | ((n144 | n210) & n315);
assign n1321 = /* CARRY 12 21  2 */ (n917 & n734) | ((n917 | n734) & n1320);
assign n388  = /* CARRY  1 23  6 */ (n381 & n379) | ((n381 | n379) & n387);
assign n486  = /* CARRY  2 22  3 */ (n169 & n103) | ((n169 | n103) & n485);
assign n1242 = /* CARRY 11 22  2 */ (n1045 & n577) | ((n1045 | n577) & n1241);
assign n402  = /* CARRY  1 24  0 */ (n221 & n401) | ((n221 | n401) & n389);
assign n798  = /* CARRY  5 26  5 */ (n774 & n81) | ((n774 | n81) & n797);
assign n297  = /* CARRY  1 18  4 */ (n102 & n170) | ((n102 | n170) & n296);
assign n479  = /* CARRY  2 21  7 */ (n155 & n274) | ((n155 | n274) & n478);
assign n1230 = /* CARRY 11 21  0 */ (n344 & n1142) | ((n344 | n1142) & n2414);
assign n1316 = /* CARRY 12 20  5 */ (n997 & n593) | ((n997 | n593) & n1315);
assign n1274 = /* CARRY 11 24  7 */ (n1078 & n737) | ((n1078 | n737) & n1273);
assign n823  = /* CARRY  5 29  1 */ (n536 & n232) | ((n536 | n232) & n822);
assign n311  = /* CARRY  1 19  3 */ (n122 & n195) | ((n122 | n195) & n310);
assign n1403 = /* CARRY 13 24  4 */ (n968 & n1356) | ((n968 | n1356) & n1402);
assign n1165 = /* CARRY 10 25  2 */ (n734 & n1059) | ((n734 | n1059) & n1164);
assign n1278 = /* CARRY 11 25  0 */ (n920 & n781) | ((n920 | n781) & n1274);
assign n1371 = /* CARRY 13 21  2 */ (n857 & n1367) | ((n857 | n1367) & n1370);
assign n1176 = /* CARRY 10 26  0 */ (n981 & n1075) | ((n981 | n1075) & n1170);
assign n1151 = /* CARRY 10 23  7 */ (n932 & n1044) | ((n932 | n1044) & n1150);
assign n1256 = /* CARRY 11 23  1 */ (n1066 & n767) | ((n1066 | n767) & n1255);
assign n425  = /* CARRY  1 25  3 */ (n249 & n248) | ((n249 | n248) & n424);
assign n803  = /* CARRY  5 27  2 */ (n103 & n595) | ((n103 | n595) & n802);
assign n1330 = /* CARRY 12 22  2 */ (n1118 & n1171) | ((n1118 | n1171) & n1329);
assign n366  = /* CARRY  1 22  2 */ (n325 & n358) | ((n325 | n358) & n365);
assign n1156 = /* CARRY 10 24  1 */ (n577 & n970) | ((n577 | n970) & n1155);
assign n282  = /* CARRY  1 17  4 */ (n80 & n152) | ((n80 | n152) & n281);
assign n509  = /* CARRY  2 24  1 */ (n211 & n144) | ((n211 | n144) & n508);
assign n1383 = /* CARRY 13 22  3 */ (n1250 & n1116) | ((n1250 | n1116) & n1382);
assign n1299 = /* CARRY 12 19  3 */ (n867 & n854) | ((n867 | n854) & n1298);
assign n815  = /* CARRY  5 28  3 */ (n778 & n122) | ((n778 | n122) & n814);
assign n500  = /* CARRY  2 23  5 */ (n197 & n247) | ((n197 | n247) & n499);
assign n1394 = /* CARRY 13 23  4 */ (n1264 & n1289) | ((n1264 | n1289) & n1393);
assign n328  = /* CARRY  1 20  1 */ (n232 & n211) | ((n232 | n211) & n327);
assign n1267 = /* CARRY 11 24  0 */ (n901 & n1075) | ((n901 | n1075) & n1262);
assign n1322 = /* CARRY 12 21  3 */ (n1287 & n852) | ((n1287 | n852) & n1321);
assign n387  = /* CARRY  1 23  5 */ (n320 & n203) | ((n320 | n203) & n386);
assign n485  = /* CARRY  2 22  2 */ (n168 & n178) | ((n168 | n178) & n484);
assign n1184 = /* CARRY 10 27  0 */ (n344 & n920) | ((n344 | n920) & n1183);
assign n1243 = /* CARRY 11 22  3 */ (n1106 & n433) | ((n1106 | n433) & n1242);
assign n403  = /* CARRY  1 24  1 */ (n222 & n353) | ((n222 | n353) & n402);
assign n799  = /* CARRY  5 26  6 */ (n672 & n274) | ((n672 | n274) & n798);
assign n298  = /* CARRY  1 18  5 */ (n97 & n171) | ((n97 | n171) & n297);
assign n476  = /* CARRY  2 21  4 */ (n152 & n79) | ((n152 | n79) & n475);
assign n1237 = /* CARRY 11 21  7 */ (n1044 & n855) | ((n1044 | n855) & n1236);
assign n1315 = /* CARRY 12 20  4 */ (n1110 & n1021) | ((n1110 | n1021) & n1314);
assign n822  = /* CARRY  5 29  0 */ (n523 & n144) | ((n523 | n144) & n819);
assign n1144 = /* CARRY 10 23  0 */ (n1142 & n979) | ((n1142 | n979) & n1143);
assign n310  = /* CARRY  1 19  2 */ (n125 & n194) | ((n125 | n194) & n309);
assign n1404 = /* CARRY 13 24  5 */ (n663 & n1355) | ((n663 | n1355) & n1403);
assign n1166 = /* CARRY 10 25  3 */ (n852 & n906) | ((n852 | n906) & n1165);
/* FF  6 19  1 */ always @(posedge clk, posedge reset) if (reset) n665 <= 1'b0; else if (n226) n665 <= n1542;
/* FF  7 24  4 */ assign n1543 = n938;
/* FF 18 20  7 */ assign n1472 = n1544;
/* FF  4 25  6 */ always @(posedge clk, posedge reset) if (reset) n239 <= 1'b0; else if (n82) n239 <= n1545;
/* FF  9 23  2 */ always @(posedge clk, posedge reset) if (reset) n965 <= 1'b0; else if (n226) n965 <= n1546;
/* FF  7 22  0 */ assign n106 = n922;
/* FF 10 22  7 */ assign n1021 = n1547;
/* FF  4 22  7 */ assign n125 = n1548;
/* FF 14 21  2 */ assign n1549 = n1426;
/* FF  5 24  5 */ always @(posedge clk) if (n157) n676 <= 1'b0 ? 1'b0 : n1550;
/* FF 10 16  7 */ always @(posedge clk, posedge reset) if (reset) n202 <= 1'b0; else if (n226) n202 <= n1551;
/* FF  5 19  4 */ always @(posedge clk, posedge reset) if (reset) n569 <= 1'b0; else if (n82) n569 <= n1552;
/* FF  2 25  3 */ assign n411 = n1553;
/* FF 10 26  7 */ assign n1064 = n1554;
/* FF 11 17  4 */ always @(posedge clk, posedge reset) if (reset) n837 <= 1'b0; else if (n51) n837 <= n1555;
/* FF 13 21  5 */ assign n1040 = n1556;
/* FF  2 19  3 */ assign n1557 = n460;
/* FF 11 23  0 */ assign n1137 = n1558;
/* FF  4 30  0 */ always @(posedge clk, posedge reset) if (reset) n262 <= 1'b0; else if (n51) n262 <= n1559;
/* FF  5 17  5 */ assign n326 = n1560;
/* FF  1 25  2 */ assign n212 = n1561;
/* FF 15 21  5 */ always @(posedge clk) if (n157) n1416 <= 1'b0 ? 1'b0 : n1562;
/* FF 10 21  3 */ assign n15 = n1133;
/* FF  6 18  6 */ always @(posedge clk) if (1'b1) n741 <= 1'b0 ? 1'b0 : n1563;
/* FF  5 27  1 */ assign n697 = n1564;
/* FF  5 22  6 */ assign n1565 = n771;
/* FF 14 22  0 */ assign n1377 = n1566;
/* FF  2 26  7 */ assign n421 = n1567;
/* FF  6 20  6 */ always @(posedge clk, posedge reset) if (reset) n744 <= 1'b0; else if (n226) n744 <= n1568;
/* FF  3 20  3 */ assign n1569 = n572;
/* FF  2 20  7 */ assign n319 = n1570;
/* FF  6 25  5 */ assign n224 = n1571;
/* FF 11 18  6 */ assign n1107 = n1572;
/* FF 12 27  5 */ assign n31 = n1344;
/* FF 14 19  2 */ always @(posedge clk) if (n53) n1353 <= n839 ? 1'b0 : n1573;
/* FF  5 30  1 */ assign n721 = n1574;
/* FF  3 22  6 */ always @(posedge clk) if (1'b1) n481 <= 1'b0 ? 1'b0 : n1575;
/* FF 13 16  0 */ always @(posedge clk) if (1'b1) n1283 <= 1'b0 ? 1'b0 : n1576;
/* FF 11 27  0 */ assign n109 = n1577;
/* FF  9 19  7 */ always @(posedge clk) if (n53) n866 <= 1'b0 ? 1'b0 : n1578;
/* FF  7 26  7 */ assign n781 = n1579;
/* FF  4 27  5 */ always @(posedge clk, posedge reset) if (reset) n537 <= 1'b0; else if (n82) n537 <= n1580;
/* FF  9 21  7 */ always @(posedge clk, posedge reset) if (reset) n416 <= 1'b0; else if (n226) n416 <= n1581;
/* FF  7 16  7 */ assign n53 = n1582;
/* FF  4 16  4 */ always @(posedge clk) if (n53) n544 <= 1'b0 ? 1'b0 : n1583;
/* FF  5 23  1 */ always @(posedge clk) if (n157) n200 <= 1'b0 ? 1'b0 : n1584;
/* FF 12 22  5 */ assign n1239 = n1585;
/* FF  1 22  3 */ assign n151 = n1586;
/* FF 13 19  6 */ assign n1294 = n1587;
/* FF 10 24  0 */ assign n1022 = n1588;
/* FF  3 27  0 */ assign n128 = n1589;
/* FF  7 25  3 */ always @(posedge clk) if (1'b1) n237 <= 1'b0 ? 1'b0 : n1590;
/* FF  4 18  5 */ always @(posedge clk, posedge reset) if (reset) n522 <= 1'b0; else if (n51) n522 <= n1591;
/* FF  7 23  3 */ always @(posedge clk, posedge reset) if (reset) n606 <= 1'b0; else if (n226) n606 <= n1592;
/* FF 14 18  5 */ always @(posedge clk) if (n53) n1212 <= 1'b0 ? 1'b0 : n1593;
/* FF  1 20  6 */ assign n119 = n1594;
/* FF  4 24  1 */ assign n1595 = n680;
/* FF  4 21  6 */ assign n576 = n1596;
/* FF 14 20  1 */ always @(posedge clk) if (n157) n1361 <= 1'b0 ? 1'b0 : n1597;
/* FF  5 25  6 */ assign n683 = n1598;
/* FF  5 20  5 */ always @(posedge clk, posedge reset) if (reset) n655 <= 1'b0; else if (n82) n655 <= n1599;
/* FF  1 17  7 */ assign n64 = n1600;
/* FF  2 24  0 */ assign n390 = n1601;
/* FF 13 22  4 */ assign n1030 = n1602;
/* FF 16 23  6 */ always @(posedge clk) if (n157) n1442 <= 1'b0 ? 1'b0 : n1603;
/* FF  2 18  4 */ assign n287 = n1604;
/* FF 11 20  1 */ assign n1605 = n1218;
/* FF  5 18  4 */ assign n100 = n1606;
/* FF 12 19  0 */ assign n1200 = n1607;
/* FF  5 28  0 */ assign n708 = n1609;
/* FF 10 20  0 */ always @(posedge clk, posedge reset) if (reset) n1006 <= 1'b0; else if (n226) n1006 <= n1610;
/* FF  6 23  7 */ always @(posedge clk) if (n157) n687 <= 1'b0 ? 1'b0 : n1611;
/* FF  3 21  4 */ assign n1612 = n582;
/* FF  4 20  1 */ always @(posedge clk) if (1'b1) n140 <= 1'b0 ? 1'b0 : n1613;
/* FF  2 23  6 */ assign n352 = n1614;
/* FF  6 24  6 */ assign n1615 = n889;
/* FF 16 25  3 */ always @(posedge clk, posedge reset) if (reset) n674 <= 1'b0; else if (n226) n674 <= n1616;
/* FF  9 27  4 */ assign n1617 = n1083;
/* FF 11 19  5 */ assign n1618 = n1209;
/* FF 17 21  5 */ always @(posedge clk, posedge reset) if (reset) n1455 <= 1'b0; else if (n1408) n1455 <= n1619;
/* FF 13 23  3 */ assign n906 = n1620;
/* FF  3 23  5 */ always @(posedge clk) if (n157) n493 <= n106 ? 1'b0 : n1621;
/* FF 15 23  2 */ always @(posedge clk) if (n157) n1425 <= 1'b0 ? 1'b0 : n1622;
/* FF  6 16  3 */ always @(posedge clk) if (n53) n728 <= 1'b0 ? 1'b0 : n1623;
/* FF  4 28  6 */ assign n529 = n1624;
/* FF 11 24  1 */ assign n1130 = n1625;
/* FF  9 22  6 */ always @(posedge clk) if (1'b1) n969 <= 1'b0 ? 1'b0 : n1626;
/* FF  4 23  5 */ always @(posedge clk) if (1'b1) n591 <= 1'b0 ? 1'b0 : n1627;
/* FF  7 15  4 */ assign n835 = n1628;
/* FF  9 24  6 */ always @(posedge clk, posedge reset) if (reset) n976 <= 1'b0; else if (n226) n976 <= n1629;
/* FF 10 17  5 */ always @(posedge clk, posedge reset) if (reset) n535 <= 1'b0; else if (n226) n535 <= n1630;
/* FF 12 21  4 */ assign n1134 = n1631;
/* FF 18 19  4 */ always @(posedge clk, posedge reset) if (reset) n1465 <= 1'b0; else if (n1408) n1465 <= n1632;
/* FF  1 23  4 */ assign n170 = n1633;
/* FF  2 22  1 */ assign n346 = n1634;
/* FF 13 20  7 */ always @(posedge clk) if (1'b1) n1309 <= 1'b0 ? 1'b0 : n1635;
/* FF 10 27  1 */ assign n811 = n1185;
/* FF 19 20  2 */ assign n1636 = n1507;
/* FF  3 24  1 */ always @(posedge clk) if (1'b1) n220 <= 1'b0 ? 1'b0 : n1637;
/* FF  7 30  2 */ always @(posedge clk, posedge reset) if (reset) n907 <= 1'b0; else if (n51) n907 <= n1638;
/* FF 11 22  0 */ assign n1123 = n1639;
/* FF  7 20  2 */ always @(posedge clk) if (1'b1) n663 <= 1'b0 ? 1'b0 : n1640;
/* FF  9 17  0 */ always @(posedge clk, posedge reset) if (reset) n945 <= 1'b0; else if (n226) n945 <= n1641;
/* FF  5 16  7 */ always @(posedge clk) if (n53) n633 <= 1'b0 ? 1'b0 : n1642;
/* FF  1 21  5 */ assign n136 = n1643;
/* FF  1 24  6 */ assign n198 = n1644;
/* FF  5 26  7 */ assign n599 = n1645;
/* FF 10 18  1 */ assign n1646 = n1111;
/* FF 14 23  0 */ assign n1388 = n1647;
/* FF  5 21  6 */ always @(posedge clk, posedge reset) if (reset) n660 <= 1'b0; else if (n82) n660 <= n1648;
/* FF  1 18  6 */ assign n75 = n1649;
/* FF 19 19  4 */ always @(posedge clk, posedge reset) if (reset) n1487 <= 1'b0; else if (n1408) n1487 <= n1650;
/* FF  6 21  2 */ assign n755 = n1651;
/* FF 16 22  5 */ assign n1652 = n1459;
/* FF  2 21  5 */ assign n159 = n1653;
/* FF 11 21  6 */ assign n1090 = n1654;
/* FF 12 20  3 */ assign n1207 = n1655;
/* FF  5 19  3 */ always @(posedge clk, posedge reset) if (reset) n645 <= 1'b0; else if (n82) n645 <= n1656;
/* FF 12 18  3 */ assign n1657 = n1291;
/* FF  5 29  3 */ assign n716 = n1658;
/* FF  3 25  6 */ always @(posedge clk, posedge reset) if (reset) n517 <= 1'b0; else if (n82) n517 <= n1659;
/* FF  2 19  4 */ assign n302 = n1660;
/* FF  6 28  4 */ assign n809 = n1661;
/* FF 10 23  1 */ assign n1025 = n1662;
/* FF  6 22  0 */ assign n187 = n1663;
/* FF  7 21  5 */ assign n873 = n1664;
/* FF  3 18  5 */ assign n80 = n1665;
/* FF  7 19  1 */ assign n853 = n1666;
/* FF  9 20  5 */ assign n356 = n1667;
/* FF  1 19  1 */ assign n88 = n1668;
/* FF 12 23  7 */ assign n1253 = n1669;
/* FF 13 24  2 */ assign n893 = n1670;
/* FF  3 20  4 */ assign n146 = n1671;
/* FF 19 22  1 */ always @(posedge clk, posedge reset) if (reset) n1499 <= 1'b0; else if (n1408) n1499 <= n1672;
/* FF  6 25  2 */ assign n218 = n1673;
/* FF 13 18  2 */ always @(posedge clk) if (n53) n1287 <= 1'b0 ? 1'b0 : n1674;
/* FF 10 25  0 */ assign n1049 = n1675;
/* FF  6 19  2 */ always @(posedge clk, posedge reset) if (reset) n742 <= 1'b0; else if (n226) n742 <= n1676;
/* FF  3 26  0 */ always @(posedge clk, posedge reset) if (reset) n526 <= 1'b0; else if (n226) n526 <= n1677;
/* FF  7 24  5 */ assign n44 = n939;
/* FF 18 20  6 */ always @(posedge clk, posedge reset) if (reset) n1471 <= 1'b0; else if (n1408) n1471 <= n1678;
/* FF  4 19  7 */ always @(posedge clk) if (1'b1) n320 <= 1'b0 ? 1'b0 : n1679;
/* FF  4 25  7 */ always @(posedge clk, posedge reset) if (reset) n603 <= 1'b0; else if (n82) n603 <= n1680;
/* FF  9 23  1 */ assign n21 = n1036;
/* FF 10 22  6 */ always @(posedge clk) if (1'b1) n974 <= 1'b0 ? 1'b0 : n1681;
/* FF  7 22  1 */ always @(posedge clk) if (1'b1) n360 <= 1'b0 ? 1'b0 : n1682;
/* FF  4 22  6 */ always @(posedge clk) if (1'b1) n586 <= 1'b0 ? 1'b0 : n1683;
/* FF 14 21  3 */ always @(posedge clk) if (n53) n1295 <= 1'b0 ? 1'b0 : n1684;
/* FF  5 24  2 */ assign n354 = n1685;
/* FF  2 25  0 */ assign n410 = n1686;
/* FF 10 26  6 */ assign n1063 = n1687;
/* FF 11 17  3 */ always @(posedge clk, posedge reset) if (reset) n190 <= 1'b0; else if (n51) n190 <= n1688;
/* FF 13 21  4 */ assign n1043 = n1689;
/* FF 19 21  5 */ assign n1496 = n1690;
/* FF  4 16  3 */ always @(posedge clk) if (n53) n543 <= 1'b0 ? 1'b0 : n1691;
/* FF 11 23  3 */ assign n1058 = n1692;
/* FF  4 30  3 */ always @(posedge clk, posedge reset) if (reset) n600 <= 1'b0; else if (n51) n600 <= n1693;
/* FF  1 22  4 */ assign n152 = n1694;
/* FF  1 25  5 */ assign n161 = n1695;
/* FF 15 21  4 */ always @(posedge clk) if (n157) n1422 <= 1'b0 ? 1'b0 : n1696;
/* FF 14 22  7 */ always @(posedge clk) if (n53) n1327 <= 1'b0 ? 1'b0 : n1697;
/* FF  5 27  0 */ assign n519 = n1698;
/* FF 10 21  0 */ assign n1699 = n1131;
/* FF  5 22  7 */ always @(posedge clk) if (n157) n668 <= 1'b0 ? 1'b0 : n1700;
/* FF  6 20  1 */ assign n162 = n871;
/* FF 11 18  7 */ assign n1095 = n1701;
/* FF 12 27  2 */ always @(posedge clk, posedge reset) if (reset) n1211 <= 1'b0; else if (n226) n1211 <= n1702;
/* FF  5 20  2 */ assign n653 = n753;
/* FF 14 19  3 */ assign n1348 = n1703;
/* FF  3 22  7 */ always @(posedge clk) if (1'b1) n482 <= 1'b0 ? 1'b0 : n1704;
/* FF  2 18  3 */ assign n1705 = n451;
/* FF 13 16  1 */ always @(posedge clk) if (1'b1) n1284 <= 1'b0 ? 1'b0 : n1706;
/* FF  3 28  7 */ always @(posedge clk) if (n157) n530 <= 1'b0 ? 1'b0 : n1707;
/* FF 11 27  3 */ assign n3 = n1708;
/* FF  6 17  1 */ assign n734 = n1709;
/* FF  7 26  4 */ assign n900 = n1710;
/* FF  3 19  6 */ assign n82 = n1711;
/* FF  9 19  6 */ assign n1712 = n1005;
/* FF  7 16  0 */ always @(posedge clk) if (n53) n551 <= 1'b0 ? 1'b0 : n1713;
/* FF 12 24  0 */ always @(posedge clk) if (1'b1) n1263 <= 1'b0 ? 1'b0 : n1714;
/* FF  9 21  6 */ always @(posedge clk, posedge reset) if (reset) n960 <= 1'b0; else if (n226) n960 <= n1715;
/* FF  5 23  0 */ always @(posedge clk) if (n157) n396 <= 1'b0 ? 1'b0 : n1716;
/* FF 12 22  4 */ assign n1215 = n1717;
/* FF 13 25  1 */ assign n1085 = n1718;
/* FF  3 21  3 */ always @(posedge clk, posedge reset) if (reset) n470 <= 1'b0; else if (n82) n470 <= n1719;
/* FF 13 19  5 */ always @(posedge clk) if (n53) n1293 <= 1'b0 ? 1'b0 : n1720;
/* FF 10 24  3 */ assign n887 = n1721;
/* FF  3 27  3 */ assign n107 = n1722;
/* FF  4 18  4 */ always @(posedge clk, posedge reset) if (reset) n556 <= 1'b0; else if (n51) n556 <= n1723;
/* FF  7 23  2 */ always @(posedge clk, posedge reset) if (reset) n881 <= 1'b0; else if (n226) n881 <= n1724;
/* FF  4 24  0 */ assign n189 = n1725;
/* FF  1 20  7 */ assign n120 = n1726;
/* FF 14 18  4 */ assign n1727 = n1410;
/* FF  4 21  7 */ always @(posedge clk) if (1'b1) n415 <= 1'b0 ? 1'b0 : n1728;
/* FF 14 20  0 */ assign n1360 = n1729;
/* FF  5 25  1 */ assign n682 = n1730;
/* FF 10 19  7 */ always @(posedge clk) if (n53) n732 <= 1'b0 ? 1'b0 : n1731;
/* FF  9 26  4 */ assign n1732 = n1073;
/* FF  1 17  6 */ assign n63 = n1733;
/* FF  2 24  3 */ assign n392 = n1734;
/* FF 13 22  5 */ assign n972 = n1735;
/* FF  4 23  2 */ assign n377 = n1736;
/* FF 11 20  2 */ always @(posedge clk) if (n53) n1119 <= 1'b0 ? 1'b0 : n1737;
/* FF  5 18  5 */ always @(posedge clk) if (1'b1) n640 <= 1'b0 ? 1'b0 : n1738;
/* FF  1 23  3 */ assign n169 = n1739;
/* FF 12 19  1 */ assign n1201 = n1740;
/* FF  1 26  4 */ assign n233 = n1741;
/* FF  5 28  1 */ assign n709 = n1742;
/* FF 10 20  3 */ assign n54 = n1127;
/* FF  6 23  0 */ always @(posedge clk) if (n157) n772 <= 1'b0 ? 1'b0 : n1743;
/* FF  4 20  0 */ always @(posedge clk) if (1'b1) n565 <= 1'b0 ? 1'b0 : n1744;
/* FF  2 23  7 */ assign n375 = n1745;
/* FF  7 18  3 */ assign n669 = n1746;
/* FF  9 27  3 */ always @(posedge clk, posedge reset) if (reset) n782 <= 1'b0; else if (n226) n782 <= n1747;
/* FF 11 19  4 */ assign n1116 = n1748;
/* FF 17 21  4 */ always @(posedge clk, posedge reset) if (reset) n1454 <= 1'b0; else if (n1408) n1454 <= n1749;
/* FF  5 21  1 */ assign n1750 = n759;
/* FF 13 23  2 */ assign n1059 = n1751;
/* FF  2 21  2 */ assign n336 = n1752;
/* FF 15 23  5 */ always @(posedge clk) if (n157) n1435 <= 1'b0 ? 1'b0 : n1753;
/* FF  4 28  5 */ assign n615 = n1754;
/* FF 11 24  2 */ assign n1096 = n1755;
/* FF  4 26  1 */ assign n1756 = n700;
/* FF  9 24  7 */ always @(posedge clk, posedge reset) if (reset) n686 <= 1'b0; else if (n226) n686 <= n1757;
/* FF 10 17  2 */ assign n1758 = n1099;
/* FF 12 21  5 */ assign n1223 = n1759;
/* FF  3 18  2 */ always @(posedge clk) if (1'b1) n325 <= 1'b0 ? 1'b0 : n1760;
/* FF  2 22  0 */ assign n307 = n1761;
/* FF 13 20  4 */ always @(posedge clk) if (1'b1) n1306 <= 1'b0 ? 1'b0 : n1762;
/* FF 10 27  2 */ assign n870 = n1763;
/* FF 19 20  3 */ assign n1764 = n1508;
/* FF  3 24  2 */ always @(posedge clk) if (1'b1) n221 <= 1'b0 ? 1'b0 : n1765;
/* FF  4 17  5 */ always @(posedge clk) if (n53) n548 <= 1'b0 ? 1'b0 : n1766;
/* FF  7 30  3 */ always @(posedge clk, posedge reset) if (reset) n261 <= 1'b0; else if (n51) n261 <= n1767;
/* FF 11 22  1 */ assign n962 = n1768;
/* FF  5 16  4 */ always @(posedge clk) if (n53) n631 <= 1'b0 ? 1'b0 : n1769;
/* FF 19 22  6 */ always @(posedge clk, posedge reset) if (reset) n1443 <= 1'b0; else if (n1408) n1443 <= n1770;
/* FF  1 24  7 */ assign n199 = n1771;
/* FF  5 26  0 */ assign n692 = n1772;
/* FF 10 18  0 */ assign n996 = n1773;
/* FF 14 23  1 */ assign n1774 = n1437;
/* FF 18 20  1 */ always @(posedge clk, posedge reset) if (reset) n1466 <= 1'b0; else if (n1408) n1466 <= n1775;
/* FF  1 18  7 */ assign n76 = n1776;
/* FF  6 21  3 */ assign n756 = n875;
/* FF  4 22  1 */ assign n226 = n1777;
/* FF 11 21  5 */ assign n1091 = n1778;
/* FF 12 20  2 */ assign n1206 = n1779;
/* FF  5 19  2 */ assign n644 = n747;
/* FF  6 26  7 */ assign n145 = n1780;
/* FF 12 18  2 */ assign n979 = n1290;
/* FF  5 29  2 */ assign n715 = n1781;
/* FF  3 25  5 */ assign n516 = n609;
/* FF  2 19  5 */ assign n303 = n461;
/* FF 10 23  2 */ assign n859 = n1782;
/* FF  6 22  7 */ assign n593 = n1783;
/* FF  7 19  0 */ assign n852 = n1784;
/* FF  9 20  2 */ assign n340 = n1785;
/* FF  1 19  0 */ assign n87 = n1786;
/* FF 12 23  4 */ assign n1251 = n1787;
/* FF 13 24  3 */ assign n894 = n1788;
/* FF  3 20  5 */ assign n464 = n573;
/* FF 13 18  3 */ assign n1789 = n1350;
/* FF 10 25  1 */ assign n1050 = n1790;
/* FF 15 20  4 */ always @(posedge clk) if (n157) n1412 <= 1'b0 ? 1'b0 : n1791;
/* FF  6 19  3 */ always @(posedge clk, posedge reset) if (reset) n175 <= 1'b0; else if (n226) n175 <= n1792;
/* FF  7 24  6 */ always @(posedge clk, posedge reset) if (reset) n883 <= 1'b0; else if (n226) n883 <= n1793;
/* FF  4 19  4 */ assign n181 = n1794;
/* FF  4 25  0 */ assign n1795 = n688;
/* FF  7 22  6 */ always @(posedge clk) if (1'b1) n179 <= 1'b0 ? 1'b0 : n1796;
/* FF 10 22  5 */ assign n344 = n1797;
/* FF  9 23  0 */ assign n1798 = n1035;
/* FF 14 21  0 */ always @(posedge clk) if (n53) n1122 <= 1'b0 ? 1'b0 : n1799;
/* FF  5 24  3 */ always @(posedge clk) if (n157) n439 <= 1'b0 ? 1'b0 : n1800;
/* FF 10 16  1 */ assign n2 = n1801;
/* FF  9 25  4 */ assign n767 = n1802;
/* FF  3 19  1 */ assign n453 = n562;
/* FF  2 25  1 */ assign n324 = n1803;
/* FF 10 26  5 */ assign n927 = n1804;
/* FF 11 17  2 */ always @(posedge clk, posedge reset) if (reset) n594 <= 1'b0; else if (n51) n594 <= n1805;
/* FF 13 21  7 */ assign n1044 = n1806;
/* FF  4 16  2 */ always @(posedge clk) if (n53) n65 <= 1'b0 ? 1'b0 : n1807;
/* FF  5 23  7 */ always @(posedge clk) if (n157) n673 <= 1'b0 ? 1'b0 : n1808;
/* FF 11 23  2 */ assign n978 = n1809;
/* FF  4 30  2 */ always @(posedge clk, posedge reset) if (reset) n98 <= 1'b0; else if (n51) n98 <= n1810;
/* FF  5 17  7 */ assign n217 = n1811;
/* FF  1 22  5 */ assign n153 = n1812;
/* FF  1 25  4 */ assign n214 = n1813;
/* FF 15 21  3 */ always @(posedge clk) if (n157) n1421 <= 1'b0 ? 1'b0 : n1814;
/* FF 10 21  1 */ assign n13 = n1815;
/* FF  6 18  4 */ always @(posedge clk) if (1'b1) n740 <= 1'b0 ? 1'b0 : n1816;
/* FF  5 27  7 */ assign n705 = n1817;
/* FF 14 22  6 */ assign n1818 = n1431;
/* FF  2 26  5 */ assign n418 = n1819;
/* FF 11 28  0 */ always @(posedge clk, posedge reset) if (reset) n671 <= 1'b0; else if (n51) n671 <= n1820;
/* FF  4 21  0 */ assign n292 = n1821;
/* FF 11 18  4 */ always @(posedge clk) if (1'b1) n1105 <= 1'b0 ? 1'b0 : n1822;
/* FF  5 20  3 */ always @(posedge clk, posedge reset) if (reset) n654 <= 1'b0; else if (n82) n654 <= n1823;
/* FF  1 17  1 */ assign n58 = n1824;
/* FF 14 19  4 */ assign n1354 = n1825;
/* FF  5 30  3 */ assign n720 = n1826;
/* FF  3 22  4 */ always @(posedge clk) if (1'b1) n480 <= 1'b0 ? 1'b0 : n1827;
/* FF 11 27  2 */ assign n1828 = n1280;
/* FF  3 15  7 */ always @(posedge clk) if (n53) n444 <= 1'b0 ? 1'b0 : n1829;
/* FF  9 19  5 */ assign n955 = n1830;
/* FF 12 19  6 */ assign n1203 = n1831;
/* FF  7 26  5 */ assign n901 = n1832;
/* FF  7 16  1 */ always @(posedge clk) if (n53) n447 <= 1'b0 ? 1'b0 : n1833;
/* FF 12 24  7 */ always @(posedge clk) if (1'b1) n1266 <= 1'b0 ? 1'b0 : n1834;
/* FF  9 21  1 */ assign n67 = n1835;
/* FF 12 22  7 */ assign n1029 = n1836;
/* FF 13 25  0 */ assign n920 = n1837;
/* FF  6 24  0 */ always @(posedge clk) if (n157) n696 <= 1'b0 ? 1'b0 : n1838;
/* FF  4 20  7 */ always @(posedge clk) if (1'b1) n250 <= 1'b0 ? 1'b0 : n1839;
/* FF  2 23  0 */ assign n372 = n1840;
/* FF  3 21  2 */ assign n469 = n581;
/* FF 13 19  4 */ assign n1841 = n1359;
/* FF 10 24  2 */ assign n1039 = n1842;
/* FF  4 18  7 */ always @(posedge clk, posedge reset) if (reset) n553 <= 1'b0; else if (n51) n553 <= n1843;
/* FF  7 23  5 */ assign n129 = n931;
/* FF  4 24  7 */ always @(posedge clk) if (n157) n520 <= 1'b0 ? 1'b0 : n1844;
/* FF  1 20  4 */ assign n117 = n1845;
/* FF 14 18  3 */ always @(posedge clk) if (n53) n1310 <= 1'b0 ? 1'b0 : n1846;
/* FF 14 20  3 */ always @(posedge clk) if (n157) n1362 <= 1'b0 ? 1'b0 : n1847;
/* FF  9 26  5 */ assign n36 = n1074;
/* FF 10 19  0 */ always @(posedge clk) if (n53) n52 <= 1'b0 ? 1'b0 : n1848;
/* FF  5 25  0 */ assign n291 = n1849;
/* FF  2 24  2 */ assign n391 = n1850;
/* FF 13 22  6 */ assign n785 = n1851;
/* FF 16 23  4 */ always @(posedge clk) if (n157) n1446 <= 1'b0 ? 1'b0 : n1852;
/* FF 11 20  3 */ assign n1853 = n1219;
/* FF  4 29  3 */ always @(posedge clk) if (n157) n624 <= 1'b0 ? 1'b0 : n1854;
/* FF  5 18  6 */ always @(posedge clk) if (1'b1) n641 <= 1'b0 ? 1'b0 : n1855;
/* FF  1 23  2 */ assign n168 = n1856;
/* FF  2 22  7 */ assign n351 = n1857;
/* FF 19 20  4 */ assign n910 = n1858;
/* FF  1 26  5 */ assign n234 = n1859;
/* FF  5 28  6 */ assign n706 = n1860;
/* FF  6 29  5 */ assign n821 = n1861;
/* FF 10 20  2 */ assign n1862 = n1126;
/* FF 11 22  6 */ assign n685 = n1863;
/* FF  6 23  1 */ assign n380 = n1864;
/* FF  7 18  0 */ always @(posedge clk) if (1'b1) n844 <= 1'b0 ? 1'b0 : n1865;
/* FF  9 27  2 */ always @(posedge clk, posedge reset) if (reset) n987 <= 1'b0; else if (n226) n987 <= n1866;
/* FF 11 19  7 */ assign n1117 = n1867;
/* FF 17 21  7 */ always @(posedge clk, posedge reset) if (reset) n1457 <= 1'b0; else if (n1408) n1457 <= n1868;
/* FF  3 17  7 */ always @(posedge clk, posedge reset) if (reset) n446 <= 1'b0; else if (n82) n446 <= n1869;
/* FF  1 18  0 */ assign n69 = n1870;
/* FF 12 16  4 */ assign n1190 = n1871;
/* FF 13 23  1 */ assign n1066 = n1872;
/* FF  3 23  7 */ assign n204 = n1873;
/* FF  2 21  3 */ assign n156 = n1874;
/* FF 15 23  4 */ always @(posedge clk) if (n157) n1434 <= 1'b0 ? 1'b0 : n1875;
/* FF  6 16  5 */ always @(posedge clk) if (n53) n729 <= 1'b0 ? 1'b0 : n1876;
/* FF  4 28  4 */ assign n613 = n1877;
/* FF  7 27  6 */ assign n905 = n1878;
/* FF 11 24  3 */ assign n1097 = n1879;
/* FF 12 18  5 */ always @(posedge clk) if (1'b1) n1195 <= 1'b0 ? 1'b0 : n1880;
/* FF  4 26  0 */ assign n610 = n1881;
/* FF  9 22  0 */ always @(posedge clk) if (1'b1) n967 <= 1'b0 ? 1'b0 : n1882;
/* FF  9 24  4 */ assign n1883 = n1047;
/* FF 10 17  3 */ assign n11 = n1100;
/* FF 12 21  6 */ assign n1224 = n1884;
/* FF 18 19  6 */ assign n1346 = n1885;
/* FF 13 20  5 */ always @(posedge clk) if (1'b1) n1307 <= 1'b0 ? 1'b0 : n1886;
/* FF 10 27  3 */ always @(posedge clk) if (1'b1) n1060 <= 1'b0 ? 1'b0 : n1887;
/* FF  3 24  3 */ always @(posedge clk) if (1'b1) n222 <= 1'b0 ? 1'b0 : n1888;
/* FF  4 17  6 */ always @(posedge clk) if (n53) n549 <= 1'b0 ? 1'b0 : n1889;
/* FF  7 30  0 */ always @(posedge clk, posedge reset) if (reset) n252 <= 1'b0; else if (n51) n252 <= n1890;
/* FF  1 19  7 */ assign n94 = n1891;
/* FF  5 16  5 */ always @(posedge clk) if (n53) n632 <= 1'b0 ? 1'b0 : n1892;
/* FF  1 21  7 */ assign n138 = n1893;
/* FF 19 22  7 */ always @(posedge clk, posedge reset) if (reset) n77 <= 1'b0; else if (n1408) n77 <= n1894;
/* FF 13 18  4 */ always @(posedge clk) if (n53) n1288 <= 1'b0 ? 1'b0 : n1895;
/* FF 10 25  6 */ assign n1055 = n1896;
/* FF  1 24  4 */ assign n196 = n1897;
/* FF  5 26  1 */ assign n617 = n1898;
/* FF 10 18  7 */ always @(posedge clk) if (n53) n649 <= 1'b0 ? 1'b0 : n1899;
/* FF 14 23  2 */ always @(posedge clk) if (n53) n1141 <= 1'b0 ? 1'b0 : n1900;
/* FF 19 19  6 */ always @(posedge clk, posedge reset) if (reset) n1489 <= 1'b0; else if (n1408) n1489 <= n1901;
/* FF  6 21  0 */ always @(posedge clk, posedge reset) if (reset) n733 <= 1'b0; else if (n82) n733 <= n1902;
/* FF  2 27  3 */ assign n420 = n1903;
/* FF  4 22  0 */ always @(posedge clk) if (1'b1) n584 <= 1'b0 ? 1'b0 : n1904;
/* FF 11 21  4 */ assign n941 = n1905;
/* FF 12 20  1 */ assign n1199 = n1906;
/* FF  5 19  1 */ assign n643 = n1907;
/* FF  6 26  6 */ always @(posedge clk) if (1'b1) n790 <= 1'b0 ? 1'b0 : n1908;
/* FF  2 25  6 */ always @(posedge clk) if (1'b1) n414 <= 1'b0 ? 1'b0 : n1909;
/* FF 19 21  3 */ assign n1495 = n1910;
/* FF  5 29  5 */ assign n699 = n1911;
/* FF  3 25  4 */ assign n434 = n1912;
/* FF  2 19  6 */ always @(posedge clk, posedge reset) if (reset) n304 <= 1'b0; else if (n82) n304 <= n1913;
/* FF  6 28  6 */ assign n810 = n1914;
/* FF 11 23  5 */ assign n1140 = n1915;
/* FF 10 23  3 */ assign n1026 = n1916;
/* FF  6 22  6 */ always @(posedge clk) if (1'b1) n765 <= 1'b0 ? 1'b0 : n1917;
/* FF 11 26  6 */ assign n1174 = n1918;
/* FF  7 19  3 */ assign n855 = n1919;
/* FF 12 25  1 */ always @(posedge clk, posedge reset) if (reset) n775 <= 1'b0; else if (n226) n775 <= n1920;
/* FF  9 20  3 */ assign n379 = n1921;
/* FF  5 22  1 */ assign n1922 = n769;
/* FF 12 23  5 */ always @(posedge clk) if (1'b1) n1252 <= 1'b0 ? 1'b0 : n1923;
/* FF 13 24  0 */ assign n1075 = n1924;
/* FF  3 20  6 */ always @(posedge clk, posedge reset) if (reset) n139 <= 1'b0; else if (n82) n139 <= n1925;
/* FF  6 25  0 */ always @(posedge clk) if (n157) n707 <= 1'b0 ? 1'b0 : n1926;
/* FF 15 20  5 */ always @(posedge clk) if (n157) n598 <= 1'b0 ? 1'b0 : n1927;
/* FF  6 19  4 */ assign n1928 = n862;
/* FF  7 24  7 */ always @(posedge clk, posedge reset) if (reset) n768 <= 1'b0; else if (n226) n768 <= n1929;
/* FF  4 19  5 */ always @(posedge clk) if (1'b1) n209 <= 1'b0 ? 1'b0 : n1930;
/* FF 12 17  4 */ always @(posedge clk) if (n53) n1192 <= 1'b0 ? 1'b0 : n1931;
/* FF  7 22  7 */ always @(posedge clk) if (1'b1) n183 <= 1'b0 ? 1'b0 : n1932;
/* FF  9 23  7 */ always @(posedge clk, posedge reset) if (reset) n884 <= 1'b0; else if (n226) n884 <= n1933;
/* FF  4 25  1 */ assign n579 = n689;
/* FF 14 21  1 */ assign n1366 = n1934;
/* FF  5 24  0 */ always @(posedge clk) if (n157) n524 <= 1'b0 ? 1'b0 : n1935;
/* FF 10 16  0 */ assign n1936 = n1092;
/* FF  3 19  0 */ assign n1937 = n561;
/* FF 10 26  4 */ assign n1012 = n1938;
/* FF 11 17  1 */ always @(posedge clk, posedge reset) if (reset) n675 <= 1'b0; else if (n51) n675 <= n1939;
/* FF 13 21  6 */ assign n1042 = n1940;
/* FF  4 16  1 */ always @(posedge clk) if (n53) n448 <= 1'b0 ? 1'b0 : n1941;
/* FF  5 23  6 */ assign n1942 = n777;
/* FF  4 30  5 */ always @(posedge clk, posedge reset) if (reset) n95 <= 1'b0; else if (n51) n95 <= n1943;
/* FF  5 17  6 */ always @(posedge clk) if (1'b1) n636 <= 1'b0 ? 1'b0 : n1944;
/* FF  1 22  6 */ assign n154 = n1945;
/* FF 10 24  5 */ assign n1032 = n1946;
/* FF 13 19  3 */ assign n1292 = n1947;
/* FF  1 25  7 */ assign n215 = n1948;
/* FF 15 21  2 */ always @(posedge clk) if (n157) n1420 <= 1'b0 ? 1'b0 : n1949;
/* FF 10 21  6 */ always @(posedge clk, posedge reset) if (reset) n1009 <= 1'b0; else if (n226) n1009 <= n1950;
/* FF  6 18  3 */ always @(posedge clk) if (1'b1) n739 <= 1'b0 ? 1'b0 : n1951;
/* FF  5 27  6 */ assign n704 = n1952;
/* FF 14 22  5 */ assign n1378 = n1953;
/* FF  2 26  4 */ always @(posedge clk) if (1'b1) n432 <= 1'b0 ? 1'b0 : n1954;
/* FF  6 20  3 */ always @(posedge clk, posedge reset) if (reset) n578 <= 1'b0; else if (n226) n578 <= n1955;
/* FF  4 21  1 */ always @(posedge clk) if (1'b1) n126 <= 1'b0 ? 1'b0 : n1956;
/* FF 11 18  5 */ assign n1106 = n1957;
/* FF  5 20  0 */ assign n1958 = n752;
/* FF  1 17  0 */ assign n57 = n1959;
/* FF  2 24  5 */ assign n394 = n1960;
/* FF 14 19  5 */ assign n1355 = n1961;
/* FF  5 30  4 */ assign n723 = n1962;
/* FF  3 22  5 */ assign n103 = n1963;
/* FF  2 18  1 */ assign n286 = n1964;
/* FF 11 20  4 */ always @(posedge clk) if (n53) n1120 <= 1'b0 ? 1'b0 : n1965;
/* FF 15 22  4 */ assign n1415 = n1966;
/* FF  6 17  7 */ always @(posedge clk) if (1'b1) n736 <= 1'b0 ? 1'b0 : n1967;
/* FF  7 26  2 */ always @(posedge clk) if (1'b1) n898 <= 1'b0 ? 1'b0 : n1968;
/* FF  3 28  1 */ assign n1969 = n622;
/* FF  9 19  4 */ assign n954 = n1970;
/* FF 11 27  5 */ assign n1971 = n1281;
/* FF 12 19  7 */ assign n1204 = n1972;
/* FF  9 21  0 */ assign n1973 = n1015;
/* FF 12 22  6 */ assign n1191 = n1974;
/* FF  3 21  1 */ assign n1975 = n580;
/* FF  4 20  6 */ assign n81 = n1976;
/* FF  2 23  1 */ assign n342 = n1977;
/* FF 13 18  1 */ assign n1978 = n1349;
/* FF  4 18  6 */ always @(posedge clk, posedge reset) if (reset) n96 <= 1'b0; else if (n51) n96 <= n1979;
/* FF  7 25  0 */ assign n890 = n1980;
/* FF  4 24  6 */ always @(posedge clk) if (n157) n595 <= 1'b0 ? 1'b0 : n1981;
/* FF 14 18  2 */ always @(posedge clk) if (n53) n1001 <= 1'b0 ? 1'b0 : n1982;
/* FF  1 20  5 */ assign n118 = n1983;
/* FF  7 23  4 */ assign n1984 = n930;
/* FF 14 20  2 */ always @(posedge clk) if (n157) n783 <= 1'b0 ? 1'b0 : n1985;
/* FF  9 26  6 */ always @(posedge clk, posedge reset) if (reset) n942 <= 1'b0; else if (n226) n942 <= n1986;
/* FF 10 19  1 */ always @(posedge clk) if (n53) n843 <= 1'b0 ? 1'b0 : n1987;
/* FF  5 25  3 */ assign n679 = n1988;
/* FF 13 22  7 */ assign n786 = n1989;
/* FF 16 23  5 */ always @(posedge clk) if (n157) n1440 <= 1'b0 ? 1'b0 : n1990;
/* FF  4 23  0 */ always @(posedge clk) if (1'b1) n589 <= 1'b0 ? 1'b0 : n1991;
/* FF  4 29  4 */ assign n248 = n1992;
/* FF  5 18  7 */ assign n97 = n1993;
/* FF  1 23  1 */ assign n167 = n1994;
/* FF  2 22  6 */ assign n350 = n1995;
/* FF 13 20  2 */ always @(posedge clk) if (1'b1) n1304 <= 1'b0 ? 1'b0 : n1996;
/* FF  1 26  6 */ assign n235 = n1997;
/* FF  5 28  7 */ assign n620 = n1998;
/* FF 10 20  5 */ always @(posedge clk, posedge reset) if (reset) n751 <= 1'b0; else if (n226) n751 <= n1999;
/* FF 11 22  7 */ assign n933 = n2000;
/* FF 16 20  1 */ assign n1439 = n2001;
/* FF  7 18  1 */ assign n845 = n2002;
/* FF  9 27  1 */ assign n38 = n1082;
/* FF 11 19  6 */ always @(posedge clk) if (n53) n1110 <= 1'b0 ? 1'b0 : n2003;
/* FF 17 21  6 */ always @(posedge clk, posedge reset) if (reset) n1456 <= 1'b0; else if (n1408) n1456 <= n2004;
/* FF  5 21  3 */ assign n658 = n760;
/* FF  3 17  6 */ always @(posedge clk, posedge reset) if (reset) n445 <= 1'b0; else if (n82) n445 <= n2005;
/* FF 19 19  1 */ always @(posedge clk, posedge reset) if (reset) n1485 <= 1'b0; else if (n1408) n1485 <= n2006;
/* FF  1 18  1 */ assign n70 = n2007;
/* FF 13 23  0 */ assign n1065 = n2008;
/* FF  2 21  0 */ assign n2009 = n2010;
/* FF 11 21  3 */ assign n985 = n2012;
/* FF 15 23  7 */ always @(posedge clk) if (n157) n1226 <= 1'b0 ? 1'b0 : n2013;
/* FF  6 16  4 */ always @(posedge clk) if (n53) n634 <= 1'b0 ? 1'b0 : n2014;
/* FF  4 28  3 */ always @(posedge clk) if (1'b1) n265 <= 1'b0 ? 1'b0 : n2015;
/* FF  7 27  1 */ always @(posedge clk) if (1'b1) n903 <= 1'b0 ? 1'b0 : n2016;
/* FF 11 24  4 */ assign n971 = n2017;
/* FF 12 18  4 */ assign n1194 = n2018;
/* FF  4 26  3 */ always @(posedge clk) if (n157) n256 <= 1'b0 ? 1'b0 : n2019;
/* FF  9 24  5 */ assign n27 = n1048;
/* FF 10 17  0 */ assign n2020 = n1098;
/* FF 12 21  7 */ assign n1225 = n2021;
/* FF  3 18  0 */ always @(posedge clk) if (1'b1) n323 <= 1'b0 ? 1'b0 : n2022;
/* FF  3 24  4 */ always @(posedge clk) if (1'b1) n399 <= 1'b0 ? 1'b0 : n2023;
/* FF  4 17  7 */ always @(posedge clk) if (n53) n550 <= 1'b0 ? 1'b0 : n2024;
/* FF  7 30  1 */ always @(posedge clk, posedge reset) if (reset) n254 <= 1'b0; else if (n51) n254 <= n2025;
/* FF  1 19  6 */ assign n93 = n2026;
/* FF 12 23  2 */ assign n1249 = n2027;
/* FF  7 20  5 */ always @(posedge clk) if (1'b1) n865 <= 1'b0 ? 1'b0 : n2028;
/* FF  9 17  5 */ always @(posedge clk, posedge reset) if (reset) n946 <= 1'b0; else if (n226) n946 <= n2029;
/* FF  1 21  6 */ assign n137 = n2030;
/* FF 19 22  4 */ always @(posedge clk, posedge reset) if (reset) n1502 <= 1'b0; else if (n1408) n1502 <= n2031;
/* FF 13 18  5 */ assign n1289 = n2032;
/* FF 10 25  7 */ assign n1056 = n2033;
/* FF  1 24  5 */ assign n197 = n2034;
/* FF  5 26  2 */ assign n693 = n2035;
/* FF 14 23  3 */ always @(posedge clk) if (n53) n1118 <= 1'b0 ? 1'b0 : n2036;
/* FF 10 18  6 */ assign n2037 = n1113;
/* FF 18 20  3 */ always @(posedge clk, posedge reset) if (reset) n1468 <= 1'b0; else if (n1408) n1468 <= n2038;
/* FF  6 21  1 */ assign n2039 = n874;
/* FF 16 22  6 */ assign n443 = n2040;
/* FF  4 22  3 */ assign n122 = n2041;
/* FF 14 21  6 */ always @(posedge clk) if (n53) n867 <= 1'b0 ? 1'b0 : n2042;
/* FF 12 20  0 */ assign n1198 = n2043;
/* FF  5 19  0 */ assign n2044 = n746;
/* FF  6 26  5 */ assign n104 = n2045;
/* FF  2 25  7 */ assign n274 = n2046;
/* FF 10 26  3 */ assign n995 = n2047;
/* FF 13 21  1 */ assign n1041 = n2048;
/* FF  5 29  4 */ assign n717 = n2049;
/* FF  3 25  3 */ assign n2050 = n608;
/* FF  2 19  7 */ always @(posedge clk, posedge reset) if (reset) n305 <= 1'b0; else if (n82) n305 <= n2051;
/* FF 10 23  4 */ assign n1027 = n2052;
/* FF 11 23  4 */ assign n1139 = n2053;
/* FF  6 22  5 */ always @(posedge clk) if (1'b1) n764 <= 1'b0 ? 1'b0 : n2054;
/* FF 11 26  7 */ assign n1175 = n2055;
/* FF  7 19  2 */ assign n854 = n2056;
/* FF  9 20  0 */ always @(posedge clk, posedge reset) if (reset) n670 <= 1'b0; else if (n226) n670 <= n2057;
/* FF  5 22  2 */ always @(posedge clk) if (n157) n666 <= 1'b0 ? 1'b0 : n2058;
/* FF 14 24  0 */ always @(posedge clk) if (1'b1) n1379 <= 1'b0 ? 1'b0 : n2059;
/* FF  2 26  3 */ always @(posedge clk) if (1'b1) n431 <= 1'b0 ? 1'b0 : n2060;
/* FF 13 24  1 */ assign n1076 = n2061;
/* FF  3 20  7 */ always @(posedge clk, posedge reset) if (reset) n465 <= 1'b0; else if (n82) n465 <= n2062;
/* FF  2 20  3 */ assign n316 = n2063;
/* FF 11 18  2 */ always @(posedge clk) if (1'b1) n1103 <= 1'b0 ? 1'b0 : n2064;
/* FF 15 20  6 */ always @(posedge clk) if (n157) n1413 <= 1'b0 ? 1'b0 : n2065;
/* FF  3 26  7 */ always @(posedge clk, posedge reset) if (reset) n251 <= 1'b0; else if (n226) n251 <= n2066;
/* FF  6 19  5 */ assign n48 = n863;
/* FF  4 19  2 */ always @(posedge clk) if (1'b1) n559 <= 1'b0 ? 1'b0 : n2067;
/* FF  7 24  0 */ assign n2068 = n936;
/* FF 12 17  5 */ always @(posedge clk) if (n53) n1108 <= 1'b0 ? 1'b0 : n2069;
/* FF  4 25  2 */ always @(posedge clk, posedge reset) if (reset) n275 <= 1'b0; else if (n82) n275 <= n2070;
/* FF  9 23  6 */ always @(posedge clk, posedge reset) if (reset) n973 <= 1'b0; else if (n226) n973 <= n2071;
/* FF 10 22  3 */ always @(posedge clk) if (1'b1) n1020 <= 1'b0 ? 1'b0 : n2072;
/* FF  7 22  4 */ assign n878 = n923;
/* FF  5 24  1 */ assign n357 = n2073;
/* FF 10 16  3 */ always @(posedge clk, posedge reset) if (reset) n521 <= 1'b0; else if (n226) n521 <= n2074;
/* FF  3 19  3 */ assign n2075 = n563;
/* FF 11 17  0 */ assign n1094 = n2076;
/* FF  4 16  0 */ always @(posedge clk) if (n53) n542 <= 1'b0 ? 1'b0 : n2077;
/* FF  5 23  5 */ assign n253 = n2078;
/* FF 12 22  1 */ assign n1229 = n2079;
/* FF  4 30  4 */ always @(posedge clk, posedge reset) if (reset) n101 <= 1'b0; else if (n51) n101 <= n2080;
/* FF  5 17  1 */ assign n160 = n2081;
/* FF  1 22  7 */ assign n155 = n2082;
/* FF 13 19  2 */ always @(posedge clk) if (n53) n1285 <= 1'b0 ? 1'b0 : n2083;
/* FF 10 24  4 */ assign n1034 = n2084;
/* FF  1 25  6 */ assign n208 = n2085;
/* FF 15 21  1 */ always @(posedge clk) if (n157) n1419 <= 1'b0 ? 1'b0 : n2086;
/* FF 10 21  7 */ always @(posedge clk, posedge reset) if (reset) n538 <= 1'b0; else if (n226) n538 <= n2087;
/* FF  6 18  2 */ always @(posedge clk) if (1'b1) n738 <= 1'b0 ? 1'b0 : n2088;
/* FF  5 27  5 */ assign n703 = n2089;
/* FF 14 22  4 */ always @(posedge clk) if (n53) n1136 <= 1'b0 ? 1'b0 : n2090;
/* FF  6 20  2 */ always @(posedge clk, posedge reset) if (reset) n749 <= 1'b0; else if (n226) n749 <= n2091;
/* FF  4 21  2 */ always @(posedge clk) if (1'b1) n227 <= 1'b0 ? 1'b0 : n2092;
/* FF 14 20  5 */ always @(posedge clk) if (n157) n1364 <= 1'b0 ? 1'b0 : n2093;
/* FF 12 27  1 */ assign n29 = n1342;
/* FF  5 20  1 */ assign n627 = n2094;
/* FF  1 17  3 */ assign n60 = n2095;
/* FF  2 24  4 */ assign n393 = n2096;
/* FF 13 22  0 */ assign n1057 = n2097;
/* FF 14 19  6 */ assign n1356 = n2098;
/* FF  5 30  5 */ assign n722 = n2099;
/* FF  3 22  2 */ always @(posedge clk) if (1'b1) n180 <= 1'b0 ? 1'b0 : n2100;
/* FF  2 18  0 */ assign n2101 = n450;
/* FF 11 20  5 */ assign n1121 = n2102;
/* FF 15 22  5 */ assign n1429 = n2103;
/* FF  3 28  2 */ always @(posedge clk) if (n157) n523 <= 1'b0 ? 1'b0 : n2104;
/* FF  7 26  3 */ always @(posedge clk) if (1'b1) n899 <= 1'b0 ? 1'b0 : n2105;
/* FF  9 19  3 */ always @(posedge clk) if (n53) n953 <= 1'b0 ? 1'b0 : n2106;
/* FF 12 19  4 */ assign n657 = n2107;
/* FF  7 16  3 */ assign n2108 = n915;
/* FF 12 24  5 */ always @(posedge clk) if (1'b1) n1265 <= 1'b0 ? 1'b0 : n2109;
/* FF  9 21  3 */ assign n85 = n1017;
/* FF  3 21  0 */ always @(posedge clk, posedge reset) if (reset) n468 <= 1'b0; else if (n82) n468 <= n2110;
/* FF  4 20  5 */ always @(posedge clk) if (1'b1) n188 <= 1'b0 ? 1'b0 : n2111;
/* FF  2 23  2 */ assign n343 = n2112;
/* FF  7 18  6 */ always @(posedge clk) if (1'b1) n848 <= 1'b0 ? 1'b0 : n2113;
/* FF  6 24  2 */ assign n216 = n2114;
/* FF 11 19  1 */ assign n1008 = n2115;
/* FF  3 27  4 */ always @(posedge clk) if (1'b1) n532 <= 1'b0 ? 1'b0 : n2116;
/* FF  4 18  1 */ always @(posedge clk, posedge reset) if (reset) n555 <= 1'b0; else if (n51) n555 <= n2117;
/* FF 12 16  2 */ always @(posedge clk) if (1'b1) n1189 <= 1'b0 ? 1'b0 : n2118;
/* FF 13 23  7 */ assign n1069 = n2119;
/* FF  7 23  7 */ always @(posedge clk, posedge reset) if (reset) n678 <= 1'b0; else if (n226) n678 <= n2120;
/* FF  4 24  5 */ always @(posedge clk) if (n157) n597 <= 1'b0 ? 1'b0 : n2121;
/* FF  1 20  2 */ assign n115 = n2122;
/* FF 14 18  1 */ assign n2123 = n1409;
/* FF  9 26  7 */ always @(posedge clk, posedge reset) if (reset) n791 <= 1'b0; else if (n226) n791 <= n2124;
/* FF 10 19  2 */ always @(posedge clk) if (n53) n914 <= 1'b0 ? 1'b0 : n2125;
/* FF 16 23  2 */ assign n1444 = n2126;
/* FF  4 23  1 */ assign n201 = n2127;
/* FF  7 15  0 */ assign n6 = n2128;
/* FF  9 24  2 */ always @(posedge clk, posedge reset) if (reset) n975 <= 1'b0; else if (n226) n975 <= n2129;
/* FF 12 21  0 */ assign n1217 = n2130;
/* FF  4 29  5 */ assign n245 = n2131;
/* FF  1 23  0 */ assign n166 = n2132;
/* FF  2 22  5 */ assign n349 = n2133;
/* FF 13 20  3 */ always @(posedge clk) if (1'b1) n1305 <= 1'b0 ? 1'b0 : n2134;
/* FF  1 26  7 */ always @(posedge clk) if (1'b1) n236 <= 1'b0 ? 1'b0 : n2135;
/* FF  5 28  4 */ assign n711 = n2136;
/* FF 10 20  4 */ always @(posedge clk, posedge reset) if (reset) n1007 <= 1'b0; else if (n226) n1007 <= n2137;
/* FF 11 22  4 */ assign n982 = n2138;
/* FF  6 23  3 */ assign n2139 = n886;
/* FF  1 24  2 */ assign n194 = n2140;
/* FF 14 23  4 */ assign n1389 = n2141;
/* FF  9 27  0 */ assign n2142 = n1081;
/* FF 17 21  1 */ always @(posedge clk, posedge reset) if (reset) n1451 <= 1'b0; else if (n1408) n1451 <= n2143;
/* FF  5 21  2 */ assign n650 = n2144;
/* FF  1 18  2 */ assign n71 = n2145;
/* FF 19 19  0 */ assign n1484 = n2146;
/* FF  6 21  6 */ assign n2147 = n876;
/* FF  3 23  1 */ always @(posedge clk) if (n157) n397 <= n106 ? 1'b0 : n2148;
/* FF  2 21  1 */ assign n335 = n2149;
/* FF 11 21  2 */ assign n860 = n2150;
/* FF 12 20  7 */ assign n1210 = n2151;
/* FF 15 23  6 */ always @(posedge clk) if (n157) n1436 <= 1'b0 ? 1'b0 : n2152;
/* FF  6 16  7 */ assign n731 = n2153;
/* FF  7 27  0 */ always @(posedge clk) if (1'b1) n902 <= 1'b0 ? 1'b0 : n2154;
/* FF 11 24  5 */ assign n926 = n2155;
/* FF 12 18  7 */ assign n1197 = n2156;
/* FF  4 26  2 */ always @(posedge clk) if (n157) n611 <= 1'b0 ? 1'b0 : n2157;
/* FF  9 22  2 */ always @(posedge clk) if (1'b1) n966 <= 1'b0 ? 1'b0 : n2158;
/* FF 13 15  4 */ always @(posedge clk, posedge reset) if (reset) ready <= 1'b1; else if (1'b1) ready <= n2159;
/* FF 10 17  1 */ assign n7 = n2160;
/* FF 18 19  0 */ always @(posedge clk, posedge reset) if (reset) n1461 <= 1'b0; else if (n1408) n1461 <= n2161;
/* FF  3 18  1 */ assign n272 = n2162;
/* FF  7 19  5 */ assign n121 = n2163;
/* FF  3 24  5 */ always @(posedge clk) if (1'b1) n417 <= 1'b0 ? 1'b0 : n2164;
/* FF  4 17  0 */ assign n545 = n2165;
/* FF  7 30  6 */ always @(posedge clk, posedge reset) if (reset) n642 <= 1'b0; else if (n51) n642 <= n2166;
/* FF  1 19  5 */ assign n92 = n2167;
/* FF 12 23  3 */ always @(posedge clk) if (1'b1) n1250 <= 1'b0 ? 1'b0 : n2168;
/* FF 13 24  6 */ assign n1077 = n2169;
/* FF  5 16  3 */ always @(posedge clk) if (n53) n630 <= 1'b0 ? 1'b0 : n2170;
/* FF  1 21  1 */ assign n133 = n2171;
/* FF 19 22  5 */ always @(posedge clk, posedge reset) if (reset) n1497 <= 1'b0; else if (n1408) n1497 <= n2172;
/* FF 10 25  4 */ assign n1053 = n2173;
/* FF 13 18  6 */ assign n2174 = n1351;
/* FF  5 26  3 */ assign n619 = n2175;
/* FF 10 18  5 */ assign n999 = n2176;
/* FF 11 25  2 */ assign n51 = n2177;
/* FF 18 20  2 */ always @(posedge clk, posedge reset) if (reset) n1467 <= 1'b0; else if (n1408) n1467 <= n2178;
/* FF  4 22  2 */ assign n178 = n2179;
/* FF 14 21  7 */ assign n1368 = n2180;
/* FF  5 24  6 */ assign n362 = n2181;
/* FF  9 25  1 */ assign n981 = n2182;
/* FF  5 19  7 */ assign n648 = n2183;
/* FF  2 25  4 */ assign n412 = n2184;
/* FF 10 26  2 */ assign n1062 = n2185;
/* FF 11 17  7 */ always @(posedge clk, posedge reset) if (reset) n588 <= 1'b0; else if (n51) n588 <= n2186;
/* FF 13 21  0 */ assign n1142 = n2187;
/* FF  5 29  7 */ assign n506 = n2189;
/* FF 10 23  5 */ assign n994 = n2190;
/* FF  2 19  0 */ assign n2191 = n458;
/* FF 11 23  7 */ assign n990 = n2192;
/* FF  6 22  4 */ always @(posedge clk) if (1'b1) n249 <= 1'b0 ? 1'b0 : n2193;
/* FF  7 21  1 */ always @(posedge clk) if (n53) n766 <= n839 ? 1'b0 : n2194;
/* FF  1 25  1 */ assign n211 = n2195;
/* FF 12 25  3 */ assign n19 = n1337;
/* FF  9 20  1 */ assign n959 = n2196;
/* FF  5 22  3 */ assign n2197 = n770;
/* FF  6 20  5 */ assign n164 = n872;
/* FF  3 20  0 */ assign n2198 = n570;
/* FF  2 20  2 */ always @(posedge clk, posedge reset) if (reset) n142 <= 1'b1; else if (1'b1) n142 <= n2199;
/* FF  6 25  6 */ assign n2200 = n896;
/* FF 11 18  3 */ always @(posedge clk) if (1'b1) n1104 <= 1'b0 ? 1'b0 : n2201;
/* FF 12 27  6 */ always @(posedge clk, posedge reset) if (reset) n1205 <= 1'b0; else if (n226) n1205 <= n2202;
/* FF  6 19  6 */ always @(posedge clk, posedge reset) if (reset) n743 <= 1'b0; else if (n226) n743 <= n2203;
/* FF  7 24  1 */ assign n35 = n937;
/* FF  4 19  3 */ always @(posedge clk) if (1'b1) n127 <= 1'b0 ? 1'b0 : n2204;
/* FF  7 22  5 */ assign n157 = n924;
/* FF  9 23  5 */ assign n23 = n1038;
/* FF  4 25  3 */ assign n2205 = n690;
/* FF 10 22  2 */ assign n1019 = n2206;
/* FF 15 22  2 */ assign n577 = n2207;
/* FF  3 19  2 */ always @(posedge clk, posedge reset) if (reset) n454 <= 1'b0; else if (n82) n454 <= n2208;
/* FF  7 16  4 */ assign n838 = n2209;
/* FF  5 23  4 */ assign n361 = n2210;
/* FF 12 22  0 */ assign n1228 = n2211;
/* FF 13 25  5 */ assign n1336 = n2212;
/* FF  4 30  7 */ always @(posedge clk, posedge reset) if (reset) n618 <= 1'b0; else if (n51) n618 <= n2213;
/* FF  5 17  0 */ always @(posedge clk) if (1'b1) n635 <= 1'b0 ? 1'b0 : n2214;
/* FF  1 22  0 */ assign n148 = n2215;
/* FF  9 18  5 */ assign n948 = n2217;
/* FF 10 24  7 */ assign n934 = n2218;
/* FF 13 19  1 */ assign n2219 = n1358;
/* FF 15 21  0 */ always @(posedge clk) if (n157) n1418 <= 1'b0 ? 1'b0 : n2220;
/* FF 10 21  4 */ always @(posedge clk, posedge reset) if (reset) n1011 <= 1'b0; else if (n226) n1011 <= n2221;
/* FF  5 27  4 */ assign n702 = n2222;
/* FF  6 18  1 */ assign n737 = n2223;
/* FF  4 21  3 */ always @(posedge clk) if (1'b1) n158 <= 1'b0 ? 1'b0 : n2224;
/* FF 14 20  4 */ always @(posedge clk) if (n157) n1363 <= 1'b0 ? 1'b0 : n2225;
/* FF  5 25  5 */ assign n363 = n2226;
/* FF  9 26  0 */ assign n2227 = n1071;
/* FF  5 20  6 */ always @(posedge clk, posedge reset) if (reset) n656 <= 1'b0; else if (n82) n656 <= n2228;
/* FF  1 17  2 */ assign n59 = n2229;
/* FF  2 24  7 */ assign n395 = n2230;
/* FF 13 22  1 */ assign n970 = n2231;
/* FF  3 22  3 */ always @(posedge clk) if (1'b1) n381 <= 1'b0 ? 1'b0 : n2232;
/* FF 11 20  6 */ assign n2233 = n1220;
/* FF  3 28  3 */ always @(posedge clk) if (n157) n536 <= 1'b0 ? 1'b0 : n2234;
/* FF 11 27  7 */ always @(posedge clk) if (1'b1) n1086 <= 1'b0 ? 1'b0 : n2235;
/* FF  7 26  0 */ always @(posedge clk) if (1'b1) n897 <= 1'b0 ? 1'b0 : n2236;
/* FF  9 19  2 */ assign n2237 = n1004;
/* FF 12 19  5 */ assign n1002 = n2238;
/* FF  1 26  0 */ assign n230 = n2239;
/* FF 12 24  4 */ always @(posedge clk) if (1'b1) n1264 <= 1'b0 ? 1'b0 : n2240;
/* FF  9 21  2 */ assign n2241 = n1016;
/* FF  6 23  4 */ always @(posedge clk) if (n157) n773 <= 1'b0 ? 1'b0 : n2242;
/* FF  6 24  5 */ assign n219 = n2243;
/* FF  2 23  3 */ assign n373 = n2244;
/* FF  3 21  7 */ assign n466 = n2245;
/* FF 11 19  0 */ always @(posedge clk) if (n53) n1114 <= 1'b0 ? 1'b0 : n2246;
/* FF  9 27  7 */ always @(posedge clk, posedge reset) if (reset) n787 <= 1'b0; else if (n226) n787 <= n2247;
/* FF 12 26  5 */ always @(posedge clk, posedge reset) if (reset) n1279 <= 1'b0; else if (n226) n1279 <= n2248;
/* FF  7 18  7 */ assign n849 = n2249;
/* FF  4 18  0 */ always @(posedge clk, posedge reset) if (reset) n554 <= 1'b0; else if (n51) n554 <= n2250;
/* FF  7 25  6 */ assign n892 = n2251;
/* FF 13 23  6 */ assign n1067 = n2252;
/* FF  7 23  6 */ always @(posedge clk, posedge reset) if (reset) n882 <= 1'b0; else if (n226) n882 <= n2253;
/* FF  4 24  4 */ assign n2254 = n681;
/* FF  1 20  3 */ assign n116 = n2255;
/* FF 14 18  0 */ assign n1347 = n2256;
/* FF 15 23  1 */ always @(posedge clk) if (n157) n1432 <= 1'b0 ? 1'b0 : n2257;
/* FF 10 19  3 */ always @(posedge clk) if (n53) n637 <= 1'b0 ? 1'b0 : n2258;
/* FF 18 21  6 */ assign n2259 = n1498;
/* FF 16 23  3 */ assign n1445 = n2260;
/* FF  4 23  6 */ always @(posedge clk) if (1'b1) n592 <= 1'b0 ? 1'b0 : n2261;
/* FF  7 15  3 */ assign n834 = n913;
/* FF  9 24  3 */ always @(posedge clk, posedge reset) if (reset) n518 <= 1'b0; else if (n226) n518 <= n2262;
/* FF 10 17  6 */ always @(posedge clk, posedge reset) if (reset) n993 <= 1'b0; else if (n226) n993 <= n2263;
/* FF 12 21  1 */ assign n1216 = n2264;
/* FF  5 18  1 */ always @(posedge clk) if (1'b1) n638 <= 1'b0 ? 1'b0 : n2265;
/* FF  1 23  7 */ assign n173 = n2266;
/* FF  2 22  4 */ assign n348 = n2267;
/* FF 10 27  6 */ assign n1010 = n2268;
/* FF  5 28  5 */ assign n712 = n2269;
/* FF 10 20  7 */ always @(posedge clk, posedge reset) if (reset) n587 <= 1'b0; else if (n226) n587 <= n2270;
/* FF 11 22  5 */ assign n983 = n2271;
/* FF  1 24  3 */ assign n195 = n2272;
/* FF  5 26  4 */ assign n694 = n2273;
/* FF 17 21  0 */ always @(posedge clk, posedge reset) if (reset) n1450 <= 1'b0; else if (n1408) n1450 <= n2274;
/* FF  5 21  5 */ assign n651 = n761;
/* FF  1 18  3 */ assign n72 = n2275;
/* FF  6 21  7 */ assign n757 = n2276;
/* FF  3 23  0 */ always @(posedge clk) if (n157) n398 <= n106 ? 1'b0 : n2277;
/* FF  2 21  6 */ assign n338 = n2278;
/* FF 11 21  1 */ assign n869 = n2279;
/* FF 12 20  6 */ assign n958 = n2280;
/* FF  6 16  6 */ always @(posedge clk) if (n53) n730 <= 1'b0 ? 1'b0 : n2281;
/* FF 11 24  6 */ assign n1152 = n2282;
/* FF 12 18  6 */ always @(posedge clk) if (1'b1) n1196 <= 1'b0 ? 1'b0 : n2283;
/* FF  9 22  3 */ always @(posedge clk) if (1'b1) n968 <= 1'b0 ? 1'b0 : n2284;
/* FF  6 22  3 */ assign n763 = n2285;
/* FF 18 19  1 */ always @(posedge clk, posedge reset) if (reset) n1462 <= 1'b0; else if (n1408) n1462 <= n2286;
/* FF  3 18  6 */ always @(posedge clk) if (1'b1) n449 <= 1'b0 ? 1'b0 : n2287;
/* FF  6 27  4 */ always @(posedge clk) if (n157) n774 <= 1'b0 ? 1'b0 : n2288;
/* FF 11 16  1 */ always @(posedge clk) if (n53) n842 <= 1'b0 ? 1'b0 : n2289;
/* FF 12 25  4 */ always @(posedge clk, posedge reset) if (reset) n1275 <= 1'b0; else if (n226) n1275 <= n2290;
/* FF  7 19  4 */ assign n102 = n2291;
/* FF  3 24  6 */ always @(posedge clk) if (1'b1) n400 <= 1'b0 ? 1'b0 : n2292;
/* FF  4 17  1 */ always @(posedge clk) if (n53) n546 <= 1'b0 ? 1'b0 : n2293;
/* FF  7 30  7 */ always @(posedge clk, posedge reset) if (reset) n238 <= 1'b0; else if (n51) n238 <= n2294;
/* FF  1 19  4 */ assign n91 = n2295;
/* FF 12 23  0 */ assign n918 = n2296;
/* FF  9 20  6 */ assign n355 = n2297;
/* FF 13 24  7 */ assign n1078 = n2298;
/* FF  5 16  0 */ assign n628 = n2299;
/* FF  1 21  0 */ assign n132 = n2300;
/* FF 19 22  2 */ always @(posedge clk, posedge reset) if (reset) n1500 <= 1'b0; else if (n1408) n1500 <= n2301;
/* FF 13 18  7 */ always @(posedge clk) if (n53) n957 <= 1'b0 ? 1'b0 : n2302;
/* FF 10 25  5 */ assign n1054 = n2303;
/* FF 15 20  0 */ assign n2304 = n1441;
/* FF 10 18  4 */ always @(posedge clk) if (n53) n998 <= 1'b0 ? 1'b0 : n2305;
/* FF 11 25  1 */ assign n861 = n2306;
/* FF 18 20  5 */ always @(posedge clk, posedge reset) if (reset) n1470 <= 1'b0; else if (n1408) n1470 <= n2307;
/* FF  7 22  2 */ always @(posedge clk) if (1'b1) n359 <= 1'b0 ? 1'b0 : n2308;
/* FF  4 25  4 */ assign n601 = n2309;
/* FF  4 22  5 */ assign n247 = n2310;
/* FF 14 21  4 */ assign n1367 = n2311;
/* FF  9 25  0 */ always @(posedge clk) if (1'b1) n788 <= 1'b0 ? 1'b0 : n2312;
/* FF 10 16  5 */ assign n8 = n2313;
/* FF  5 24  7 */ always @(posedge clk) if (n157) n534 <= 1'b0 ? 1'b0 : n2314;
/* FF  5 19  6 */ always @(posedge clk, posedge reset) if (reset) n647 <= 1'b0; else if (n82) n647 <= n2315;
/* FF  6 26  3 */ always @(posedge clk) if (1'b1) n789 <= 1'b0 ? 1'b0 : n2316;
/* FF  2 25  5 */ always @(posedge clk) if (1'b1) n413 <= 1'b0 ? 1'b0 : n2317;
/* FF 10 26  1 */ assign n1023 = n2318;
/* FF 11 17  6 */ always @(posedge clk, posedge reset) if (reset) n467 <= 1'b0; else if (n51) n467 <= n2319;
/* FF 13 21  3 */ assign n1031 = n2320;
/* FF  5 29  6 */ assign n437 = n2321;
/* FF  3 25  1 */ assign n242 = n2322;
/* FF  2 19  1 */ assign n301 = n459;
/* FF  6 28  3 */ assign n604 = n2323;
/* FF 10 23  6 */ assign n1000 = n2324;
/* FF 11 23  6 */ assign n989 = n2325;
/* FF 11 26  5 */ always @(posedge clk) if (1'b1) n1173 <= 1'b0 ? 1'b0 : n2326;
/* FF  7 21  0 */ assign n2327 = n921;
/* FF  1 25  0 */ assign n210 = n2328;
/* FF 15 21  7 */ always @(posedge clk) if (n157) n1417 <= 1'b0 ? 1'b0 : n2329;
/* FF  5 27  3 */ assign n701 = n2330;
/* FF 14 22  2 */ always @(posedge clk) if (n53) n1135 <= 1'b0 ? 1'b0 : n2331;
/* FF  5 22  4 */ always @(posedge clk) if (n157) n667 <= 1'b0 ? 1'b0 : n2332;
/* FF 14 24  2 */ assign n1398 = n2333;
/* FF  2 26  1 */ assign n430 = n2334;
/* FF  6 20  4 */ always @(posedge clk, posedge reset) if (reset) n662 <= 1'b0; else if (n226) n662 <= n2335;
/* FF  6 25  7 */ always @(posedge clk) if (n157) n621 <= 1'b0 ? 1'b0 : n2336;
/* FF  2 20  5 */ assign n318 = n2337;
/* FF  3 20  1 */ assign n462 = n571;
/* FF 11 18  0 */ assign n1101 = n2338;
/* FF 12 27  7 */ always @(posedge clk, posedge reset) if (reset) n174 <= 1'b0; else if (n226) n174 <= n2339;
/* FF  6 19  7 */ always @(posedge clk, posedge reset) if (reset) n568 <= 1'b0; else if (n226) n568 <= n2340;
/* FF  7 24  2 */ always @(posedge clk, posedge reset) if (reset) n868 <= 1'b0; else if (n226) n868 <= n2341;
/* FF  4 19  0 */ always @(posedge clk) if (1'b1) n560 <= 1'b0 ? 1'b0 : n2342;
/* FF 14 19  0 */ always @(posedge clk) if (n53) n1227 <= n839 ? 1'b0 : n2343;
/* FF  9 23  4 */ assign n2344 = n1037;
/* FF 10 22  1 */ always @(posedge clk) if (1'b1) n1018 <= 1'b0 ? 1'b0 : n2345;
/* FF 15 22  3 */ always @(posedge clk) if (1'b1) n1428 <= 1'b0 ? 1'b0 : n2346;
/* FF  3 19  5 */ always @(posedge clk, posedge reset) if (reset) n455 <= 1'b0; else if (n82) n455 <= n2347;
/* FF  7 16  5 */ assign n839 = n2348;
/* FF  9 21  5 */ always @(posedge clk, posedge reset) if (reset) n718 <= 1'b0; else if (n226) n718 <= n2349;
/* FF  5 23  3 */ always @(posedge clk) if (n157) n672 <= 1'b0 ? 1'b0 : n2350;
/* FF 12 22  3 */ assign n1213 = n2351;
/* FF 13 25  4 */ assign n290 = n2352;
/* FF  4 30  6 */ always @(posedge clk, posedge reset) if (reset) n456 <= 1'b0; else if (n51) n456 <= n2353;
/* FF  5 17  3 */ assign n79 = n2354;
/* FF  1 22  1 */ assign n149 = n2355;
/* FF  9 18  6 */ assign n947 = n2356;
/* FF 10 24  6 */ assign n935 = n2357;
/* FF  7 23  1 */ assign n123 = n929;
/* FF 14 18  7 */ always @(posedge clk) if (n53) n1214 <= 1'b0 ? 1'b0 : n2358;
/* FF  4 21  4 */ assign n574 = n2359;
/* FF  9 26  1 */ assign n33 = n1072;
/* FF 10 19  4 */ always @(posedge clk) if (n53) n916 <= 1'b0 ? 1'b0 : n2360;
/* FF  5 25  4 */ assign n207 = n2361;
/* FF  1 17  5 */ assign n62 = n2362;
/* FF  2 24  6 */ assign n186 = n2363;
/* FF 13 22  2 */ assign n1045 = n2364;
/* FF  3 22  0 */ assign n177 = n2365;
/* FF  2 18  6 */ always @(posedge clk, posedge reset) if (reset) n289 <= 1'b0; else if (n82) n289 <= n2366;
/* FF 11 20  7 */ always @(posedge clk) if (n53) n917 <= 1'b0 ? 1'b0 : n2367;
/* FF 11 27  6 */ assign n111 = n1282;
/* FF  9 19  1 */ always @(posedge clk) if (n53) n952 <= 1'b0 ? 1'b0 : n2368;
/* FF 12 19  2 */ assign n1202 = n2369;
/* FF  1 26  1 */ assign n231 = n2370;
/* FF  5 28  2 */ assign n710 = n2371;
/* FF 15 16  6 */ assign n911 = n1438;
/* FF  6 23  5 */ assign n203 = n2372;
/* FF  3 21  6 */ always @(posedge clk, posedge reset) if (reset) n471 <= 1'b0; else if (n82) n471 <= n2373;
/* FF  4 20  3 */ always @(posedge clk) if (1'b1) n566 <= 1'b0 ? 1'b0 : n2374;
/* FF  2 23  4 */ assign n374 = n2375;
/* FF  7 18  4 */ always @(posedge clk) if (1'b1) n846 <= 1'b0 ? 1'b0 : n2376;
/* FF  9 27  6 */ always @(posedge clk, posedge reset) if (reset) n988 <= 1'b0; else if (n226) n988 <= n2377;
/* FF  6 24  4 */ always @(posedge clk) if (n157) n778 <= 1'b0 ? 1'b0 : n2378;
/* FF  3 27  6 */ always @(posedge clk) if (1'b1) n533 <= 1'b0 ? 1'b0 : n2379;
/* FF  7 25  5 */ always @(posedge clk) if (1'b1) n891 <= 1'b0 ? 1'b0 : n2380;
/* FF  4 18  3 */ always @(posedge clk, posedge reset) if (reset) n99 <= 1'b0; else if (n51) n99 <= n2381;
/* FF 11 19  3 */ always @(posedge clk) if (n53) n1115 <= 1'b0 ? 1'b0 : n2382;
/* FF 13 23  5 */ assign n1070 = n2383;
/* FF  1 20  0 */ assign n113 = n2384;
/* FF 15 23  0 */ always @(posedge clk) if (n157) n1424 <= 1'b0 ? 1'b0 : n2385;
/* FF 18 21  7 */ assign n1474 = n2386;
/* FF  4 26  4 */ assign n246 = n2387;
/* FF  4 23  7 */ assign n277 = n2388;
/* FF  7 15  2 */ assign n2389 = n912;
/* FF 12 21  2 */ assign n1221 = n2390;
/* FF 10 17  7 */ always @(posedge clk, posedge reset) if (reset) n719 <= 1'b0; else if (n226) n719 <= n2391;
/* FF  4 29  7 */ always @(posedge clk) if (n157) n257 <= 1'b0 ? 1'b0 : n2392;
/* FF  5 18  2 */ always @(posedge clk) if (1'b1) n639 <= 1'b0 ? 1'b0 : n2393;
/* FF  1 23  6 */ assign n172 = n2394;
/* FF  2 22  3 */ assign n347 = n2395;
/* FF 10 27  7 */ assign n616 = n2396;
/* FF  6 29  1 */ assign n820 = n2397;
/* FF 11 22  2 */ assign n858 = n2398;
/* FF  7 20  0 */ always @(posedge clk) if (1'b1) n857 <= 1'b0 ? 1'b0 : n2399;
/* FF 10 15  7 */ always @(posedge clk, posedge reset) if (reset) n50 <= 1'b1; else if (1'b1) n50 <= n2400;
/* FF  1 24  0 */ assign n193 = n2401;
/* FF  5 26  5 */ assign n695 = n2402;
/* FF 10 18  3 */ assign n2403 = n1112;
/* FF 17 21  3 */ always @(posedge clk, posedge reset) if (reset) n1453 <= 1'b0; else if (n1408) n1453 <= n2404;
/* FF  5 21  4 */ always @(posedge clk, posedge reset) if (reset) n659 <= 1'b0; else if (n82) n659 <= n2405;
/* FF  1 18  4 */ assign n73 = n2406;
/* FF 19 19  2 */ always @(posedge clk, posedge reset) if (reset) n1486 <= 1'b0; else if (n1408) n1486 <= n2407;
/* FF  6 21  4 */ always @(posedge clk, posedge reset) if (reset) n558 <= 1'b0; else if (n82) n558 <= n2408;
/* FF  2 27  7 */ assign n185 = n2409;
/* FF  3 23  3 */ always @(posedge clk) if (n157) n492 <= n106 ? 1'b0 : n2410;
/* FF  2 21  7 */ assign n339 = n2411;
/* FF 11 21  0 */ assign n2412 = n2413;
/* FF 12 20  5 */ assign n1109 = n2415;
/* FF  7 27  2 */ assign n144 = n2416;
/* FF  4 28  0 */ assign n614 = n2417;
/* FF 11 24  7 */ assign n1153 = n2418;
/* FF  5 29  1 */ assign n713 = n2419;
/* FF 13 15  2 */ always @(posedge clk, posedge reset) if (reset) n49 <= 1'b0; else if (1'b1) n49 <= n2420;
/* FF 11 26  2 */ assign n1171 = n2421;
/* FF 18 19  2 */ always @(posedge clk, posedge reset) if (reset) n1463 <= 1'b0; else if (n1408) n1463 <= n2422;
/* FF  3 18  7 */ always @(posedge clk) if (1'b1) n205 <= 1'b0 ? 1'b0 : n2423;
/* FF  7 19  7 */ assign n850 = n2424;
/* FF 12 25  5 */ assign n17 = n1338;
/* FF  3 24  7 */ always @(posedge clk) if (1'b1) n223 <= 1'b0 ? 1'b0 : n2425;
/* FF  4 17  2 */ always @(posedge clk) if (n53) n78 <= 1'b0 ? 1'b0 : n2426;
/* FF  7 30  4 */ always @(posedge clk, posedge reset) if (reset) n557 <= 1'b0; else if (n51) n557 <= n2427;
/* FF  1 19  3 */ assign n90 = n2428;
/* FF 12 23  1 */ always @(posedge clk) if (1'b1) n1248 <= 1'b0 ? 1'b0 : n2429;
/* FF 13 24  4 */ assign n1014 = n2430;
/* FF  5 16  1 */ always @(posedge clk) if (n53) n629 <= 1'b0 ? 1'b0 : n2431;
/* FF  1 21  3 */ assign n135 = n2432;
/* FF 19 22  3 */ always @(posedge clk, posedge reset) if (reset) n1501 <= 1'b0; else if (n1408) n1501 <= n2433;
/* FF 13 18  0 */ assign n1286 = n2434;
/* FF 10 25  2 */ assign n1051 = n2435;
/* FF 15 20  1 */ assign n141 = n2436;
/* FF 11 25  0 */ assign n919 = n2437;
/* FF 18 20  4 */ always @(posedge clk, posedge reset) if (reset) n1469 <= 1'b0; else if (n1408) n1469 <= n2438;
/* FF  7 22  3 */ always @(posedge clk) if (1'b1) n877 <= 1'b0 ? 1'b0 : n2439;
/* FF  9 23  3 */ always @(posedge clk, posedge reset) if (reset) n503 <= 1'b0; else if (n226) n503 <= n2440;
/* FF  4 25  5 */ assign n602 = n691;
/* FF  4 22  4 */ assign n585 = n2441;
/* FF 14 21  5 */ assign n2442 = n1427;
/* FF  5 24  4 */ assign n358 = n2443;
/* FF  9 25  3 */ assign n984 = n2444;
/* FF 10 16  4 */ assign n2445 = n1093;
/* FF 13 27  2 */ always @(posedge clk) if (n53) n1340 <= n839 ? 1'b0 : n2446;
/* FF  5 19  5 */ assign n646 = n748;
/* FF  6 26  2 */ always @(posedge clk) if (1'b1) n494 <= 1'b0 ? 1'b0 : n2447;
/* FF  2 25  2 */ assign n322 = n2448;
/* FF 13 21  2 */ assign n745 = n2449;
/* FF 11 17  5 */ always @(posedge clk, posedge reset) if (reset) n176 <= 1'b0; else if (n51) n176 <= n2450;
/* FF 10 26  0 */ assign n1061 = n2451;
/* FF  3 25  0 */ assign n2452 = n607;
/* FF  2 19  2 */ always @(posedge clk, posedge reset) if (reset) n66 <= 1'b0; else if (n82) n66 <= n2453;
/* FF 10 23  7 */ assign n1028 = n2454;
/* FF 11 23  1 */ assign n1138 = n2455;
/* FF  4 30  1 */ always @(posedge clk, posedge reset) if (reset) n438 <= 1'b0; else if (n51) n438 <= n2456;
/* FF  1 25  3 */ assign n213 = n2457;
/* FF 15 21  6 */ always @(posedge clk) if (n157) n1423 <= 1'b0 ? 1'b0 : n2458;
/* FF  5 27  2 */ assign n505 = n2459;
/* FF 10 21  2 */ assign n2460 = n1132;
/* FF 14 22  1 */ assign n2461 = n1430;
/* FF  5 22  5 */ assign n401 = n2462;
/* FF  2 26  0 */ assign n419 = n2463;
/* FF  6 20  7 */ always @(posedge clk, posedge reset) if (reset) n341 <= 1'b0; else if (n226) n341 <= n2464;
/* FF  3 20  2 */ always @(posedge clk, posedge reset) if (reset) n463 <= 1'b0; else if (n82) n463 <= n2465;
/* FF  2 20  4 */ assign n317 = n2466;
/* FF  6 25  4 */ always @(posedge clk) if (n157) n784 <= 1'b0 ? 1'b0 : n2467;
/* FF 11 18  1 */ always @(posedge clk) if (1'b1) n1102 <= 1'b0 ? 1'b0 : n2468;
/* FF 12 27  4 */ assign n2469 = n1343;
/* FF  7 24  3 */ always @(posedge clk, posedge reset) if (reset) n885 <= 1'b0; else if (n226) n885 <= n2470;
/* FF  4 19  1 */ always @(posedge clk) if (1'b1) n244 <= 1'b0 ? 1'b0 : n2471;
/* FF 14 19  1 */ assign n1352 = n2472;
/* FF  5 30  0 */ assign n507 = n2473;
/* FF 10 22  0 */ assign n932 = n2474;
/* FF  6 17  3 */ assign n735 = n2475;
/* FF  7 26  6 */ assign n684 = n2476;
/* FF  3 19  4 */ assign n321 = n564;
/* FF  9 21  4 */ always @(posedge clk, posedge reset) if (reset) n963 <= 1'b0; else if (n226) n963 <= n2477;
/* FF 12 24  2 */ always @(posedge clk) if (1'b1) n1254 <= 1'b0 ? 1'b0 : n2478;
/* FF  5 23  2 */ assign n2479 = n776;
/* FF 12 22  2 */ assign n1238 = n2480;
/* FF 13 25  7 */ always @(posedge clk) if (1'b1) n1079 <= 1'b0 ? 1'b0 : n2481;
/* FF  9 18  7 */ assign n949 = n2482;
/* FF  1 22  2 */ assign n150 = n2483;
/* FF 10 24  1 */ assign n1013 = n2484;
/* FF  3 27  1 */ always @(posedge clk) if (1'b1) n531 <= 1'b0 ? 1'b0 : n2485;
/* FF  4 24  2 */ always @(posedge clk) if (n157) n596 <= 1'b0 ? 1'b0 : n2486;
/* FF  7 23  0 */ assign n2487 = n928;
/* FF 14 18  6 */ assign n2488 = n1411;
/* FF  4 21  5 */ assign n575 = n2489;
/* FF 14 20  6 */ always @(posedge clk) if (n157) n1365 <= 1'b0 ? 1'b0 : n2490;
/* FF  9 26  2 */ always @(posedge clk, posedge reset) if (reset) n980 <= 1'b0; else if (n226) n980 <= n2491;
/* FF 10 19  5 */ always @(posedge clk) if (n53) n841 <= 1'b0 ? 1'b0 : n2492;
/* FF  5 25  7 */ always @(posedge clk) if (1'b1) n527 <= 1'b0 ? 1'b0 : n2493;
/* FF  5 20  4 */ assign n652 = n754;
/* FF  1 17  4 */ assign n61 = n2494;
/* FF  2 24  1 */ assign n376 = n2495;
/* FF 13 22  3 */ assign n433 = n2496;
/* FF  3 22  1 */ always @(posedge clk) if (1'b1) n184 <= 1'b0 ? 1'b0 : n2497;
/* FF  2 18  5 */ assign n288 = n452;
/* FF  4 29  0 */ always @(posedge clk) if (n157) n623 <= 1'b0 ? 1'b0 : n2498;
/* FF  9 19  0 */ assign n2499 = n1003;
/* FF 12 19  3 */ assign n750 = n2500;
/* FF  1 26  2 */ assign n232 = n2501;
/* FF  5 28  3 */ assign n698 = n2502;
/* FF 10 20  1 */ assign n46 = n2503;
/* FF  6 29  6 */ assign n780 = n2504;
/* FF 15 16  7 */ assign n1408 = n2505;
/* FF  6 24  7 */ always @(posedge clk) if (n157) n605 <= 1'b0 ? 1'b0 : n2506;
/* FF  4 20  2 */ always @(posedge clk) if (1'b1) n225 <= 1'b0 ? 1'b0 : n2507;
/* FF  2 23  5 */ assign n206 = n2508;
/* FF  7 18  5 */ always @(posedge clk) if (1'b1) n847 <= 1'b0 ? 1'b0 : n2509;
/* FF  9 27  5 */ assign n40 = n1084;
/* FF  3 21  5 */ assign n457 = n583;
/* FF 11 19  2 */ assign n2510 = n1208;
/* FF  4 18  2 */ always @(posedge clk, posedge reset) if (reset) n306 <= 1'b0; else if (n51) n306 <= n2511;
/* FF 13 23  4 */ assign n1068 = n2512;
/* FF  1 20  1 */ assign n114 = n2513;
/* FF 15 23  3 */ always @(posedge clk) if (n157) n1433 <= 1'b0 ? 1'b0 : n2514;
/* FF  6 16  0 */ assign n727 = n2515;
/* FF  7 27  5 */ always @(posedge clk) if (1'b1) n904 <= 1'b0 ? 1'b0 : n2516;
/* FF 11 24  0 */ assign n1129 = n2517;
/* FF 18 21  4 */ assign n1473 = n2518;
/* FF  4 26  7 */ always @(posedge clk) if (n157) n612 <= 1'b0 ? 1'b0 : n2519;
/* FF  9 22  5 */ always @(posedge clk) if (1'b1) n758 <= 1'b0 ? 1'b0 : n2520;
/* FF  4 23  4 */ always @(posedge clk) if (1'b1) n590 <= 1'b0 ? 1'b0 : n2521;
/* FF  9 24  1 */ assign n25 = n1046;
/* FF 10 17  4 */ always @(posedge clk, posedge reset) if (reset) n992 <= 1'b0; else if (n226) n992 <= n2522;
/* FF 12 21  3 */ assign n1222 = n2523;
/* FF  5 18  3 */ always @(posedge clk) if (1'b1) n378 <= 1'b0 ? 1'b0 : n2524;
/* FF  1 23  5 */ assign n171 = n2525;
/* FF  2 22  2 */ assign n124 = n2526;
/* FF 13 20  6 */ always @(posedge clk) if (1'b1) n1308 <= 1'b0 ? 1'b0 : n2527;
/* FF 10 27  0 */ assign n880 = n2528;
/* FF  3 24  0 */ assign n83 = n2529;
/* FF 11 22  3 */ assign n925 = n2530;
/* FF  7 20  1 */ always @(posedge clk) if (1'b1) n864 <= 1'b0 ? 1'b0 : n2531;
/* FF  1 24  1 */ assign n182 = n2532;
/* FF  5 26  6 */ assign n504 = n2533;
/* FF 10 18  2 */ always @(posedge clk) if (n53) n997 <= 1'b0 ? 1'b0 : n2534;
/* FF 17 21  2 */ always @(posedge clk, posedge reset) if (reset) n1452 <= 1'b0; else if (n1408) n1452 <= n2535;
/* FF  5 21  7 */ always @(posedge clk, posedge reset) if (reset) n661 <= 1'b0; else if (n82) n661 <= n2536;
/* FF  1 18  5 */ assign n74 = n2537;
/* FF  2 27  0 */ always @(posedge clk) if (1'b1) n435 <= 1'b0 ? 1'b0 : n2538;
/* FF 19 19  5 */ always @(posedge clk, posedge reset) if (reset) n1488 <= 1'b0; else if (n1408) n1488 <= n2539;
/* FF  6 21  5 */ always @(posedge clk, posedge reset) if (reset) n552 <= 1'b0; else if (n82) n552 <= n2540;
/* FF  3 23  2 */ assign n491 = n2541;
/* FF  5 14  6 */ always @(posedge clk, posedge reset) if (reset) n541 <= 1'b0; else if (n226) n541 <= n2542;
/* FF  2 21  4 */ assign n337 = n2543;
/* FF 11 21  7 */ assign n1125 = n2544;
/* FF 12 20  4 */ assign n956 = n2545;
/* FF 12 18  0 */ always @(posedge clk) if (1'b1) n1193 <= 1'b0 ? 1'b0 : n2546;
/* FF  5 29  0 */ assign n714 = n2547;
/* FF  3 25  7 */ always @(posedge clk, posedge reset) if (reset) n240 <= 1'b0; else if (n82) n240 <= n2548;
/* FF 10 23  0 */ assign n1024 = n2549;
/* FF  6 22  1 */ always @(posedge clk) if (1'b1) n762 <= 1'b0 ? 1'b0 : n2550;
/* FF 11 26  3 */ assign n1172 = n2551;
/* FF 18 19  3 */ always @(posedge clk, posedge reset) if (reset) n1464 <= 1'b0; else if (n1408) n1464 <= n2552;
/* FF  3 18  4 */ always @(posedge clk) if (1'b1) n243 <= 1'b0 ? 1'b0 : n2553;
/* FF  7 19  6 */ always @(posedge clk) if (1'b1) n856 <= 1'b0 ? 1'b0 : n2554;
/* FF 12 25  6 */ always @(posedge clk, posedge reset) if (reset) n1276 <= 1'b0; else if (n226) n1276 <= n2555;
/* FF  9 20  4 */ assign n353 = n2556;
/* FF  4 17  3 */ always @(posedge clk) if (n53) n547 <= 1'b0 ? 1'b0 : n2557;
/* FF  7 30  5 */ always @(posedge clk, posedge reset) if (reset) n255 <= 1'b0; else if (n51) n255 <= n2558;
/* FF  1 19  2 */ assign n89 = n2559;
/* FF 12 23  6 */ assign n1154 = n2560;
/* FF 13 24  5 */ assign n779 = n2561;
/* FF  1 21  2 */ always @(posedge clk) if (1'b1) n134 <= 1'b0 ? 1'b0 : n2562;
/* FF 10 25  3 */ assign n1052 = n2563;

endmodule

