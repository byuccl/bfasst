`ifndef LUCONST
`define LUCONST

localparam[3:0] AND = 4'b0000;
localparam[3:0] OR = 4'b0001;
localparam[3:0] ADD = 4'b0010;
localparam[3:0] SUB = 4'b0011;
localparam[3:0] LESS_THAN = 4'b0111;
localparam[3:0] SRL = 4'b1000;
localparam[3:0] SLL = 4'b1001;
localparam[3:0] SRA = 4'b1010;
localparam[3:0] XOR = 4'b1101;


`endif 