
module chip (input clk, input rst, output \data_out[7] , output \data_out[5] , output \data_out[6] , output \data_out[0] , output read_e, output \data_out[2] , output \data_out[3] , output \data_out[1] , output \data_out[4] , output write_e, output \port_addr[6] , output \port_addr[7] , output \port_addr[4] , output \port_addr[5] , output \port_addr[3] , output \port_addr[2] , output \port_addr[0] , output \port_addr[1] , input \data_in[7] , input \data_in[6] , input \data_in[0] , input \data_in[5] , input \data_in[4] , input \data_in[3] , input \data_in[1] , input \data_in[2] );

wire n1, clk, rst, \data_out[7] , \data_out[5] , \data_out[6] , \data_out[0] , \data_out[2] , \data_out[3] , \data_out[1] ;
wire \data_out[4] , \port_addr[6] , \port_addr[7] , \port_addr[4] , n18, n20, \port_addr[5] , \port_addr[3] , \port_addr[2] , n24;
wire \port_addr[0] , \port_addr[1] , n28, n33, n35, n38, n39, n40, n42, n43;
wire n44, n45, n47, n48, n49, n50, n51, n52, n53, n54;
wire n57, n58, n59, n60, n61, n62, n63, n64, n65, n66;
wire n67, n69, n72, n73, n75, n76, n77, n78, n79, n80;
wire n81, n82, n83, n84, n85, n86, n87, n88, n92, n93;
wire n94, n97, n98, n99, n100, n102, n103, n104, n107, n108;
wire n112, n113, n114, n115, n116, n117, n118, n119, n120, n121;
wire n122, n123, n124, n125, n126, n127, n128, n129, n130, n131;
wire n132, n134, n135, n136, n137, n138, n139, n140, n141, n142;
wire n143, n144, n145, n146, n147, n148, n149, n150, n151, n152;
wire n153, n154, n155, n158, n159, n160, n161, n162, n163, n164;
wire n165, n166, n167, n168, n169, n172, n173, n174, n175, n176;
wire n177, n178, n179, n180, n182, n183, n184, n185, n186, n187;
wire n188, n189, n190, n191, n192, n193, n194, n196, n197, n198;
wire n199, n201, n202, n203, n204, n205, n206, n207, n208, n209;
wire n210, n211, n212, n213, n214, n215, n216, n217, n218, n219;
wire n220, n221, n222, n223, n224, n225, n226, n227, n228, n229;
wire n230, n231, n232, n235, n236, n237, n238, n239, n240, n241;
wire n242, n243, n244, n245, n246, n247, n248, n249, n250, n251;
wire n254, n261, n262, n263, n264, n265, n269, n270, n271, n272;
wire n276, n277, n278, n279, n280, n281, n282, n283, n284, n285;
wire n286, n287, n288, n289, n294, n295, n297, n298, n299, open_0;
wire open_1, open_2, open_3, open_4, open_5, open_6, open_7, open_8, open_9, open_10;
wire open_11, open_12, open_13, open_14, open_15, open_16, open_17, open_18, open_19, open_20;
wire open_21, open_22, open_23, open_24, open_25, open_26, open_27, open_28, open_29, open_30;
wire open_31, open_32, open_33, open_34, open_35, open_36, open_37, open_38, open_39, open_40;
wire open_41, open_42, open_43, open_44, open_45, open_46, open_47, open_48, open_49, open_50;
wire open_51, open_52, open_53, open_54, open_55, open_56, open_57, open_58, open_59, open_60;
wire open_61, open_62, open_63, open_64, open_65, open_66, open_67, open_68, open_69, open_70;
wire open_71, open_72, open_73, open_74, open_75, open_76, open_77, open_78, open_79, open_80;
wire open_81, open_82, open_83, open_84, open_85, open_86, open_87, open_88, open_89, open_90;
wire open_91, open_92, open_93, open_94, open_95, open_96, open_97, open_98, open_99, open_100;
wire open_101, open_102, open_103, open_104, open_105, open_106, open_107, open_108, open_109, open_110;
wire open_111, open_112, open_113, open_114, open_115, open_116, open_117, open_118, open_119, open_120;
wire open_121, open_122, open_123, open_124, open_125, open_126, open_127, open_128, open_129, open_130;
wire open_131, open_132, n300, n301, n302, n303, n304, n305, n306, n307;
wire n308, n309, n310, n311, n312, n313, n314, n315, n316, n317;
wire n318, n319, n320, n321, n322, n323, n324, n325, n326, n327;
wire n328, n329, n330, n331, n332, n333, n334, n335, n336, n337;
wire n338, n339, n340, n341, n342, n343, n344, n345, n346, n347;
wire n348, n349, n350, n351, n352, n353, n354, n355, n356, n357;
wire n358, n359, n360, n361, n362, n363, n364, n365, n366, n367;
wire n368, n369, n370, n371, n372, n373, n374, n375, n376, n377;
wire n378, n379, n380, n381, n382, n383, n384, n385, n386, n387;
wire n388, n389, n390, n391, n392, n393, n394, n395, n396, n397;
wire n398, n399, n400, n401, n402, n403, n404, n405, n406, n407;
wire n408, n409, n410, n411, n412, n413, n414, n415, n416, n417;
wire n418, n419, n420, n421, n422, n423, n424, n425, n426, n427;
wire n428, n429, n430, n431, n432, n433, n434, n435, n436, n437;
wire n438, n439, n440, n441, n442, n443, n444, n445, n446, n447;
wire n448, n449, n450, n451, n452, n453, n454, n455, n456, n457;
wire n458, n459, n460, n461, n462, n463, n464, n465, n466, n467;
wire n468, n469, n470, n471, n472, n473, n474, n475, n476, n477;
wire n478, n479, n480, n481, n482, n483, n484, n485, n486, n487;
wire n488, n489, n490, n491, n492, n493, n494, n495, n496, n497;
wire n498, n499, n500, n501, n502, n503, n504, n505, n506, n507;
wire n508, n509, n510, n511, n512, n513, n514, n515, n516, n517;
wire n518, n519, n520, n521, n522, n523, n524, n525, n526, n527;
wire n528, n529, n530, n531, n532, n533, n534, n535, n536, n537;
wire n538, n539, n540, n541, n542, n543, n544, n545, n546, n547;
wire n548, n549, n550, n551, n552, n553, n554, n555, n556, n557;
wire n558, n559, n560, n561, n562, n563, n564, n565, n566, n567;
wire n568, n569, n570, n571, n572, n573, n574, n575, n576, n577;
wire n578, n579, n580, n581, n582, n583, n584, n585, n586, n587;
wire n588, n589, n590, n591, n592, n593;
reg read_e = 0, n10 = 0, write_e = 0, n19 = 0, n27 = 0, n29 = 0, n30 = 0, n31 = 0, n32 = 0, n34 = 0;
reg n36 = 0, n37 = 0, n41 = 0, n46 = 0, n55 = 0, n56 = 0, n68 = 0, n70 = 0, n71 = 0, n74 = 0;
reg n89 = 0, n90 = 0, n91 = 0, n95 = 0, n96 = 0, n101 = 0, n105 = 0, n106 = 0, n109 = 0, n110 = 0;
reg n111 = 0, n133 = 0, n156 = 0, n157 = 0, n170 = 0, n171 = 0, n181 = 0, n195 = 0, n200 = 0, n233 = 0;
reg n234 = 0, n252 = 0, n253 = 0, n255 = 0, n256 = 0, n257 = 0, n258 = 0, n259 = 0, n260 = 0, n266 = 0;
reg n267 = 0, n268 = 0, n273 = 0, n274 = 0, n275 = 0, n290 = 0, n291 = 0, n292 = 0, n293 = 0, n296 = 0;
assign n356 = 1;
assign n419 = 1;
assign n425 = 1;
assign n443 = 1;
assign n482 = 1;
assign n514 = 1;
assign n552 = 1;

SB_RAM40_4K #(
  .READ_MODE(0),
  .WRITE_MODE(0),
  .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
) ram40_8_25 (
  .WADDR({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n101, n19, n74, n34}),
  .RADDR({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n97, n20, n98, n73}),
  .MASK({n38, n38, n38, n38, n38, n66, n66, n66, n66, n66, n66, n66, n66, n66, n66, n66}),
  .WDATA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n56, n32, n29, n55, n36, n37, n27, n89, n30, n31, n10}),
  .RDATA({open_0, open_1, open_2, open_3, open_4, n18, n72, n63, n82, n83, n84, n85, n86, n87, n81, n75}),
  .WE(n38),
  .WCLKE(n43),
  .WCLK(clk),
  .RE(n38),
  .RCLKE(1'b1),
  .RCLK(clk)
);

SB_RAM40_4K #(
  .READ_MODE(3),
  .WRITE_MODE(3),
  .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
) ram40_8_23 (
  .WADDR({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RADDR({n56, n32, n29, n55, n36, n37, n27, n89, n30, n31, n10}),
  .MASK({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .WDATA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RDATA({open_13, open_14, open_15, open_16, n65, open_17, open_18, open_19, open_20, open_21, open_22, open_23, n61, open_25, open_26, open_27}),
  .WE(n38),
  .WCLKE(n79),
  .WCLK(1'b0),
  .RE(n38),
  .RCLKE(1'b1),
  .RCLK(clk)
);

SB_RAM40_4K #(
  .READ_MODE(3),
  .WRITE_MODE(3),
  .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
) ram40_8_21 (
  .WADDR({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RADDR({n56, n32, n29, n55, n36, n37, n27, n89, n30, n31, n10}),
  .MASK({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .WDATA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RDATA({open_28, open_29, open_30, open_31, n57, open_32, open_33, open_34, open_35, open_36, open_37, open_38, n58, open_40, open_41, open_42}),
  .WE(n38),
  .WCLKE(n79),
  .WCLK(1'b0),
  .RE(n38),
  .RCLKE(1'b1),
  .RCLK(clk)
);

SB_RAM40_4K #(
  .READ_MODE(3),
  .WRITE_MODE(3),
  .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
) ram40_25_25 (
  .WADDR({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RADDR({n56, n32, n29, n55, n36, n37, n27, n89, n30, n31, n10}),
  .MASK({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .WDATA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RDATA({open_43, open_44, open_45, open_46, n62, open_47, open_48, open_49, open_50, open_51, open_52, open_53, n245, open_55, open_56, open_57}),
  .WE(n38),
  .WCLKE(n79),
  .WCLK(1'b0),
  .RE(n38),
  .RCLKE(1'b1),
  .RCLK(clk)
);

SB_RAM40_4K #(
  .READ_MODE(3),
  .WRITE_MODE(3),
  .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
) ram40_8_19 (
  .WADDR({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RADDR({n56, n32, n29, n55, n36, n37, n27, n89, n30, n31, n10}),
  .MASK({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .WDATA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RDATA({open_58, open_59, open_60, open_61, n76, open_62, open_63, open_64, open_65, open_66, open_67, open_68, n77, open_70, open_71, open_72}),
  .WE(n38),
  .WCLKE(n79),
  .WCLK(1'b0),
  .RE(n38),
  .RCLKE(1'b1),
  .RCLK(clk)
);

SB_RAM40_4K #(
  .READ_MODE(3),
  .WRITE_MODE(3),
  .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
) ram40_25_21 (
  .WADDR({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RADDR({n56, n32, n29, n55, n36, n37, n27, n89, n30, n31, n10}),
  .MASK({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .WDATA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RDATA({open_73, open_74, open_75, open_76, n54, open_77, open_78, open_79, open_80, open_81, open_82, open_83, n297, open_85, open_86, open_87}),
  .WE(n38),
  .WCLKE(n79),
  .WCLK(1'b0),
  .RE(n38),
  .RCLKE(1'b1),
  .RCLK(clk)
);

SB_RAM40_4K #(
  .READ_MODE(3),
  .WRITE_MODE(3),
  .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
) ram40_25_23 (
  .WADDR({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RADDR({n56, n32, n29, n55, n36, n37, n27, n89, n30, n31, n10}),
  .MASK({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .WDATA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RDATA({open_88, open_89, open_90, open_91, n298, open_92, open_93, open_94, open_95, open_96, open_97, open_98, n59, open_100, open_101, open_102}),
  .WE(n38),
  .WCLKE(n79),
  .WCLK(1'b0),
  .RE(n38),
  .RCLKE(1'b1),
  .RCLK(clk)
);

SB_RAM40_4K #(
  .READ_MODE(3),
  .WRITE_MODE(3),
  .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
) ram40_25_19 (
  .WADDR({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RADDR({n56, n32, n29, n55, n36, n37, n27, n89, n30, n31, n10}),
  .MASK({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .WDATA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RDATA({open_103, open_104, open_105, open_106, n299, open_107, open_108, open_109, open_110, open_111, open_112, open_113, n53, open_115, open_116, open_117}),
  .WE(n38),
  .WCLKE(n79),
  .WCLK(1'b0),
  .RE(n38),
  .RCLKE(1'b1),
  .RCLK(clk)
);

SB_RAM40_4K #(
  .READ_MODE(3),
  .WRITE_MODE(3),
  .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
) ram40_8_27 (
  .WADDR({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RADDR({n56, n32, n29, n55, n36, n37, n27, n89, n30, n31, n10}),
  .MASK({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .WDATA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RDATA({open_118, open_119, open_120, open_121, n67, open_122, open_123, open_124, open_125, open_126, open_127, open_128, n24, open_130, open_131, open_132}),
  .WE(n38),
  .WCLKE(n79),
  .WCLK(1'b0),
  .RE(n38),
  .RCLKE(1'b1),
  .RCLK(clk)
);

assign n338 = /* LUT   15 28  1 */ 1'b0;
assign n345 = /* LUT   15 28  3 */ 1'b0;
assign n355 = /* LUT   11 27  0 */ 1'b0;
assign n361 = /* LUT   12 24  1 */ 1'b0;
assign n406 = /* LUT   13 20  1 */ 1'b0;
assign n410 = /* LUT   14 26  2 */ 1'b0;
assign n418 = /* LUT   14 26  0 */ 1'b0;
assign n424 = /* LUT   14 23  0 */ 1'b0;
assign n442 = /* LUT   11 26  0 */ 1'b0;
assign n481 = /* LUT   15 28  0 */ 1'b0;
assign n488 = /* LUT   15 28  2 */ 1'b0;
assign n496 = /* LUT   11 27  1 */ 1'b0;
assign n513 = /* LUT   12 24  0 */ 1'b0;
assign n545 = /* LUT   20 22  7 */ 1'b0;
assign n551 = /* LUT   13 20  0 */ 1'b0;
assign n558 = /* LUT   14 26  3 */ 1'b0;
assign n564 = /* LUT   14 26  1 */ 1'b0;
assign n574 = /* LUT   14 23  1 */ 1'b0;
assign n590 = /* LUT   11 26  1 */ 1'b0;
assign n311 = /* LUT   14 21  4 */ (n228 ? (n41 ? 1'b0 : !n156) : 1'b0);
assign n312 = /* LUT   15 20  2 */ (n53 ? (n123 ? (n269 ? !n54 : 1'b0) : 1'b0) : 1'b0);
assign n313 = /* LUT    9 25  0 */ (n71 ? n96 : n87);
assign n314 = /* LUT   17 22  5 */ (n298 ? !n297 : 1'b0);
assign n315 = /* LUT   12 23  4 */ (n69 ? (n92 ? n133 : 1'b1) : !n24);
assign n316 = /* LUT   11 26  7 */ (n114 ? (n66 ? n130 : n19) : n19);
assign n317 = /* LUT    7 21  2 */ (n77 ? n41 : 1'b0);
assign n318 = /* LUT   12 25  2 */ (n210 ? !n50 : n50);
assign n319 = /* LUT   14 21  2 */ (n267 ? 1'b0 : (n41 ? 1'b0 : !n156));
assign n320 = /* LUT   15 20  4 */ (n53 ? (n54 ? (n269 ? n123 : 1'b0) : 1'b0) : 1'b0);
assign n321 = /* LUT   14 24  0 */ (n283 ? !n29 : n29);
assign n322 = /* LUT   13 24  1 */ (n57 ? (n69 ? (n165 ? !n133 : 1'b1) : 1'b0) : (n165 ? !n133 : 1'b1));
assign n323 = /* LUT   11 26  5 */ (n114 ? (n66 ? n129 : n101) : n101);
assign n324 = /* LUT   15 25  1 */ (n64 ? (n196 ? n244 : 1'b0) : 1'b0);
assign n325 = /* LUT   15 21  7 */ (n254 ? (n231 ? (n217 ? !n263 : 1'b1) : 1'b1) : 1'b1);
assign n326 = /* LUT   15 20  6 */ (n53 ? (n244 ? (n269 ? !n54 : 1'b0) : 1'b0) : 1'b0);
assign n327 = /* LUT   14 21  0 */ (n229 ? (n230 ? !n228 : 1'b0) : 1'b0);
assign n328 = /* LUT   14 24  2 */ (n285 ? !n56 : n56);
assign n329 = /* LUT   15 19  7 */ (n53 ? (n64 ? (n102 ? !n54 : 1'b0) : 1'b0) : 1'b0);
assign n330 = /* LUT   10 26  5 */ (rst ? !n74 : !n51);
assign n331 = /* LUT   13 21  7 */ (n192 ? !n193 : 1'b1);
assign n332 = /* LUT   15 21  5 */ (n64 ? (n54 ? (n102 ? !n53 : 1'b0) : 1'b0) : 1'b0);
assign n333 = /* LUT    9 25  6 */ n55;
assign n334 = /* LUT   17 22  3 */ (n297 ? n298 : 1'b0);
assign n335 = /* LUT   14 24  4 */ (n59 ? (n69 ? (n167 ? !n133 : 1'b1) : 1'b0) : (n167 ? !n133 : 1'b1));
assign n336 = /* LUT   15 19  1 */ (n53 ? (n64 ? (n161 ? !n54 : 1'b0) : 1'b0) : 1'b0);
assign n339 = /* LUT   14 19  0 */ (n251 ? !n252 : 1'b0);
assign n340 = /* LUT   14 22  6 */ n276;
assign n341 = /* LUT   11 18  6 */ (n39 ? !n115 : 1'b0);
assign n342 = /* LUT   15 21  3 */ (n90 ? (n291 ? 1'b0 : !n233) : (n291 ? 1'b0 : !n266));
assign n343 = /* LUT   15 22  3 */ (n233 ? 1'b0 : (n275 ? 1'b0 : (read_e ? 1'b0 : !n274)));
assign n346 = /* LUT   14 19  2 */ (n214 ? (n121 ? 1'b0 : !n212) : 1'b0);
assign n347 = /* LUT   10 24  4 */ n27;
assign n348 = /* LUT   13 19  2 */ (n46 ? n211 : (n212 ? 1'b0 : (n211 ? 1'b1 : !n181)));
assign n349 = /* LUT   14 22  4 */ n239;
assign n350 = /* LUT   16 21  5 */ (n53 ? (n54 ? (n64 ? n244 : 1'b0) : 1'b0) : 1'b0);
assign n351 = /* LUT   12 24  3 */ (n203 ? !n169 : n169);
assign n352 = /* LUT   15 21  1 */ (n292 ? 1'b0 : (n290 ? 1'b0 : (n133 ? 1'b0 : !n195)));
assign n353 = /* LUT   15 22  1 */ (n264 ? (n157 ? !n274 : !n293) : 1'b0);
assign n357 = /* LUT    7 26  7 */ n43;
assign n358 = /* LUT   14 19  4 */ (n251 ? (n252 ? 1'b1 : (n46 ? 1'b0 : !n253)) : (n252 ? 1'b1 : (n46 ? 1'b1 : n253)));
assign n359 = /* LUT   10 24  6 */ n36;
assign n362 = /* LUT   15 27  4 */ !n34;
assign n363 = /* LUT   16 21  7 */ (n53 ? (n54 ? (n102 ? n269 : 1'b0) : 1'b0) : 1'b0);
assign n364 = /* LUT   13 19  0 */ (n185 ? (n154 ? !n182 : 1'b1) : 1'b0);
assign n365 = /* LUT   14 20  5 */ (n229 ? (n232 ? 1'b0 : !n195) : 1'b0);
assign n366 = /* LUT   15 22  7 */ (n53 ? (n54 ? (n269 ? n244 : 1'b0) : 1'b0) : 1'b0);
assign n367 = /* LUT   12 22  5 */ (n61 ? !n41 : 1'b1);
assign n368 = /* LUT   11 27  2 */ (n179 ? !n19 : n19);
assign n369 = /* LUT   15 28  7 */ !n19;
assign n370 = /* LUT   14 19  6 */ (n214 ? (n212 ? n255 : 1'b1) : 1'b0);
assign n371 = /* LUT   16 21  1 */ (n269 ? (n54 ? (n102 ? !n53 : 1'b0) : 1'b0) : 1'b0);
assign n372 = /* LUT   12 24  7 */ (n207 ? !n94 : n94);
assign n373 = /* LUT   14 20  7 */ (n230 ? !n232 : 1'b0);
assign n374 = /* LUT    9 26  1 */ (n100 ? !rst : 1'b0);
assign n375 = /* LUT   15 22  5 */ (n53 ? (n54 ? (n161 ? n269 : 1'b0) : 1'b0) : 1'b0);
assign n376 = /* LUT   12 19  4 */ (n143 ? 1'b0 : (n40 ? n47 : 1'b1));
assign n377 = /* LUT   13 19  4 */ (n143 ? 1'b0 : (n40 ? n194 : 1'b1));
assign n378 = /* LUT   10 24  2 */ (n71 ? n105 : n85);
assign n379 = /* LUT   12 24  5 */ (n205 ? !n80 : n80);
assign n380 = /* LUT   14 20  1 */ !n220;
assign n381 = /* LUT    7 25  1 */ 1'b1;
assign n382 = /* LUT   13 25  2 */ (n248 ? (n166 ? n133 : 1'b0) : 1'b1);
assign n383 = /* LUT   11 27  6 */ (n173 ? n135 : n131);
assign n384 = /* LUT   12 19  2 */ (n52 ? (n151 ? (n39 ? n149 : 1'b1) : 1'b0) : (n39 ? n149 : 1'b1));
assign n385 = /* LUT   11 19  1 */ (n118 ? (n39 ? !n138 : 1'b0) : 1'b1);
assign n386 = /* LUT   14 20  3 */ n28;
assign n387 = /* LUT    9 26  5 */ (n99 ? (n112 ? (n19 ? !n20 : n20) : 1'b1) : 1'b1);
assign n388 = /* LUT   13 23  7 */ (n199 ? (n163 ? n133 : 1'b0) : 1'b1);
assign n389 = /* LUT   12 19  0 */ (n35 ? (n142 ? (n115 ? n121 : 1'b0) : 1'b0) : 1'b0);
assign n390 = /* LUT   13 22  6 */ (n57 ? !n41 : 1'b1);
assign n391 = /* LUT   11 19  3 */ (n119 ? (n52 ? !n142 : 1'b0) : 1'b1);
assign n392 = /* LUT   12 26  4 */ (n34 ? (n66 ? 1'b0 : n178) : (n66 ? n114 : 1'b0));
assign n393 = /* LUT    9 26  7 */ n100;
assign n394 = /* LUT    6 24  6 */ (n61 ? !n45 : 1'b0);
assign n395 = /* LUT   11 19  5 */ (n52 ? (n144 ? (n39 ? n35 : 1'b1) : 1'b0) : (n39 ? n35 : 1'b1));
assign n396 = /* LUT   12 26  6 */ !n34;
assign n397 = /* LUT   17 21  5 */ (n296 ? n299 : 1'b0);
assign n398 = /* LUT   13 23  3 */ (n69 ? (n236 ? n133 : 1'b1) : !n61);
assign n399 = /* LUT   13 20  3 */ (n223 ? !n194 : n194);
assign n400 = /* LUT   11 19  7 */ (n117 ? (n52 ? !n121 : 1'b0) : 1'b1);
assign n401 = /* LUT   12 26  0 */ (n114 ? (n66 ? n174 : n34) : n34);
assign n402 = /* LUT   14 26  4 */ (n286 ? 1'b0 : (n64 ? (n196 ? !n244 : 1'b1) : 1'b1));
assign n403 = /* LUT   17 21  7 */ n268;
assign n404 = /* LUT   14 25  2 */ (n62 ? (n69 ? (n88 ? !n133 : 1'b1) : 1'b0) : (n88 ? !n133 : 1'b1));
assign n407 = /* LUT   14 23  4 */ (n279 ? !n27 : n27);
assign n408 = /* LUT   12 26  2 */ (n173 ? (rst ? 1'b0 : n175) : (rst ? 1'b0 : n172));
assign n411 = /* LUT    9 24  6 */ (n71 ? n91 : n84);
assign n412 = /* LUT   11 24  3 */ (n69 ? (n31 ? 1'b1 : n133) : !n76);
assign n413 = /* LUT   12 18  5 */ (n137 ? (n39 ? !n151 : 1'b0) : 1'b1);
assign n414 = /* LUT   13 20  7 */ (n227 ? !n122 : n122);
assign n415 = /* LUT   14 23  6 */ (n281 ? !n36 : n36);
assign n416 = /* LUT   12 20  7 */ (n145 ? (n154 ? !n189 : 1'b1) : 1'b0);
assign n420 = /* LUT   12 21  6 */ (n58 ? !n41 : 1'b1);
assign n421 = /* LUT   14 25  6 */ (n69 ? (n240 ? n133 : 1'b1) : !n245);
assign n422 = /* LUT   13 20  5 */ (n225 ? !n191 : n191);
assign n426 = /* LUT   12 20  5 */ (n147 ? (n154 ? !n190 : 1'b1) : 1'b0);
assign n427 = /* LUT   11 25  6 */ (n125 ? (n127 ? n133 : 1'b0) : 1'b1);
assign n428 = /* LUT   14 25  4 */ (n69 ? !n133 : 1'b0);
assign n429 = /* LUT   10 25  6 */ n10;
assign n430 = /* LUT   16 22  5 */ (n53 ? 1'b0 : !n54);
assign n431 = /* LUT   14 23  2 */ (n277 ? !n30 : n30);
assign n432 = /* LUT   12 20  3 */ (n143 ? 1'b0 : (n40 ? n122 : 1'b1));
assign n433 = /* LUT   11 26  2 */ n176;
assign n434 = /* LUT    7 21  7 */ (n76 ? !n41 : 1'b1);
assign n435 = /* LUT   13 24  6 */ (n201 ? (n238 ? n246 : 1'b0) : 1'b1);
assign n436 = /* LUT   10 25  4 */ n56;
assign n437 = /* LUT    6 28  4 */ (n67 ? !n45 : 1'b0);
assign n438 = /* LUT   12 25  5 */ n89;
assign n439 = /* LUT   12 20  1 */ (n146 ? (n154 ? !n186 : 1'b1) : 1'b0);
assign n440 = /* LUT   11 25  2 */ !n108;
assign n444 = /* LUT   13 24  4 */ (n197 ? (n60 ? n133 : 1'b0) : 1'b1);
assign n445 = /* LUT   10 25  2 */ (n71 ? n109 : n18);
assign n446 = /* LUT   12 25  7 */ n29;
assign n447 = /* LUT   16 22  1 */ (n269 ? (n123 ? n196 : 1'b0) : 1'b0);
assign n448 = /* LUT   14 21  7 */ (n102 ? (n64 ? n196 : 1'b0) : 1'b0);
assign n449 = /* LUT   15 20  1 */ (n123 ? (n54 ? (n269 ? !n53 : 1'b0) : 1'b0) : 1'b0);
assign n450 = /* LUT   11 25  0 */ (n69 ? (n126 ? n133 : 1'b1) : !n77);
assign n451 = /* LUT   17 22  4 */ (n297 ? !n298 : 1'b0);
assign n452 = /* LUT   12 23  7 */ (n159 ? (n162 ? n133 : 1'b0) : 1'b1);
assign n453 = /* LUT   11 26  6 */ (n173 ? n134 : n132);
assign n454 = /* LUT   10 26  2 */ (n113 ? (n34 ? n73 : !n73) : 1'b0);
assign n455 = /* LUT   10 25  0 */ (n71 ? n110 : n72);
assign n456 = /* LUT   12 25  1 */ (n209 ? !n107 : n107);
assign n457 = /* LUT   15 26  2 */ (n244 ? (n64 ? (n196 ? !n288 : 1'b0) : 1'b0) : 1'b0);
assign n458 = /* LUT   14 21  5 */ (n68 ? 1'b0 : (n41 ? 1'b0 : (n156 ? 1'b0 : !n256)));
assign n459 = /* LUT   15 20  3 */ (n53 ? (n64 ? (n123 ? !n54 : 1'b0) : 1'b0) : 1'b0);
assign n460 = /* LUT   14 24  1 */ (n284 ? !n32 : n32);
assign n461 = /* LUT   12 23  5 */ (n69 ? (n48 ? n133 : 1'b1) : !n58);
assign n462 = /* LUT   13 24  0 */ (n1 ? (n246 ? n10 : 1'b1) : 1'b0);
assign n463 = /* LUT   11 26  4 */ (n128 ? n19 : !n19);
assign n464 = /* LUT    6 26  2 */ (n65 ? !n45 : 1'b0);
assign n465 = /* LUT   13 21  2 */ (n152 ? (n153 ? (n155 ? !n28 : 1'b0) : 1'b0) : 1'b0);
assign n466 = /* LUT   14 22  3 */ (write_e ? 1'b0 : (read_e ? 1'b0 : (n239 ? 1'b0 : !n276)));
assign n467 = /* LUT   12 25  3 */ (n71 ? n171 : n63);
assign n468 = /* LUT   15 20  5 */ (n64 ? (n54 ? (n123 ? !n53 : 1'b0) : 1'b0) : 1'b0);
assign n469 = /* LUT   14 21  3 */ (n260 ? 1'b0 : (n68 ? 1'b0 : (n195 ? 1'b0 : !n256)));
assign n470 = /* LUT    9 25  5 */ (n71 ? n95 : n82);
assign n471 = /* LUT   15 19  4 */ (n53 ? (n244 ? (n64 ? !n54 : 1'b0) : 1'b0) : 1'b0);
assign n472 = /* LUT   10 26  6 */ n33;
assign n473 = /* LUT   13 21  4 */ (n139 ? n148 : 1'b0);
assign n474 = /* LUT   15 21  6 */ (n53 ? (n269 ? (n161 ? !n54 : 1'b0) : 1'b0) : 1'b0);
assign n475 = /* LUT   15 20  7 */ (n53 ? (n269 ? (n102 ? !n54 : 1'b0) : 1'b0) : 1'b0);
assign n476 = /* LUT    9 25  7 */ n30;
assign n477 = /* LUT   17 22  2 */ (n297 ? 1'b0 : !n298);
assign n478 = /* LUT   14 24  5 */ (n247 ? (n241 ? n246 : 1'b0) : 1'b1);
assign n479 = /* LUT   14 21  1 */ (n267 ? 1'b0 : !n234);
assign n483 = /* LUT   15 21  4 */ (n270 ? (n68 ? 1'b0 : (n291 ? 1'b0 : !write_e)) : 1'b0);
assign n484 = /* LUT   15 22  2 */ (n261 ? (n157 ? !n200 : !n275) : 1'b0);
assign n485 = /* LUT   14 24  7 */ (n243 ? (n242 ? n246 : 1'b0) : 1'b1);
assign n486 = /* LUT   15 19  0 */ (n181 ? 1'b0 : !n258);
assign n489 = /* LUT   14 19  1 */ (n253 ? 1'b0 : !n252);
assign n490 = /* LUT   13 19  3 */ (n212 ? (n181 ? !n46 : 1'b0) : 1'b0);
assign n491 = /* LUT   15 21  2 */ (n272 ? (n262 ? n265 : 1'b0) : 1'b0);
assign n492 = /* LUT   15 22  0 */ (n293 ? 1'b0 : (n200 ? 1'b0 : (n273 ? 1'b0 : !n266)));
assign n493 = /* LUT    7 26  6 */ (n77 ? !n45 : 1'b0);
assign n494 = /* LUT   15 19  2 */ (n53 ? (n54 ? (n161 ? n64 : 1'b0) : 1'b0) : 1'b0);
assign n497 = /* LUT   15 28  4 */ n294;
assign n498 = /* LUT   14 19  3 */ (n46 ? 1'b0 : !n181);
assign n499 = /* LUT   13 19  1 */ (n140 ? (n211 ? n46 : n213) : 1'b1);
assign n500 = /* LUT   16 21  6 */ (n244 ? (n54 ? (n269 ? !n53 : 1'b0) : 1'b0) : 1'b0);
assign n501 = /* LUT   12 24  2 */ (n202 ? !n93 : n93);
assign n502 = /* LUT   11 18  5 */ (n116 ? 1'b1 : (n136 ? 1'b1 : (n138 ? 1'b0 : n52)));
assign n503 = /* LUT   15 21  0 */ (n90 ? (n257 ? 1'b0 : !n292) : (n257 ? 1'b0 : !n259));
assign n504 = /* LUT   15 22  6 */ (n123 ? (n64 ? n196 : 1'b0) : 1'b0);
assign n505 = /* LUT    7 26  4 */ (n33 ? !rst : 1'b0);
assign n506 = /* LUT   11 27  3 */ (n180 ? !n101 : n101);
assign n507 = /* LUT   14 19  5 */ (n212 ? (n46 ? 1'b0 : (n181 ? 1'b0 : !n251)) : 1'b0);
assign n508 = /* LUT   13 19  7 */ (n184 ? (n154 ? !n187 : 1'b1) : 1'b0);
assign n509 = /* LUT   16 21  0 */ (n161 ? (n64 ? n196 : 1'b0) : 1'b0);
assign n510 = /* LUT   10 24  1 */ (n71 ? n106 : n83);
assign n511 = /* LUT   14 20  4 */ !n28;
assign n515 = /* LUT   15 22  4 */ (n102 ? (n269 ? n196 : 1'b0) : 1'b0);
assign n516 = /* LUT   11 27  5 */ (n173 ? (rst ? 1'b0 : n135) : (rst ? 1'b0 : n131));
assign n517 = /* LUT   14 19  7 */ (n215 ? !n216 : 1'b0);
assign n518 = /* LUT   13 19  5 */ (n143 ? 1'b0 : (n40 ? n191 : 1'b1));
assign n519 = /* LUT   16 21  2 */ (n244 ? (n54 ? (n64 ? !n53 : 1'b0) : 1'b0) : 1'b0);
assign n520 = /* LUT   12 24  6 */ (n206 ? !n103 : n103);
assign n521 = /* LUT   14 20  6 */ (n229 ? (n230 ? (n218 ? 1'b0 : !n219) : !n218) : (n230 ? !n219 : 1'b0));
assign n522 = /* LUT    9 26  2 */ !n66;
assign n523 = /* LUT    7 25  2 */ n31;
assign n524 = /* LUT   13 22  3 */ (n65 ? !n41 : 1'b1);
assign n525 = /* LUT    6 24  3 */ (n57 ? !n45 : 1'b0);
assign n526 = /* LUT   12 19  5 */ (n150 ? !n143 : 1'b0);
assign n527 = /* LUT   12 24  4 */ (n204 ? !n104 : n104);
assign n528 = /* LUT   14 20  0 */ (n214 ? (n212 ? (n260 ? 1'b0 : !n256) : 1'b0) : 1'b0);
assign n529 = /* LUT    9 26  4 */ (n101 ? n97 : !n97);
assign n530 = /* LUT    7 25  0 */ (n71 ? n70 : n81);
assign n531 = /* LUT   14 27  2 */ !n101;
assign n532 = /* LUT   12 19  3 */ (n39 ? (n121 ? (n78 ? n142 : 1'b1) : 1'b0) : (n78 ? n142 : 1'b1));
assign n533 = /* LUT   13 22  5 */ (n67 ? !n41 : 1'b1);
assign n534 = /* LUT   11 19  0 */ (n78 ? (n144 ? (n39 ? n142 : 1'b1) : 1'b0) : (n39 ? n142 : 1'b1));
assign n535 = /* LUT   12 26  5 */ !n34;
assign n536 = /* LUT   14 20  2 */ (n143 ? 1'b0 : (n232 ? 1'b1 : (n221 ? !n195 : 1'b0)));
assign n537 = /* LUT    9 26  6 */ (n74 ? !n51 : n51);
assign n538 = /* LUT   13 23  6 */ (n69 ? (n237 ? n133 : 1'b1) : !n65);
assign n539 = /* LUT   12 19  1 */ (n141 ? (n183 ? 1'b1 : (n149 ? 1'b0 : n52)) : 1'b1);
assign n540 = /* LUT   11 19  2 */ (n78 ? (n115 ? (n52 ? n35 : 1'b1) : 1'b0) : (n52 ? n35 : 1'b1));
assign n541 = /* LUT    7 28  2 */ (n24 ? !n45 : 1'b0);
assign n542 = /* LUT   12 26  7 */ (n173 ? n175 : n172);
assign n543 = /* LUT   14 28  7 */ !n74;
assign n544 = /* LUT   13 20  2 */ (n222 ? !n153 : n153);
assign n546 = /* LUT   11 19  4 */ (n39 ? (n144 ? (n78 ? n35 : 1'b1) : 1'b0) : (n78 ? n35 : 1'b1));
assign n547 = /* LUT   17 21  4 */ (n296 ? !n299 : 1'b0);
assign n548 = /* LUT    7 27  5 */ (n76 ? !n45 : 1'b0);
assign n549 = /* LUT    6 23  2 */ (n58 ? !n45 : 1'b0);
assign n553 = /* LUT   11 19  6 */ (n120 ? (n78 ? !n138 : 1'b0) : 1'b1);
assign n554 = /* LUT   12 26  3 */ (n178 ? !n66 : 1'b0);
assign n555 = /* LUT   15 23  5 */ (n66 ? n271 : 1'b0);
assign n556 = /* LUT   12 21  3 */ (n24 ? !n41 : 1'b1);
assign n559 = /* LUT   17 21  6 */ (n296 ? n295 : 1'b0);
assign n560 = /* LUT   13 23  0 */ (n69 ? (n235 ? n133 : 1'b1) : !n67);
assign n561 = /* LUT   13 20  6 */ (n226 ? !n152 : n152);
assign n562 = /* LUT   14 23  5 */ (n280 ? !n37 : n37);
assign n565 = /* LUT   17 21  0 */ (n296 ? 1'b0 : !n268);
assign n566 = /* LUT    9 24  7 */ n37;
assign n567 = /* LUT   12 18  4 */ (n52 ? (n115 ? (n78 ? n149 : 1'b1) : 1'b0) : (n78 ? n149 : 1'b1));
assign n568 = /* LUT   13 20  4 */ (n224 ? !n155 : n155);
assign n569 = /* LUT   14 23  7 */ (n282 ? !n55 : n55);
assign n570 = /* LUT   12 20  6 */ (n188 ? (n154 ? 1'b0 : (n40 ? n155 : 1'b1)) : (n40 ? n155 : 1'b1));
assign n571 = /* LUT   17 21  2 */ (n53 ? (n297 ? (n54 ? n299 : 1'b0) : 1'b0) : (n297 ? 1'b0 : (n54 ? 1'b0 : !n299)));
assign n572 = /* LUT   11 24  6 */ (n133 ? (n108 ? (n42 ? !n124 : 1'b1) : (n42 ? 1'b1 : !n124)) : !n124);
assign n575 = /* LUT   12 20  4 */ (n144 ? (n149 ? (n150 ? n151 : 1'b0) : 1'b0) : 1'b0);
assign n576 = /* LUT   16 22  4 */ (n269 ? (n54 ? (n161 ? !n53 : 1'b0) : 1'b0) : 1'b0);
assign n577 = /* LUT   12 25  4 */ (n71 ? n170 : n86);
assign n578 = /* LUT   14 23  3 */ (n278 ? !n89 : n89);
assign n579 = /* LUT   12 20  2 */ (n143 ? 1'b0 : (n40 ? n153 : 1'b1));
assign n580 = /* LUT   13 24  7 */ (n198 ? (n49 ? n133 : 1'b0) : 1'b1);
assign n581 = /* LUT   11 26  3 */ (n177 ? n101 : !n101);
assign n582 = /* LUT   12 18  2 */ (n78 ? !n151 : 1'b0);
assign n583 = /* LUT   10 25  5 */ n32;
assign n584 = /* LUT   16 22  6 */ (n64 ? (n54 ? (n161 ? !n53 : 1'b0) : 1'b0) : 1'b0);
assign n585 = /* LUT   15 20  0 */ (n257 ? 1'b0 : (n258 ? 1'b0 : (n255 ? 1'b0 : !n259)));
assign n586 = /* LUT   12 20  0 */ (n143 ? 1'b0 : (n40 ? n152 : 1'b1));
assign n587 = /* LUT   11 25  1 */ !n10;
assign n588 = /* LUT   12 23  6 */ (n160 ? (n164 ? n133 : 1'b0) : 1'b1);
assign n591 = /* LUT   13 21  1 */ (n122 ? (n191 ? (n47 ? n194 : 1'b0) : 1'b0) : 1'b0);
assign n592 = /* LUT   10 25  3 */ (n71 ? n111 : n75);
assign n593 = /* LUT   12 25  0 */ (n208 ? !n168 : n168);
assign n284 = /* CARRY 14 24  0 */ (1'b0 & n29) | ((1'b0 | n29) & n283);
assign n300 = /* CARRY 15 28  1 */ (1'b0 & n250) | ((1'b0 | n250) & n306);
assign n294 = /* CARRY 15 28  3 */ (1'b0 & n249) | ((1'b0 | n249) & n307);
assign n204 = /* CARRY 12 24  3 */ (1'b0 & n169) | ((1'b0 | n169) & n203);
assign n301 = /* CARRY 11 27  0 */ (n34 & 1'b0) | ((n34 | 1'b0) & n356);
assign n202 = /* CARRY 12 24  1 */ (1'b0 & n42) | ((1'b0 | n42) & n308);
assign n180 = /* CARRY 11 27  2 */ (1'b0 & n19) | ((1'b0 | n19) & n179);
assign n208 = /* CARRY 12 24  7 */ (1'b0 & n94) | ((1'b0 | n94) & n207);
assign n206 = /* CARRY 12 24  5 */ (1'b0 & n80) | ((1'b0 | n80) & n205);
assign n224 = /* CARRY 13 20  3 */ (1'b0 & n194) | ((1'b0 | n194) & n223);
assign n222 = /* CARRY 13 20  1 */ (1'b0 & n47) | ((1'b0 | n47) & n309);
assign n280 = /* CARRY 14 23  4 */ (1'b0 & n27) | ((1'b0 | n27) & n279);
assign n302 = /* CARRY 14 26  2 */ (n19 & 1'b0) | ((n19 | 1'b0) & n310);
assign n282 = /* CARRY 14 23  6 */ (1'b0 & n36) | ((1'b0 | n36) & n281);
assign n303 = /* CARRY 14 26  0 */ (n34 & 1'b0) | ((n34 | 1'b0) & n419);
assign n226 = /* CARRY 13 20  5 */ (1'b0 & n191) | ((1'b0 | n191) & n225);
assign n304 = /* CARRY 14 23  0 */ (n10 & 1'b0) | ((n10 | 1'b0) & n425);
assign n278 = /* CARRY 14 23  2 */ (1'b0 & n30) | ((1'b0 | n30) & n277);
assign n177 = /* CARRY 11 26  2 */ (n19 & n38) | ((n19 | n38) & n176);
assign n305 = /* CARRY 11 26  0 */ (n34 & 1'b0) | ((n34 | 1'b0) & n443);
assign n210 = /* CARRY 12 25  1 */ (1'b0 & n107) | ((1'b0 | n107) & n209);
assign n285 = /* CARRY 14 24  1 */ (1'b0 & n32) | ((1'b0 | n32) & n284);
assign n306 = /* CARRY 15 28  0 */ (n287 & 1'b0) | ((n287 | 1'b0) & n482);
assign n307 = /* CARRY 15 28  2 */ (1'b0 & n289) | ((1'b0 | n289) & n300);
assign n179 = /* CARRY 11 27  1 */ (1'b0 & n74) | ((1'b0 | n74) & n301);
assign n203 = /* CARRY 12 24  2 */ (1'b0 & n93) | ((1'b0 | n93) & n202);
assign n308 = /* CARRY 12 24  0 */ (n108 & 1'b0) | ((n108 | 1'b0) & n514);
assign n207 = /* CARRY 12 24  6 */ (1'b0 & n103) | ((1'b0 | n103) & n206);
assign n205 = /* CARRY 12 24  4 */ (1'b0 & n104) | ((1'b0 | n104) & n204);
assign n223 = /* CARRY 13 20  2 */ (1'b0 & n153) | ((1'b0 | n153) & n222);
assign n309 = /* CARRY 13 20  0 */ (n220 & 1'b0) | ((n220 | 1'b0) & n552);
assign n286 = /* CARRY 14 26  3 */ (n101 & 1'b0) | ((n101 | 1'b0) & n302);
assign n227 = /* CARRY 13 20  6 */ (1'b0 & n152) | ((1'b0 | n152) & n226);
assign n281 = /* CARRY 14 23  5 */ (1'b0 & n37) | ((1'b0 | n37) & n280);
assign n310 = /* CARRY 14 26  1 */ (n74 & 1'b0) | ((n74 | 1'b0) & n303);
assign n225 = /* CARRY 13 20  4 */ (1'b0 & n155) | ((1'b0 | n155) & n224);
assign n283 = /* CARRY 14 23  7 */ (1'b0 & n55) | ((1'b0 | n55) & n282);
assign n277 = /* CARRY 14 23  1 */ (1'b0 & n31) | ((1'b0 | n31) & n304);
assign n279 = /* CARRY 14 23  3 */ (1'b0 & n89) | ((1'b0 | n89) & n278);
assign n176 = /* CARRY 11 26  1 */ (n74 & n38) | ((n74 | n38) & n305);
assign n209 = /* CARRY 12 25  0 */ (1'b0 & n168) | ((1'b0 | n168) & n208);
/* FF 14 21  4 */ assign n231 = n311;
/* FF 15 20  2 */ always @(posedge clk, posedge rst) if (rst) n257 <= 1'b0; else if (1'b1) n257 <= n312;
/* FF  9 25  0 */ assign n93 = n313;
/* FF 17 22  5 */ assign n244 = n314;
/* FF 12 23  4 */ assign n159 = n315;
/* FF 11 26  7 */ assign n132 = n316;
/* FF  7 21  2 */ assign n28 = n317;
/* FF 12 25  2 */ assign n167 = n318;
/* FF 14 21  2 */ assign n229 = n319;
/* FF 15 20  4 */ always @(posedge clk, posedge rst) if (rst) n259 <= 1'b0; else if (1'b1) n259 <= n320;
/* FF 14 24  0 */ assign n240 = n321;
/* FF 13 24  1 */ assign n201 = n322;
/* FF 11 26  5 */ assign n131 = n323;
/* FF 15 25  1 */ always @(posedge clk, posedge rst) if (rst) n133 <= 1'b0; else if (1'b1) n133 <= n324;
/* FF 15 21  7 */ always @(posedge clk, posedge rst) if (rst) n268 <= 1'b0; else if (1'b1) n268 <= n325;
/* FF 15 20  6 */ always @(posedge clk, posedge rst) if (rst) n195 <= 1'b0; else if (1'b1) n195 <= n326;
/* FF 14 21  0 */ assign n143 = n327;
/* FF 14 24  2 */ assign n242 = n328;
/* FF 15 19  7 */ always @(posedge clk, posedge rst) if (rst) n46 <= 1'b0; else if (1'b1) n46 <= n329;
/* FF 10 26  5 */ assign n113 = n330;
/* FF 13 21  7 */ always @(posedge clk, posedge rst) if (rst) n90 <= 1'b0; else if (n68) n90 <= n331;
/* FF 15 21  5 */ always @(posedge clk, posedge rst) if (rst) n266 <= 1'b0; else if (1'b1) n266 <= n332;
/* FF  9 25  6 */ always @(posedge clk) if (1'b1) n95 <= 1'b0 ? 1'b0 : n333;
/* FF 17 22  3 */ assign n123 = n334;
/* FF 14 24  4 */ assign n243 = n335;
/* FF 15 19  1 */ always @(posedge clk, posedge rst) if (rst) n181 <= 1'b0; else if (1'b1) n181 <= n336;
/* FF 15 28  1 */ assign n337 = n338;
/* FF 14 19  0 */ assign n211 = n339;
/* FF 14 22  6 */ always @(posedge clk, posedge rst) if (rst) read_e <= 1'b0; else if (1'b1) read_e <= n340;
/* FF 11 18  6 */ assign n116 = n341;
/* FF 15 21  3 */ assign n264 = n342;
/* FF 15 22  3 */ assign n272 = n343;
/* FF 15 28  3 */ assign n344 = n345;
/* FF 14 19  2 */ assign n213 = n346;
/* FF 10 24  4 */ always @(posedge clk) if (1'b1) n105 <= 1'b0 ? 1'b0 : n347;
/* FF 13 19  2 */ assign n78 = n348;
/* FF 14 22  4 */ always @(posedge clk, posedge rst) if (rst) write_e <= 1'b0; else if (1'b1) write_e <= n349;
/* FF 16 21  5 */ always @(posedge clk, posedge rst) if (rst) n234 <= 1'b0; else if (1'b1) n234 <= n350;
/* FF 12 24  3 */ assign n60 = n351;
/* FF 15 21  1 */ assign n262 = n352;
/* FF 15 22  1 */ assign n66 = n353;
/* FF 11 27  0 */ assign n354 = n355;
/* FF  7 26  7 */ always @(posedge clk) if (1'b1) n71 <= n44 ? 1'b0 : n357;
/* FF 14 19  4 */ assign n215 = n358;
/* FF 10 24  6 */ always @(posedge clk) if (1'b1) n106 <= 1'b0 ? 1'b0 : n359;
/* FF 12 24  1 */ assign n360 = n361;
/* FF 15 27  4 */ assign n287 = n362;
/* FF 16 21  7 */ always @(posedge clk, posedge rst) if (rst) n292 <= 1'b0; else if (1'b1) n292 <= n363;
/* FF 13 19  0 */ assign n115 = n364;
/* FF 14 20  5 */ assign n154 = n365;
/* FF 15 22  7 */ always @(posedge clk, posedge rst) if (rst) n275 <= 1'b0; else if (1'b1) n275 <= n366;
/* FF 12 22  5 */ assign n155 = n367;
/* FF 11 27  2 */ assign n134 = n368;
/* FF 15 28  7 */ assign n289 = n369;
/* FF 14 19  6 */ assign n216 = n370;
/* FF 16 21  1 */ always @(posedge clk, posedge rst) if (rst) n156 <= 1'b0; else if (1'b1) n156 <= n371;
/* FF 12 24  7 */ assign n165 = n372;
/* FF 14 20  7 */ assign n40 = n373;
/* FF  9 26  1 */ assign n98 = n374;
/* FF 15 22  5 */ always @(posedge clk, posedge rst) if (rst) n200 <= 1'b0; else if (1'b1) n200 <= n375;
/* FF 12 19  4 */ assign n142 = n376;
/* FF 13 19  4 */ assign n184 = n377;
/* FF 10 24  2 */ assign n104 = n378;
/* FF 12 24  5 */ assign n163 = n379;
/* FF 14 20  1 */ assign n218 = n380;
/* FF  7 25  1 */ assign n38 = n381;
/* FF 13 25  2 */ always @(posedge clk, posedge rst) if (rst) n29 <= 1'b0; else if (n1) n29 <= n382;
/* FF 11 27  6 */ always @(posedge clk) if (1'b1) n101 <= rst ? 1'b0 : n383;
/* FF 12 19  2 */ assign n140 = n384;
/* FF 11 19  1 */ assign \data_out[4]  = n385;
/* FF 14 20  3 */ assign n219 = n386;
/* FF  9 26  5 */ assign n44 = n387;
/* FF 13 23  7 */ always @(posedge clk, posedge rst) if (rst) n37 <= 1'b0; else if (n1) n37 <= n388;
/* FF 12 19  0 */ assign n139 = n389;
/* FF 13 22  6 */ assign n122 = n390;
/* FF 11 19  3 */ assign \data_out[2]  = n391;
/* FF 12 26  4 */ assign n51 = n392;
/* FF  9 26  7 */ always @(posedge clk) if (1'b1) n74 <= rst ? 1'b0 : n393;
/* FF  6 24  6 */ assign \port_addr[4]  = n394;
/* FF 11 19  5 */ assign n120 = n395;
/* FF 12 26  6 */ assign n175 = n396;
/* FF 17 21  5 */ assign n64 = n397;
/* FF 13 23  3 */ assign n198 = n398;
/* FF 13 20  3 */ assign n187 = n399;
/* FF 11 19  7 */ assign \data_out[1]  = n400;
/* FF 12 26  0 */ assign n172 = n401;
/* FF 14 26  4 */ assign n178 = n402;
/* FF 17 21  7 */ always @(posedge clk, posedge rst) if (rst) n296 <= 1'b1; else if (1'b1) n296 <= n403;
/* FF 14 25  2 */ assign n247 = n404;
/* FF 13 20  1 */ assign n405 = n406;
/* FF 14 23  4 */ assign n236 = n407;
/* FF 12 26  2 */ assign n73 = n408;
/* FF 14 26  2 */ assign n409 = n410;
/* FF  9 24  6 */ assign n80 = n411;
/* FF 11 24  3 */ assign n124 = n412;
/* FF 12 18  5 */ assign \data_out[6]  = n413;
/* FF 13 20  7 */ assign n190 = n414;
/* FF 14 23  6 */ assign n48 = n415;
/* FF 12 20  7 */ assign n151 = n416;
/* FF 14 26  0 */ assign n417 = n418;
/* FF 12 21  6 */ assign n152 = n420;
/* FF 14 25  6 */ assign n248 = n421;
/* FF 13 20  5 */ assign n182 = n422;
/* FF 14 23  0 */ assign n423 = n424;
/* FF 12 20  5 */ assign n149 = n426;
/* FF 11 25  6 */ always @(posedge clk, posedge rst) if (rst) n10 <= 1'b0; else if (n1) n10 <= n427;
/* FF 14 25  4 */ assign n246 = n428;
/* FF 10 25  6 */ always @(posedge clk) if (1'b1) n111 <= 1'b0 ? 1'b0 : n429;
/* FF 16 22  5 */ assign n196 = n430;
/* FF 14 23  2 */ assign n92 = n431;
/* FF 12 20  3 */ assign n147 = n432;
/* FF 11 26  2 */ assign n128 = n433;
/* FF  7 21  7 */ assign n47 = n434;
/* FF 13 24  6 */ always @(posedge clk, posedge rst) if (rst) n55 <= 1'b0; else if (n1) n55 <= n435;
/* FF 10 25  4 */ always @(posedge clk) if (1'b1) n109 <= 1'b0 ? 1'b0 : n436;
/* FF  6 28  4 */ assign \port_addr[3]  = n437;
/* FF 12 25  5 */ always @(posedge clk) if (1'b1) n170 <= 1'b0 ? 1'b0 : n438;
/* FF 12 20  1 */ assign n144 = n439;
/* FF 11 25  2 */ assign n127 = n440;
/* FF 11 26  0 */ assign n441 = n442;
/* FF 13 24  4 */ always @(posedge clk, posedge rst) if (rst) n89 <= 1'b0; else if (n1) n89 <= n444;
/* FF 10 25  2 */ assign n50 = n445;
/* FF 12 25  7 */ always @(posedge clk) if (1'b1) n171 <= 1'b0 ? 1'b0 : n446;
/* FF 16 22  1 */ assign n276 = n447;
/* FF 14 21  7 */ always @(posedge clk, posedge rst) if (rst) n41 <= 1'b0; else if (1'b1) n41 <= n448;
/* FF 15 20  1 */ always @(posedge clk, posedge rst) if (rst) n256 <= 1'b0; else if (1'b1) n256 <= n449;
/* FF 11 25  0 */ assign n125 = n450;
/* FF 17 22  4 */ assign n102 = n451;
/* FF 12 23  7 */ always @(posedge clk, posedge rst) if (rst) n30 <= 1'b0; else if (n1) n30 <= n452;
/* FF 11 26  6 */ assign n33 = n453;
/* FF 10 26  2 */ assign n112 = n454;
/* FF 10 25  0 */ assign n107 = n455;
/* FF 12 25  1 */ assign n88 = n456;
/* FF 15 26  2 */ assign n114 = n457;
/* FF 14 21  5 */ assign n232 = n458;
/* FF 15 20  3 */ always @(posedge clk, posedge rst) if (rst) n258 <= 1'b0; else if (1'b1) n258 <= n459;
/* FF 14 24  1 */ assign n241 = n460;
/* FF 12 23  5 */ assign n160 = n461;
/* FF 13 24  0 */ assign n158 = n462;
/* FF 11 26  4 */ assign n130 = n463;
/* FF  6 26  2 */ assign \port_addr[5]  = n464;
/* FF 13 21  2 */ assign n193 = n465;
/* FF 14 22  3 */ assign n45 = n466;
/* FF 12 25  3 */ assign n168 = n467;
/* FF 15 20  5 */ always @(posedge clk, posedge rst) if (rst) n255 <= 1'b0; else if (1'b1) n255 <= n468;
/* FF 14 21  3 */ assign n230 = n469;
/* FF  9 25  5 */ assign n94 = n470;
/* FF 15 19  4 */ always @(posedge clk, posedge rst) if (rst) n253 <= 1'b0; else if (1'b1) n253 <= n471;
/* FF 10 26  6 */ always @(posedge clk) if (1'b1) n19 <= rst ? 1'b0 : n472;
/* FF 13 21  4 */ always @(posedge clk, posedge rst) if (rst) n157 <= 1'b0; else if (n68) n157 <= n473;
/* FF 15 21  6 */ always @(posedge clk, posedge rst) if (rst) n267 <= 1'b0; else if (1'b1) n267 <= n474;
/* FF 15 20  7 */ always @(posedge clk, posedge rst) if (rst) n260 <= 1'b0; else if (1'b1) n260 <= n475;
/* FF  9 25  7 */ always @(posedge clk) if (1'b1) n96 <= 1'b0 ? 1'b0 : n476;
/* FF 17 22  2 */ assign n161 = n477;
/* FF 14 24  5 */ always @(posedge clk, posedge rst) if (rst) n32 <= 1'b0; else if (n1) n32 <= n478;
/* FF 14 21  1 */ assign n228 = n479;
/* FF 15 28  0 */ assign n480 = n481;
/* FF 15 21  4 */ assign n265 = n483;
/* FF 15 22  2 */ assign n271 = n484;
/* FF 14 24  7 */ always @(posedge clk, posedge rst) if (rst) n56 <= 1'b0; else if (n1) n56 <= n485;
/* FF 15 19  0 */ assign n251 = n486;
/* FF 15 28  2 */ assign n487 = n488;
/* FF 14 19  1 */ assign n212 = n489;
/* FF 13 19  3 */ assign n183 = n490;
/* FF 15 21  2 */ assign n263 = n491;
/* FF 15 22  0 */ assign n270 = n492;
/* FF  7 26  6 */ assign \port_addr[0]  = n493;
/* FF 15 19  2 */ always @(posedge clk, posedge rst) if (rst) n252 <= 1'b0; else if (1'b1) n252 <= n494;
/* FF 11 27  1 */ assign n495 = n496;
/* FF 15 28  4 */ assign n288 = n497;
/* FF 14 19  3 */ assign n214 = n498;
/* FF 13 19  1 */ assign \data_out[7]  = n499;
/* FF 16 21  6 */ always @(posedge clk, posedge rst) if (rst) n68 <= 1'b0; else if (1'b1) n68 <= n500;
/* FF 12 24  2 */ assign n162 = n501;
/* FF 11 18  5 */ assign \data_out[5]  = n502;
/* FF 15 21  0 */ assign n261 = n503;
/* FF 15 22  6 */ always @(posedge clk, posedge rst) if (rst) n274 <= 1'b0; else if (1'b1) n274 <= n504;
/* FF  7 26  4 */ assign n20 = n505;
/* FF 11 27  3 */ assign n135 = n506;
/* FF 14 19  5 */ assign n52 = n507;
/* FF 13 19  7 */ assign n35 = n508;
/* FF 16 21  0 */ always @(posedge clk, posedge rst) if (rst) n291 <= 1'b0; else if (1'b1) n291 <= n509;
/* FF 10 24  1 */ assign n103 = n510;
/* FF 14 20  4 */ assign n220 = n511;
/* FF 12 24  0 */ assign n512 = n513;
/* FF 15 22  4 */ always @(posedge clk, posedge rst) if (rst) n273 <= 1'b0; else if (1'b1) n273 <= n515;
/* FF 11 27  5 */ assign n97 = n516;
/* FF 14 19  7 */ assign n39 = n517;
/* FF 13 19  5 */ assign n185 = n518;
/* FF 16 21  2 */ always @(posedge clk, posedge rst) if (rst) n233 <= 1'b0; else if (1'b1) n233 <= n519;
/* FF 12 24  6 */ assign n164 = n520;
/* FF 14 20  6 */ assign n221 = n521;
/* FF  9 26  2 */ assign n43 = n522;
/* FF  7 25  2 */ always @(posedge clk) if (1'b1) n70 <= 1'b0 ? 1'b0 : n523;
/* FF 13 22  3 */ assign n191 = n524;
/* FF  6 24  3 */ assign \port_addr[7]  = n525;
/* FF 12 19  5 */ assign n138 = n526;
/* FF 12 24  4 */ assign n49 = n527;
/* FF 14 20  0 */ assign n217 = n528;
/* FF  9 26  4 */ assign n99 = n529;
/* FF  7 25  0 */ assign n42 = n530;
/* FF 14 27  2 */ assign n249 = n531;
/* FF 12 19  3 */ assign n141 = n532;
/* FF 13 22  5 */ assign n194 = n533;
/* FF 11 19  0 */ assign n117 = n534;
/* FF 12 26  5 */ assign n174 = n535;
/* FF 14 20  2 */ assign n121 = n536;
/* FF  9 26  6 */ assign n100 = n537;
/* FF 13 23  6 */ assign n199 = n538;
/* FF 12 19  1 */ assign \data_out[0]  = n539;
/* FF 11 19  2 */ assign n118 = n540;
/* FF  7 28  2 */ assign \port_addr[2]  = n541;
/* FF 12 26  7 */ always @(posedge clk) if (1'b1) n34 <= rst ? 1'b0 : n542;
/* FF 14 28  7 */ assign n250 = n543;
/* FF 13 20  2 */ assign n186 = n544;
/* FF 20 22  7 */ assign n79 = n545;
/* FF 11 19  4 */ assign n119 = n546;
/* FF 17 21  4 */ assign n269 = n547;
/* FF  7 27  5 */ assign \port_addr[1]  = n548;
/* FF  6 23  2 */ assign \port_addr[6]  = n549;
/* FF 13 20  0 */ assign n550 = n551;
/* FF 11 19  6 */ assign \data_out[3]  = n553;
/* FF 12 26  3 */ assign n173 = n554;
/* FF 15 23  5 */ assign n69 = n555;
/* FF 12 21  3 */ assign n153 = n556;
/* FF 14 26  3 */ assign n557 = n558;
/* FF 17 21  6 */ always @(posedge clk, posedge rst) if (rst) n290 <= 1'b0; else if (1'b1) n290 <= n559;
/* FF 13 23  0 */ assign n197 = n560;
/* FF 13 20  6 */ assign n189 = n561;
/* FF 14 23  5 */ assign n237 = n562;
/* FF 14 26  1 */ assign n563 = n564;
/* FF 17 21  0 */ assign n1 = n565;
/* FF  9 24  7 */ always @(posedge clk) if (1'b1) n91 <= 1'b0 ? 1'b0 : n566;
/* FF 12 18  4 */ assign n137 = n567;
/* FF 13 20  4 */ assign n188 = n568;
/* FF 14 23  7 */ assign n238 = n569;
/* FF 12 20  6 */ assign n150 = n570;
/* FF 17 21  2 */ assign n295 = n571;
/* FF 11 24  6 */ always @(posedge clk, posedge rst) if (rst) n31 <= 1'b0; else if (n158) n31 <= n572;
/* FF 14 23  1 */ assign n573 = n574;
/* FF 12 20  4 */ assign n148 = n575;
/* FF 16 22  4 */ assign n239 = n576;
/* FF 12 25  4 */ assign n169 = n577;
/* FF 14 23  3 */ assign n235 = n578;
/* FF 12 20  2 */ assign n146 = n579;
/* FF 13 24  7 */ always @(posedge clk, posedge rst) if (rst) n27 <= 1'b0; else if (n1) n27 <= n580;
/* FF 11 26  3 */ assign n129 = n581;
/* FF 12 18  2 */ assign n136 = n582;
/* FF 10 25  5 */ always @(posedge clk) if (1'b1) n110 <= 1'b0 ? 1'b0 : n583;
/* FF 16 22  6 */ always @(posedge clk, posedge rst) if (rst) n293 <= 1'b0; else if (1'b1) n293 <= n584;
/* FF 15 20  0 */ assign n254 = n585;
/* FF 12 20  0 */ assign n145 = n586;
/* FF 11 25  1 */ assign n126 = n587;
/* FF 12 23  6 */ always @(posedge clk, posedge rst) if (rst) n36 <= 1'b0; else if (n1) n36 <= n588;
/* FF 11 26  1 */ assign n589 = n590;
/* FF 13 21  1 */ assign n192 = n591;
/* FF 10 25  3 */ assign n108 = n592;
/* FF 12 25  0 */ assign n166 = n593;

// Warning: unmatched port '\data_in[7] '
// Warning: unmatched port '\data_in[6] '
// Warning: unmatched port '\data_in[0] '
// Warning: unmatched port '\data_in[5] '
// Warning: unmatched port '\data_in[4] '
// Warning: unmatched port '\data_in[3] '
// Warning: unmatched port '\data_in[1] '
// Warning: unmatched port '\data_in[2] '

endmodule

