// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 12 2017 08:25:46

// File Generated:     Dec 6 2018 15:12:25

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "uart" view "INTERFACE"

module uart (
    output_axis_tdata,
    input_axis_tdata,
    txd,
    tx_busy,
    rxd,
    rx_overrun_error,
    rx_frame_error,
    rx_busy,
    rst,
    output_axis_tvalid,
    output_axis_tready,
    input_axis_tvalid,
    input_axis_tready,
    clk);

    output [7:0] output_axis_tdata;
    input [7:0] input_axis_tdata;
    output txd;
    output tx_busy;
    input rxd;
    output rx_overrun_error;
    output rx_frame_error;
    output rx_busy;
    input rst;
    output output_axis_tvalid;
    input output_axis_tready;
    input input_axis_tvalid;
    output input_axis_tready;
    input clk;

    wire N__9136;
    wire N__9135;
    wire N__9134;
    wire N__9125;
    wire N__9124;
    wire N__9123;
    wire N__9116;
    wire N__9115;
    wire N__9114;
    wire N__9107;
    wire N__9106;
    wire N__9105;
    wire N__9098;
    wire N__9097;
    wire N__9096;
    wire N__9089;
    wire N__9088;
    wire N__9087;
    wire N__9080;
    wire N__9079;
    wire N__9078;
    wire N__9071;
    wire N__9070;
    wire N__9069;
    wire N__9062;
    wire N__9061;
    wire N__9060;
    wire N__9053;
    wire N__9052;
    wire N__9051;
    wire N__9044;
    wire N__9043;
    wire N__9042;
    wire N__9035;
    wire N__9034;
    wire N__9033;
    wire N__9026;
    wire N__9025;
    wire N__9024;
    wire N__9017;
    wire N__9016;
    wire N__9015;
    wire N__9008;
    wire N__9007;
    wire N__9006;
    wire N__8999;
    wire N__8998;
    wire N__8997;
    wire N__8990;
    wire N__8989;
    wire N__8988;
    wire N__8981;
    wire N__8980;
    wire N__8979;
    wire N__8972;
    wire N__8971;
    wire N__8970;
    wire N__8963;
    wire N__8962;
    wire N__8961;
    wire N__8954;
    wire N__8953;
    wire N__8952;
    wire N__8945;
    wire N__8944;
    wire N__8943;
    wire N__8936;
    wire N__8935;
    wire N__8934;
    wire N__8927;
    wire N__8926;
    wire N__8925;
    wire N__8918;
    wire N__8917;
    wire N__8916;
    wire N__8909;
    wire N__8908;
    wire N__8907;
    wire N__8900;
    wire N__8899;
    wire N__8898;
    wire N__8891;
    wire N__8890;
    wire N__8889;
    wire N__8872;
    wire N__8871;
    wire N__8868;
    wire N__8867;
    wire N__8862;
    wire N__8859;
    wire N__8858;
    wire N__8855;
    wire N__8852;
    wire N__8849;
    wire N__8848;
    wire N__8847;
    wire N__8842;
    wire N__8839;
    wire N__8836;
    wire N__8835;
    wire N__8832;
    wire N__8827;
    wire N__8824;
    wire N__8821;
    wire N__8818;
    wire N__8813;
    wire N__8810;
    wire N__8803;
    wire N__8800;
    wire N__8799;
    wire N__8796;
    wire N__8793;
    wire N__8790;
    wire N__8787;
    wire N__8782;
    wire N__8779;
    wire N__8776;
    wire N__8775;
    wire N__8772;
    wire N__8771;
    wire N__8770;
    wire N__8767;
    wire N__8764;
    wire N__8761;
    wire N__8758;
    wire N__8757;
    wire N__8754;
    wire N__8753;
    wire N__8748;
    wire N__8745;
    wire N__8742;
    wire N__8741;
    wire N__8738;
    wire N__8735;
    wire N__8730;
    wire N__8727;
    wire N__8724;
    wire N__8721;
    wire N__8718;
    wire N__8713;
    wire N__8710;
    wire N__8701;
    wire N__8698;
    wire N__8697;
    wire N__8694;
    wire N__8691;
    wire N__8688;
    wire N__8685;
    wire N__8680;
    wire N__8677;
    wire N__8674;
    wire N__8673;
    wire N__8670;
    wire N__8669;
    wire N__8668;
    wire N__8667;
    wire N__8664;
    wire N__8663;
    wire N__8660;
    wire N__8657;
    wire N__8654;
    wire N__8651;
    wire N__8648;
    wire N__8645;
    wire N__8642;
    wire N__8639;
    wire N__8636;
    wire N__8633;
    wire N__8630;
    wire N__8627;
    wire N__8626;
    wire N__8619;
    wire N__8612;
    wire N__8609;
    wire N__8604;
    wire N__8601;
    wire N__8596;
    wire N__8595;
    wire N__8592;
    wire N__8589;
    wire N__8586;
    wire N__8583;
    wire N__8578;
    wire N__8575;
    wire N__8572;
    wire N__8571;
    wire N__8570;
    wire N__8567;
    wire N__8566;
    wire N__8565;
    wire N__8564;
    wire N__8561;
    wire N__8558;
    wire N__8555;
    wire N__8552;
    wire N__8549;
    wire N__8546;
    wire N__8543;
    wire N__8538;
    wire N__8535;
    wire N__8532;
    wire N__8529;
    wire N__8528;
    wire N__8525;
    wire N__8518;
    wire N__8515;
    wire N__8512;
    wire N__8509;
    wire N__8506;
    wire N__8503;
    wire N__8500;
    wire N__8491;
    wire N__8488;
    wire N__8487;
    wire N__8484;
    wire N__8481;
    wire N__8478;
    wire N__8475;
    wire N__8470;
    wire N__8467;
    wire N__8464;
    wire N__8463;
    wire N__8462;
    wire N__8459;
    wire N__8458;
    wire N__8455;
    wire N__8454;
    wire N__8453;
    wire N__8450;
    wire N__8447;
    wire N__8444;
    wire N__8441;
    wire N__8438;
    wire N__8435;
    wire N__8434;
    wire N__8429;
    wire N__8426;
    wire N__8423;
    wire N__8420;
    wire N__8417;
    wire N__8414;
    wire N__8411;
    wire N__8404;
    wire N__8399;
    wire N__8396;
    wire N__8393;
    wire N__8390;
    wire N__8383;
    wire N__8382;
    wire N__8381;
    wire N__8380;
    wire N__8379;
    wire N__8378;
    wire N__8377;
    wire N__8376;
    wire N__8375;
    wire N__8374;
    wire N__8371;
    wire N__8370;
    wire N__8367;
    wire N__8366;
    wire N__8363;
    wire N__8360;
    wire N__8359;
    wire N__8356;
    wire N__8355;
    wire N__8352;
    wire N__8351;
    wire N__8348;
    wire N__8347;
    wire N__8344;
    wire N__8343;
    wire N__8342;
    wire N__8339;
    wire N__8336;
    wire N__8335;
    wire N__8334;
    wire N__8333;
    wire N__8332;
    wire N__8331;
    wire N__8330;
    wire N__8329;
    wire N__8328;
    wire N__8315;
    wire N__8298;
    wire N__8291;
    wire N__8288;
    wire N__8279;
    wire N__8270;
    wire N__8269;
    wire N__8268;
    wire N__8267;
    wire N__8266;
    wire N__8265;
    wire N__8264;
    wire N__8263;
    wire N__8262;
    wire N__8261;
    wire N__8260;
    wire N__8259;
    wire N__8258;
    wire N__8257;
    wire N__8256;
    wire N__8255;
    wire N__8248;
    wire N__8247;
    wire N__8246;
    wire N__8245;
    wire N__8244;
    wire N__8243;
    wire N__8242;
    wire N__8241;
    wire N__8238;
    wire N__8233;
    wire N__8224;
    wire N__8215;
    wire N__8208;
    wire N__8199;
    wire N__8196;
    wire N__8189;
    wire N__8180;
    wire N__8175;
    wire N__8170;
    wire N__8169;
    wire N__8158;
    wire N__8153;
    wire N__8150;
    wire N__8147;
    wire N__8144;
    wire N__8141;
    wire N__8134;
    wire N__8131;
    wire N__8130;
    wire N__8127;
    wire N__8124;
    wire N__8121;
    wire N__8118;
    wire N__8113;
    wire N__8110;
    wire N__8107;
    wire N__8106;
    wire N__8103;
    wire N__8100;
    wire N__8097;
    wire N__8094;
    wire N__8091;
    wire N__8088;
    wire N__8083;
    wire N__8080;
    wire N__8079;
    wire N__8076;
    wire N__8073;
    wire N__8070;
    wire N__8067;
    wire N__8062;
    wire N__8059;
    wire N__8056;
    wire N__8055;
    wire N__8052;
    wire N__8049;
    wire N__8046;
    wire N__8043;
    wire N__8040;
    wire N__8037;
    wire N__8032;
    wire N__8029;
    wire N__8028;
    wire N__8025;
    wire N__8022;
    wire N__8019;
    wire N__8016;
    wire N__8013;
    wire N__8010;
    wire N__8005;
    wire N__8002;
    wire N__7999;
    wire N__7998;
    wire N__7995;
    wire N__7992;
    wire N__7989;
    wire N__7986;
    wire N__7983;
    wire N__7980;
    wire N__7975;
    wire N__7972;
    wire N__7971;
    wire N__7970;
    wire N__7969;
    wire N__7966;
    wire N__7963;
    wire N__7960;
    wire N__7959;
    wire N__7958;
    wire N__7955;
    wire N__7952;
    wire N__7949;
    wire N__7946;
    wire N__7943;
    wire N__7940;
    wire N__7939;
    wire N__7936;
    wire N__7925;
    wire N__7922;
    wire N__7917;
    wire N__7914;
    wire N__7909;
    wire N__7906;
    wire N__7905;
    wire N__7902;
    wire N__7899;
    wire N__7894;
    wire N__7891;
    wire N__7888;
    wire N__7885;
    wire N__7884;
    wire N__7883;
    wire N__7882;
    wire N__7881;
    wire N__7878;
    wire N__7877;
    wire N__7874;
    wire N__7871;
    wire N__7868;
    wire N__7865;
    wire N__7862;
    wire N__7859;
    wire N__7856;
    wire N__7853;
    wire N__7850;
    wire N__7847;
    wire N__7846;
    wire N__7843;
    wire N__7838;
    wire N__7831;
    wire N__7828;
    wire N__7821;
    wire N__7818;
    wire N__7813;
    wire N__7810;
    wire N__7809;
    wire N__7806;
    wire N__7803;
    wire N__7800;
    wire N__7797;
    wire N__7792;
    wire N__7789;
    wire N__7788;
    wire N__7787;
    wire N__7786;
    wire N__7785;
    wire N__7784;
    wire N__7781;
    wire N__7778;
    wire N__7775;
    wire N__7772;
    wire N__7769;
    wire N__7766;
    wire N__7763;
    wire N__7760;
    wire N__7757;
    wire N__7754;
    wire N__7751;
    wire N__7750;
    wire N__7747;
    wire N__7744;
    wire N__7735;
    wire N__7732;
    wire N__7729;
    wire N__7724;
    wire N__7721;
    wire N__7714;
    wire N__7711;
    wire N__7708;
    wire N__7707;
    wire N__7704;
    wire N__7701;
    wire N__7696;
    wire N__7693;
    wire N__7690;
    wire N__7687;
    wire N__7684;
    wire N__7681;
    wire N__7678;
    wire N__7675;
    wire N__7672;
    wire N__7669;
    wire N__7666;
    wire N__7663;
    wire N__7660;
    wire N__7659;
    wire N__7658;
    wire N__7657;
    wire N__7656;
    wire N__7655;
    wire N__7654;
    wire N__7653;
    wire N__7652;
    wire N__7651;
    wire N__7650;
    wire N__7649;
    wire N__7646;
    wire N__7645;
    wire N__7642;
    wire N__7639;
    wire N__7622;
    wire N__7619;
    wire N__7616;
    wire N__7613;
    wire N__7608;
    wire N__7607;
    wire N__7606;
    wire N__7605;
    wire N__7602;
    wire N__7595;
    wire N__7592;
    wire N__7585;
    wire N__7580;
    wire N__7575;
    wire N__7570;
    wire N__7567;
    wire N__7564;
    wire N__7563;
    wire N__7560;
    wire N__7557;
    wire N__7552;
    wire N__7549;
    wire N__7546;
    wire N__7543;
    wire N__7540;
    wire N__7537;
    wire N__7534;
    wire N__7531;
    wire N__7528;
    wire N__7527;
    wire N__7526;
    wire N__7525;
    wire N__7524;
    wire N__7523;
    wire N__7522;
    wire N__7521;
    wire N__7520;
    wire N__7519;
    wire N__7518;
    wire N__7515;
    wire N__7498;
    wire N__7493;
    wire N__7490;
    wire N__7487;
    wire N__7486;
    wire N__7485;
    wire N__7484;
    wire N__7483;
    wire N__7482;
    wire N__7481;
    wire N__7478;
    wire N__7475;
    wire N__7472;
    wire N__7469;
    wire N__7466;
    wire N__7463;
    wire N__7456;
    wire N__7441;
    wire N__7438;
    wire N__7437;
    wire N__7436;
    wire N__7433;
    wire N__7432;
    wire N__7431;
    wire N__7430;
    wire N__7425;
    wire N__7422;
    wire N__7419;
    wire N__7414;
    wire N__7405;
    wire N__7402;
    wire N__7399;
    wire N__7396;
    wire N__7393;
    wire N__7390;
    wire N__7387;
    wire N__7384;
    wire N__7383;
    wire N__7382;
    wire N__7381;
    wire N__7380;
    wire N__7379;
    wire N__7378;
    wire N__7377;
    wire N__7376;
    wire N__7375;
    wire N__7374;
    wire N__7373;
    wire N__7372;
    wire N__7371;
    wire N__7370;
    wire N__7369;
    wire N__7368;
    wire N__7367;
    wire N__7366;
    wire N__7365;
    wire N__7364;
    wire N__7363;
    wire N__7362;
    wire N__7361;
    wire N__7360;
    wire N__7359;
    wire N__7358;
    wire N__7357;
    wire N__7356;
    wire N__7355;
    wire N__7354;
    wire N__7353;
    wire N__7352;
    wire N__7285;
    wire N__7282;
    wire N__7279;
    wire N__7276;
    wire N__7273;
    wire N__7270;
    wire N__7267;
    wire N__7266;
    wire N__7265;
    wire N__7264;
    wire N__7263;
    wire N__7262;
    wire N__7259;
    wire N__7256;
    wire N__7255;
    wire N__7254;
    wire N__7253;
    wire N__7252;
    wire N__7249;
    wire N__7246;
    wire N__7245;
    wire N__7244;
    wire N__7243;
    wire N__7242;
    wire N__7241;
    wire N__7240;
    wire N__7239;
    wire N__7238;
    wire N__7237;
    wire N__7236;
    wire N__7233;
    wire N__7232;
    wire N__7231;
    wire N__7228;
    wire N__7227;
    wire N__7224;
    wire N__7221;
    wire N__7218;
    wire N__7215;
    wire N__7212;
    wire N__7209;
    wire N__7206;
    wire N__7203;
    wire N__7200;
    wire N__7197;
    wire N__7192;
    wire N__7189;
    wire N__7188;
    wire N__7187;
    wire N__7186;
    wire N__7185;
    wire N__7182;
    wire N__7181;
    wire N__7178;
    wire N__7177;
    wire N__7176;
    wire N__7175;
    wire N__7172;
    wire N__7169;
    wire N__7164;
    wire N__7163;
    wire N__7162;
    wire N__7161;
    wire N__7158;
    wire N__7155;
    wire N__7152;
    wire N__7149;
    wire N__7140;
    wire N__7137;
    wire N__7134;
    wire N__7133;
    wire N__7132;
    wire N__7123;
    wire N__7118;
    wire N__7115;
    wire N__7108;
    wire N__7105;
    wire N__7102;
    wire N__7099;
    wire N__7096;
    wire N__7093;
    wire N__7090;
    wire N__7087;
    wire N__7082;
    wire N__7079;
    wire N__7074;
    wire N__7073;
    wire N__7072;
    wire N__7069;
    wire N__7066;
    wire N__7061;
    wire N__7054;
    wire N__7051;
    wire N__7048;
    wire N__7043;
    wire N__7040;
    wire N__7037;
    wire N__7032;
    wire N__7023;
    wire N__7016;
    wire N__7013;
    wire N__7008;
    wire N__7005;
    wire N__7002;
    wire N__6999;
    wire N__6992;
    wire N__6981;
    wire N__6974;
    wire N__6961;
    wire N__6960;
    wire N__6957;
    wire N__6954;
    wire N__6951;
    wire N__6948;
    wire N__6945;
    wire N__6942;
    wire N__6937;
    wire N__6934;
    wire N__6931;
    wire N__6930;
    wire N__6927;
    wire N__6924;
    wire N__6921;
    wire N__6918;
    wire N__6915;
    wire N__6912;
    wire N__6907;
    wire N__6904;
    wire N__6901;
    wire N__6898;
    wire N__6897;
    wire N__6894;
    wire N__6891;
    wire N__6888;
    wire N__6885;
    wire N__6880;
    wire N__6877;
    wire N__6874;
    wire N__6873;
    wire N__6870;
    wire N__6867;
    wire N__6862;
    wire N__6859;
    wire N__6856;
    wire N__6853;
    wire N__6850;
    wire N__6849;
    wire N__6846;
    wire N__6843;
    wire N__6838;
    wire N__6837;
    wire N__6836;
    wire N__6835;
    wire N__6834;
    wire N__6833;
    wire N__6832;
    wire N__6827;
    wire N__6824;
    wire N__6821;
    wire N__6816;
    wire N__6813;
    wire N__6812;
    wire N__6811;
    wire N__6810;
    wire N__6809;
    wire N__6808;
    wire N__6807;
    wire N__6806;
    wire N__6805;
    wire N__6804;
    wire N__6799;
    wire N__6794;
    wire N__6787;
    wire N__6778;
    wire N__6777;
    wire N__6776;
    wire N__6775;
    wire N__6774;
    wire N__6767;
    wire N__6764;
    wire N__6761;
    wire N__6756;
    wire N__6747;
    wire N__6736;
    wire N__6733;
    wire N__6730;
    wire N__6727;
    wire N__6726;
    wire N__6725;
    wire N__6724;
    wire N__6723;
    wire N__6722;
    wire N__6721;
    wire N__6714;
    wire N__6713;
    wire N__6712;
    wire N__6711;
    wire N__6710;
    wire N__6709;
    wire N__6708;
    wire N__6707;
    wire N__6700;
    wire N__6699;
    wire N__6698;
    wire N__6697;
    wire N__6696;
    wire N__6693;
    wire N__6692;
    wire N__6691;
    wire N__6690;
    wire N__6689;
    wire N__6686;
    wire N__6677;
    wire N__6670;
    wire N__6669;
    wire N__6668;
    wire N__6667;
    wire N__6664;
    wire N__6655;
    wire N__6652;
    wire N__6643;
    wire N__6638;
    wire N__6635;
    wire N__6632;
    wire N__6629;
    wire N__6626;
    wire N__6607;
    wire N__6604;
    wire N__6603;
    wire N__6598;
    wire N__6597;
    wire N__6596;
    wire N__6595;
    wire N__6594;
    wire N__6593;
    wire N__6592;
    wire N__6589;
    wire N__6586;
    wire N__6577;
    wire N__6576;
    wire N__6575;
    wire N__6574;
    wire N__6573;
    wire N__6572;
    wire N__6571;
    wire N__6570;
    wire N__6569;
    wire N__6568;
    wire N__6567;
    wire N__6566;
    wire N__6563;
    wire N__6560;
    wire N__6555;
    wire N__6554;
    wire N__6551;
    wire N__6544;
    wire N__6539;
    wire N__6536;
    wire N__6533;
    wire N__6524;
    wire N__6519;
    wire N__6516;
    wire N__6499;
    wire N__6498;
    wire N__6495;
    wire N__6492;
    wire N__6489;
    wire N__6486;
    wire N__6481;
    wire N__6478;
    wire N__6477;
    wire N__6476;
    wire N__6475;
    wire N__6472;
    wire N__6469;
    wire N__6466;
    wire N__6465;
    wire N__6464;
    wire N__6461;
    wire N__6454;
    wire N__6451;
    wire N__6448;
    wire N__6445;
    wire N__6442;
    wire N__6439;
    wire N__6436;
    wire N__6431;
    wire N__6424;
    wire N__6421;
    wire N__6418;
    wire N__6415;
    wire N__6412;
    wire N__6409;
    wire N__6406;
    wire N__6403;
    wire N__6400;
    wire N__6397;
    wire N__6394;
    wire N__6391;
    wire N__6388;
    wire N__6385;
    wire N__6382;
    wire N__6379;
    wire N__6376;
    wire N__6373;
    wire N__6370;
    wire N__6367;
    wire N__6364;
    wire N__6361;
    wire N__6358;
    wire N__6355;
    wire N__6352;
    wire N__6349;
    wire N__6346;
    wire N__6343;
    wire N__6340;
    wire N__6337;
    wire N__6334;
    wire N__6331;
    wire N__6328;
    wire N__6325;
    wire N__6322;
    wire N__6321;
    wire N__6320;
    wire N__6315;
    wire N__6314;
    wire N__6313;
    wire N__6312;
    wire N__6311;
    wire N__6308;
    wire N__6305;
    wire N__6304;
    wire N__6303;
    wire N__6302;
    wire N__6301;
    wire N__6300;
    wire N__6299;
    wire N__6298;
    wire N__6297;
    wire N__6296;
    wire N__6295;
    wire N__6294;
    wire N__6293;
    wire N__6292;
    wire N__6289;
    wire N__6288;
    wire N__6287;
    wire N__6282;
    wire N__6279;
    wire N__6276;
    wire N__6273;
    wire N__6262;
    wire N__6245;
    wire N__6242;
    wire N__6237;
    wire N__6220;
    wire N__6217;
    wire N__6214;
    wire N__6211;
    wire N__6208;
    wire N__6207;
    wire N__6204;
    wire N__6201;
    wire N__6196;
    wire N__6193;
    wire N__6190;
    wire N__6187;
    wire N__6184;
    wire N__6181;
    wire N__6178;
    wire N__6175;
    wire N__6172;
    wire N__6169;
    wire N__6166;
    wire N__6163;
    wire N__6160;
    wire N__6157;
    wire N__6154;
    wire N__6151;
    wire N__6148;
    wire N__6145;
    wire N__6142;
    wire N__6139;
    wire N__6136;
    wire N__6133;
    wire N__6130;
    wire N__6127;
    wire N__6124;
    wire N__6121;
    wire N__6118;
    wire N__6115;
    wire N__6112;
    wire N__6109;
    wire N__6106;
    wire N__6103;
    wire N__6100;
    wire N__6097;
    wire N__6094;
    wire N__6091;
    wire N__6088;
    wire N__6085;
    wire N__6082;
    wire N__6079;
    wire N__6076;
    wire N__6073;
    wire N__6070;
    wire N__6067;
    wire N__6064;
    wire N__6063;
    wire N__6060;
    wire N__6057;
    wire N__6052;
    wire N__6049;
    wire N__6046;
    wire N__6043;
    wire N__6040;
    wire N__6037;
    wire N__6034;
    wire N__6031;
    wire N__6028;
    wire N__6027;
    wire N__6024;
    wire N__6021;
    wire N__6016;
    wire N__6013;
    wire N__6010;
    wire N__6007;
    wire N__6004;
    wire N__6001;
    wire N__6000;
    wire N__5997;
    wire N__5994;
    wire N__5991;
    wire N__5988;
    wire N__5985;
    wire N__5982;
    wire N__5977;
    wire N__5974;
    wire N__5971;
    wire N__5968;
    wire N__5965;
    wire N__5962;
    wire N__5959;
    wire N__5956;
    wire N__5955;
    wire N__5952;
    wire N__5949;
    wire N__5944;
    wire N__5941;
    wire N__5938;
    wire N__5935;
    wire N__5932;
    wire N__5929;
    wire N__5928;
    wire N__5925;
    wire N__5922;
    wire N__5919;
    wire N__5916;
    wire N__5913;
    wire N__5910;
    wire N__5905;
    wire N__5902;
    wire N__5899;
    wire N__5896;
    wire N__5893;
    wire N__5890;
    wire N__5887;
    wire N__5884;
    wire N__5881;
    wire N__5878;
    wire N__5875;
    wire N__5872;
    wire N__5869;
    wire N__5866;
    wire N__5863;
    wire N__5860;
    wire N__5857;
    wire N__5854;
    wire N__5851;
    wire N__5850;
    wire N__5847;
    wire N__5844;
    wire N__5841;
    wire N__5836;
    wire N__5833;
    wire N__5830;
    wire N__5827;
    wire N__5824;
    wire N__5823;
    wire N__5820;
    wire N__5817;
    wire N__5814;
    wire N__5809;
    wire N__5806;
    wire N__5803;
    wire N__5800;
    wire N__5797;
    wire N__5794;
    wire N__5791;
    wire N__5790;
    wire N__5787;
    wire N__5784;
    wire N__5781;
    wire N__5778;
    wire N__5773;
    wire N__5770;
    wire N__5767;
    wire N__5764;
    wire N__5761;
    wire N__5758;
    wire N__5755;
    wire N__5754;
    wire N__5751;
    wire N__5748;
    wire N__5743;
    wire N__5740;
    wire N__5737;
    wire N__5734;
    wire N__5731;
    wire N__5728;
    wire N__5725;
    wire N__5724;
    wire N__5721;
    wire N__5718;
    wire N__5715;
    wire N__5712;
    wire N__5707;
    wire N__5704;
    wire N__5701;
    wire N__5698;
    wire N__5695;
    wire N__5692;
    wire N__5691;
    wire N__5688;
    wire N__5685;
    wire N__5680;
    wire N__5677;
    wire N__5674;
    wire N__5671;
    wire N__5668;
    wire N__5665;
    wire N__5662;
    wire N__5659;
    wire N__5658;
    wire N__5655;
    wire N__5652;
    wire N__5647;
    wire N__5644;
    wire N__5641;
    wire N__5638;
    wire N__5635;
    wire N__5632;
    wire N__5629;
    wire N__5626;
    wire N__5625;
    wire N__5622;
    wire N__5619;
    wire N__5614;
    wire N__5611;
    wire N__5610;
    wire N__5607;
    wire N__5604;
    wire N__5599;
    wire N__5596;
    wire N__5593;
    wire N__5590;
    wire N__5587;
    wire N__5586;
    wire N__5583;
    wire N__5580;
    wire N__5577;
    wire N__5572;
    wire N__5569;
    wire N__5566;
    wire N__5563;
    wire N__5560;
    wire N__5557;
    wire N__5554;
    wire N__5553;
    wire N__5552;
    wire N__5549;
    wire N__5544;
    wire N__5539;
    wire N__5536;
    wire N__5533;
    wire N__5530;
    wire N__5527;
    wire N__5526;
    wire N__5523;
    wire N__5520;
    wire N__5519;
    wire N__5516;
    wire N__5511;
    wire N__5506;
    wire N__5503;
    wire N__5500;
    wire N__5497;
    wire N__5494;
    wire N__5493;
    wire N__5490;
    wire N__5487;
    wire N__5484;
    wire N__5483;
    wire N__5480;
    wire N__5477;
    wire N__5474;
    wire N__5467;
    wire N__5464;
    wire N__5461;
    wire N__5458;
    wire N__5455;
    wire N__5454;
    wire N__5453;
    wire N__5450;
    wire N__5447;
    wire N__5444;
    wire N__5441;
    wire N__5438;
    wire N__5431;
    wire N__5428;
    wire N__5425;
    wire N__5422;
    wire N__5419;
    wire N__5418;
    wire N__5415;
    wire N__5412;
    wire N__5409;
    wire N__5408;
    wire N__5405;
    wire N__5402;
    wire N__5399;
    wire N__5396;
    wire N__5393;
    wire N__5390;
    wire N__5387;
    wire N__5380;
    wire N__5377;
    wire N__5374;
    wire N__5371;
    wire N__5368;
    wire N__5365;
    wire N__5364;
    wire N__5363;
    wire N__5362;
    wire N__5361;
    wire N__5360;
    wire N__5359;
    wire N__5356;
    wire N__5355;
    wire N__5348;
    wire N__5341;
    wire N__5338;
    wire N__5335;
    wire N__5326;
    wire N__5325;
    wire N__5324;
    wire N__5323;
    wire N__5322;
    wire N__5321;
    wire N__5320;
    wire N__5317;
    wire N__5304;
    wire N__5301;
    wire N__5296;
    wire N__5295;
    wire N__5294;
    wire N__5293;
    wire N__5292;
    wire N__5291;
    wire N__5286;
    wire N__5283;
    wire N__5282;
    wire N__5279;
    wire N__5276;
    wire N__5273;
    wire N__5272;
    wire N__5271;
    wire N__5270;
    wire N__5269;
    wire N__5266;
    wire N__5263;
    wire N__5260;
    wire N__5257;
    wire N__5254;
    wire N__5251;
    wire N__5242;
    wire N__5233;
    wire N__5230;
    wire N__5225;
    wire N__5218;
    wire N__5215;
    wire N__5212;
    wire N__5209;
    wire N__5206;
    wire N__5203;
    wire N__5200;
    wire N__5197;
    wire N__5194;
    wire N__5193;
    wire N__5190;
    wire N__5187;
    wire N__5186;
    wire N__5183;
    wire N__5178;
    wire N__5173;
    wire N__5170;
    wire N__5167;
    wire N__5164;
    wire N__5163;
    wire N__5162;
    wire N__5159;
    wire N__5156;
    wire N__5153;
    wire N__5150;
    wire N__5147;
    wire N__5144;
    wire N__5137;
    wire N__5134;
    wire N__5131;
    wire N__5128;
    wire N__5125;
    wire N__5122;
    wire N__5119;
    wire N__5118;
    wire N__5115;
    wire N__5112;
    wire N__5111;
    wire N__5108;
    wire N__5105;
    wire N__5102;
    wire N__5095;
    wire N__5092;
    wire N__5089;
    wire N__5086;
    wire N__5083;
    wire N__5080;
    wire N__5077;
    wire N__5074;
    wire N__5071;
    wire N__5068;
    wire N__5065;
    wire N__5062;
    wire N__5059;
    wire N__5056;
    wire N__5053;
    wire N__5050;
    wire N__5047;
    wire N__5044;
    wire N__5041;
    wire N__5038;
    wire N__5035;
    wire N__5032;
    wire N__5029;
    wire N__5026;
    wire N__5023;
    wire N__5020;
    wire N__5017;
    wire N__5014;
    wire N__5013;
    wire N__5010;
    wire N__5007;
    wire N__5002;
    wire N__4999;
    wire N__4996;
    wire N__4993;
    wire N__4992;
    wire N__4989;
    wire N__4986;
    wire N__4983;
    wire N__4978;
    wire N__4975;
    wire N__4972;
    wire N__4969;
    wire N__4966;
    wire N__4963;
    wire N__4962;
    wire N__4959;
    wire N__4956;
    wire N__4951;
    wire N__4948;
    wire N__4945;
    wire N__4942;
    wire N__4941;
    wire N__4940;
    wire N__4939;
    wire N__4938;
    wire N__4937;
    wire N__4936;
    wire N__4935;
    wire N__4934;
    wire N__4933;
    wire N__4932;
    wire N__4929;
    wire N__4928;
    wire N__4925;
    wire N__4924;
    wire N__4921;
    wire N__4920;
    wire N__4917;
    wire N__4916;
    wire N__4913;
    wire N__4910;
    wire N__4909;
    wire N__4906;
    wire N__4905;
    wire N__4902;
    wire N__4901;
    wire N__4898;
    wire N__4891;
    wire N__4874;
    wire N__4859;
    wire N__4852;
    wire N__4849;
    wire N__4848;
    wire N__4845;
    wire N__4842;
    wire N__4837;
    wire N__4834;
    wire N__4831;
    wire N__4828;
    wire N__4825;
    wire N__4822;
    wire N__4819;
    wire N__4816;
    wire N__4813;
    wire N__4810;
    wire N__4807;
    wire N__4804;
    wire N__4801;
    wire N__4798;
    wire N__4795;
    wire N__4792;
    wire N__4791;
    wire N__4788;
    wire N__4785;
    wire N__4782;
    wire N__4779;
    wire N__4774;
    wire N__4771;
    wire N__4768;
    wire N__4765;
    wire N__4762;
    wire N__4759;
    wire N__4758;
    wire N__4755;
    wire N__4752;
    wire N__4749;
    wire N__4746;
    wire N__4743;
    wire N__4738;
    wire N__4735;
    wire N__4732;
    wire N__4729;
    wire N__4726;
    wire N__4723;
    wire N__4720;
    wire N__4717;
    wire N__4716;
    wire N__4713;
    wire N__4710;
    wire N__4707;
    wire N__4702;
    wire N__4699;
    wire N__4696;
    wire N__4693;
    wire N__4690;
    wire N__4689;
    wire N__4686;
    wire N__4683;
    wire N__4678;
    wire N__4675;
    wire N__4672;
    wire N__4669;
    wire N__4668;
    wire N__4665;
    wire N__4662;
    wire N__4657;
    wire N__4654;
    wire N__4651;
    wire N__4648;
    wire N__4645;
    wire N__4642;
    wire N__4641;
    wire N__4638;
    wire N__4635;
    wire N__4630;
    wire N__4627;
    wire N__4624;
    wire N__4621;
    wire N__4618;
    wire N__4617;
    wire N__4614;
    wire N__4611;
    wire N__4606;
    wire N__4603;
    wire N__4600;
    wire N__4597;
    wire N__4596;
    wire N__4595;
    wire N__4594;
    wire N__4591;
    wire N__4586;
    wire N__4583;
    wire N__4576;
    wire N__4575;
    wire N__4572;
    wire N__4569;
    wire N__4566;
    wire N__4563;
    wire N__4558;
    wire N__4555;
    wire N__4552;
    wire N__4549;
    wire N__4546;
    wire N__4543;
    wire N__4540;
    wire N__4537;
    wire N__4534;
    wire N__4531;
    wire N__4528;
    wire N__4525;
    wire N__4522;
    wire N__4521;
    wire N__4518;
    wire N__4515;
    wire N__4510;
    wire N__4507;
    wire N__4504;
    wire N__4501;
    wire N__4498;
    wire N__4495;
    wire N__4492;
    wire N__4489;
    wire N__4488;
    wire N__4485;
    wire N__4482;
    wire N__4477;
    wire N__4474;
    wire N__4471;
    wire N__4468;
    wire N__4465;
    wire N__4462;
    wire N__4461;
    wire N__4458;
    wire N__4455;
    wire N__4450;
    wire N__4447;
    wire N__4444;
    wire N__4441;
    wire N__4438;
    wire N__4435;
    wire N__4434;
    wire N__4431;
    wire N__4428;
    wire N__4423;
    wire N__4420;
    wire N__4417;
    wire N__4414;
    wire N__4411;
    wire N__4408;
    wire N__4405;
    wire N__4402;
    wire N__4399;
    wire N__4396;
    wire N__4395;
    wire N__4392;
    wire N__4389;
    wire N__4384;
    wire N__4381;
    wire N__4378;
    wire N__4375;
    wire N__4372;
    wire N__4369;
    wire N__4368;
    wire N__4365;
    wire N__4362;
    wire N__4357;
    wire N__4354;
    wire N__4351;
    wire N__4348;
    wire N__4347;
    wire N__4344;
    wire N__4341;
    wire N__4336;
    wire N__4333;
    wire N__4330;
    wire N__4327;
    wire N__4324;
    wire N__4321;
    wire N__4318;
    wire N__4315;
    wire N__4312;
    wire N__4309;
    wire N__4306;
    wire N__4303;
    wire N__4300;
    wire N__4297;
    wire N__4294;
    wire N__4291;
    wire N__4288;
    wire N__4285;
    wire N__4282;
    wire N__4279;
    wire N__4276;
    wire N__4273;
    wire N__4272;
    wire N__4271;
    wire N__4270;
    wire N__4265;
    wire N__4264;
    wire N__4263;
    wire N__4262;
    wire N__4261;
    wire N__4258;
    wire N__4257;
    wire N__4254;
    wire N__4253;
    wire N__4250;
    wire N__4247;
    wire N__4242;
    wire N__4239;
    wire N__4236;
    wire N__4229;
    wire N__4226;
    wire N__4213;
    wire N__4212;
    wire N__4211;
    wire N__4210;
    wire N__4207;
    wire N__4206;
    wire N__4201;
    wire N__4198;
    wire N__4195;
    wire N__4192;
    wire N__4189;
    wire N__4180;
    wire N__4177;
    wire N__4174;
    wire N__4173;
    wire N__4170;
    wire N__4167;
    wire N__4162;
    wire N__4161;
    wire N__4160;
    wire N__4159;
    wire N__4156;
    wire N__4149;
    wire N__4144;
    wire N__4141;
    wire N__4138;
    wire N__4135;
    wire N__4134;
    wire N__4131;
    wire N__4128;
    wire N__4127;
    wire N__4126;
    wire N__4125;
    wire N__4120;
    wire N__4117;
    wire N__4114;
    wire N__4111;
    wire N__4104;
    wire N__4099;
    wire N__4098;
    wire N__4095;
    wire N__4092;
    wire N__4091;
    wire N__4086;
    wire N__4083;
    wire N__4080;
    wire N__4075;
    wire N__4074;
    wire N__4071;
    wire N__4068;
    wire N__4065;
    wire N__4062;
    wire N__4057;
    wire N__4054;
    wire N__4051;
    wire N__4048;
    wire N__4045;
    wire N__4042;
    wire N__4039;
    wire N__4036;
    wire N__4033;
    wire N__4030;
    wire N__4029;
    wire N__4028;
    wire N__4027;
    wire N__4024;
    wire N__4019;
    wire N__4016;
    wire N__4013;
    wire N__4006;
    wire N__4003;
    wire N__4000;
    wire N__3999;
    wire N__3998;
    wire N__3997;
    wire N__3994;
    wire N__3989;
    wire N__3986;
    wire N__3979;
    wire N__3976;
    wire N__3973;
    wire N__3972;
    wire N__3969;
    wire N__3966;
    wire N__3961;
    wire N__3960;
    wire N__3957;
    wire N__3954;
    wire N__3949;
    wire N__3946;
    wire N__3943;
    wire N__3942;
    wire N__3939;
    wire N__3936;
    wire N__3931;
    wire N__3930;
    wire N__3927;
    wire N__3926;
    wire N__3925;
    wire N__3924;
    wire N__3923;
    wire N__3920;
    wire N__3917;
    wire N__3912;
    wire N__3909;
    wire N__3906;
    wire N__3895;
    wire N__3894;
    wire N__3893;
    wire N__3892;
    wire N__3891;
    wire N__3888;
    wire N__3885;
    wire N__3880;
    wire N__3877;
    wire N__3868;
    wire N__3867;
    wire N__3864;
    wire N__3861;
    wire N__3858;
    wire N__3855;
    wire N__3854;
    wire N__3851;
    wire N__3848;
    wire N__3845;
    wire N__3838;
    wire N__3835;
    wire N__3832;
    wire N__3829;
    wire N__3826;
    wire N__3823;
    wire N__3822;
    wire N__3821;
    wire N__3820;
    wire N__3819;
    wire N__3818;
    wire N__3817;
    wire N__3816;
    wire N__3815;
    wire N__3814;
    wire N__3813;
    wire N__3812;
    wire N__3811;
    wire N__3810;
    wire N__3809;
    wire N__3808;
    wire N__3807;
    wire N__3806;
    wire N__3805;
    wire N__3804;
    wire N__3803;
    wire N__3800;
    wire N__3799;
    wire N__3796;
    wire N__3779;
    wire N__3766;
    wire N__3761;
    wire N__3750;
    wire N__3739;
    wire N__3738;
    wire N__3735;
    wire N__3734;
    wire N__3733;
    wire N__3730;
    wire N__3727;
    wire N__3724;
    wire N__3721;
    wire N__3712;
    wire N__3709;
    wire N__3706;
    wire N__3703;
    wire N__3700;
    wire N__3697;
    wire N__3696;
    wire N__3695;
    wire N__3694;
    wire N__3691;
    wire N__3690;
    wire N__3689;
    wire N__3686;
    wire N__3683;
    wire N__3682;
    wire N__3675;
    wire N__3666;
    wire N__3661;
    wire N__3660;
    wire N__3659;
    wire N__3658;
    wire N__3657;
    wire N__3656;
    wire N__3649;
    wire N__3642;
    wire N__3637;
    wire N__3634;
    wire N__3631;
    wire N__3628;
    wire N__3625;
    wire N__3622;
    wire N__3619;
    wire N__3616;
    wire N__3613;
    wire N__3610;
    wire N__3607;
    wire N__3604;
    wire N__3601;
    wire N__3600;
    wire N__3599;
    wire N__3596;
    wire N__3593;
    wire N__3590;
    wire N__3583;
    wire N__3582;
    wire N__3579;
    wire N__3576;
    wire N__3573;
    wire N__3568;
    wire N__3565;
    wire N__3562;
    wire N__3559;
    wire N__3556;
    wire N__3555;
    wire N__3552;
    wire N__3551;
    wire N__3550;
    wire N__3549;
    wire N__3548;
    wire N__3545;
    wire N__3542;
    wire N__3539;
    wire N__3536;
    wire N__3533;
    wire N__3528;
    wire N__3517;
    wire N__3514;
    wire N__3511;
    wire N__3508;
    wire N__3507;
    wire N__3506;
    wire N__3505;
    wire N__3504;
    wire N__3503;
    wire N__3502;
    wire N__3499;
    wire N__3494;
    wire N__3485;
    wire N__3478;
    wire N__3475;
    wire N__3472;
    wire N__3469;
    wire N__3466;
    wire N__3463;
    wire N__3460;
    wire N__3457;
    wire N__3454;
    wire N__3451;
    wire N__3448;
    wire N__3445;
    wire N__3442;
    wire N__3439;
    wire N__3436;
    wire N__3435;
    wire N__3432;
    wire N__3429;
    wire N__3424;
    wire N__3421;
    wire N__3418;
    wire N__3415;
    wire N__3412;
    wire N__3409;
    wire N__3406;
    wire N__3405;
    wire N__3402;
    wire N__3399;
    wire N__3394;
    wire N__3393;
    wire N__3390;
    wire N__3387;
    wire N__3382;
    wire N__3379;
    wire N__3376;
    wire N__3373;
    wire N__3370;
    wire N__3367;
    wire N__3364;
    wire N__3361;
    wire N__3358;
    wire N__3355;
    wire N__3352;
    wire N__3351;
    wire N__3348;
    wire N__3345;
    wire N__3340;
    wire N__3337;
    wire N__3334;
    wire N__3331;
    wire N__3328;
    wire N__3325;
    wire N__3322;
    wire N__3319;
    wire N__3316;
    wire N__3313;
    wire N__3310;
    wire N__3307;
    wire N__3304;
    wire N__3301;
    wire VCCG0;
    wire GNDG0;
    wire tx_busy_c;
    wire \uart_tx_inst.n721 ;
    wire input_axis_tready_c;
    wire \uart_tx_inst.n701 ;
    wire \uart_tx_inst.n535 ;
    wire rx_busy_c;
    wire n588_cascade_;
    wire n707_cascade_;
    wire \uart_tx_inst.n7_cascade_ ;
    wire n1165;
    wire n4;
    wire \uart_tx_inst.n613 ;
    wire n707;
    wire rx_overrun_error_c;
    wire \uart_rx_inst.n984 ;
    wire n705_cascade_;
    wire n1167_cascade_;
    wire n1698;
    wire \uart_rx_inst.n677_cascade_ ;
    wire \uart_rx_inst.n607_cascade_ ;
    wire \uart_rx_inst.n603_cascade_ ;
    wire n1471;
    wire \uart_tx_inst.n485_cascade_ ;
    wire \uart_tx_inst.n30_adj_196_cascade_ ;
    wire \uart_tx_inst.n34_cascade_ ;
    wire \uart_tx_inst.n189_cascade_ ;
    wire \uart_tx_inst.bit_cnt_0 ;
    wire \uart_tx_inst.n7_adj_195 ;
    wire \uart_tx_inst.bit_cnt_1 ;
    wire \uart_tx_inst.n15_cascade_ ;
    wire bit_cnt_2;
    wire \uart_tx_inst.bit_cnt_3 ;
    wire \uart_tx_inst.n1723_cascade_ ;
    wire \uart_rx_inst.n681 ;
    wire \uart_tx_inst.n13 ;
    wire output_axis_tready_c;
    wire output_axis_tvalid_c;
    wire \uart_rx_inst.n30_cascade_ ;
    wire \uart_rx_inst.n32_cascade_ ;
    wire \uart_rx_inst.n34 ;
    wire output_axis_tvalid_N_175_cascade_;
    wire \uart_rx_inst.n509_cascade_ ;
    wire \uart_rx_inst.n31 ;
    wire \uart_rx_inst.n33 ;
    wire \uart_rx_inst.n1479 ;
    wire \uart_rx_inst.n1045 ;
    wire \uart_rx_inst.output_axis_tvalid_N_174 ;
    wire n1711_cascade_;
    wire n1220_cascade_;
    wire \uart_rx_inst.bit_cnt_3 ;
    wire \uart_rx_inst.output_axis_tvalid_N_172_cascade_ ;
    wire \uart_rx_inst.n232_cascade_ ;
    wire \uart_rx_inst.n1468 ;
    wire \uart_rx_inst.n1502 ;
    wire \uart_rx_inst.n235 ;
    wire \uart_rx_inst.bit_cnt_1 ;
    wire \uart_rx_inst.bit_cnt_2 ;
    wire n705;
    wire n1167;
    wire bit_cnt_0;
    wire \uart_rx_inst.n677 ;
    wire \uart_rx_inst.output_axis_tvalid_N_172 ;
    wire \uart_rx_inst.output_axis_tvalid_N_173 ;
    wire n695_cascade_;
    wire n695;
    wire output_axis_tvalid_N_175;
    wire n680;
    wire data_reg_0;
    wire output_axis_tdata_c_0;
    wire rxd_c;
    wire \uart_tx_inst.n910_cascade_ ;
    wire \uart_tx_inst.n920_cascade_ ;
    wire \uart_tx_inst.n930_cascade_ ;
    wire \uart_tx_inst.n31_adj_199 ;
    wire \uart_tx_inst.n915 ;
    wire \uart_tx_inst.n875_cascade_ ;
    wire \uart_tx_inst.n880_cascade_ ;
    wire \uart_tx_inst.n895_cascade_ ;
    wire \uart_tx_inst.n900_cascade_ ;
    wire \uart_tx_inst.n925 ;
    wire \uart_tx_inst.n935 ;
    wire \uart_rx_inst.n509 ;
    wire \uart_rx_inst.prescale_reg_0 ;
    wire bfn_9_5_0_;
    wire \uart_rx_inst.n1648 ;
    wire \uart_rx_inst.n1141 ;
    wire \uart_rx_inst.prescale_reg_1 ;
    wire \uart_rx_inst.n819 ;
    wire \uart_rx_inst.n1564 ;
    wire \uart_rx_inst.prescale_reg_2 ;
    wire \uart_rx_inst.n814 ;
    wire \uart_rx_inst.n1565 ;
    wire \uart_rx_inst.prescale_reg_3 ;
    wire \uart_rx_inst.n809 ;
    wire \uart_rx_inst.n1566 ;
    wire \uart_rx_inst.prescale_reg_4 ;
    wire \uart_rx_inst.n804 ;
    wire \uart_rx_inst.n1567 ;
    wire \uart_rx_inst.n1756 ;
    wire \uart_rx_inst.prescale_reg_5 ;
    wire \uart_rx_inst.n799 ;
    wire \uart_rx_inst.n1568 ;
    wire \uart_rx_inst.prescale_reg_6 ;
    wire \uart_rx_inst.n794 ;
    wire \uart_rx_inst.n1569 ;
    wire \uart_rx_inst.prescale_reg_7 ;
    wire \uart_rx_inst.n789 ;
    wire \uart_rx_inst.n1570 ;
    wire \uart_rx_inst.n1571 ;
    wire \uart_rx_inst.prescale_reg_8 ;
    wire \uart_rx_inst.n784 ;
    wire bfn_9_6_0_;
    wire \uart_rx_inst.prescale_reg_9 ;
    wire \uart_rx_inst.n779 ;
    wire \uart_rx_inst.n1572 ;
    wire \uart_rx_inst.n1744 ;
    wire \uart_rx_inst.prescale_reg_10 ;
    wire \uart_rx_inst.n774 ;
    wire \uart_rx_inst.n1573 ;
    wire \uart_rx_inst.prescale_reg_11 ;
    wire \uart_rx_inst.n769 ;
    wire \uart_rx_inst.n1574 ;
    wire \uart_rx_inst.prescale_reg_12 ;
    wire \uart_rx_inst.n764 ;
    wire \uart_rx_inst.n1575 ;
    wire \uart_rx_inst.prescale_reg_13 ;
    wire \uart_rx_inst.n759 ;
    wire \uart_rx_inst.n1576 ;
    wire \uart_rx_inst.prescale_reg_14 ;
    wire \uart_rx_inst.n754 ;
    wire \uart_rx_inst.n1577 ;
    wire \uart_rx_inst.prescale_reg_15 ;
    wire \uart_rx_inst.n749 ;
    wire \uart_rx_inst.n1578 ;
    wire \uart_rx_inst.n1579 ;
    wire \uart_rx_inst.prescale_reg_16 ;
    wire \uart_rx_inst.n744 ;
    wire bfn_9_7_0_;
    wire \uart_rx_inst.prescale_reg_17 ;
    wire \uart_rx_inst.n739 ;
    wire \uart_rx_inst.n1580 ;
    wire \uart_rx_inst.n712 ;
    wire \uart_rx_inst.prescale_reg_18 ;
    wire \uart_rx_inst.n1581 ;
    wire \uart_rx_inst.n729 ;
    wire \uart_rx_inst.n1743 ;
    wire \uart_rx_inst.n1740 ;
    wire \uart_rx_inst.n1741 ;
    wire \uart_rx_inst.n1747 ;
    wire \uart_rx_inst.n1745 ;
    wire \uart_rx_inst.n1750 ;
    wire \uart_rx_inst.n1755 ;
    wire \uart_rx_inst.n1754 ;
    wire \uart_rx_inst.n1751 ;
    wire \uart_rx_inst.n1758 ;
    wire \uart_rx_inst.n1742 ;
    wire \uart_rx_inst.n1739 ;
    wire \uart_rx_inst.n1757 ;
    wire n1711;
    wire n1220;
    wire rxd_reg;
    wire rx_frame_error_c;
    wire n697;
    wire data_reg_6;
    wire output_axis_tdata_c_6;
    wire data_reg_2;
    wire output_axis_tdata_c_2;
    wire data_reg_7;
    wire output_axis_tdata_c_7;
    wire data_reg_4;
    wire output_axis_tdata_c_4;
    wire data_reg_5;
    wire output_axis_tdata_c_5;
    wire data_reg_1;
    wire output_axis_tdata_c_1;
    wire data_reg_3;
    wire output_axis_tdata_c_3;
    wire n703;
    wire \uart_tx_inst.n905_cascade_ ;
    wire \uart_tx_inst.n890_cascade_ ;
    wire \uart_tx_inst.n33_adj_198 ;
    wire \uart_tx_inst.n860_cascade_ ;
    wire bfn_11_2_0_;
    wire \uart_tx_inst.prescale_reg_1 ;
    wire \uart_tx_inst.n1546 ;
    wire \uart_tx_inst.prescale_reg_2 ;
    wire \uart_tx_inst.n1547 ;
    wire \uart_tx_inst.n1170 ;
    wire \uart_tx_inst.prescale_reg_3 ;
    wire \uart_tx_inst.n33 ;
    wire \uart_tx_inst.n1548 ;
    wire \uart_tx_inst.n1549 ;
    wire \uart_tx_inst.n1550 ;
    wire \uart_tx_inst.prescale_reg_6 ;
    wire \uart_tx_inst.n30 ;
    wire \uart_tx_inst.n1551 ;
    wire \uart_tx_inst.prescale_reg_7 ;
    wire \uart_tx_inst.n29 ;
    wire \uart_tx_inst.n1552 ;
    wire \uart_tx_inst.n1553 ;
    wire bfn_11_3_0_;
    wire \uart_tx_inst.prescale_reg_9 ;
    wire \uart_tx_inst.n27 ;
    wire \uart_tx_inst.n1554 ;
    wire \uart_tx_inst.prescale_reg_10 ;
    wire \uart_tx_inst.n26 ;
    wire \uart_tx_inst.n1555 ;
    wire \uart_tx_inst.prescale_reg_11 ;
    wire \uart_tx_inst.n25 ;
    wire \uart_tx_inst.n1556 ;
    wire \uart_tx_inst.prescale_reg_12 ;
    wire \uart_tx_inst.n24 ;
    wire \uart_tx_inst.n1557 ;
    wire \uart_tx_inst.prescale_reg_13 ;
    wire \uart_tx_inst.n23 ;
    wire \uart_tx_inst.n1558 ;
    wire \uart_tx_inst.prescale_reg_14 ;
    wire \uart_tx_inst.n22 ;
    wire \uart_tx_inst.n1559 ;
    wire \uart_tx_inst.prescale_reg_15 ;
    wire \uart_tx_inst.n21 ;
    wire \uart_tx_inst.n1560 ;
    wire \uart_tx_inst.n1561 ;
    wire \uart_tx_inst.prescale_reg_16 ;
    wire \uart_tx_inst.n20 ;
    wire bfn_11_4_0_;
    wire \uart_tx_inst.prescale_reg_17 ;
    wire \uart_tx_inst.n19 ;
    wire \uart_tx_inst.n1562 ;
    wire \uart_tx_inst.prescale_reg_18 ;
    wire \uart_tx_inst.n1563 ;
    wire \uart_tx_inst.n18 ;
    wire \uart_rx_inst.n328 ;
    wire bfn_11_5_0_;
    wire \uart_rx_inst.n327 ;
    wire \uart_rx_inst.n1530 ;
    wire \uart_rx_inst.n326 ;
    wire \uart_rx_inst.n1531 ;
    wire \uart_rx_inst.n325 ;
    wire \uart_rx_inst.n1532 ;
    wire \uart_rx_inst.n324 ;
    wire \uart_rx_inst.n1533 ;
    wire \uart_rx_inst.n323 ;
    wire \uart_rx_inst.n1534 ;
    wire \uart_rx_inst.n322 ;
    wire \uart_rx_inst.n1535 ;
    wire \uart_rx_inst.n321 ;
    wire \uart_rx_inst.n1536 ;
    wire \uart_rx_inst.n1537 ;
    wire \uart_rx_inst.n320 ;
    wire bfn_11_6_0_;
    wire \uart_rx_inst.n319 ;
    wire \uart_rx_inst.n1538 ;
    wire \uart_rx_inst.n318 ;
    wire \uart_rx_inst.n1539 ;
    wire \uart_rx_inst.n317 ;
    wire \uart_rx_inst.n1540 ;
    wire \uart_rx_inst.n316 ;
    wire \uart_rx_inst.n1541 ;
    wire \uart_rx_inst.n315 ;
    wire \uart_rx_inst.n1542 ;
    wire \uart_rx_inst.n314 ;
    wire \uart_rx_inst.n1543 ;
    wire \uart_rx_inst.n313 ;
    wire \uart_rx_inst.n1544 ;
    wire \uart_rx_inst.n1545 ;
    wire bfn_11_7_0_;
    wire \uart_rx_inst.n312 ;
    wire \uart_rx_inst.n232 ;
    wire \uart_rx_inst.n1746 ;
    wire \uart_tx_inst.prescale_reg_0 ;
    wire \uart_tx_inst.n32_adj_197 ;
    wire \uart_tx_inst.n32 ;
    wire \uart_tx_inst.n865_cascade_ ;
    wire \uart_tx_inst.prescale_reg_4 ;
    wire \uart_tx_inst.n31 ;
    wire \uart_tx_inst.n870_cascade_ ;
    wire \uart_tx_inst.prescale_reg_5 ;
    wire \uart_tx_inst.n485 ;
    wire \uart_tx_inst.n28 ;
    wire input_axis_tready_N_72;
    wire \uart_tx_inst.n885_cascade_ ;
    wire \uart_tx_inst.n165 ;
    wire \uart_tx_inst.prescale_reg_8 ;
    wire \uart_tx_inst.n873 ;
    wire \uart_tx_inst.data_reg_1 ;
    wire \uart_tx_inst.data_reg_2 ;
    wire \uart_tx_inst.data_reg_3 ;
    wire \uart_tx_inst.data_reg_4 ;
    wire \uart_tx_inst.data_reg_5 ;
    wire \uart_tx_inst.data_reg_6 ;
    wire input_axis_tvalid_c;
    wire \uart_tx_inst.data_reg_8 ;
    wire \uart_tx_inst.data_reg_7 ;
    wire \uart_tx_inst.n189 ;
    wire \uart_tx_inst.data_reg_0 ;
    wire \uart_tx_inst.n7 ;
    wire \uart_tx_inst.n15 ;
    wire txd_c;
    wire clk_c;
    wire \uart_tx_inst.n719 ;
    wire rst_c;
    wire n108;
    wire bfn_12_5_0_;
    wire n107;
    wire \uart_tx_inst.n1582 ;
    wire n106;
    wire \uart_tx_inst.n1583 ;
    wire n105;
    wire \uart_tx_inst.n1584 ;
    wire n104;
    wire \uart_tx_inst.n1585 ;
    wire n103;
    wire \uart_tx_inst.n1586 ;
    wire n102;
    wire \uart_tx_inst.n1587 ;
    wire n101;
    wire \uart_tx_inst.n1588 ;
    wire \uart_tx_inst.n1589 ;
    wire input_axis_tdata_c_0;
    wire n100;
    wire bfn_12_6_0_;
    wire input_axis_tdata_c_1;
    wire n99;
    wire \uart_tx_inst.n1590 ;
    wire input_axis_tdata_c_2;
    wire n98;
    wire \uart_tx_inst.n1591 ;
    wire input_axis_tdata_c_3;
    wire n97;
    wire \uart_tx_inst.n1592 ;
    wire input_axis_tdata_c_4;
    wire n96;
    wire \uart_tx_inst.n1593 ;
    wire input_axis_tdata_c_5;
    wire n95;
    wire \uart_tx_inst.n1594 ;
    wire input_axis_tdata_c_6;
    wire n94;
    wire \uart_tx_inst.n1595 ;
    wire input_axis_tdata_c_7;
    wire CONSTANT_ONE_NET;
    wire \uart_tx_inst.n1596 ;
    wire n93;
    wire _gnd_net_;

    PRE_IO_GBUF clk_pad_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__9134),
            .GLOBALBUFFEROUTPUT(clk_c));
    defparam clk_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam clk_pad_iopad.PULLUP=1'b0;
    IO_PAD clk_pad_iopad (
            .OE(N__9136),
            .DIN(N__9135),
            .DOUT(N__9134),
            .PACKAGEPIN(clk));
    defparam clk_pad_preio.PIN_TYPE=6'b000001;
    defparam clk_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO clk_pad_preio (
            .PADOEN(N__9136),
            .PADOUT(N__9135),
            .PADIN(N__9134),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam input_axis_tdata_pad_0_iopad.IO_STANDARD="SB_LVCMOS";
    defparam input_axis_tdata_pad_0_iopad.PULLUP=1'b0;
    IO_PAD input_axis_tdata_pad_0_iopad (
            .OE(N__9125),
            .DIN(N__9124),
            .DOUT(N__9123),
            .PACKAGEPIN(input_axis_tdata[0]));
    defparam input_axis_tdata_pad_0_preio.PIN_TYPE=6'b000001;
    defparam input_axis_tdata_pad_0_preio.NEG_TRIGGER=1'b0;
    PRE_IO input_axis_tdata_pad_0_preio (
            .PADOEN(N__9125),
            .PADOUT(N__9124),
            .PADIN(N__9123),
            .CLOCKENABLE(),
            .DIN0(input_axis_tdata_c_0),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam input_axis_tdata_pad_1_iopad.IO_STANDARD="SB_LVCMOS";
    defparam input_axis_tdata_pad_1_iopad.PULLUP=1'b0;
    IO_PAD input_axis_tdata_pad_1_iopad (
            .OE(N__9116),
            .DIN(N__9115),
            .DOUT(N__9114),
            .PACKAGEPIN(input_axis_tdata[1]));
    defparam input_axis_tdata_pad_1_preio.PIN_TYPE=6'b000001;
    defparam input_axis_tdata_pad_1_preio.NEG_TRIGGER=1'b0;
    PRE_IO input_axis_tdata_pad_1_preio (
            .PADOEN(N__9116),
            .PADOUT(N__9115),
            .PADIN(N__9114),
            .CLOCKENABLE(),
            .DIN0(input_axis_tdata_c_1),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam input_axis_tdata_pad_2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam input_axis_tdata_pad_2_iopad.PULLUP=1'b0;
    IO_PAD input_axis_tdata_pad_2_iopad (
            .OE(N__9107),
            .DIN(N__9106),
            .DOUT(N__9105),
            .PACKAGEPIN(input_axis_tdata[2]));
    defparam input_axis_tdata_pad_2_preio.PIN_TYPE=6'b000001;
    defparam input_axis_tdata_pad_2_preio.NEG_TRIGGER=1'b0;
    PRE_IO input_axis_tdata_pad_2_preio (
            .PADOEN(N__9107),
            .PADOUT(N__9106),
            .PADIN(N__9105),
            .CLOCKENABLE(),
            .DIN0(input_axis_tdata_c_2),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam input_axis_tdata_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam input_axis_tdata_pad_3_iopad.PULLUP=1'b0;
    IO_PAD input_axis_tdata_pad_3_iopad (
            .OE(N__9098),
            .DIN(N__9097),
            .DOUT(N__9096),
            .PACKAGEPIN(input_axis_tdata[3]));
    defparam input_axis_tdata_pad_3_preio.PIN_TYPE=6'b000001;
    defparam input_axis_tdata_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO input_axis_tdata_pad_3_preio (
            .PADOEN(N__9098),
            .PADOUT(N__9097),
            .PADIN(N__9096),
            .CLOCKENABLE(),
            .DIN0(input_axis_tdata_c_3),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam input_axis_tdata_pad_4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam input_axis_tdata_pad_4_iopad.PULLUP=1'b0;
    IO_PAD input_axis_tdata_pad_4_iopad (
            .OE(N__9089),
            .DIN(N__9088),
            .DOUT(N__9087),
            .PACKAGEPIN(input_axis_tdata[4]));
    defparam input_axis_tdata_pad_4_preio.PIN_TYPE=6'b000001;
    defparam input_axis_tdata_pad_4_preio.NEG_TRIGGER=1'b0;
    PRE_IO input_axis_tdata_pad_4_preio (
            .PADOEN(N__9089),
            .PADOUT(N__9088),
            .PADIN(N__9087),
            .CLOCKENABLE(),
            .DIN0(input_axis_tdata_c_4),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam input_axis_tdata_pad_5_iopad.IO_STANDARD="SB_LVCMOS";
    defparam input_axis_tdata_pad_5_iopad.PULLUP=1'b0;
    IO_PAD input_axis_tdata_pad_5_iopad (
            .OE(N__9080),
            .DIN(N__9079),
            .DOUT(N__9078),
            .PACKAGEPIN(input_axis_tdata[5]));
    defparam input_axis_tdata_pad_5_preio.PIN_TYPE=6'b000001;
    defparam input_axis_tdata_pad_5_preio.NEG_TRIGGER=1'b0;
    PRE_IO input_axis_tdata_pad_5_preio (
            .PADOEN(N__9080),
            .PADOUT(N__9079),
            .PADIN(N__9078),
            .CLOCKENABLE(),
            .DIN0(input_axis_tdata_c_5),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam input_axis_tdata_pad_6_iopad.IO_STANDARD="SB_LVCMOS";
    defparam input_axis_tdata_pad_6_iopad.PULLUP=1'b0;
    IO_PAD input_axis_tdata_pad_6_iopad (
            .OE(N__9071),
            .DIN(N__9070),
            .DOUT(N__9069),
            .PACKAGEPIN(input_axis_tdata[6]));
    defparam input_axis_tdata_pad_6_preio.PIN_TYPE=6'b000001;
    defparam input_axis_tdata_pad_6_preio.NEG_TRIGGER=1'b0;
    PRE_IO input_axis_tdata_pad_6_preio (
            .PADOEN(N__9071),
            .PADOUT(N__9070),
            .PADIN(N__9069),
            .CLOCKENABLE(),
            .DIN0(input_axis_tdata_c_6),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam input_axis_tdata_pad_7_iopad.IO_STANDARD="SB_LVCMOS";
    defparam input_axis_tdata_pad_7_iopad.PULLUP=1'b0;
    IO_PAD input_axis_tdata_pad_7_iopad (
            .OE(N__9062),
            .DIN(N__9061),
            .DOUT(N__9060),
            .PACKAGEPIN(input_axis_tdata[7]));
    defparam input_axis_tdata_pad_7_preio.PIN_TYPE=6'b000001;
    defparam input_axis_tdata_pad_7_preio.NEG_TRIGGER=1'b0;
    PRE_IO input_axis_tdata_pad_7_preio (
            .PADOEN(N__9062),
            .PADOUT(N__9061),
            .PADIN(N__9060),
            .CLOCKENABLE(),
            .DIN0(input_axis_tdata_c_7),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam input_axis_tready_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam input_axis_tready_pad_iopad.PULLUP=1'b0;
    IO_PAD input_axis_tready_pad_iopad (
            .OE(N__9053),
            .DIN(N__9052),
            .DOUT(N__9051),
            .PACKAGEPIN(input_axis_tready));
    defparam input_axis_tready_pad_preio.PIN_TYPE=6'b011001;
    defparam input_axis_tready_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO input_axis_tready_pad_preio (
            .PADOEN(N__9053),
            .PADOUT(N__9052),
            .PADIN(N__9051),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__3358),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam input_axis_tvalid_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam input_axis_tvalid_pad_iopad.PULLUP=1'b0;
    IO_PAD input_axis_tvalid_pad_iopad (
            .OE(N__9044),
            .DIN(N__9043),
            .DOUT(N__9042),
            .PACKAGEPIN(input_axis_tvalid));
    defparam input_axis_tvalid_pad_preio.PIN_TYPE=6'b000001;
    defparam input_axis_tvalid_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO input_axis_tvalid_pad_preio (
            .PADOEN(N__9044),
            .PADOUT(N__9043),
            .PADIN(N__9042),
            .CLOCKENABLE(),
            .DIN0(input_axis_tvalid_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam output_axis_tdata_pad_0_iopad.IO_STANDARD="SB_LVCMOS";
    defparam output_axis_tdata_pad_0_iopad.PULLUP=1'b0;
    IO_PAD output_axis_tdata_pad_0_iopad (
            .OE(N__9035),
            .DIN(N__9034),
            .DOUT(N__9033),
            .PACKAGEPIN(output_axis_tdata[0]));
    defparam output_axis_tdata_pad_0_preio.PIN_TYPE=6'b011001;
    defparam output_axis_tdata_pad_0_preio.NEG_TRIGGER=1'b0;
    PRE_IO output_axis_tdata_pad_0_preio (
            .PADOEN(N__9035),
            .PADOUT(N__9034),
            .PADIN(N__9033),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__4057),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam output_axis_tdata_pad_1_iopad.IO_STANDARD="SB_LVCMOS";
    defparam output_axis_tdata_pad_1_iopad.PULLUP=1'b0;
    IO_PAD output_axis_tdata_pad_1_iopad (
            .OE(N__9026),
            .DIN(N__9025),
            .DOUT(N__9024),
            .PACKAGEPIN(output_axis_tdata[1]));
    defparam output_axis_tdata_pad_1_preio.PIN_TYPE=6'b011001;
    defparam output_axis_tdata_pad_1_preio.NEG_TRIGGER=1'b0;
    PRE_IO output_axis_tdata_pad_1_preio (
            .PADOEN(N__9026),
            .PADOUT(N__9025),
            .PADIN(N__9024),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__5467),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam output_axis_tdata_pad_2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam output_axis_tdata_pad_2_iopad.PULLUP=1'b0;
    IO_PAD output_axis_tdata_pad_2_iopad (
            .OE(N__9017),
            .DIN(N__9016),
            .DOUT(N__9015),
            .PACKAGEPIN(output_axis_tdata[2]));
    defparam output_axis_tdata_pad_2_preio.PIN_TYPE=6'b011001;
    defparam output_axis_tdata_pad_2_preio.NEG_TRIGGER=1'b0;
    PRE_IO output_axis_tdata_pad_2_preio (
            .PADOEN(N__9017),
            .PADOUT(N__9016),
            .PADIN(N__9015),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__5137),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam output_axis_tdata_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam output_axis_tdata_pad_3_iopad.PULLUP=1'b0;
    IO_PAD output_axis_tdata_pad_3_iopad (
            .OE(N__9008),
            .DIN(N__9007),
            .DOUT(N__9006),
            .PACKAGEPIN(output_axis_tdata[3]));
    defparam output_axis_tdata_pad_3_preio.PIN_TYPE=6'b011001;
    defparam output_axis_tdata_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO output_axis_tdata_pad_3_preio (
            .PADOEN(N__9008),
            .PADOUT(N__9007),
            .PADIN(N__9006),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__5431),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam output_axis_tdata_pad_4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam output_axis_tdata_pad_4_iopad.PULLUP=1'b0;
    IO_PAD output_axis_tdata_pad_4_iopad (
            .OE(N__8999),
            .DIN(N__8998),
            .DOUT(N__8997),
            .PACKAGEPIN(output_axis_tdata[4]));
    defparam output_axis_tdata_pad_4_preio.PIN_TYPE=6'b011001;
    defparam output_axis_tdata_pad_4_preio.NEG_TRIGGER=1'b0;
    PRE_IO output_axis_tdata_pad_4_preio (
            .PADOEN(N__8999),
            .PADOUT(N__8998),
            .PADIN(N__8997),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__5539),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam output_axis_tdata_pad_5_iopad.IO_STANDARD="SB_LVCMOS";
    defparam output_axis_tdata_pad_5_iopad.PULLUP=1'b0;
    IO_PAD output_axis_tdata_pad_5_iopad (
            .OE(N__8990),
            .DIN(N__8989),
            .DOUT(N__8988),
            .PACKAGEPIN(output_axis_tdata[5]));
    defparam output_axis_tdata_pad_5_preio.PIN_TYPE=6'b011001;
    defparam output_axis_tdata_pad_5_preio.NEG_TRIGGER=1'b0;
    PRE_IO output_axis_tdata_pad_5_preio (
            .PADOEN(N__8990),
            .PADOUT(N__8989),
            .PADIN(N__8988),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__5506),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam output_axis_tdata_pad_6_iopad.IO_STANDARD="SB_LVCMOS";
    defparam output_axis_tdata_pad_6_iopad.PULLUP=1'b0;
    IO_PAD output_axis_tdata_pad_6_iopad (
            .OE(N__8981),
            .DIN(N__8980),
            .DOUT(N__8979),
            .PACKAGEPIN(output_axis_tdata[6]));
    defparam output_axis_tdata_pad_6_preio.PIN_TYPE=6'b011001;
    defparam output_axis_tdata_pad_6_preio.NEG_TRIGGER=1'b0;
    PRE_IO output_axis_tdata_pad_6_preio (
            .PADOEN(N__8981),
            .PADOUT(N__8980),
            .PADIN(N__8979),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__5173),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam output_axis_tdata_pad_7_iopad.IO_STANDARD="SB_LVCMOS";
    defparam output_axis_tdata_pad_7_iopad.PULLUP=1'b0;
    IO_PAD output_axis_tdata_pad_7_iopad (
            .OE(N__8972),
            .DIN(N__8971),
            .DOUT(N__8970),
            .PACKAGEPIN(output_axis_tdata[7]));
    defparam output_axis_tdata_pad_7_preio.PIN_TYPE=6'b011001;
    defparam output_axis_tdata_pad_7_preio.NEG_TRIGGER=1'b0;
    PRE_IO output_axis_tdata_pad_7_preio (
            .PADOEN(N__8972),
            .PADOUT(N__8971),
            .PADIN(N__8970),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__5095),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam output_axis_tready_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam output_axis_tready_pad_iopad.PULLUP=1'b0;
    IO_PAD output_axis_tready_pad_iopad (
            .OE(N__8963),
            .DIN(N__8962),
            .DOUT(N__8961),
            .PACKAGEPIN(output_axis_tready));
    defparam output_axis_tready_pad_preio.PIN_TYPE=6'b000001;
    defparam output_axis_tready_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO output_axis_tready_pad_preio (
            .PADOEN(N__8963),
            .PADOUT(N__8962),
            .PADIN(N__8961),
            .CLOCKENABLE(),
            .DIN0(output_axis_tready_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam output_axis_tvalid_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam output_axis_tvalid_pad_iopad.PULLUP=1'b0;
    IO_PAD output_axis_tvalid_pad_iopad (
            .OE(N__8954),
            .DIN(N__8953),
            .DOUT(N__8952),
            .PACKAGEPIN(output_axis_tvalid));
    defparam output_axis_tvalid_pad_preio.PIN_TYPE=6'b011001;
    defparam output_axis_tvalid_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO output_axis_tvalid_pad_preio (
            .PADOEN(N__8954),
            .PADOUT(N__8953),
            .PADIN(N__8952),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__3607),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam rst_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam rst_pad_iopad.PULLUP=1'b0;
    IO_PAD rst_pad_iopad (
            .OE(N__8945),
            .DIN(N__8944),
            .DOUT(N__8943),
            .PACKAGEPIN(rst));
    defparam rst_pad_preio.PIN_TYPE=6'b000001;
    defparam rst_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO rst_pad_preio (
            .PADOEN(N__8945),
            .PADOUT(N__8944),
            .PADIN(N__8943),
            .CLOCKENABLE(),
            .DIN0(rst_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam rx_busy_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam rx_busy_pad_iopad.PULLUP=1'b0;
    IO_PAD rx_busy_pad_iopad (
            .OE(N__8936),
            .DIN(N__8935),
            .DOUT(N__8934),
            .PACKAGEPIN(rx_busy));
    defparam rx_busy_pad_preio.PIN_TYPE=6'b011001;
    defparam rx_busy_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO rx_busy_pad_preio (
            .PADOEN(N__8936),
            .PADOUT(N__8935),
            .PADIN(N__8934),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__3322),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam rx_frame_error_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam rx_frame_error_pad_iopad.PULLUP=1'b0;
    IO_PAD rx_frame_error_pad_iopad (
            .OE(N__8927),
            .DIN(N__8926),
            .DOUT(N__8925),
            .PACKAGEPIN(rx_frame_error));
    defparam rx_frame_error_pad_preio.PIN_TYPE=6'b011001;
    defparam rx_frame_error_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO rx_frame_error_pad_preio (
            .PADOEN(N__8927),
            .PADOUT(N__8926),
            .PADIN(N__8925),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__5218),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam rx_overrun_error_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam rx_overrun_error_pad_iopad.PULLUP=1'b0;
    IO_PAD rx_overrun_error_pad_iopad (
            .OE(N__8918),
            .DIN(N__8917),
            .DOUT(N__8916),
            .PACKAGEPIN(rx_overrun_error));
    defparam rx_overrun_error_pad_preio.PIN_TYPE=6'b011001;
    defparam rx_overrun_error_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO rx_overrun_error_pad_preio (
            .PADOEN(N__8918),
            .PADOUT(N__8917),
            .PADIN(N__8916),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__3382),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam rxd_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam rxd_pad_iopad.PULLUP=1'b0;
    IO_PAD rxd_pad_iopad (
            .OE(N__8909),
            .DIN(N__8908),
            .DOUT(N__8907),
            .PACKAGEPIN(rxd));
    defparam rxd_pad_preio.PIN_TYPE=6'b000001;
    defparam rxd_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO rxd_pad_preio (
            .PADOEN(N__8909),
            .PADOUT(N__8908),
            .PADIN(N__8907),
            .CLOCKENABLE(),
            .DIN0(rxd_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam tx_busy_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam tx_busy_pad_iopad.PULLUP=1'b0;
    IO_PAD tx_busy_pad_iopad (
            .OE(N__8900),
            .DIN(N__8899),
            .DOUT(N__8898),
            .PACKAGEPIN(tx_busy));
    defparam tx_busy_pad_preio.PIN_TYPE=6'b011001;
    defparam tx_busy_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO tx_busy_pad_preio (
            .PADOEN(N__8900),
            .PADOUT(N__8899),
            .PADIN(N__8898),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__3304),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam txd_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam txd_pad_iopad.PULLUP=1'b0;
    IO_PAD txd_pad_iopad (
            .OE(N__8891),
            .DIN(N__8890),
            .DOUT(N__8889),
            .PACKAGEPIN(txd));
    defparam txd_pad_preio.PIN_TYPE=6'b011001;
    defparam txd_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO txd_pad_preio (
            .PADOEN(N__8891),
            .PADOUT(N__8890),
            .PADIN(N__8889),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7405),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    CascadeMux I__2137 (
            .O(N__8872),
            .I(N__8868));
    InMux I__2136 (
            .O(N__8871),
            .I(N__8862));
    InMux I__2135 (
            .O(N__8868),
            .I(N__8862));
    CascadeMux I__2134 (
            .O(N__8867),
            .I(N__8859));
    LocalMux I__2133 (
            .O(N__8862),
            .I(N__8855));
    InMux I__2132 (
            .O(N__8859),
            .I(N__8852));
    CascadeMux I__2131 (
            .O(N__8858),
            .I(N__8849));
    Span4Mux_h I__2130 (
            .O(N__8855),
            .I(N__8842));
    LocalMux I__2129 (
            .O(N__8852),
            .I(N__8842));
    InMux I__2128 (
            .O(N__8849),
            .I(N__8839));
    CascadeMux I__2127 (
            .O(N__8848),
            .I(N__8836));
    CascadeMux I__2126 (
            .O(N__8847),
            .I(N__8832));
    Span4Mux_s1_h I__2125 (
            .O(N__8842),
            .I(N__8827));
    LocalMux I__2124 (
            .O(N__8839),
            .I(N__8827));
    InMux I__2123 (
            .O(N__8836),
            .I(N__8824));
    CascadeMux I__2122 (
            .O(N__8835),
            .I(N__8821));
    InMux I__2121 (
            .O(N__8832),
            .I(N__8818));
    Span4Mux_v I__2120 (
            .O(N__8827),
            .I(N__8813));
    LocalMux I__2119 (
            .O(N__8824),
            .I(N__8813));
    InMux I__2118 (
            .O(N__8821),
            .I(N__8810));
    LocalMux I__2117 (
            .O(N__8818),
            .I(input_axis_tdata_c_3));
    Odrv4 I__2116 (
            .O(N__8813),
            .I(input_axis_tdata_c_3));
    LocalMux I__2115 (
            .O(N__8810),
            .I(input_axis_tdata_c_3));
    InMux I__2114 (
            .O(N__8803),
            .I(N__8800));
    LocalMux I__2113 (
            .O(N__8800),
            .I(N__8796));
    InMux I__2112 (
            .O(N__8799),
            .I(N__8793));
    Span4Mux_s1_v I__2111 (
            .O(N__8796),
            .I(N__8790));
    LocalMux I__2110 (
            .O(N__8793),
            .I(N__8787));
    Span4Mux_v I__2109 (
            .O(N__8790),
            .I(N__8782));
    Span4Mux_v I__2108 (
            .O(N__8787),
            .I(N__8782));
    Odrv4 I__2107 (
            .O(N__8782),
            .I(n97));
    InMux I__2106 (
            .O(N__8779),
            .I(\uart_tx_inst.n1592 ));
    InMux I__2105 (
            .O(N__8776),
            .I(N__8772));
    InMux I__2104 (
            .O(N__8775),
            .I(N__8767));
    LocalMux I__2103 (
            .O(N__8772),
            .I(N__8764));
    InMux I__2102 (
            .O(N__8771),
            .I(N__8761));
    CascadeMux I__2101 (
            .O(N__8770),
            .I(N__8758));
    LocalMux I__2100 (
            .O(N__8767),
            .I(N__8754));
    Span4Mux_h I__2099 (
            .O(N__8764),
            .I(N__8748));
    LocalMux I__2098 (
            .O(N__8761),
            .I(N__8748));
    InMux I__2097 (
            .O(N__8758),
            .I(N__8745));
    CascadeMux I__2096 (
            .O(N__8757),
            .I(N__8742));
    Span4Mux_s3_v I__2095 (
            .O(N__8754),
            .I(N__8738));
    CascadeMux I__2094 (
            .O(N__8753),
            .I(N__8735));
    Span4Mux_s1_h I__2093 (
            .O(N__8748),
            .I(N__8730));
    LocalMux I__2092 (
            .O(N__8745),
            .I(N__8730));
    InMux I__2091 (
            .O(N__8742),
            .I(N__8727));
    CascadeMux I__2090 (
            .O(N__8741),
            .I(N__8724));
    IoSpan4Mux I__2089 (
            .O(N__8738),
            .I(N__8721));
    InMux I__2088 (
            .O(N__8735),
            .I(N__8718));
    Span4Mux_v I__2087 (
            .O(N__8730),
            .I(N__8713));
    LocalMux I__2086 (
            .O(N__8727),
            .I(N__8713));
    InMux I__2085 (
            .O(N__8724),
            .I(N__8710));
    Odrv4 I__2084 (
            .O(N__8721),
            .I(input_axis_tdata_c_4));
    LocalMux I__2083 (
            .O(N__8718),
            .I(input_axis_tdata_c_4));
    Odrv4 I__2082 (
            .O(N__8713),
            .I(input_axis_tdata_c_4));
    LocalMux I__2081 (
            .O(N__8710),
            .I(input_axis_tdata_c_4));
    InMux I__2080 (
            .O(N__8701),
            .I(N__8698));
    LocalMux I__2079 (
            .O(N__8698),
            .I(N__8694));
    InMux I__2078 (
            .O(N__8697),
            .I(N__8691));
    Span4Mux_s1_v I__2077 (
            .O(N__8694),
            .I(N__8688));
    LocalMux I__2076 (
            .O(N__8691),
            .I(N__8685));
    Span4Mux_v I__2075 (
            .O(N__8688),
            .I(N__8680));
    Span4Mux_v I__2074 (
            .O(N__8685),
            .I(N__8680));
    Odrv4 I__2073 (
            .O(N__8680),
            .I(n96));
    InMux I__2072 (
            .O(N__8677),
            .I(\uart_tx_inst.n1593 ));
    CascadeMux I__2071 (
            .O(N__8674),
            .I(N__8670));
    CascadeMux I__2070 (
            .O(N__8673),
            .I(N__8664));
    InMux I__2069 (
            .O(N__8670),
            .I(N__8660));
    CascadeMux I__2068 (
            .O(N__8669),
            .I(N__8657));
    CascadeMux I__2067 (
            .O(N__8668),
            .I(N__8654));
    InMux I__2066 (
            .O(N__8667),
            .I(N__8651));
    InMux I__2065 (
            .O(N__8664),
            .I(N__8648));
    CascadeMux I__2064 (
            .O(N__8663),
            .I(N__8645));
    LocalMux I__2063 (
            .O(N__8660),
            .I(N__8642));
    InMux I__2062 (
            .O(N__8657),
            .I(N__8639));
    InMux I__2061 (
            .O(N__8654),
            .I(N__8636));
    LocalMux I__2060 (
            .O(N__8651),
            .I(N__8633));
    LocalMux I__2059 (
            .O(N__8648),
            .I(N__8630));
    InMux I__2058 (
            .O(N__8645),
            .I(N__8627));
    Span4Mux_h I__2057 (
            .O(N__8642),
            .I(N__8619));
    LocalMux I__2056 (
            .O(N__8639),
            .I(N__8619));
    LocalMux I__2055 (
            .O(N__8636),
            .I(N__8619));
    Span4Mux_s2_v I__2054 (
            .O(N__8633),
            .I(N__8612));
    Span4Mux_s2_v I__2053 (
            .O(N__8630),
            .I(N__8612));
    LocalMux I__2052 (
            .O(N__8627),
            .I(N__8612));
    CascadeMux I__2051 (
            .O(N__8626),
            .I(N__8609));
    Span4Mux_v I__2050 (
            .O(N__8619),
            .I(N__8604));
    Span4Mux_v I__2049 (
            .O(N__8612),
            .I(N__8604));
    InMux I__2048 (
            .O(N__8609),
            .I(N__8601));
    Odrv4 I__2047 (
            .O(N__8604),
            .I(input_axis_tdata_c_5));
    LocalMux I__2046 (
            .O(N__8601),
            .I(input_axis_tdata_c_5));
    InMux I__2045 (
            .O(N__8596),
            .I(N__8592));
    InMux I__2044 (
            .O(N__8595),
            .I(N__8589));
    LocalMux I__2043 (
            .O(N__8592),
            .I(N__8586));
    LocalMux I__2042 (
            .O(N__8589),
            .I(N__8583));
    Span4Mux_v I__2041 (
            .O(N__8586),
            .I(N__8578));
    Span4Mux_v I__2040 (
            .O(N__8583),
            .I(N__8578));
    Odrv4 I__2039 (
            .O(N__8578),
            .I(n95));
    InMux I__2038 (
            .O(N__8575),
            .I(\uart_tx_inst.n1594 ));
    CascadeMux I__2037 (
            .O(N__8572),
            .I(N__8567));
    InMux I__2036 (
            .O(N__8571),
            .I(N__8561));
    InMux I__2035 (
            .O(N__8570),
            .I(N__8558));
    InMux I__2034 (
            .O(N__8567),
            .I(N__8555));
    CascadeMux I__2033 (
            .O(N__8566),
            .I(N__8552));
    CascadeMux I__2032 (
            .O(N__8565),
            .I(N__8549));
    CascadeMux I__2031 (
            .O(N__8564),
            .I(N__8546));
    LocalMux I__2030 (
            .O(N__8561),
            .I(N__8543));
    LocalMux I__2029 (
            .O(N__8558),
            .I(N__8538));
    LocalMux I__2028 (
            .O(N__8555),
            .I(N__8538));
    InMux I__2027 (
            .O(N__8552),
            .I(N__8535));
    InMux I__2026 (
            .O(N__8549),
            .I(N__8532));
    InMux I__2025 (
            .O(N__8546),
            .I(N__8529));
    Span4Mux_s2_v I__2024 (
            .O(N__8543),
            .I(N__8525));
    Span4Mux_s2_v I__2023 (
            .O(N__8538),
            .I(N__8518));
    LocalMux I__2022 (
            .O(N__8535),
            .I(N__8518));
    LocalMux I__2021 (
            .O(N__8532),
            .I(N__8518));
    LocalMux I__2020 (
            .O(N__8529),
            .I(N__8515));
    CascadeMux I__2019 (
            .O(N__8528),
            .I(N__8512));
    Span4Mux_v I__2018 (
            .O(N__8525),
            .I(N__8509));
    Span4Mux_v I__2017 (
            .O(N__8518),
            .I(N__8506));
    Span4Mux_v I__2016 (
            .O(N__8515),
            .I(N__8503));
    InMux I__2015 (
            .O(N__8512),
            .I(N__8500));
    Odrv4 I__2014 (
            .O(N__8509),
            .I(input_axis_tdata_c_6));
    Odrv4 I__2013 (
            .O(N__8506),
            .I(input_axis_tdata_c_6));
    Odrv4 I__2012 (
            .O(N__8503),
            .I(input_axis_tdata_c_6));
    LocalMux I__2011 (
            .O(N__8500),
            .I(input_axis_tdata_c_6));
    InMux I__2010 (
            .O(N__8491),
            .I(N__8488));
    LocalMux I__2009 (
            .O(N__8488),
            .I(N__8484));
    InMux I__2008 (
            .O(N__8487),
            .I(N__8481));
    Span4Mux_s1_v I__2007 (
            .O(N__8484),
            .I(N__8478));
    LocalMux I__2006 (
            .O(N__8481),
            .I(N__8475));
    Span4Mux_v I__2005 (
            .O(N__8478),
            .I(N__8470));
    Span4Mux_v I__2004 (
            .O(N__8475),
            .I(N__8470));
    Odrv4 I__2003 (
            .O(N__8470),
            .I(n94));
    InMux I__2002 (
            .O(N__8467),
            .I(\uart_tx_inst.n1595 ));
    CascadeMux I__2001 (
            .O(N__8464),
            .I(N__8459));
    CascadeMux I__2000 (
            .O(N__8463),
            .I(N__8455));
    InMux I__1999 (
            .O(N__8462),
            .I(N__8450));
    InMux I__1998 (
            .O(N__8459),
            .I(N__8447));
    CascadeMux I__1997 (
            .O(N__8458),
            .I(N__8444));
    InMux I__1996 (
            .O(N__8455),
            .I(N__8441));
    CascadeMux I__1995 (
            .O(N__8454),
            .I(N__8438));
    CascadeMux I__1994 (
            .O(N__8453),
            .I(N__8435));
    LocalMux I__1993 (
            .O(N__8450),
            .I(N__8429));
    LocalMux I__1992 (
            .O(N__8447),
            .I(N__8429));
    InMux I__1991 (
            .O(N__8444),
            .I(N__8426));
    LocalMux I__1990 (
            .O(N__8441),
            .I(N__8423));
    InMux I__1989 (
            .O(N__8438),
            .I(N__8420));
    InMux I__1988 (
            .O(N__8435),
            .I(N__8417));
    InMux I__1987 (
            .O(N__8434),
            .I(N__8414));
    Span4Mux_s3_v I__1986 (
            .O(N__8429),
            .I(N__8411));
    LocalMux I__1985 (
            .O(N__8426),
            .I(N__8404));
    Sp12to4 I__1984 (
            .O(N__8423),
            .I(N__8404));
    LocalMux I__1983 (
            .O(N__8420),
            .I(N__8404));
    LocalMux I__1982 (
            .O(N__8417),
            .I(N__8399));
    LocalMux I__1981 (
            .O(N__8414),
            .I(N__8399));
    Span4Mux_v I__1980 (
            .O(N__8411),
            .I(N__8396));
    Span12Mux_s7_v I__1979 (
            .O(N__8404),
            .I(N__8393));
    Span4Mux_v I__1978 (
            .O(N__8399),
            .I(N__8390));
    Odrv4 I__1977 (
            .O(N__8396),
            .I(input_axis_tdata_c_7));
    Odrv12 I__1976 (
            .O(N__8393),
            .I(input_axis_tdata_c_7));
    Odrv4 I__1975 (
            .O(N__8390),
            .I(input_axis_tdata_c_7));
    CascadeMux I__1974 (
            .O(N__8383),
            .I(N__8371));
    CascadeMux I__1973 (
            .O(N__8382),
            .I(N__8367));
    CascadeMux I__1972 (
            .O(N__8381),
            .I(N__8363));
    CascadeMux I__1971 (
            .O(N__8380),
            .I(N__8360));
    CascadeMux I__1970 (
            .O(N__8379),
            .I(N__8356));
    CascadeMux I__1969 (
            .O(N__8378),
            .I(N__8352));
    CascadeMux I__1968 (
            .O(N__8377),
            .I(N__8348));
    CascadeMux I__1967 (
            .O(N__8376),
            .I(N__8344));
    CascadeMux I__1966 (
            .O(N__8375),
            .I(N__8339));
    CascadeMux I__1965 (
            .O(N__8374),
            .I(N__8336));
    InMux I__1964 (
            .O(N__8371),
            .I(N__8315));
    InMux I__1963 (
            .O(N__8370),
            .I(N__8315));
    InMux I__1962 (
            .O(N__8367),
            .I(N__8315));
    InMux I__1961 (
            .O(N__8366),
            .I(N__8315));
    InMux I__1960 (
            .O(N__8363),
            .I(N__8315));
    InMux I__1959 (
            .O(N__8360),
            .I(N__8315));
    InMux I__1958 (
            .O(N__8359),
            .I(N__8298));
    InMux I__1957 (
            .O(N__8356),
            .I(N__8298));
    InMux I__1956 (
            .O(N__8355),
            .I(N__8298));
    InMux I__1955 (
            .O(N__8352),
            .I(N__8298));
    InMux I__1954 (
            .O(N__8351),
            .I(N__8298));
    InMux I__1953 (
            .O(N__8348),
            .I(N__8298));
    InMux I__1952 (
            .O(N__8347),
            .I(N__8298));
    InMux I__1951 (
            .O(N__8344),
            .I(N__8298));
    InMux I__1950 (
            .O(N__8343),
            .I(N__8291));
    InMux I__1949 (
            .O(N__8342),
            .I(N__8291));
    InMux I__1948 (
            .O(N__8339),
            .I(N__8291));
    InMux I__1947 (
            .O(N__8336),
            .I(N__8288));
    InMux I__1946 (
            .O(N__8335),
            .I(N__8279));
    InMux I__1945 (
            .O(N__8334),
            .I(N__8279));
    InMux I__1944 (
            .O(N__8333),
            .I(N__8279));
    InMux I__1943 (
            .O(N__8332),
            .I(N__8279));
    InMux I__1942 (
            .O(N__8331),
            .I(N__8270));
    InMux I__1941 (
            .O(N__8330),
            .I(N__8270));
    InMux I__1940 (
            .O(N__8329),
            .I(N__8270));
    InMux I__1939 (
            .O(N__8328),
            .I(N__8270));
    LocalMux I__1938 (
            .O(N__8315),
            .I(N__8248));
    LocalMux I__1937 (
            .O(N__8298),
            .I(N__8248));
    LocalMux I__1936 (
            .O(N__8291),
            .I(N__8248));
    LocalMux I__1935 (
            .O(N__8288),
            .I(N__8238));
    LocalMux I__1934 (
            .O(N__8279),
            .I(N__8233));
    LocalMux I__1933 (
            .O(N__8270),
            .I(N__8233));
    InMux I__1932 (
            .O(N__8269),
            .I(N__8224));
    InMux I__1931 (
            .O(N__8268),
            .I(N__8224));
    InMux I__1930 (
            .O(N__8267),
            .I(N__8224));
    InMux I__1929 (
            .O(N__8266),
            .I(N__8224));
    InMux I__1928 (
            .O(N__8265),
            .I(N__8215));
    InMux I__1927 (
            .O(N__8264),
            .I(N__8215));
    InMux I__1926 (
            .O(N__8263),
            .I(N__8215));
    InMux I__1925 (
            .O(N__8262),
            .I(N__8215));
    InMux I__1924 (
            .O(N__8261),
            .I(N__8208));
    InMux I__1923 (
            .O(N__8260),
            .I(N__8208));
    InMux I__1922 (
            .O(N__8259),
            .I(N__8208));
    InMux I__1921 (
            .O(N__8258),
            .I(N__8199));
    InMux I__1920 (
            .O(N__8257),
            .I(N__8199));
    InMux I__1919 (
            .O(N__8256),
            .I(N__8199));
    InMux I__1918 (
            .O(N__8255),
            .I(N__8199));
    Span4Mux_v I__1917 (
            .O(N__8248),
            .I(N__8196));
    InMux I__1916 (
            .O(N__8247),
            .I(N__8189));
    InMux I__1915 (
            .O(N__8246),
            .I(N__8189));
    InMux I__1914 (
            .O(N__8245),
            .I(N__8189));
    InMux I__1913 (
            .O(N__8244),
            .I(N__8180));
    InMux I__1912 (
            .O(N__8243),
            .I(N__8180));
    InMux I__1911 (
            .O(N__8242),
            .I(N__8180));
    InMux I__1910 (
            .O(N__8241),
            .I(N__8180));
    Span4Mux_s2_h I__1909 (
            .O(N__8238),
            .I(N__8175));
    Span4Mux_s2_h I__1908 (
            .O(N__8233),
            .I(N__8175));
    LocalMux I__1907 (
            .O(N__8224),
            .I(N__8170));
    LocalMux I__1906 (
            .O(N__8215),
            .I(N__8170));
    LocalMux I__1905 (
            .O(N__8208),
            .I(N__8158));
    LocalMux I__1904 (
            .O(N__8199),
            .I(N__8158));
    Sp12to4 I__1903 (
            .O(N__8196),
            .I(N__8158));
    LocalMux I__1902 (
            .O(N__8189),
            .I(N__8158));
    LocalMux I__1901 (
            .O(N__8180),
            .I(N__8158));
    Span4Mux_v I__1900 (
            .O(N__8175),
            .I(N__8153));
    Span4Mux_s2_h I__1899 (
            .O(N__8170),
            .I(N__8153));
    InMux I__1898 (
            .O(N__8169),
            .I(N__8150));
    Span12Mux_s6_h I__1897 (
            .O(N__8158),
            .I(N__8147));
    Span4Mux_h I__1896 (
            .O(N__8153),
            .I(N__8144));
    LocalMux I__1895 (
            .O(N__8150),
            .I(N__8141));
    Odrv12 I__1894 (
            .O(N__8147),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__1893 (
            .O(N__8144),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__1892 (
            .O(N__8141),
            .I(CONSTANT_ONE_NET));
    InMux I__1891 (
            .O(N__8134),
            .I(\uart_tx_inst.n1596 ));
    InMux I__1890 (
            .O(N__8131),
            .I(N__8127));
    InMux I__1889 (
            .O(N__8130),
            .I(N__8124));
    LocalMux I__1888 (
            .O(N__8127),
            .I(N__8121));
    LocalMux I__1887 (
            .O(N__8124),
            .I(N__8118));
    Span4Mux_v I__1886 (
            .O(N__8121),
            .I(N__8113));
    Span4Mux_v I__1885 (
            .O(N__8118),
            .I(N__8113));
    Odrv4 I__1884 (
            .O(N__8113),
            .I(n93));
    InMux I__1883 (
            .O(N__8110),
            .I(\uart_tx_inst.n1583 ));
    InMux I__1882 (
            .O(N__8107),
            .I(N__8103));
    InMux I__1881 (
            .O(N__8106),
            .I(N__8100));
    LocalMux I__1880 (
            .O(N__8103),
            .I(N__8097));
    LocalMux I__1879 (
            .O(N__8100),
            .I(N__8094));
    Span4Mux_h I__1878 (
            .O(N__8097),
            .I(N__8091));
    Span4Mux_h I__1877 (
            .O(N__8094),
            .I(N__8088));
    Odrv4 I__1876 (
            .O(N__8091),
            .I(n105));
    Odrv4 I__1875 (
            .O(N__8088),
            .I(n105));
    InMux I__1874 (
            .O(N__8083),
            .I(\uart_tx_inst.n1584 ));
    InMux I__1873 (
            .O(N__8080),
            .I(N__8076));
    InMux I__1872 (
            .O(N__8079),
            .I(N__8073));
    LocalMux I__1871 (
            .O(N__8076),
            .I(N__8070));
    LocalMux I__1870 (
            .O(N__8073),
            .I(N__8067));
    Span4Mux_v I__1869 (
            .O(N__8070),
            .I(N__8062));
    Span4Mux_v I__1868 (
            .O(N__8067),
            .I(N__8062));
    Odrv4 I__1867 (
            .O(N__8062),
            .I(n104));
    InMux I__1866 (
            .O(N__8059),
            .I(\uart_tx_inst.n1585 ));
    InMux I__1865 (
            .O(N__8056),
            .I(N__8052));
    InMux I__1864 (
            .O(N__8055),
            .I(N__8049));
    LocalMux I__1863 (
            .O(N__8052),
            .I(N__8046));
    LocalMux I__1862 (
            .O(N__8049),
            .I(N__8043));
    Span4Mux_v I__1861 (
            .O(N__8046),
            .I(N__8040));
    Span4Mux_s3_v I__1860 (
            .O(N__8043),
            .I(N__8037));
    Odrv4 I__1859 (
            .O(N__8040),
            .I(n103));
    Odrv4 I__1858 (
            .O(N__8037),
            .I(n103));
    InMux I__1857 (
            .O(N__8032),
            .I(\uart_tx_inst.n1586 ));
    InMux I__1856 (
            .O(N__8029),
            .I(N__8025));
    InMux I__1855 (
            .O(N__8028),
            .I(N__8022));
    LocalMux I__1854 (
            .O(N__8025),
            .I(N__8019));
    LocalMux I__1853 (
            .O(N__8022),
            .I(N__8016));
    Span4Mux_s3_v I__1852 (
            .O(N__8019),
            .I(N__8013));
    Span4Mux_v I__1851 (
            .O(N__8016),
            .I(N__8010));
    Odrv4 I__1850 (
            .O(N__8013),
            .I(n102));
    Odrv4 I__1849 (
            .O(N__8010),
            .I(n102));
    InMux I__1848 (
            .O(N__8005),
            .I(\uart_tx_inst.n1587 ));
    InMux I__1847 (
            .O(N__8002),
            .I(N__7999));
    LocalMux I__1846 (
            .O(N__7999),
            .I(N__7995));
    InMux I__1845 (
            .O(N__7998),
            .I(N__7992));
    Span4Mux_v I__1844 (
            .O(N__7995),
            .I(N__7989));
    LocalMux I__1843 (
            .O(N__7992),
            .I(N__7986));
    Span4Mux_h I__1842 (
            .O(N__7989),
            .I(N__7983));
    Span12Mux_s4_v I__1841 (
            .O(N__7986),
            .I(N__7980));
    Odrv4 I__1840 (
            .O(N__7983),
            .I(n101));
    Odrv12 I__1839 (
            .O(N__7980),
            .I(n101));
    InMux I__1838 (
            .O(N__7975),
            .I(\uart_tx_inst.n1588 ));
    CascadeMux I__1837 (
            .O(N__7972),
            .I(N__7966));
    CascadeMux I__1836 (
            .O(N__7971),
            .I(N__7963));
    InMux I__1835 (
            .O(N__7970),
            .I(N__7960));
    InMux I__1834 (
            .O(N__7969),
            .I(N__7955));
    InMux I__1833 (
            .O(N__7966),
            .I(N__7952));
    InMux I__1832 (
            .O(N__7963),
            .I(N__7949));
    LocalMux I__1831 (
            .O(N__7960),
            .I(N__7946));
    InMux I__1830 (
            .O(N__7959),
            .I(N__7943));
    InMux I__1829 (
            .O(N__7958),
            .I(N__7940));
    LocalMux I__1828 (
            .O(N__7955),
            .I(N__7936));
    LocalMux I__1827 (
            .O(N__7952),
            .I(N__7925));
    LocalMux I__1826 (
            .O(N__7949),
            .I(N__7925));
    Span4Mux_s2_v I__1825 (
            .O(N__7946),
            .I(N__7925));
    LocalMux I__1824 (
            .O(N__7943),
            .I(N__7925));
    LocalMux I__1823 (
            .O(N__7940),
            .I(N__7925));
    CascadeMux I__1822 (
            .O(N__7939),
            .I(N__7922));
    Span4Mux_h I__1821 (
            .O(N__7936),
            .I(N__7917));
    Span4Mux_v I__1820 (
            .O(N__7925),
            .I(N__7917));
    InMux I__1819 (
            .O(N__7922),
            .I(N__7914));
    Odrv4 I__1818 (
            .O(N__7917),
            .I(input_axis_tdata_c_0));
    LocalMux I__1817 (
            .O(N__7914),
            .I(input_axis_tdata_c_0));
    InMux I__1816 (
            .O(N__7909),
            .I(N__7906));
    LocalMux I__1815 (
            .O(N__7906),
            .I(N__7902));
    InMux I__1814 (
            .O(N__7905),
            .I(N__7899));
    Span4Mux_v I__1813 (
            .O(N__7902),
            .I(N__7894));
    LocalMux I__1812 (
            .O(N__7899),
            .I(N__7894));
    Span4Mux_v I__1811 (
            .O(N__7894),
            .I(N__7891));
    Odrv4 I__1810 (
            .O(N__7891),
            .I(n100));
    InMux I__1809 (
            .O(N__7888),
            .I(bfn_12_6_0_));
    CascadeMux I__1808 (
            .O(N__7885),
            .I(N__7878));
    CascadeMux I__1807 (
            .O(N__7884),
            .I(N__7874));
    InMux I__1806 (
            .O(N__7883),
            .I(N__7871));
    CascadeMux I__1805 (
            .O(N__7882),
            .I(N__7868));
    CascadeMux I__1804 (
            .O(N__7881),
            .I(N__7865));
    InMux I__1803 (
            .O(N__7878),
            .I(N__7862));
    InMux I__1802 (
            .O(N__7877),
            .I(N__7859));
    InMux I__1801 (
            .O(N__7874),
            .I(N__7856));
    LocalMux I__1800 (
            .O(N__7871),
            .I(N__7853));
    InMux I__1799 (
            .O(N__7868),
            .I(N__7850));
    InMux I__1798 (
            .O(N__7865),
            .I(N__7847));
    LocalMux I__1797 (
            .O(N__7862),
            .I(N__7843));
    LocalMux I__1796 (
            .O(N__7859),
            .I(N__7838));
    LocalMux I__1795 (
            .O(N__7856),
            .I(N__7838));
    Span4Mux_s3_v I__1794 (
            .O(N__7853),
            .I(N__7831));
    LocalMux I__1793 (
            .O(N__7850),
            .I(N__7831));
    LocalMux I__1792 (
            .O(N__7847),
            .I(N__7831));
    CascadeMux I__1791 (
            .O(N__7846),
            .I(N__7828));
    Span4Mux_v I__1790 (
            .O(N__7843),
            .I(N__7821));
    Span4Mux_s3_v I__1789 (
            .O(N__7838),
            .I(N__7821));
    Span4Mux_v I__1788 (
            .O(N__7831),
            .I(N__7821));
    InMux I__1787 (
            .O(N__7828),
            .I(N__7818));
    Odrv4 I__1786 (
            .O(N__7821),
            .I(input_axis_tdata_c_1));
    LocalMux I__1785 (
            .O(N__7818),
            .I(input_axis_tdata_c_1));
    InMux I__1784 (
            .O(N__7813),
            .I(N__7810));
    LocalMux I__1783 (
            .O(N__7810),
            .I(N__7806));
    InMux I__1782 (
            .O(N__7809),
            .I(N__7803));
    Span4Mux_s2_v I__1781 (
            .O(N__7806),
            .I(N__7800));
    LocalMux I__1780 (
            .O(N__7803),
            .I(N__7797));
    Odrv4 I__1779 (
            .O(N__7800),
            .I(n99));
    Odrv4 I__1778 (
            .O(N__7797),
            .I(n99));
    InMux I__1777 (
            .O(N__7792),
            .I(\uart_tx_inst.n1590 ));
    CascadeMux I__1776 (
            .O(N__7789),
            .I(N__7781));
    InMux I__1775 (
            .O(N__7788),
            .I(N__7778));
    CascadeMux I__1774 (
            .O(N__7787),
            .I(N__7775));
    CascadeMux I__1773 (
            .O(N__7786),
            .I(N__7772));
    CascadeMux I__1772 (
            .O(N__7785),
            .I(N__7769));
    InMux I__1771 (
            .O(N__7784),
            .I(N__7766));
    InMux I__1770 (
            .O(N__7781),
            .I(N__7763));
    LocalMux I__1769 (
            .O(N__7778),
            .I(N__7760));
    InMux I__1768 (
            .O(N__7775),
            .I(N__7757));
    InMux I__1767 (
            .O(N__7772),
            .I(N__7754));
    InMux I__1766 (
            .O(N__7769),
            .I(N__7751));
    LocalMux I__1765 (
            .O(N__7766),
            .I(N__7747));
    LocalMux I__1764 (
            .O(N__7763),
            .I(N__7744));
    Span4Mux_s3_v I__1763 (
            .O(N__7760),
            .I(N__7735));
    LocalMux I__1762 (
            .O(N__7757),
            .I(N__7735));
    LocalMux I__1761 (
            .O(N__7754),
            .I(N__7735));
    LocalMux I__1760 (
            .O(N__7751),
            .I(N__7735));
    CascadeMux I__1759 (
            .O(N__7750),
            .I(N__7732));
    IoSpan4Mux I__1758 (
            .O(N__7747),
            .I(N__7729));
    Span4Mux_s3_v I__1757 (
            .O(N__7744),
            .I(N__7724));
    Span4Mux_v I__1756 (
            .O(N__7735),
            .I(N__7724));
    InMux I__1755 (
            .O(N__7732),
            .I(N__7721));
    Odrv4 I__1754 (
            .O(N__7729),
            .I(input_axis_tdata_c_2));
    Odrv4 I__1753 (
            .O(N__7724),
            .I(input_axis_tdata_c_2));
    LocalMux I__1752 (
            .O(N__7721),
            .I(input_axis_tdata_c_2));
    InMux I__1751 (
            .O(N__7714),
            .I(N__7711));
    LocalMux I__1750 (
            .O(N__7711),
            .I(N__7708));
    Span4Mux_s1_v I__1749 (
            .O(N__7708),
            .I(N__7704));
    InMux I__1748 (
            .O(N__7707),
            .I(N__7701));
    Span4Mux_v I__1747 (
            .O(N__7704),
            .I(N__7696));
    LocalMux I__1746 (
            .O(N__7701),
            .I(N__7696));
    Span4Mux_v I__1745 (
            .O(N__7696),
            .I(N__7693));
    Odrv4 I__1744 (
            .O(N__7693),
            .I(n98));
    InMux I__1743 (
            .O(N__7690),
            .I(\uart_tx_inst.n1591 ));
    InMux I__1742 (
            .O(N__7687),
            .I(N__7684));
    LocalMux I__1741 (
            .O(N__7684),
            .I(\uart_tx_inst.data_reg_3 ));
    InMux I__1740 (
            .O(N__7681),
            .I(N__7678));
    LocalMux I__1739 (
            .O(N__7678),
            .I(\uart_tx_inst.data_reg_4 ));
    CascadeMux I__1738 (
            .O(N__7675),
            .I(N__7672));
    InMux I__1737 (
            .O(N__7672),
            .I(N__7669));
    LocalMux I__1736 (
            .O(N__7669),
            .I(\uart_tx_inst.data_reg_5 ));
    InMux I__1735 (
            .O(N__7666),
            .I(N__7663));
    LocalMux I__1734 (
            .O(N__7663),
            .I(\uart_tx_inst.data_reg_6 ));
    InMux I__1733 (
            .O(N__7660),
            .I(N__7646));
    CascadeMux I__1732 (
            .O(N__7659),
            .I(N__7642));
    CascadeMux I__1731 (
            .O(N__7658),
            .I(N__7639));
    InMux I__1730 (
            .O(N__7657),
            .I(N__7622));
    InMux I__1729 (
            .O(N__7656),
            .I(N__7622));
    InMux I__1728 (
            .O(N__7655),
            .I(N__7622));
    InMux I__1727 (
            .O(N__7654),
            .I(N__7622));
    InMux I__1726 (
            .O(N__7653),
            .I(N__7622));
    InMux I__1725 (
            .O(N__7652),
            .I(N__7622));
    InMux I__1724 (
            .O(N__7651),
            .I(N__7622));
    InMux I__1723 (
            .O(N__7650),
            .I(N__7622));
    InMux I__1722 (
            .O(N__7649),
            .I(N__7619));
    LocalMux I__1721 (
            .O(N__7646),
            .I(N__7616));
    InMux I__1720 (
            .O(N__7645),
            .I(N__7613));
    InMux I__1719 (
            .O(N__7642),
            .I(N__7608));
    InMux I__1718 (
            .O(N__7639),
            .I(N__7608));
    LocalMux I__1717 (
            .O(N__7622),
            .I(N__7602));
    LocalMux I__1716 (
            .O(N__7619),
            .I(N__7595));
    Span4Mux_s1_v I__1715 (
            .O(N__7616),
            .I(N__7595));
    LocalMux I__1714 (
            .O(N__7613),
            .I(N__7595));
    LocalMux I__1713 (
            .O(N__7608),
            .I(N__7592));
    InMux I__1712 (
            .O(N__7607),
            .I(N__7585));
    InMux I__1711 (
            .O(N__7606),
            .I(N__7585));
    InMux I__1710 (
            .O(N__7605),
            .I(N__7585));
    Span4Mux_s3_h I__1709 (
            .O(N__7602),
            .I(N__7580));
    Span4Mux_h I__1708 (
            .O(N__7595),
            .I(N__7580));
    Span4Mux_h I__1707 (
            .O(N__7592),
            .I(N__7575));
    LocalMux I__1706 (
            .O(N__7585),
            .I(N__7575));
    Odrv4 I__1705 (
            .O(N__7580),
            .I(input_axis_tvalid_c));
    Odrv4 I__1704 (
            .O(N__7575),
            .I(input_axis_tvalid_c));
    InMux I__1703 (
            .O(N__7570),
            .I(N__7567));
    LocalMux I__1702 (
            .O(N__7567),
            .I(N__7564));
    Span4Mux_s0_h I__1701 (
            .O(N__7564),
            .I(N__7560));
    InMux I__1700 (
            .O(N__7563),
            .I(N__7557));
    Odrv4 I__1699 (
            .O(N__7560),
            .I(\uart_tx_inst.data_reg_8 ));
    LocalMux I__1698 (
            .O(N__7557),
            .I(\uart_tx_inst.data_reg_8 ));
    InMux I__1697 (
            .O(N__7552),
            .I(N__7549));
    LocalMux I__1696 (
            .O(N__7549),
            .I(\uart_tx_inst.data_reg_7 ));
    CEMux I__1695 (
            .O(N__7546),
            .I(N__7543));
    LocalMux I__1694 (
            .O(N__7543),
            .I(N__7540));
    Span4Mux_s0_h I__1693 (
            .O(N__7540),
            .I(N__7537));
    Odrv4 I__1692 (
            .O(N__7537),
            .I(\uart_tx_inst.n189 ));
    InMux I__1691 (
            .O(N__7534),
            .I(N__7531));
    LocalMux I__1690 (
            .O(N__7531),
            .I(\uart_tx_inst.data_reg_0 ));
    InMux I__1689 (
            .O(N__7528),
            .I(N__7515));
    InMux I__1688 (
            .O(N__7527),
            .I(N__7498));
    InMux I__1687 (
            .O(N__7526),
            .I(N__7498));
    InMux I__1686 (
            .O(N__7525),
            .I(N__7498));
    InMux I__1685 (
            .O(N__7524),
            .I(N__7498));
    InMux I__1684 (
            .O(N__7523),
            .I(N__7498));
    InMux I__1683 (
            .O(N__7522),
            .I(N__7498));
    InMux I__1682 (
            .O(N__7521),
            .I(N__7498));
    InMux I__1681 (
            .O(N__7520),
            .I(N__7498));
    InMux I__1680 (
            .O(N__7519),
            .I(N__7493));
    InMux I__1679 (
            .O(N__7518),
            .I(N__7493));
    LocalMux I__1678 (
            .O(N__7515),
            .I(N__7490));
    LocalMux I__1677 (
            .O(N__7498),
            .I(N__7487));
    LocalMux I__1676 (
            .O(N__7493),
            .I(N__7478));
    Span12Mux_v I__1675 (
            .O(N__7490),
            .I(N__7475));
    Span4Mux_s1_h I__1674 (
            .O(N__7487),
            .I(N__7472));
    InMux I__1673 (
            .O(N__7486),
            .I(N__7469));
    InMux I__1672 (
            .O(N__7485),
            .I(N__7466));
    InMux I__1671 (
            .O(N__7484),
            .I(N__7463));
    InMux I__1670 (
            .O(N__7483),
            .I(N__7456));
    InMux I__1669 (
            .O(N__7482),
            .I(N__7456));
    InMux I__1668 (
            .O(N__7481),
            .I(N__7456));
    Odrv4 I__1667 (
            .O(N__7478),
            .I(\uart_tx_inst.n7 ));
    Odrv12 I__1666 (
            .O(N__7475),
            .I(\uart_tx_inst.n7 ));
    Odrv4 I__1665 (
            .O(N__7472),
            .I(\uart_tx_inst.n7 ));
    LocalMux I__1664 (
            .O(N__7469),
            .I(\uart_tx_inst.n7 ));
    LocalMux I__1663 (
            .O(N__7466),
            .I(\uart_tx_inst.n7 ));
    LocalMux I__1662 (
            .O(N__7463),
            .I(\uart_tx_inst.n7 ));
    LocalMux I__1661 (
            .O(N__7456),
            .I(\uart_tx_inst.n7 ));
    InMux I__1660 (
            .O(N__7441),
            .I(N__7438));
    LocalMux I__1659 (
            .O(N__7438),
            .I(N__7433));
    InMux I__1658 (
            .O(N__7437),
            .I(N__7425));
    InMux I__1657 (
            .O(N__7436),
            .I(N__7425));
    Span4Mux_s3_h I__1656 (
            .O(N__7433),
            .I(N__7422));
    InMux I__1655 (
            .O(N__7432),
            .I(N__7419));
    InMux I__1654 (
            .O(N__7431),
            .I(N__7414));
    InMux I__1653 (
            .O(N__7430),
            .I(N__7414));
    LocalMux I__1652 (
            .O(N__7425),
            .I(\uart_tx_inst.n15 ));
    Odrv4 I__1651 (
            .O(N__7422),
            .I(\uart_tx_inst.n15 ));
    LocalMux I__1650 (
            .O(N__7419),
            .I(\uart_tx_inst.n15 ));
    LocalMux I__1649 (
            .O(N__7414),
            .I(\uart_tx_inst.n15 ));
    IoInMux I__1648 (
            .O(N__7405),
            .I(N__7402));
    LocalMux I__1647 (
            .O(N__7402),
            .I(N__7399));
    IoSpan4Mux I__1646 (
            .O(N__7399),
            .I(N__7396));
    Span4Mux_s3_v I__1645 (
            .O(N__7396),
            .I(N__7393));
    Span4Mux_v I__1644 (
            .O(N__7393),
            .I(N__7390));
    Span4Mux_v I__1643 (
            .O(N__7390),
            .I(N__7387));
    Odrv4 I__1642 (
            .O(N__7387),
            .I(txd_c));
    ClkMux I__1641 (
            .O(N__7384),
            .I(N__7285));
    ClkMux I__1640 (
            .O(N__7383),
            .I(N__7285));
    ClkMux I__1639 (
            .O(N__7382),
            .I(N__7285));
    ClkMux I__1638 (
            .O(N__7381),
            .I(N__7285));
    ClkMux I__1637 (
            .O(N__7380),
            .I(N__7285));
    ClkMux I__1636 (
            .O(N__7379),
            .I(N__7285));
    ClkMux I__1635 (
            .O(N__7378),
            .I(N__7285));
    ClkMux I__1634 (
            .O(N__7377),
            .I(N__7285));
    ClkMux I__1633 (
            .O(N__7376),
            .I(N__7285));
    ClkMux I__1632 (
            .O(N__7375),
            .I(N__7285));
    ClkMux I__1631 (
            .O(N__7374),
            .I(N__7285));
    ClkMux I__1630 (
            .O(N__7373),
            .I(N__7285));
    ClkMux I__1629 (
            .O(N__7372),
            .I(N__7285));
    ClkMux I__1628 (
            .O(N__7371),
            .I(N__7285));
    ClkMux I__1627 (
            .O(N__7370),
            .I(N__7285));
    ClkMux I__1626 (
            .O(N__7369),
            .I(N__7285));
    ClkMux I__1625 (
            .O(N__7368),
            .I(N__7285));
    ClkMux I__1624 (
            .O(N__7367),
            .I(N__7285));
    ClkMux I__1623 (
            .O(N__7366),
            .I(N__7285));
    ClkMux I__1622 (
            .O(N__7365),
            .I(N__7285));
    ClkMux I__1621 (
            .O(N__7364),
            .I(N__7285));
    ClkMux I__1620 (
            .O(N__7363),
            .I(N__7285));
    ClkMux I__1619 (
            .O(N__7362),
            .I(N__7285));
    ClkMux I__1618 (
            .O(N__7361),
            .I(N__7285));
    ClkMux I__1617 (
            .O(N__7360),
            .I(N__7285));
    ClkMux I__1616 (
            .O(N__7359),
            .I(N__7285));
    ClkMux I__1615 (
            .O(N__7358),
            .I(N__7285));
    ClkMux I__1614 (
            .O(N__7357),
            .I(N__7285));
    ClkMux I__1613 (
            .O(N__7356),
            .I(N__7285));
    ClkMux I__1612 (
            .O(N__7355),
            .I(N__7285));
    ClkMux I__1611 (
            .O(N__7354),
            .I(N__7285));
    ClkMux I__1610 (
            .O(N__7353),
            .I(N__7285));
    ClkMux I__1609 (
            .O(N__7352),
            .I(N__7285));
    GlobalMux I__1608 (
            .O(N__7285),
            .I(N__7282));
    gio2CtrlBuf I__1607 (
            .O(N__7282),
            .I(clk_c));
    CEMux I__1606 (
            .O(N__7279),
            .I(N__7276));
    LocalMux I__1605 (
            .O(N__7276),
            .I(N__7273));
    Sp12to4 I__1604 (
            .O(N__7273),
            .I(N__7270));
    Odrv12 I__1603 (
            .O(N__7270),
            .I(\uart_tx_inst.n719 ));
    SRMux I__1602 (
            .O(N__7267),
            .I(N__7259));
    SRMux I__1601 (
            .O(N__7266),
            .I(N__7256));
    SRMux I__1600 (
            .O(N__7265),
            .I(N__7249));
    SRMux I__1599 (
            .O(N__7264),
            .I(N__7246));
    CascadeMux I__1598 (
            .O(N__7263),
            .I(N__7233));
    SRMux I__1597 (
            .O(N__7262),
            .I(N__7228));
    LocalMux I__1596 (
            .O(N__7259),
            .I(N__7224));
    LocalMux I__1595 (
            .O(N__7256),
            .I(N__7221));
    InMux I__1594 (
            .O(N__7255),
            .I(N__7218));
    SRMux I__1593 (
            .O(N__7254),
            .I(N__7215));
    InMux I__1592 (
            .O(N__7253),
            .I(N__7212));
    InMux I__1591 (
            .O(N__7252),
            .I(N__7209));
    LocalMux I__1590 (
            .O(N__7249),
            .I(N__7206));
    LocalMux I__1589 (
            .O(N__7246),
            .I(N__7203));
    InMux I__1588 (
            .O(N__7245),
            .I(N__7200));
    SRMux I__1587 (
            .O(N__7244),
            .I(N__7197));
    InMux I__1586 (
            .O(N__7243),
            .I(N__7192));
    InMux I__1585 (
            .O(N__7242),
            .I(N__7192));
    SRMux I__1584 (
            .O(N__7241),
            .I(N__7189));
    CascadeMux I__1583 (
            .O(N__7240),
            .I(N__7182));
    SRMux I__1582 (
            .O(N__7239),
            .I(N__7178));
    InMux I__1581 (
            .O(N__7238),
            .I(N__7172));
    SRMux I__1580 (
            .O(N__7237),
            .I(N__7169));
    InMux I__1579 (
            .O(N__7236),
            .I(N__7164));
    InMux I__1578 (
            .O(N__7233),
            .I(N__7164));
    SRMux I__1577 (
            .O(N__7232),
            .I(N__7158));
    SRMux I__1576 (
            .O(N__7231),
            .I(N__7155));
    LocalMux I__1575 (
            .O(N__7228),
            .I(N__7152));
    SRMux I__1574 (
            .O(N__7227),
            .I(N__7149));
    Span4Mux_v I__1573 (
            .O(N__7224),
            .I(N__7140));
    Span4Mux_v I__1572 (
            .O(N__7221),
            .I(N__7140));
    LocalMux I__1571 (
            .O(N__7218),
            .I(N__7140));
    LocalMux I__1570 (
            .O(N__7215),
            .I(N__7140));
    LocalMux I__1569 (
            .O(N__7212),
            .I(N__7137));
    LocalMux I__1568 (
            .O(N__7209),
            .I(N__7134));
    Span4Mux_v I__1567 (
            .O(N__7206),
            .I(N__7123));
    Span4Mux_h I__1566 (
            .O(N__7203),
            .I(N__7123));
    LocalMux I__1565 (
            .O(N__7200),
            .I(N__7123));
    LocalMux I__1564 (
            .O(N__7197),
            .I(N__7123));
    LocalMux I__1563 (
            .O(N__7192),
            .I(N__7118));
    LocalMux I__1562 (
            .O(N__7189),
            .I(N__7118));
    SRMux I__1561 (
            .O(N__7188),
            .I(N__7115));
    InMux I__1560 (
            .O(N__7187),
            .I(N__7108));
    InMux I__1559 (
            .O(N__7186),
            .I(N__7108));
    InMux I__1558 (
            .O(N__7185),
            .I(N__7108));
    InMux I__1557 (
            .O(N__7182),
            .I(N__7105));
    SRMux I__1556 (
            .O(N__7181),
            .I(N__7102));
    LocalMux I__1555 (
            .O(N__7178),
            .I(N__7099));
    InMux I__1554 (
            .O(N__7177),
            .I(N__7096));
    InMux I__1553 (
            .O(N__7176),
            .I(N__7093));
    SRMux I__1552 (
            .O(N__7175),
            .I(N__7090));
    LocalMux I__1551 (
            .O(N__7172),
            .I(N__7087));
    LocalMux I__1550 (
            .O(N__7169),
            .I(N__7082));
    LocalMux I__1549 (
            .O(N__7164),
            .I(N__7082));
    SRMux I__1548 (
            .O(N__7163),
            .I(N__7079));
    InMux I__1547 (
            .O(N__7162),
            .I(N__7074));
    InMux I__1546 (
            .O(N__7161),
            .I(N__7074));
    LocalMux I__1545 (
            .O(N__7158),
            .I(N__7069));
    LocalMux I__1544 (
            .O(N__7155),
            .I(N__7066));
    Span4Mux_v I__1543 (
            .O(N__7152),
            .I(N__7061));
    LocalMux I__1542 (
            .O(N__7149),
            .I(N__7061));
    Span4Mux_v I__1541 (
            .O(N__7140),
            .I(N__7054));
    Span4Mux_h I__1540 (
            .O(N__7137),
            .I(N__7054));
    Span4Mux_h I__1539 (
            .O(N__7134),
            .I(N__7054));
    InMux I__1538 (
            .O(N__7133),
            .I(N__7051));
    SRMux I__1537 (
            .O(N__7132),
            .I(N__7048));
    Span4Mux_v I__1536 (
            .O(N__7123),
            .I(N__7043));
    Span4Mux_h I__1535 (
            .O(N__7118),
            .I(N__7043));
    LocalMux I__1534 (
            .O(N__7115),
            .I(N__7040));
    LocalMux I__1533 (
            .O(N__7108),
            .I(N__7037));
    LocalMux I__1532 (
            .O(N__7105),
            .I(N__7032));
    LocalMux I__1531 (
            .O(N__7102),
            .I(N__7032));
    Span4Mux_h I__1530 (
            .O(N__7099),
            .I(N__7023));
    LocalMux I__1529 (
            .O(N__7096),
            .I(N__7023));
    LocalMux I__1528 (
            .O(N__7093),
            .I(N__7023));
    LocalMux I__1527 (
            .O(N__7090),
            .I(N__7023));
    Span4Mux_v I__1526 (
            .O(N__7087),
            .I(N__7016));
    Span4Mux_h I__1525 (
            .O(N__7082),
            .I(N__7016));
    LocalMux I__1524 (
            .O(N__7079),
            .I(N__7016));
    LocalMux I__1523 (
            .O(N__7074),
            .I(N__7013));
    InMux I__1522 (
            .O(N__7073),
            .I(N__7008));
    SRMux I__1521 (
            .O(N__7072),
            .I(N__7008));
    Span12Mux_s8_h I__1520 (
            .O(N__7069),
            .I(N__7005));
    Span12Mux_s8_h I__1519 (
            .O(N__7066),
            .I(N__7002));
    IoSpan4Mux I__1518 (
            .O(N__7061),
            .I(N__6999));
    Span4Mux_v I__1517 (
            .O(N__7054),
            .I(N__6992));
    LocalMux I__1516 (
            .O(N__7051),
            .I(N__6992));
    LocalMux I__1515 (
            .O(N__7048),
            .I(N__6992));
    Span4Mux_v I__1514 (
            .O(N__7043),
            .I(N__6981));
    Span4Mux_h I__1513 (
            .O(N__7040),
            .I(N__6981));
    Span4Mux_h I__1512 (
            .O(N__7037),
            .I(N__6981));
    Span4Mux_s3_h I__1511 (
            .O(N__7032),
            .I(N__6981));
    Span4Mux_v I__1510 (
            .O(N__7023),
            .I(N__6981));
    Span4Mux_v I__1509 (
            .O(N__7016),
            .I(N__6974));
    Span4Mux_h I__1508 (
            .O(N__7013),
            .I(N__6974));
    LocalMux I__1507 (
            .O(N__7008),
            .I(N__6974));
    Odrv12 I__1506 (
            .O(N__7005),
            .I(rst_c));
    Odrv12 I__1505 (
            .O(N__7002),
            .I(rst_c));
    Odrv4 I__1504 (
            .O(N__6999),
            .I(rst_c));
    Odrv4 I__1503 (
            .O(N__6992),
            .I(rst_c));
    Odrv4 I__1502 (
            .O(N__6981),
            .I(rst_c));
    Odrv4 I__1501 (
            .O(N__6974),
            .I(rst_c));
    InMux I__1500 (
            .O(N__6961),
            .I(N__6957));
    InMux I__1499 (
            .O(N__6960),
            .I(N__6954));
    LocalMux I__1498 (
            .O(N__6957),
            .I(N__6951));
    LocalMux I__1497 (
            .O(N__6954),
            .I(N__6948));
    Span4Mux_v I__1496 (
            .O(N__6951),
            .I(N__6945));
    Span4Mux_s2_v I__1495 (
            .O(N__6948),
            .I(N__6942));
    Odrv4 I__1494 (
            .O(N__6945),
            .I(n108));
    Odrv4 I__1493 (
            .O(N__6942),
            .I(n108));
    InMux I__1492 (
            .O(N__6937),
            .I(bfn_12_5_0_));
    InMux I__1491 (
            .O(N__6934),
            .I(N__6931));
    LocalMux I__1490 (
            .O(N__6931),
            .I(N__6927));
    InMux I__1489 (
            .O(N__6930),
            .I(N__6924));
    Span4Mux_v I__1488 (
            .O(N__6927),
            .I(N__6921));
    LocalMux I__1487 (
            .O(N__6924),
            .I(N__6918));
    Span4Mux_h I__1486 (
            .O(N__6921),
            .I(N__6915));
    Span4Mux_s1_v I__1485 (
            .O(N__6918),
            .I(N__6912));
    Odrv4 I__1484 (
            .O(N__6915),
            .I(n107));
    Odrv4 I__1483 (
            .O(N__6912),
            .I(n107));
    InMux I__1482 (
            .O(N__6907),
            .I(\uart_tx_inst.n1582 ));
    InMux I__1481 (
            .O(N__6904),
            .I(N__6901));
    LocalMux I__1480 (
            .O(N__6901),
            .I(N__6898));
    Span4Mux_v I__1479 (
            .O(N__6898),
            .I(N__6894));
    InMux I__1478 (
            .O(N__6897),
            .I(N__6891));
    Span4Mux_h I__1477 (
            .O(N__6894),
            .I(N__6888));
    LocalMux I__1476 (
            .O(N__6891),
            .I(N__6885));
    Odrv4 I__1475 (
            .O(N__6888),
            .I(n106));
    Odrv12 I__1474 (
            .O(N__6885),
            .I(n106));
    CascadeMux I__1473 (
            .O(N__6880),
            .I(\uart_tx_inst.n865_cascade_ ));
    CascadeMux I__1472 (
            .O(N__6877),
            .I(N__6874));
    InMux I__1471 (
            .O(N__6874),
            .I(N__6870));
    InMux I__1470 (
            .O(N__6873),
            .I(N__6867));
    LocalMux I__1469 (
            .O(N__6870),
            .I(\uart_tx_inst.prescale_reg_4 ));
    LocalMux I__1468 (
            .O(N__6867),
            .I(\uart_tx_inst.prescale_reg_4 ));
    CascadeMux I__1467 (
            .O(N__6862),
            .I(N__6859));
    InMux I__1466 (
            .O(N__6859),
            .I(N__6856));
    LocalMux I__1465 (
            .O(N__6856),
            .I(\uart_tx_inst.n31 ));
    CascadeMux I__1464 (
            .O(N__6853),
            .I(\uart_tx_inst.n870_cascade_ ));
    InMux I__1463 (
            .O(N__6850),
            .I(N__6846));
    InMux I__1462 (
            .O(N__6849),
            .I(N__6843));
    LocalMux I__1461 (
            .O(N__6846),
            .I(\uart_tx_inst.prescale_reg_5 ));
    LocalMux I__1460 (
            .O(N__6843),
            .I(\uart_tx_inst.prescale_reg_5 ));
    InMux I__1459 (
            .O(N__6838),
            .I(N__6827));
    InMux I__1458 (
            .O(N__6837),
            .I(N__6827));
    InMux I__1457 (
            .O(N__6836),
            .I(N__6824));
    InMux I__1456 (
            .O(N__6835),
            .I(N__6821));
    InMux I__1455 (
            .O(N__6834),
            .I(N__6816));
    InMux I__1454 (
            .O(N__6833),
            .I(N__6816));
    CascadeMux I__1453 (
            .O(N__6832),
            .I(N__6813));
    LocalMux I__1452 (
            .O(N__6827),
            .I(N__6799));
    LocalMux I__1451 (
            .O(N__6824),
            .I(N__6799));
    LocalMux I__1450 (
            .O(N__6821),
            .I(N__6794));
    LocalMux I__1449 (
            .O(N__6816),
            .I(N__6794));
    InMux I__1448 (
            .O(N__6813),
            .I(N__6787));
    InMux I__1447 (
            .O(N__6812),
            .I(N__6787));
    InMux I__1446 (
            .O(N__6811),
            .I(N__6787));
    InMux I__1445 (
            .O(N__6810),
            .I(N__6778));
    InMux I__1444 (
            .O(N__6809),
            .I(N__6778));
    InMux I__1443 (
            .O(N__6808),
            .I(N__6778));
    InMux I__1442 (
            .O(N__6807),
            .I(N__6778));
    InMux I__1441 (
            .O(N__6806),
            .I(N__6767));
    InMux I__1440 (
            .O(N__6805),
            .I(N__6767));
    InMux I__1439 (
            .O(N__6804),
            .I(N__6767));
    Span4Mux_s3_h I__1438 (
            .O(N__6799),
            .I(N__6764));
    Span4Mux_v I__1437 (
            .O(N__6794),
            .I(N__6761));
    LocalMux I__1436 (
            .O(N__6787),
            .I(N__6756));
    LocalMux I__1435 (
            .O(N__6778),
            .I(N__6756));
    InMux I__1434 (
            .O(N__6777),
            .I(N__6747));
    InMux I__1433 (
            .O(N__6776),
            .I(N__6747));
    InMux I__1432 (
            .O(N__6775),
            .I(N__6747));
    InMux I__1431 (
            .O(N__6774),
            .I(N__6747));
    LocalMux I__1430 (
            .O(N__6767),
            .I(\uart_tx_inst.n485 ));
    Odrv4 I__1429 (
            .O(N__6764),
            .I(\uart_tx_inst.n485 ));
    Odrv4 I__1428 (
            .O(N__6761),
            .I(\uart_tx_inst.n485 ));
    Odrv12 I__1427 (
            .O(N__6756),
            .I(\uart_tx_inst.n485 ));
    LocalMux I__1426 (
            .O(N__6747),
            .I(\uart_tx_inst.n485 ));
    InMux I__1425 (
            .O(N__6736),
            .I(N__6733));
    LocalMux I__1424 (
            .O(N__6733),
            .I(N__6730));
    Odrv4 I__1423 (
            .O(N__6730),
            .I(\uart_tx_inst.n28 ));
    InMux I__1422 (
            .O(N__6727),
            .I(N__6714));
    InMux I__1421 (
            .O(N__6726),
            .I(N__6714));
    InMux I__1420 (
            .O(N__6725),
            .I(N__6714));
    InMux I__1419 (
            .O(N__6724),
            .I(N__6700));
    InMux I__1418 (
            .O(N__6723),
            .I(N__6700));
    InMux I__1417 (
            .O(N__6722),
            .I(N__6700));
    InMux I__1416 (
            .O(N__6721),
            .I(N__6693));
    LocalMux I__1415 (
            .O(N__6714),
            .I(N__6686));
    InMux I__1414 (
            .O(N__6713),
            .I(N__6677));
    InMux I__1413 (
            .O(N__6712),
            .I(N__6677));
    InMux I__1412 (
            .O(N__6711),
            .I(N__6677));
    InMux I__1411 (
            .O(N__6710),
            .I(N__6677));
    InMux I__1410 (
            .O(N__6709),
            .I(N__6670));
    InMux I__1409 (
            .O(N__6708),
            .I(N__6670));
    InMux I__1408 (
            .O(N__6707),
            .I(N__6670));
    LocalMux I__1407 (
            .O(N__6700),
            .I(N__6664));
    InMux I__1406 (
            .O(N__6699),
            .I(N__6655));
    InMux I__1405 (
            .O(N__6698),
            .I(N__6655));
    InMux I__1404 (
            .O(N__6697),
            .I(N__6655));
    InMux I__1403 (
            .O(N__6696),
            .I(N__6655));
    LocalMux I__1402 (
            .O(N__6693),
            .I(N__6652));
    InMux I__1401 (
            .O(N__6692),
            .I(N__6643));
    InMux I__1400 (
            .O(N__6691),
            .I(N__6643));
    InMux I__1399 (
            .O(N__6690),
            .I(N__6643));
    InMux I__1398 (
            .O(N__6689),
            .I(N__6643));
    Span4Mux_s0_h I__1397 (
            .O(N__6686),
            .I(N__6638));
    LocalMux I__1396 (
            .O(N__6677),
            .I(N__6638));
    LocalMux I__1395 (
            .O(N__6670),
            .I(N__6635));
    InMux I__1394 (
            .O(N__6669),
            .I(N__6632));
    InMux I__1393 (
            .O(N__6668),
            .I(N__6629));
    InMux I__1392 (
            .O(N__6667),
            .I(N__6626));
    Odrv4 I__1391 (
            .O(N__6664),
            .I(input_axis_tready_N_72));
    LocalMux I__1390 (
            .O(N__6655),
            .I(input_axis_tready_N_72));
    Odrv4 I__1389 (
            .O(N__6652),
            .I(input_axis_tready_N_72));
    LocalMux I__1388 (
            .O(N__6643),
            .I(input_axis_tready_N_72));
    Odrv4 I__1387 (
            .O(N__6638),
            .I(input_axis_tready_N_72));
    Odrv4 I__1386 (
            .O(N__6635),
            .I(input_axis_tready_N_72));
    LocalMux I__1385 (
            .O(N__6632),
            .I(input_axis_tready_N_72));
    LocalMux I__1384 (
            .O(N__6629),
            .I(input_axis_tready_N_72));
    LocalMux I__1383 (
            .O(N__6626),
            .I(input_axis_tready_N_72));
    CascadeMux I__1382 (
            .O(N__6607),
            .I(\uart_tx_inst.n885_cascade_ ));
    InMux I__1381 (
            .O(N__6604),
            .I(N__6598));
    InMux I__1380 (
            .O(N__6603),
            .I(N__6598));
    LocalMux I__1379 (
            .O(N__6598),
            .I(N__6589));
    InMux I__1378 (
            .O(N__6597),
            .I(N__6586));
    InMux I__1377 (
            .O(N__6596),
            .I(N__6577));
    InMux I__1376 (
            .O(N__6595),
            .I(N__6577));
    InMux I__1375 (
            .O(N__6594),
            .I(N__6577));
    InMux I__1374 (
            .O(N__6593),
            .I(N__6577));
    CascadeMux I__1373 (
            .O(N__6592),
            .I(N__6563));
    Span4Mux_s1_v I__1372 (
            .O(N__6589),
            .I(N__6560));
    LocalMux I__1371 (
            .O(N__6586),
            .I(N__6555));
    LocalMux I__1370 (
            .O(N__6577),
            .I(N__6555));
    InMux I__1369 (
            .O(N__6576),
            .I(N__6551));
    InMux I__1368 (
            .O(N__6575),
            .I(N__6544));
    InMux I__1367 (
            .O(N__6574),
            .I(N__6544));
    InMux I__1366 (
            .O(N__6573),
            .I(N__6544));
    InMux I__1365 (
            .O(N__6572),
            .I(N__6539));
    InMux I__1364 (
            .O(N__6571),
            .I(N__6539));
    InMux I__1363 (
            .O(N__6570),
            .I(N__6536));
    InMux I__1362 (
            .O(N__6569),
            .I(N__6533));
    InMux I__1361 (
            .O(N__6568),
            .I(N__6524));
    InMux I__1360 (
            .O(N__6567),
            .I(N__6524));
    InMux I__1359 (
            .O(N__6566),
            .I(N__6524));
    InMux I__1358 (
            .O(N__6563),
            .I(N__6524));
    Span4Mux_s0_h I__1357 (
            .O(N__6560),
            .I(N__6519));
    Span4Mux_s1_v I__1356 (
            .O(N__6555),
            .I(N__6519));
    InMux I__1355 (
            .O(N__6554),
            .I(N__6516));
    LocalMux I__1354 (
            .O(N__6551),
            .I(\uart_tx_inst.n165 ));
    LocalMux I__1353 (
            .O(N__6544),
            .I(\uart_tx_inst.n165 ));
    LocalMux I__1352 (
            .O(N__6539),
            .I(\uart_tx_inst.n165 ));
    LocalMux I__1351 (
            .O(N__6536),
            .I(\uart_tx_inst.n165 ));
    LocalMux I__1350 (
            .O(N__6533),
            .I(\uart_tx_inst.n165 ));
    LocalMux I__1349 (
            .O(N__6524),
            .I(\uart_tx_inst.n165 ));
    Odrv4 I__1348 (
            .O(N__6519),
            .I(\uart_tx_inst.n165 ));
    LocalMux I__1347 (
            .O(N__6516),
            .I(\uart_tx_inst.n165 ));
    InMux I__1346 (
            .O(N__6499),
            .I(N__6495));
    CascadeMux I__1345 (
            .O(N__6498),
            .I(N__6492));
    LocalMux I__1344 (
            .O(N__6495),
            .I(N__6489));
    InMux I__1343 (
            .O(N__6492),
            .I(N__6486));
    Odrv4 I__1342 (
            .O(N__6489),
            .I(\uart_tx_inst.prescale_reg_8 ));
    LocalMux I__1341 (
            .O(N__6486),
            .I(\uart_tx_inst.prescale_reg_8 ));
    CEMux I__1340 (
            .O(N__6481),
            .I(N__6478));
    LocalMux I__1339 (
            .O(N__6478),
            .I(N__6472));
    CEMux I__1338 (
            .O(N__6477),
            .I(N__6469));
    CEMux I__1337 (
            .O(N__6476),
            .I(N__6466));
    CEMux I__1336 (
            .O(N__6475),
            .I(N__6461));
    Span4Mux_v I__1335 (
            .O(N__6472),
            .I(N__6454));
    LocalMux I__1334 (
            .O(N__6469),
            .I(N__6454));
    LocalMux I__1333 (
            .O(N__6466),
            .I(N__6454));
    CEMux I__1332 (
            .O(N__6465),
            .I(N__6451));
    CEMux I__1331 (
            .O(N__6464),
            .I(N__6448));
    LocalMux I__1330 (
            .O(N__6461),
            .I(N__6445));
    Span4Mux_h I__1329 (
            .O(N__6454),
            .I(N__6442));
    LocalMux I__1328 (
            .O(N__6451),
            .I(N__6439));
    LocalMux I__1327 (
            .O(N__6448),
            .I(N__6436));
    Span4Mux_s0_v I__1326 (
            .O(N__6445),
            .I(N__6431));
    Span4Mux_s0_h I__1325 (
            .O(N__6442),
            .I(N__6431));
    Odrv12 I__1324 (
            .O(N__6439),
            .I(\uart_tx_inst.n873 ));
    Odrv4 I__1323 (
            .O(N__6436),
            .I(\uart_tx_inst.n873 ));
    Odrv4 I__1322 (
            .O(N__6431),
            .I(\uart_tx_inst.n873 ));
    InMux I__1321 (
            .O(N__6424),
            .I(N__6421));
    LocalMux I__1320 (
            .O(N__6421),
            .I(\uart_tx_inst.data_reg_1 ));
    InMux I__1319 (
            .O(N__6418),
            .I(N__6415));
    LocalMux I__1318 (
            .O(N__6415),
            .I(\uart_tx_inst.data_reg_2 ));
    InMux I__1317 (
            .O(N__6412),
            .I(N__6409));
    LocalMux I__1316 (
            .O(N__6409),
            .I(N__6406));
    Span4Mux_v I__1315 (
            .O(N__6406),
            .I(N__6403));
    Odrv4 I__1314 (
            .O(N__6403),
            .I(\uart_rx_inst.n317 ));
    InMux I__1313 (
            .O(N__6400),
            .I(\uart_rx_inst.n1540 ));
    InMux I__1312 (
            .O(N__6397),
            .I(N__6394));
    LocalMux I__1311 (
            .O(N__6394),
            .I(N__6391));
    Span4Mux_h I__1310 (
            .O(N__6391),
            .I(N__6388));
    Odrv4 I__1309 (
            .O(N__6388),
            .I(\uart_rx_inst.n316 ));
    InMux I__1308 (
            .O(N__6385),
            .I(\uart_rx_inst.n1541 ));
    InMux I__1307 (
            .O(N__6382),
            .I(N__6379));
    LocalMux I__1306 (
            .O(N__6379),
            .I(N__6376));
    Span4Mux_v I__1305 (
            .O(N__6376),
            .I(N__6373));
    Odrv4 I__1304 (
            .O(N__6373),
            .I(\uart_rx_inst.n315 ));
    InMux I__1303 (
            .O(N__6370),
            .I(\uart_rx_inst.n1542 ));
    InMux I__1302 (
            .O(N__6367),
            .I(N__6364));
    LocalMux I__1301 (
            .O(N__6364),
            .I(N__6361));
    Span4Mux_h I__1300 (
            .O(N__6361),
            .I(N__6358));
    Odrv4 I__1299 (
            .O(N__6358),
            .I(\uart_rx_inst.n314 ));
    InMux I__1298 (
            .O(N__6355),
            .I(\uart_rx_inst.n1543 ));
    InMux I__1297 (
            .O(N__6352),
            .I(N__6349));
    LocalMux I__1296 (
            .O(N__6349),
            .I(N__6346));
    Span4Mux_v I__1295 (
            .O(N__6346),
            .I(N__6343));
    Odrv4 I__1294 (
            .O(N__6343),
            .I(\uart_rx_inst.n313 ));
    InMux I__1293 (
            .O(N__6340),
            .I(\uart_rx_inst.n1544 ));
    InMux I__1292 (
            .O(N__6337),
            .I(bfn_11_7_0_));
    InMux I__1291 (
            .O(N__6334),
            .I(N__6331));
    LocalMux I__1290 (
            .O(N__6331),
            .I(N__6328));
    Span4Mux_v I__1289 (
            .O(N__6328),
            .I(N__6325));
    Odrv4 I__1288 (
            .O(N__6325),
            .I(\uart_rx_inst.n312 ));
    InMux I__1287 (
            .O(N__6322),
            .I(N__6315));
    InMux I__1286 (
            .O(N__6321),
            .I(N__6315));
    InMux I__1285 (
            .O(N__6320),
            .I(N__6308));
    LocalMux I__1284 (
            .O(N__6315),
            .I(N__6305));
    InMux I__1283 (
            .O(N__6314),
            .I(N__6289));
    InMux I__1282 (
            .O(N__6313),
            .I(N__6282));
    InMux I__1281 (
            .O(N__6312),
            .I(N__6282));
    InMux I__1280 (
            .O(N__6311),
            .I(N__6279));
    LocalMux I__1279 (
            .O(N__6308),
            .I(N__6276));
    Span4Mux_v I__1278 (
            .O(N__6305),
            .I(N__6273));
    InMux I__1277 (
            .O(N__6304),
            .I(N__6262));
    InMux I__1276 (
            .O(N__6303),
            .I(N__6262));
    InMux I__1275 (
            .O(N__6302),
            .I(N__6262));
    InMux I__1274 (
            .O(N__6301),
            .I(N__6262));
    InMux I__1273 (
            .O(N__6300),
            .I(N__6262));
    InMux I__1272 (
            .O(N__6299),
            .I(N__6245));
    InMux I__1271 (
            .O(N__6298),
            .I(N__6245));
    InMux I__1270 (
            .O(N__6297),
            .I(N__6245));
    InMux I__1269 (
            .O(N__6296),
            .I(N__6245));
    InMux I__1268 (
            .O(N__6295),
            .I(N__6245));
    InMux I__1267 (
            .O(N__6294),
            .I(N__6245));
    InMux I__1266 (
            .O(N__6293),
            .I(N__6245));
    InMux I__1265 (
            .O(N__6292),
            .I(N__6245));
    LocalMux I__1264 (
            .O(N__6289),
            .I(N__6242));
    InMux I__1263 (
            .O(N__6288),
            .I(N__6237));
    InMux I__1262 (
            .O(N__6287),
            .I(N__6237));
    LocalMux I__1261 (
            .O(N__6282),
            .I(\uart_rx_inst.n232 ));
    LocalMux I__1260 (
            .O(N__6279),
            .I(\uart_rx_inst.n232 ));
    Odrv4 I__1259 (
            .O(N__6276),
            .I(\uart_rx_inst.n232 ));
    Odrv4 I__1258 (
            .O(N__6273),
            .I(\uart_rx_inst.n232 ));
    LocalMux I__1257 (
            .O(N__6262),
            .I(\uart_rx_inst.n232 ));
    LocalMux I__1256 (
            .O(N__6245),
            .I(\uart_rx_inst.n232 ));
    Odrv4 I__1255 (
            .O(N__6242),
            .I(\uart_rx_inst.n232 ));
    LocalMux I__1254 (
            .O(N__6237),
            .I(\uart_rx_inst.n232 ));
    InMux I__1253 (
            .O(N__6220),
            .I(N__6217));
    LocalMux I__1252 (
            .O(N__6217),
            .I(N__6214));
    Span4Mux_h I__1251 (
            .O(N__6214),
            .I(N__6211));
    Odrv4 I__1250 (
            .O(N__6211),
            .I(\uart_rx_inst.n1746 ));
    InMux I__1249 (
            .O(N__6208),
            .I(N__6204));
    InMux I__1248 (
            .O(N__6207),
            .I(N__6201));
    LocalMux I__1247 (
            .O(N__6204),
            .I(\uart_tx_inst.prescale_reg_0 ));
    LocalMux I__1246 (
            .O(N__6201),
            .I(\uart_tx_inst.prescale_reg_0 ));
    InMux I__1245 (
            .O(N__6196),
            .I(N__6193));
    LocalMux I__1244 (
            .O(N__6193),
            .I(N__6190));
    Odrv12 I__1243 (
            .O(N__6190),
            .I(\uart_tx_inst.n32_adj_197 ));
    InMux I__1242 (
            .O(N__6187),
            .I(N__6184));
    LocalMux I__1241 (
            .O(N__6184),
            .I(\uart_tx_inst.n32 ));
    InMux I__1240 (
            .O(N__6181),
            .I(N__6178));
    LocalMux I__1239 (
            .O(N__6178),
            .I(N__6175));
    Odrv12 I__1238 (
            .O(N__6175),
            .I(\uart_rx_inst.n325 ));
    InMux I__1237 (
            .O(N__6172),
            .I(\uart_rx_inst.n1532 ));
    CascadeMux I__1236 (
            .O(N__6169),
            .I(N__6166));
    InMux I__1235 (
            .O(N__6166),
            .I(N__6163));
    LocalMux I__1234 (
            .O(N__6163),
            .I(N__6160));
    Odrv4 I__1233 (
            .O(N__6160),
            .I(\uart_rx_inst.n324 ));
    InMux I__1232 (
            .O(N__6157),
            .I(\uart_rx_inst.n1533 ));
    InMux I__1231 (
            .O(N__6154),
            .I(N__6151));
    LocalMux I__1230 (
            .O(N__6151),
            .I(N__6148));
    Odrv4 I__1229 (
            .O(N__6148),
            .I(\uart_rx_inst.n323 ));
    InMux I__1228 (
            .O(N__6145),
            .I(\uart_rx_inst.n1534 ));
    InMux I__1227 (
            .O(N__6142),
            .I(N__6139));
    LocalMux I__1226 (
            .O(N__6139),
            .I(N__6136));
    Span4Mux_h I__1225 (
            .O(N__6136),
            .I(N__6133));
    Odrv4 I__1224 (
            .O(N__6133),
            .I(\uart_rx_inst.n322 ));
    InMux I__1223 (
            .O(N__6130),
            .I(\uart_rx_inst.n1535 ));
    InMux I__1222 (
            .O(N__6127),
            .I(N__6124));
    LocalMux I__1221 (
            .O(N__6124),
            .I(N__6121));
    Odrv4 I__1220 (
            .O(N__6121),
            .I(\uart_rx_inst.n321 ));
    InMux I__1219 (
            .O(N__6118),
            .I(\uart_rx_inst.n1536 ));
    InMux I__1218 (
            .O(N__6115),
            .I(N__6112));
    LocalMux I__1217 (
            .O(N__6112),
            .I(N__6109));
    Span4Mux_v I__1216 (
            .O(N__6109),
            .I(N__6106));
    Odrv4 I__1215 (
            .O(N__6106),
            .I(\uart_rx_inst.n320 ));
    InMux I__1214 (
            .O(N__6103),
            .I(bfn_11_6_0_));
    InMux I__1213 (
            .O(N__6100),
            .I(N__6097));
    LocalMux I__1212 (
            .O(N__6097),
            .I(N__6094));
    Span4Mux_v I__1211 (
            .O(N__6094),
            .I(N__6091));
    Odrv4 I__1210 (
            .O(N__6091),
            .I(\uart_rx_inst.n319 ));
    InMux I__1209 (
            .O(N__6088),
            .I(\uart_rx_inst.n1538 ));
    InMux I__1208 (
            .O(N__6085),
            .I(N__6082));
    LocalMux I__1207 (
            .O(N__6082),
            .I(N__6079));
    Span4Mux_h I__1206 (
            .O(N__6079),
            .I(N__6076));
    Odrv4 I__1205 (
            .O(N__6076),
            .I(\uart_rx_inst.n318 ));
    InMux I__1204 (
            .O(N__6073),
            .I(\uart_rx_inst.n1539 ));
    InMux I__1203 (
            .O(N__6070),
            .I(N__6067));
    LocalMux I__1202 (
            .O(N__6067),
            .I(N__6064));
    Span4Mux_s2_h I__1201 (
            .O(N__6064),
            .I(N__6060));
    InMux I__1200 (
            .O(N__6063),
            .I(N__6057));
    Odrv4 I__1199 (
            .O(N__6060),
            .I(\uart_tx_inst.prescale_reg_14 ));
    LocalMux I__1198 (
            .O(N__6057),
            .I(\uart_tx_inst.prescale_reg_14 ));
    InMux I__1197 (
            .O(N__6052),
            .I(N__6049));
    LocalMux I__1196 (
            .O(N__6049),
            .I(N__6046));
    Span4Mux_s2_v I__1195 (
            .O(N__6046),
            .I(N__6043));
    Odrv4 I__1194 (
            .O(N__6043),
            .I(\uart_tx_inst.n22 ));
    InMux I__1193 (
            .O(N__6040),
            .I(\uart_tx_inst.n1559 ));
    CascadeMux I__1192 (
            .O(N__6037),
            .I(N__6034));
    InMux I__1191 (
            .O(N__6034),
            .I(N__6031));
    LocalMux I__1190 (
            .O(N__6031),
            .I(N__6028));
    Span4Mux_v I__1189 (
            .O(N__6028),
            .I(N__6024));
    InMux I__1188 (
            .O(N__6027),
            .I(N__6021));
    Odrv4 I__1187 (
            .O(N__6024),
            .I(\uart_tx_inst.prescale_reg_15 ));
    LocalMux I__1186 (
            .O(N__6021),
            .I(\uart_tx_inst.prescale_reg_15 ));
    InMux I__1185 (
            .O(N__6016),
            .I(N__6013));
    LocalMux I__1184 (
            .O(N__6013),
            .I(N__6010));
    Span4Mux_s2_v I__1183 (
            .O(N__6010),
            .I(N__6007));
    Odrv4 I__1182 (
            .O(N__6007),
            .I(\uart_tx_inst.n21 ));
    InMux I__1181 (
            .O(N__6004),
            .I(\uart_tx_inst.n1560 ));
    InMux I__1180 (
            .O(N__6001),
            .I(N__5997));
    CascadeMux I__1179 (
            .O(N__6000),
            .I(N__5994));
    LocalMux I__1178 (
            .O(N__5997),
            .I(N__5991));
    InMux I__1177 (
            .O(N__5994),
            .I(N__5988));
    Span4Mux_s2_h I__1176 (
            .O(N__5991),
            .I(N__5985));
    LocalMux I__1175 (
            .O(N__5988),
            .I(N__5982));
    Odrv4 I__1174 (
            .O(N__5985),
            .I(\uart_tx_inst.prescale_reg_16 ));
    Odrv4 I__1173 (
            .O(N__5982),
            .I(\uart_tx_inst.prescale_reg_16 ));
    InMux I__1172 (
            .O(N__5977),
            .I(N__5974));
    LocalMux I__1171 (
            .O(N__5974),
            .I(N__5971));
    Odrv4 I__1170 (
            .O(N__5971),
            .I(\uart_tx_inst.n20 ));
    InMux I__1169 (
            .O(N__5968),
            .I(bfn_11_4_0_));
    CascadeMux I__1168 (
            .O(N__5965),
            .I(N__5962));
    InMux I__1167 (
            .O(N__5962),
            .I(N__5959));
    LocalMux I__1166 (
            .O(N__5959),
            .I(N__5956));
    Span4Mux_s2_h I__1165 (
            .O(N__5956),
            .I(N__5952));
    InMux I__1164 (
            .O(N__5955),
            .I(N__5949));
    Odrv4 I__1163 (
            .O(N__5952),
            .I(\uart_tx_inst.prescale_reg_17 ));
    LocalMux I__1162 (
            .O(N__5949),
            .I(\uart_tx_inst.prescale_reg_17 ));
    InMux I__1161 (
            .O(N__5944),
            .I(N__5941));
    LocalMux I__1160 (
            .O(N__5941),
            .I(N__5938));
    Span4Mux_h I__1159 (
            .O(N__5938),
            .I(N__5935));
    Odrv4 I__1158 (
            .O(N__5935),
            .I(\uart_tx_inst.n19 ));
    InMux I__1157 (
            .O(N__5932),
            .I(\uart_tx_inst.n1562 ));
    InMux I__1156 (
            .O(N__5929),
            .I(N__5925));
    CascadeMux I__1155 (
            .O(N__5928),
            .I(N__5922));
    LocalMux I__1154 (
            .O(N__5925),
            .I(N__5919));
    InMux I__1153 (
            .O(N__5922),
            .I(N__5916));
    Span4Mux_v I__1152 (
            .O(N__5919),
            .I(N__5913));
    LocalMux I__1151 (
            .O(N__5916),
            .I(N__5910));
    Odrv4 I__1150 (
            .O(N__5913),
            .I(\uart_tx_inst.prescale_reg_18 ));
    Odrv4 I__1149 (
            .O(N__5910),
            .I(\uart_tx_inst.prescale_reg_18 ));
    InMux I__1148 (
            .O(N__5905),
            .I(\uart_tx_inst.n1563 ));
    InMux I__1147 (
            .O(N__5902),
            .I(N__5899));
    LocalMux I__1146 (
            .O(N__5899),
            .I(N__5896));
    Odrv4 I__1145 (
            .O(N__5896),
            .I(\uart_tx_inst.n18 ));
    InMux I__1144 (
            .O(N__5893),
            .I(N__5890));
    LocalMux I__1143 (
            .O(N__5890),
            .I(N__5887));
    Span4Mux_h I__1142 (
            .O(N__5887),
            .I(N__5884));
    Odrv4 I__1141 (
            .O(N__5884),
            .I(\uart_rx_inst.n328 ));
    InMux I__1140 (
            .O(N__5881),
            .I(bfn_11_5_0_));
    InMux I__1139 (
            .O(N__5878),
            .I(N__5875));
    LocalMux I__1138 (
            .O(N__5875),
            .I(N__5872));
    Odrv12 I__1137 (
            .O(N__5872),
            .I(\uart_rx_inst.n327 ));
    InMux I__1136 (
            .O(N__5869),
            .I(\uart_rx_inst.n1530 ));
    InMux I__1135 (
            .O(N__5866),
            .I(N__5863));
    LocalMux I__1134 (
            .O(N__5863),
            .I(N__5860));
    Odrv12 I__1133 (
            .O(N__5860),
            .I(\uart_rx_inst.n326 ));
    InMux I__1132 (
            .O(N__5857),
            .I(\uart_rx_inst.n1531 ));
    CascadeMux I__1131 (
            .O(N__5854),
            .I(N__5851));
    InMux I__1130 (
            .O(N__5851),
            .I(N__5847));
    InMux I__1129 (
            .O(N__5850),
            .I(N__5844));
    LocalMux I__1128 (
            .O(N__5847),
            .I(N__5841));
    LocalMux I__1127 (
            .O(N__5844),
            .I(\uart_tx_inst.prescale_reg_6 ));
    Odrv4 I__1126 (
            .O(N__5841),
            .I(\uart_tx_inst.prescale_reg_6 ));
    InMux I__1125 (
            .O(N__5836),
            .I(N__5833));
    LocalMux I__1124 (
            .O(N__5833),
            .I(N__5830));
    Odrv12 I__1123 (
            .O(N__5830),
            .I(\uart_tx_inst.n30 ));
    InMux I__1122 (
            .O(N__5827),
            .I(\uart_tx_inst.n1551 ));
    InMux I__1121 (
            .O(N__5824),
            .I(N__5820));
    InMux I__1120 (
            .O(N__5823),
            .I(N__5817));
    LocalMux I__1119 (
            .O(N__5820),
            .I(N__5814));
    LocalMux I__1118 (
            .O(N__5817),
            .I(\uart_tx_inst.prescale_reg_7 ));
    Odrv4 I__1117 (
            .O(N__5814),
            .I(\uart_tx_inst.prescale_reg_7 ));
    InMux I__1116 (
            .O(N__5809),
            .I(N__5806));
    LocalMux I__1115 (
            .O(N__5806),
            .I(N__5803));
    Odrv4 I__1114 (
            .O(N__5803),
            .I(\uart_tx_inst.n29 ));
    InMux I__1113 (
            .O(N__5800),
            .I(\uart_tx_inst.n1552 ));
    InMux I__1112 (
            .O(N__5797),
            .I(bfn_11_3_0_));
    CascadeMux I__1111 (
            .O(N__5794),
            .I(N__5791));
    InMux I__1110 (
            .O(N__5791),
            .I(N__5787));
    CascadeMux I__1109 (
            .O(N__5790),
            .I(N__5784));
    LocalMux I__1108 (
            .O(N__5787),
            .I(N__5781));
    InMux I__1107 (
            .O(N__5784),
            .I(N__5778));
    Odrv4 I__1106 (
            .O(N__5781),
            .I(\uart_tx_inst.prescale_reg_9 ));
    LocalMux I__1105 (
            .O(N__5778),
            .I(\uart_tx_inst.prescale_reg_9 ));
    InMux I__1104 (
            .O(N__5773),
            .I(N__5770));
    LocalMux I__1103 (
            .O(N__5770),
            .I(N__5767));
    Odrv4 I__1102 (
            .O(N__5767),
            .I(\uart_tx_inst.n27 ));
    InMux I__1101 (
            .O(N__5764),
            .I(\uart_tx_inst.n1554 ));
    InMux I__1100 (
            .O(N__5761),
            .I(N__5758));
    LocalMux I__1099 (
            .O(N__5758),
            .I(N__5755));
    Span4Mux_s2_h I__1098 (
            .O(N__5755),
            .I(N__5751));
    InMux I__1097 (
            .O(N__5754),
            .I(N__5748));
    Odrv4 I__1096 (
            .O(N__5751),
            .I(\uart_tx_inst.prescale_reg_10 ));
    LocalMux I__1095 (
            .O(N__5748),
            .I(\uart_tx_inst.prescale_reg_10 ));
    InMux I__1094 (
            .O(N__5743),
            .I(N__5740));
    LocalMux I__1093 (
            .O(N__5740),
            .I(N__5737));
    Span4Mux_s2_v I__1092 (
            .O(N__5737),
            .I(N__5734));
    Odrv4 I__1091 (
            .O(N__5734),
            .I(\uart_tx_inst.n26 ));
    InMux I__1090 (
            .O(N__5731),
            .I(\uart_tx_inst.n1555 ));
    CascadeMux I__1089 (
            .O(N__5728),
            .I(N__5725));
    InMux I__1088 (
            .O(N__5725),
            .I(N__5721));
    InMux I__1087 (
            .O(N__5724),
            .I(N__5718));
    LocalMux I__1086 (
            .O(N__5721),
            .I(N__5715));
    LocalMux I__1085 (
            .O(N__5718),
            .I(N__5712));
    Odrv4 I__1084 (
            .O(N__5715),
            .I(\uart_tx_inst.prescale_reg_11 ));
    Odrv4 I__1083 (
            .O(N__5712),
            .I(\uart_tx_inst.prescale_reg_11 ));
    InMux I__1082 (
            .O(N__5707),
            .I(N__5704));
    LocalMux I__1081 (
            .O(N__5704),
            .I(N__5701));
    Odrv4 I__1080 (
            .O(N__5701),
            .I(\uart_tx_inst.n25 ));
    InMux I__1079 (
            .O(N__5698),
            .I(\uart_tx_inst.n1556 ));
    InMux I__1078 (
            .O(N__5695),
            .I(N__5692));
    LocalMux I__1077 (
            .O(N__5692),
            .I(N__5688));
    InMux I__1076 (
            .O(N__5691),
            .I(N__5685));
    Odrv4 I__1075 (
            .O(N__5688),
            .I(\uart_tx_inst.prescale_reg_12 ));
    LocalMux I__1074 (
            .O(N__5685),
            .I(\uart_tx_inst.prescale_reg_12 ));
    InMux I__1073 (
            .O(N__5680),
            .I(N__5677));
    LocalMux I__1072 (
            .O(N__5677),
            .I(N__5674));
    Odrv4 I__1071 (
            .O(N__5674),
            .I(\uart_tx_inst.n24 ));
    InMux I__1070 (
            .O(N__5671),
            .I(\uart_tx_inst.n1557 ));
    CascadeMux I__1069 (
            .O(N__5668),
            .I(N__5665));
    InMux I__1068 (
            .O(N__5665),
            .I(N__5662));
    LocalMux I__1067 (
            .O(N__5662),
            .I(N__5659));
    Span4Mux_s2_h I__1066 (
            .O(N__5659),
            .I(N__5655));
    InMux I__1065 (
            .O(N__5658),
            .I(N__5652));
    Odrv4 I__1064 (
            .O(N__5655),
            .I(\uart_tx_inst.prescale_reg_13 ));
    LocalMux I__1063 (
            .O(N__5652),
            .I(\uart_tx_inst.prescale_reg_13 ));
    InMux I__1062 (
            .O(N__5647),
            .I(N__5644));
    LocalMux I__1061 (
            .O(N__5644),
            .I(N__5641));
    Span4Mux_s2_v I__1060 (
            .O(N__5641),
            .I(N__5638));
    Odrv4 I__1059 (
            .O(N__5638),
            .I(\uart_tx_inst.n23 ));
    InMux I__1058 (
            .O(N__5635),
            .I(\uart_tx_inst.n1558 ));
    CascadeMux I__1057 (
            .O(N__5632),
            .I(\uart_tx_inst.n860_cascade_ ));
    InMux I__1056 (
            .O(N__5629),
            .I(bfn_11_2_0_));
    InMux I__1055 (
            .O(N__5626),
            .I(N__5622));
    InMux I__1054 (
            .O(N__5625),
            .I(N__5619));
    LocalMux I__1053 (
            .O(N__5622),
            .I(\uart_tx_inst.prescale_reg_1 ));
    LocalMux I__1052 (
            .O(N__5619),
            .I(\uart_tx_inst.prescale_reg_1 ));
    InMux I__1051 (
            .O(N__5614),
            .I(\uart_tx_inst.n1546 ));
    InMux I__1050 (
            .O(N__5611),
            .I(N__5607));
    InMux I__1049 (
            .O(N__5610),
            .I(N__5604));
    LocalMux I__1048 (
            .O(N__5607),
            .I(\uart_tx_inst.prescale_reg_2 ));
    LocalMux I__1047 (
            .O(N__5604),
            .I(\uart_tx_inst.prescale_reg_2 ));
    InMux I__1046 (
            .O(N__5599),
            .I(\uart_tx_inst.n1547 ));
    SRMux I__1045 (
            .O(N__5596),
            .I(N__5593));
    LocalMux I__1044 (
            .O(N__5593),
            .I(N__5590));
    Odrv12 I__1043 (
            .O(N__5590),
            .I(\uart_tx_inst.n1170 ));
    InMux I__1042 (
            .O(N__5587),
            .I(N__5583));
    InMux I__1041 (
            .O(N__5586),
            .I(N__5580));
    LocalMux I__1040 (
            .O(N__5583),
            .I(N__5577));
    LocalMux I__1039 (
            .O(N__5580),
            .I(\uart_tx_inst.prescale_reg_3 ));
    Odrv4 I__1038 (
            .O(N__5577),
            .I(\uart_tx_inst.prescale_reg_3 ));
    InMux I__1037 (
            .O(N__5572),
            .I(N__5569));
    LocalMux I__1036 (
            .O(N__5569),
            .I(\uart_tx_inst.n33 ));
    InMux I__1035 (
            .O(N__5566),
            .I(\uart_tx_inst.n1548 ));
    InMux I__1034 (
            .O(N__5563),
            .I(\uart_tx_inst.n1549 ));
    InMux I__1033 (
            .O(N__5560),
            .I(\uart_tx_inst.n1550 ));
    InMux I__1032 (
            .O(N__5557),
            .I(N__5554));
    LocalMux I__1031 (
            .O(N__5554),
            .I(N__5549));
    InMux I__1030 (
            .O(N__5553),
            .I(N__5544));
    InMux I__1029 (
            .O(N__5552),
            .I(N__5544));
    Odrv4 I__1028 (
            .O(N__5549),
            .I(data_reg_4));
    LocalMux I__1027 (
            .O(N__5544),
            .I(data_reg_4));
    IoInMux I__1026 (
            .O(N__5539),
            .I(N__5536));
    LocalMux I__1025 (
            .O(N__5536),
            .I(N__5533));
    Span4Mux_s1_v I__1024 (
            .O(N__5533),
            .I(N__5530));
    Odrv4 I__1023 (
            .O(N__5530),
            .I(output_axis_tdata_c_4));
    InMux I__1022 (
            .O(N__5527),
            .I(N__5523));
    CascadeMux I__1021 (
            .O(N__5526),
            .I(N__5520));
    LocalMux I__1020 (
            .O(N__5523),
            .I(N__5516));
    InMux I__1019 (
            .O(N__5520),
            .I(N__5511));
    InMux I__1018 (
            .O(N__5519),
            .I(N__5511));
    Odrv12 I__1017 (
            .O(N__5516),
            .I(data_reg_5));
    LocalMux I__1016 (
            .O(N__5511),
            .I(data_reg_5));
    IoInMux I__1015 (
            .O(N__5506),
            .I(N__5503));
    LocalMux I__1014 (
            .O(N__5503),
            .I(N__5500));
    Span4Mux_s1_v I__1013 (
            .O(N__5500),
            .I(N__5497));
    Odrv4 I__1012 (
            .O(N__5497),
            .I(output_axis_tdata_c_5));
    CascadeMux I__1011 (
            .O(N__5494),
            .I(N__5490));
    InMux I__1010 (
            .O(N__5493),
            .I(N__5487));
    InMux I__1009 (
            .O(N__5490),
            .I(N__5484));
    LocalMux I__1008 (
            .O(N__5487),
            .I(N__5480));
    LocalMux I__1007 (
            .O(N__5484),
            .I(N__5477));
    InMux I__1006 (
            .O(N__5483),
            .I(N__5474));
    Odrv12 I__1005 (
            .O(N__5480),
            .I(data_reg_1));
    Odrv4 I__1004 (
            .O(N__5477),
            .I(data_reg_1));
    LocalMux I__1003 (
            .O(N__5474),
            .I(data_reg_1));
    IoInMux I__1002 (
            .O(N__5467),
            .I(N__5464));
    LocalMux I__1001 (
            .O(N__5464),
            .I(N__5461));
    Span4Mux_s3_v I__1000 (
            .O(N__5461),
            .I(N__5458));
    Odrv4 I__999 (
            .O(N__5458),
            .I(output_axis_tdata_c_1));
    CascadeMux I__998 (
            .O(N__5455),
            .I(N__5450));
    InMux I__997 (
            .O(N__5454),
            .I(N__5447));
    InMux I__996 (
            .O(N__5453),
            .I(N__5444));
    InMux I__995 (
            .O(N__5450),
            .I(N__5441));
    LocalMux I__994 (
            .O(N__5447),
            .I(N__5438));
    LocalMux I__993 (
            .O(N__5444),
            .I(data_reg_3));
    LocalMux I__992 (
            .O(N__5441),
            .I(data_reg_3));
    Odrv12 I__991 (
            .O(N__5438),
            .I(data_reg_3));
    IoInMux I__990 (
            .O(N__5431),
            .I(N__5428));
    LocalMux I__989 (
            .O(N__5428),
            .I(N__5425));
    Span4Mux_s3_v I__988 (
            .O(N__5425),
            .I(N__5422));
    Odrv4 I__987 (
            .O(N__5422),
            .I(output_axis_tdata_c_3));
    CEMux I__986 (
            .O(N__5419),
            .I(N__5415));
    CEMux I__985 (
            .O(N__5418),
            .I(N__5412));
    LocalMux I__984 (
            .O(N__5415),
            .I(N__5409));
    LocalMux I__983 (
            .O(N__5412),
            .I(N__5405));
    Span4Mux_v I__982 (
            .O(N__5409),
            .I(N__5402));
    CEMux I__981 (
            .O(N__5408),
            .I(N__5399));
    Span4Mux_v I__980 (
            .O(N__5405),
            .I(N__5396));
    Span4Mux_s1_v I__979 (
            .O(N__5402),
            .I(N__5393));
    LocalMux I__978 (
            .O(N__5399),
            .I(N__5390));
    Span4Mux_s1_v I__977 (
            .O(N__5396),
            .I(N__5387));
    Odrv4 I__976 (
            .O(N__5393),
            .I(n703));
    Odrv12 I__975 (
            .O(N__5390),
            .I(n703));
    Odrv4 I__974 (
            .O(N__5387),
            .I(n703));
    CascadeMux I__973 (
            .O(N__5380),
            .I(\uart_tx_inst.n905_cascade_ ));
    CascadeMux I__972 (
            .O(N__5377),
            .I(\uart_tx_inst.n890_cascade_ ));
    InMux I__971 (
            .O(N__5374),
            .I(N__5371));
    LocalMux I__970 (
            .O(N__5371),
            .I(N__5368));
    Odrv4 I__969 (
            .O(N__5368),
            .I(\uart_tx_inst.n33_adj_198 ));
    InMux I__968 (
            .O(N__5365),
            .I(N__5356));
    InMux I__967 (
            .O(N__5364),
            .I(N__5348));
    InMux I__966 (
            .O(N__5363),
            .I(N__5348));
    InMux I__965 (
            .O(N__5362),
            .I(N__5348));
    InMux I__964 (
            .O(N__5361),
            .I(N__5341));
    InMux I__963 (
            .O(N__5360),
            .I(N__5341));
    InMux I__962 (
            .O(N__5359),
            .I(N__5341));
    LocalMux I__961 (
            .O(N__5356),
            .I(N__5338));
    InMux I__960 (
            .O(N__5355),
            .I(N__5335));
    LocalMux I__959 (
            .O(N__5348),
            .I(n1711));
    LocalMux I__958 (
            .O(N__5341),
            .I(n1711));
    Odrv4 I__957 (
            .O(N__5338),
            .I(n1711));
    LocalMux I__956 (
            .O(N__5335),
            .I(n1711));
    InMux I__955 (
            .O(N__5326),
            .I(N__5317));
    InMux I__954 (
            .O(N__5325),
            .I(N__5304));
    InMux I__953 (
            .O(N__5324),
            .I(N__5304));
    InMux I__952 (
            .O(N__5323),
            .I(N__5304));
    InMux I__951 (
            .O(N__5322),
            .I(N__5304));
    InMux I__950 (
            .O(N__5321),
            .I(N__5304));
    InMux I__949 (
            .O(N__5320),
            .I(N__5304));
    LocalMux I__948 (
            .O(N__5317),
            .I(N__5301));
    LocalMux I__947 (
            .O(N__5304),
            .I(n1220));
    Odrv4 I__946 (
            .O(N__5301),
            .I(n1220));
    InMux I__945 (
            .O(N__5296),
            .I(N__5286));
    InMux I__944 (
            .O(N__5295),
            .I(N__5286));
    InMux I__943 (
            .O(N__5294),
            .I(N__5283));
    InMux I__942 (
            .O(N__5293),
            .I(N__5279));
    InMux I__941 (
            .O(N__5292),
            .I(N__5276));
    InMux I__940 (
            .O(N__5291),
            .I(N__5273));
    LocalMux I__939 (
            .O(N__5286),
            .I(N__5266));
    LocalMux I__938 (
            .O(N__5283),
            .I(N__5263));
    InMux I__937 (
            .O(N__5282),
            .I(N__5260));
    LocalMux I__936 (
            .O(N__5279),
            .I(N__5257));
    LocalMux I__935 (
            .O(N__5276),
            .I(N__5254));
    LocalMux I__934 (
            .O(N__5273),
            .I(N__5251));
    InMux I__933 (
            .O(N__5272),
            .I(N__5242));
    InMux I__932 (
            .O(N__5271),
            .I(N__5242));
    InMux I__931 (
            .O(N__5270),
            .I(N__5242));
    InMux I__930 (
            .O(N__5269),
            .I(N__5242));
    Span4Mux_v I__929 (
            .O(N__5266),
            .I(N__5233));
    Span4Mux_h I__928 (
            .O(N__5263),
            .I(N__5233));
    LocalMux I__927 (
            .O(N__5260),
            .I(N__5233));
    Span4Mux_v I__926 (
            .O(N__5257),
            .I(N__5233));
    Span12Mux_v I__925 (
            .O(N__5254),
            .I(N__5230));
    Span12Mux_s7_h I__924 (
            .O(N__5251),
            .I(N__5225));
    LocalMux I__923 (
            .O(N__5242),
            .I(N__5225));
    Odrv4 I__922 (
            .O(N__5233),
            .I(rxd_reg));
    Odrv12 I__921 (
            .O(N__5230),
            .I(rxd_reg));
    Odrv12 I__920 (
            .O(N__5225),
            .I(rxd_reg));
    IoInMux I__919 (
            .O(N__5218),
            .I(N__5215));
    LocalMux I__918 (
            .O(N__5215),
            .I(N__5212));
    Span4Mux_s3_h I__917 (
            .O(N__5212),
            .I(N__5209));
    Odrv4 I__916 (
            .O(N__5209),
            .I(rx_frame_error_c));
    SRMux I__915 (
            .O(N__5206),
            .I(N__5203));
    LocalMux I__914 (
            .O(N__5203),
            .I(N__5200));
    Span4Mux_h I__913 (
            .O(N__5200),
            .I(N__5197));
    Odrv4 I__912 (
            .O(N__5197),
            .I(n697));
    InMux I__911 (
            .O(N__5194),
            .I(N__5190));
    CascadeMux I__910 (
            .O(N__5193),
            .I(N__5187));
    LocalMux I__909 (
            .O(N__5190),
            .I(N__5183));
    InMux I__908 (
            .O(N__5187),
            .I(N__5178));
    InMux I__907 (
            .O(N__5186),
            .I(N__5178));
    Odrv4 I__906 (
            .O(N__5183),
            .I(data_reg_6));
    LocalMux I__905 (
            .O(N__5178),
            .I(data_reg_6));
    IoInMux I__904 (
            .O(N__5173),
            .I(N__5170));
    LocalMux I__903 (
            .O(N__5170),
            .I(N__5167));
    Odrv12 I__902 (
            .O(N__5167),
            .I(output_axis_tdata_c_6));
    CascadeMux I__901 (
            .O(N__5164),
            .I(N__5159));
    CascadeMux I__900 (
            .O(N__5163),
            .I(N__5156));
    InMux I__899 (
            .O(N__5162),
            .I(N__5153));
    InMux I__898 (
            .O(N__5159),
            .I(N__5150));
    InMux I__897 (
            .O(N__5156),
            .I(N__5147));
    LocalMux I__896 (
            .O(N__5153),
            .I(N__5144));
    LocalMux I__895 (
            .O(N__5150),
            .I(data_reg_2));
    LocalMux I__894 (
            .O(N__5147),
            .I(data_reg_2));
    Odrv12 I__893 (
            .O(N__5144),
            .I(data_reg_2));
    IoInMux I__892 (
            .O(N__5137),
            .I(N__5134));
    LocalMux I__891 (
            .O(N__5134),
            .I(N__5131));
    IoSpan4Mux I__890 (
            .O(N__5131),
            .I(N__5128));
    Span4Mux_s1_v I__889 (
            .O(N__5128),
            .I(N__5125));
    Odrv4 I__888 (
            .O(N__5125),
            .I(output_axis_tdata_c_2));
    InMux I__887 (
            .O(N__5122),
            .I(N__5119));
    LocalMux I__886 (
            .O(N__5119),
            .I(N__5115));
    CascadeMux I__885 (
            .O(N__5118),
            .I(N__5112));
    Span4Mux_v I__884 (
            .O(N__5115),
            .I(N__5108));
    InMux I__883 (
            .O(N__5112),
            .I(N__5105));
    InMux I__882 (
            .O(N__5111),
            .I(N__5102));
    Odrv4 I__881 (
            .O(N__5108),
            .I(data_reg_7));
    LocalMux I__880 (
            .O(N__5105),
            .I(data_reg_7));
    LocalMux I__879 (
            .O(N__5102),
            .I(data_reg_7));
    IoInMux I__878 (
            .O(N__5095),
            .I(N__5092));
    LocalMux I__877 (
            .O(N__5092),
            .I(N__5089));
    Odrv12 I__876 (
            .O(N__5089),
            .I(output_axis_tdata_c_7));
    InMux I__875 (
            .O(N__5086),
            .I(N__5083));
    LocalMux I__874 (
            .O(N__5083),
            .I(N__5080));
    Odrv4 I__873 (
            .O(N__5080),
            .I(\uart_rx_inst.n1750 ));
    InMux I__872 (
            .O(N__5077),
            .I(N__5074));
    LocalMux I__871 (
            .O(N__5074),
            .I(N__5071));
    Odrv4 I__870 (
            .O(N__5071),
            .I(\uart_rx_inst.n1755 ));
    CascadeMux I__869 (
            .O(N__5068),
            .I(N__5065));
    InMux I__868 (
            .O(N__5065),
            .I(N__5062));
    LocalMux I__867 (
            .O(N__5062),
            .I(\uart_rx_inst.n1754 ));
    InMux I__866 (
            .O(N__5059),
            .I(N__5056));
    LocalMux I__865 (
            .O(N__5056),
            .I(N__5053));
    Odrv4 I__864 (
            .O(N__5053),
            .I(\uart_rx_inst.n1751 ));
    InMux I__863 (
            .O(N__5050),
            .I(N__5047));
    LocalMux I__862 (
            .O(N__5047),
            .I(N__5044));
    Odrv4 I__861 (
            .O(N__5044),
            .I(\uart_rx_inst.n1758 ));
    InMux I__860 (
            .O(N__5041),
            .I(N__5038));
    LocalMux I__859 (
            .O(N__5038),
            .I(\uart_rx_inst.n1742 ));
    InMux I__858 (
            .O(N__5035),
            .I(N__5032));
    LocalMux I__857 (
            .O(N__5032),
            .I(N__5029));
    Odrv12 I__856 (
            .O(N__5029),
            .I(\uart_rx_inst.n1739 ));
    InMux I__855 (
            .O(N__5026),
            .I(N__5023));
    LocalMux I__854 (
            .O(N__5023),
            .I(N__5020));
    Odrv12 I__853 (
            .O(N__5020),
            .I(\uart_rx_inst.n1757 ));
    CascadeMux I__852 (
            .O(N__5017),
            .I(N__5014));
    InMux I__851 (
            .O(N__5014),
            .I(N__5010));
    InMux I__850 (
            .O(N__5013),
            .I(N__5007));
    LocalMux I__849 (
            .O(N__5010),
            .I(\uart_rx_inst.prescale_reg_15 ));
    LocalMux I__848 (
            .O(N__5007),
            .I(\uart_rx_inst.prescale_reg_15 ));
    InMux I__847 (
            .O(N__5002),
            .I(N__4999));
    LocalMux I__846 (
            .O(N__4999),
            .I(\uart_rx_inst.n749 ));
    InMux I__845 (
            .O(N__4996),
            .I(\uart_rx_inst.n1578 ));
    CascadeMux I__844 (
            .O(N__4993),
            .I(N__4989));
    InMux I__843 (
            .O(N__4992),
            .I(N__4986));
    InMux I__842 (
            .O(N__4989),
            .I(N__4983));
    LocalMux I__841 (
            .O(N__4986),
            .I(\uart_rx_inst.prescale_reg_16 ));
    LocalMux I__840 (
            .O(N__4983),
            .I(\uart_rx_inst.prescale_reg_16 ));
    InMux I__839 (
            .O(N__4978),
            .I(N__4975));
    LocalMux I__838 (
            .O(N__4975),
            .I(\uart_rx_inst.n744 ));
    InMux I__837 (
            .O(N__4972),
            .I(bfn_9_7_0_));
    CascadeMux I__836 (
            .O(N__4969),
            .I(N__4966));
    InMux I__835 (
            .O(N__4966),
            .I(N__4963));
    LocalMux I__834 (
            .O(N__4963),
            .I(N__4959));
    InMux I__833 (
            .O(N__4962),
            .I(N__4956));
    Odrv4 I__832 (
            .O(N__4959),
            .I(\uart_rx_inst.prescale_reg_17 ));
    LocalMux I__831 (
            .O(N__4956),
            .I(\uart_rx_inst.prescale_reg_17 ));
    InMux I__830 (
            .O(N__4951),
            .I(N__4948));
    LocalMux I__829 (
            .O(N__4948),
            .I(\uart_rx_inst.n739 ));
    InMux I__828 (
            .O(N__4945),
            .I(\uart_rx_inst.n1580 ));
    CascadeMux I__827 (
            .O(N__4942),
            .I(N__4929));
    CascadeMux I__826 (
            .O(N__4941),
            .I(N__4925));
    CascadeMux I__825 (
            .O(N__4940),
            .I(N__4921));
    CascadeMux I__824 (
            .O(N__4939),
            .I(N__4917));
    CascadeMux I__823 (
            .O(N__4938),
            .I(N__4913));
    CascadeMux I__822 (
            .O(N__4937),
            .I(N__4910));
    CascadeMux I__821 (
            .O(N__4936),
            .I(N__4906));
    CascadeMux I__820 (
            .O(N__4935),
            .I(N__4902));
    CascadeMux I__819 (
            .O(N__4934),
            .I(N__4898));
    InMux I__818 (
            .O(N__4933),
            .I(N__4891));
    InMux I__817 (
            .O(N__4932),
            .I(N__4891));
    InMux I__816 (
            .O(N__4929),
            .I(N__4891));
    InMux I__815 (
            .O(N__4928),
            .I(N__4874));
    InMux I__814 (
            .O(N__4925),
            .I(N__4874));
    InMux I__813 (
            .O(N__4924),
            .I(N__4874));
    InMux I__812 (
            .O(N__4921),
            .I(N__4874));
    InMux I__811 (
            .O(N__4920),
            .I(N__4874));
    InMux I__810 (
            .O(N__4917),
            .I(N__4874));
    InMux I__809 (
            .O(N__4916),
            .I(N__4874));
    InMux I__808 (
            .O(N__4913),
            .I(N__4874));
    InMux I__807 (
            .O(N__4910),
            .I(N__4859));
    InMux I__806 (
            .O(N__4909),
            .I(N__4859));
    InMux I__805 (
            .O(N__4906),
            .I(N__4859));
    InMux I__804 (
            .O(N__4905),
            .I(N__4859));
    InMux I__803 (
            .O(N__4902),
            .I(N__4859));
    InMux I__802 (
            .O(N__4901),
            .I(N__4859));
    InMux I__801 (
            .O(N__4898),
            .I(N__4859));
    LocalMux I__800 (
            .O(N__4891),
            .I(\uart_rx_inst.n712 ));
    LocalMux I__799 (
            .O(N__4874),
            .I(\uart_rx_inst.n712 ));
    LocalMux I__798 (
            .O(N__4859),
            .I(\uart_rx_inst.n712 ));
    InMux I__797 (
            .O(N__4852),
            .I(N__4849));
    LocalMux I__796 (
            .O(N__4849),
            .I(N__4845));
    InMux I__795 (
            .O(N__4848),
            .I(N__4842));
    Odrv4 I__794 (
            .O(N__4845),
            .I(\uart_rx_inst.prescale_reg_18 ));
    LocalMux I__793 (
            .O(N__4842),
            .I(\uart_rx_inst.prescale_reg_18 ));
    InMux I__792 (
            .O(N__4837),
            .I(\uart_rx_inst.n1581 ));
    InMux I__791 (
            .O(N__4834),
            .I(N__4831));
    LocalMux I__790 (
            .O(N__4831),
            .I(N__4828));
    Odrv4 I__789 (
            .O(N__4828),
            .I(\uart_rx_inst.n729 ));
    InMux I__788 (
            .O(N__4825),
            .I(N__4822));
    LocalMux I__787 (
            .O(N__4822),
            .I(\uart_rx_inst.n1743 ));
    InMux I__786 (
            .O(N__4819),
            .I(N__4816));
    LocalMux I__785 (
            .O(N__4816),
            .I(\uart_rx_inst.n1740 ));
    InMux I__784 (
            .O(N__4813),
            .I(N__4810));
    LocalMux I__783 (
            .O(N__4810),
            .I(\uart_rx_inst.n1741 ));
    InMux I__782 (
            .O(N__4807),
            .I(N__4804));
    LocalMux I__781 (
            .O(N__4804),
            .I(\uart_rx_inst.n1747 ));
    InMux I__780 (
            .O(N__4801),
            .I(N__4798));
    LocalMux I__779 (
            .O(N__4798),
            .I(\uart_rx_inst.n1745 ));
    InMux I__778 (
            .O(N__4795),
            .I(N__4792));
    LocalMux I__777 (
            .O(N__4792),
            .I(N__4788));
    CascadeMux I__776 (
            .O(N__4791),
            .I(N__4785));
    Span4Mux_v I__775 (
            .O(N__4788),
            .I(N__4782));
    InMux I__774 (
            .O(N__4785),
            .I(N__4779));
    Odrv4 I__773 (
            .O(N__4782),
            .I(\uart_rx_inst.prescale_reg_8 ));
    LocalMux I__772 (
            .O(N__4779),
            .I(\uart_rx_inst.prescale_reg_8 ));
    InMux I__771 (
            .O(N__4774),
            .I(N__4771));
    LocalMux I__770 (
            .O(N__4771),
            .I(N__4768));
    Span4Mux_v I__769 (
            .O(N__4768),
            .I(N__4765));
    Odrv4 I__768 (
            .O(N__4765),
            .I(\uart_rx_inst.n784 ));
    InMux I__767 (
            .O(N__4762),
            .I(bfn_9_6_0_));
    CascadeMux I__766 (
            .O(N__4759),
            .I(N__4755));
    CascadeMux I__765 (
            .O(N__4758),
            .I(N__4752));
    InMux I__764 (
            .O(N__4755),
            .I(N__4749));
    InMux I__763 (
            .O(N__4752),
            .I(N__4746));
    LocalMux I__762 (
            .O(N__4749),
            .I(N__4743));
    LocalMux I__761 (
            .O(N__4746),
            .I(\uart_rx_inst.prescale_reg_9 ));
    Odrv4 I__760 (
            .O(N__4743),
            .I(\uart_rx_inst.prescale_reg_9 ));
    InMux I__759 (
            .O(N__4738),
            .I(N__4735));
    LocalMux I__758 (
            .O(N__4735),
            .I(\uart_rx_inst.n779 ));
    InMux I__757 (
            .O(N__4732),
            .I(\uart_rx_inst.n1572 ));
    InMux I__756 (
            .O(N__4729),
            .I(N__4726));
    LocalMux I__755 (
            .O(N__4726),
            .I(N__4723));
    Span4Mux_h I__754 (
            .O(N__4723),
            .I(N__4720));
    Odrv4 I__753 (
            .O(N__4720),
            .I(\uart_rx_inst.n1744 ));
    CascadeMux I__752 (
            .O(N__4717),
            .I(N__4713));
    InMux I__751 (
            .O(N__4716),
            .I(N__4710));
    InMux I__750 (
            .O(N__4713),
            .I(N__4707));
    LocalMux I__749 (
            .O(N__4710),
            .I(\uart_rx_inst.prescale_reg_10 ));
    LocalMux I__748 (
            .O(N__4707),
            .I(\uart_rx_inst.prescale_reg_10 ));
    InMux I__747 (
            .O(N__4702),
            .I(N__4699));
    LocalMux I__746 (
            .O(N__4699),
            .I(\uart_rx_inst.n774 ));
    InMux I__745 (
            .O(N__4696),
            .I(\uart_rx_inst.n1573 ));
    CascadeMux I__744 (
            .O(N__4693),
            .I(N__4690));
    InMux I__743 (
            .O(N__4690),
            .I(N__4686));
    InMux I__742 (
            .O(N__4689),
            .I(N__4683));
    LocalMux I__741 (
            .O(N__4686),
            .I(\uart_rx_inst.prescale_reg_11 ));
    LocalMux I__740 (
            .O(N__4683),
            .I(\uart_rx_inst.prescale_reg_11 ));
    InMux I__739 (
            .O(N__4678),
            .I(N__4675));
    LocalMux I__738 (
            .O(N__4675),
            .I(\uart_rx_inst.n769 ));
    InMux I__737 (
            .O(N__4672),
            .I(\uart_rx_inst.n1574 ));
    InMux I__736 (
            .O(N__4669),
            .I(N__4665));
    InMux I__735 (
            .O(N__4668),
            .I(N__4662));
    LocalMux I__734 (
            .O(N__4665),
            .I(\uart_rx_inst.prescale_reg_12 ));
    LocalMux I__733 (
            .O(N__4662),
            .I(\uart_rx_inst.prescale_reg_12 ));
    CascadeMux I__732 (
            .O(N__4657),
            .I(N__4654));
    InMux I__731 (
            .O(N__4654),
            .I(N__4651));
    LocalMux I__730 (
            .O(N__4651),
            .I(\uart_rx_inst.n764 ));
    InMux I__729 (
            .O(N__4648),
            .I(\uart_rx_inst.n1575 ));
    CascadeMux I__728 (
            .O(N__4645),
            .I(N__4642));
    InMux I__727 (
            .O(N__4642),
            .I(N__4638));
    InMux I__726 (
            .O(N__4641),
            .I(N__4635));
    LocalMux I__725 (
            .O(N__4638),
            .I(\uart_rx_inst.prescale_reg_13 ));
    LocalMux I__724 (
            .O(N__4635),
            .I(\uart_rx_inst.prescale_reg_13 ));
    InMux I__723 (
            .O(N__4630),
            .I(N__4627));
    LocalMux I__722 (
            .O(N__4627),
            .I(\uart_rx_inst.n759 ));
    InMux I__721 (
            .O(N__4624),
            .I(\uart_rx_inst.n1576 ));
    InMux I__720 (
            .O(N__4621),
            .I(N__4618));
    LocalMux I__719 (
            .O(N__4618),
            .I(N__4614));
    InMux I__718 (
            .O(N__4617),
            .I(N__4611));
    Odrv4 I__717 (
            .O(N__4614),
            .I(\uart_rx_inst.prescale_reg_14 ));
    LocalMux I__716 (
            .O(N__4611),
            .I(\uart_rx_inst.prescale_reg_14 ));
    InMux I__715 (
            .O(N__4606),
            .I(N__4603));
    LocalMux I__714 (
            .O(N__4603),
            .I(\uart_rx_inst.n754 ));
    InMux I__713 (
            .O(N__4600),
            .I(\uart_rx_inst.n1577 ));
    InMux I__712 (
            .O(N__4597),
            .I(N__4591));
    InMux I__711 (
            .O(N__4596),
            .I(N__4586));
    InMux I__710 (
            .O(N__4595),
            .I(N__4586));
    InMux I__709 (
            .O(N__4594),
            .I(N__4583));
    LocalMux I__708 (
            .O(N__4591),
            .I(\uart_rx_inst.n509 ));
    LocalMux I__707 (
            .O(N__4586),
            .I(\uart_rx_inst.n509 ));
    LocalMux I__706 (
            .O(N__4583),
            .I(\uart_rx_inst.n509 ));
    CascadeMux I__705 (
            .O(N__4576),
            .I(N__4572));
    InMux I__704 (
            .O(N__4575),
            .I(N__4569));
    InMux I__703 (
            .O(N__4572),
            .I(N__4566));
    LocalMux I__702 (
            .O(N__4569),
            .I(N__4563));
    LocalMux I__701 (
            .O(N__4566),
            .I(\uart_rx_inst.prescale_reg_0 ));
    Odrv4 I__700 (
            .O(N__4563),
            .I(\uart_rx_inst.prescale_reg_0 ));
    InMux I__699 (
            .O(N__4558),
            .I(bfn_9_5_0_));
    CEMux I__698 (
            .O(N__4555),
            .I(N__4552));
    LocalMux I__697 (
            .O(N__4552),
            .I(N__4549));
    Span4Mux_v I__696 (
            .O(N__4549),
            .I(N__4546));
    Odrv4 I__695 (
            .O(N__4546),
            .I(\uart_rx_inst.n1648 ));
    SRMux I__694 (
            .O(N__4543),
            .I(N__4540));
    LocalMux I__693 (
            .O(N__4540),
            .I(N__4537));
    Span4Mux_s3_h I__692 (
            .O(N__4537),
            .I(N__4534));
    Span4Mux_v I__691 (
            .O(N__4534),
            .I(N__4531));
    Odrv4 I__690 (
            .O(N__4531),
            .I(\uart_rx_inst.n1141 ));
    InMux I__689 (
            .O(N__4528),
            .I(N__4525));
    LocalMux I__688 (
            .O(N__4525),
            .I(N__4522));
    Span4Mux_s3_h I__687 (
            .O(N__4522),
            .I(N__4518));
    InMux I__686 (
            .O(N__4521),
            .I(N__4515));
    Odrv4 I__685 (
            .O(N__4518),
            .I(\uart_rx_inst.prescale_reg_1 ));
    LocalMux I__684 (
            .O(N__4515),
            .I(\uart_rx_inst.prescale_reg_1 ));
    InMux I__683 (
            .O(N__4510),
            .I(N__4507));
    LocalMux I__682 (
            .O(N__4507),
            .I(N__4504));
    Odrv4 I__681 (
            .O(N__4504),
            .I(\uart_rx_inst.n819 ));
    InMux I__680 (
            .O(N__4501),
            .I(\uart_rx_inst.n1564 ));
    CascadeMux I__679 (
            .O(N__4498),
            .I(N__4495));
    InMux I__678 (
            .O(N__4495),
            .I(N__4492));
    LocalMux I__677 (
            .O(N__4492),
            .I(N__4489));
    Span4Mux_h I__676 (
            .O(N__4489),
            .I(N__4485));
    InMux I__675 (
            .O(N__4488),
            .I(N__4482));
    Odrv4 I__674 (
            .O(N__4485),
            .I(\uart_rx_inst.prescale_reg_2 ));
    LocalMux I__673 (
            .O(N__4482),
            .I(\uart_rx_inst.prescale_reg_2 ));
    InMux I__672 (
            .O(N__4477),
            .I(N__4474));
    LocalMux I__671 (
            .O(N__4474),
            .I(N__4471));
    Span4Mux_v I__670 (
            .O(N__4471),
            .I(N__4468));
    Odrv4 I__669 (
            .O(N__4468),
            .I(\uart_rx_inst.n814 ));
    InMux I__668 (
            .O(N__4465),
            .I(\uart_rx_inst.n1565 ));
    InMux I__667 (
            .O(N__4462),
            .I(N__4458));
    InMux I__666 (
            .O(N__4461),
            .I(N__4455));
    LocalMux I__665 (
            .O(N__4458),
            .I(\uart_rx_inst.prescale_reg_3 ));
    LocalMux I__664 (
            .O(N__4455),
            .I(\uart_rx_inst.prescale_reg_3 ));
    InMux I__663 (
            .O(N__4450),
            .I(N__4447));
    LocalMux I__662 (
            .O(N__4447),
            .I(\uart_rx_inst.n809 ));
    InMux I__661 (
            .O(N__4444),
            .I(\uart_rx_inst.n1566 ));
    CascadeMux I__660 (
            .O(N__4441),
            .I(N__4438));
    InMux I__659 (
            .O(N__4438),
            .I(N__4435));
    LocalMux I__658 (
            .O(N__4435),
            .I(N__4431));
    InMux I__657 (
            .O(N__4434),
            .I(N__4428));
    Odrv4 I__656 (
            .O(N__4431),
            .I(\uart_rx_inst.prescale_reg_4 ));
    LocalMux I__655 (
            .O(N__4428),
            .I(\uart_rx_inst.prescale_reg_4 ));
    InMux I__654 (
            .O(N__4423),
            .I(N__4420));
    LocalMux I__653 (
            .O(N__4420),
            .I(N__4417));
    Odrv4 I__652 (
            .O(N__4417),
            .I(\uart_rx_inst.n804 ));
    InMux I__651 (
            .O(N__4414),
            .I(\uart_rx_inst.n1567 ));
    InMux I__650 (
            .O(N__4411),
            .I(N__4408));
    LocalMux I__649 (
            .O(N__4408),
            .I(N__4405));
    Span4Mux_h I__648 (
            .O(N__4405),
            .I(N__4402));
    Odrv4 I__647 (
            .O(N__4402),
            .I(\uart_rx_inst.n1756 ));
    InMux I__646 (
            .O(N__4399),
            .I(N__4396));
    LocalMux I__645 (
            .O(N__4396),
            .I(N__4392));
    InMux I__644 (
            .O(N__4395),
            .I(N__4389));
    Odrv4 I__643 (
            .O(N__4392),
            .I(\uart_rx_inst.prescale_reg_5 ));
    LocalMux I__642 (
            .O(N__4389),
            .I(\uart_rx_inst.prescale_reg_5 ));
    InMux I__641 (
            .O(N__4384),
            .I(N__4381));
    LocalMux I__640 (
            .O(N__4381),
            .I(N__4378));
    Odrv4 I__639 (
            .O(N__4378),
            .I(\uart_rx_inst.n799 ));
    InMux I__638 (
            .O(N__4375),
            .I(\uart_rx_inst.n1568 ));
    CascadeMux I__637 (
            .O(N__4372),
            .I(N__4369));
    InMux I__636 (
            .O(N__4369),
            .I(N__4365));
    InMux I__635 (
            .O(N__4368),
            .I(N__4362));
    LocalMux I__634 (
            .O(N__4365),
            .I(\uart_rx_inst.prescale_reg_6 ));
    LocalMux I__633 (
            .O(N__4362),
            .I(\uart_rx_inst.prescale_reg_6 ));
    InMux I__632 (
            .O(N__4357),
            .I(N__4354));
    LocalMux I__631 (
            .O(N__4354),
            .I(\uart_rx_inst.n794 ));
    InMux I__630 (
            .O(N__4351),
            .I(\uart_rx_inst.n1569 ));
    InMux I__629 (
            .O(N__4348),
            .I(N__4344));
    InMux I__628 (
            .O(N__4347),
            .I(N__4341));
    LocalMux I__627 (
            .O(N__4344),
            .I(\uart_rx_inst.prescale_reg_7 ));
    LocalMux I__626 (
            .O(N__4341),
            .I(\uart_rx_inst.prescale_reg_7 ));
    InMux I__625 (
            .O(N__4336),
            .I(N__4333));
    LocalMux I__624 (
            .O(N__4333),
            .I(\uart_rx_inst.n789 ));
    InMux I__623 (
            .O(N__4330),
            .I(\uart_rx_inst.n1570 ));
    CascadeMux I__622 (
            .O(N__4327),
            .I(\uart_tx_inst.n880_cascade_ ));
    CascadeMux I__621 (
            .O(N__4324),
            .I(\uart_tx_inst.n895_cascade_ ));
    CascadeMux I__620 (
            .O(N__4321),
            .I(\uart_tx_inst.n900_cascade_ ));
    InMux I__619 (
            .O(N__4318),
            .I(N__4315));
    LocalMux I__618 (
            .O(N__4315),
            .I(\uart_tx_inst.n925 ));
    InMux I__617 (
            .O(N__4312),
            .I(N__4309));
    LocalMux I__616 (
            .O(N__4309),
            .I(\uart_tx_inst.n935 ));
    CascadeMux I__615 (
            .O(N__4306),
            .I(\uart_tx_inst.n920_cascade_ ));
    CascadeMux I__614 (
            .O(N__4303),
            .I(\uart_tx_inst.n930_cascade_ ));
    InMux I__613 (
            .O(N__4300),
            .I(N__4297));
    LocalMux I__612 (
            .O(N__4297),
            .I(\uart_tx_inst.n31_adj_199 ));
    InMux I__611 (
            .O(N__4294),
            .I(N__4291));
    LocalMux I__610 (
            .O(N__4291),
            .I(\uart_tx_inst.n915 ));
    CascadeMux I__609 (
            .O(N__4288),
            .I(\uart_tx_inst.n875_cascade_ ));
    SRMux I__608 (
            .O(N__4285),
            .I(N__4282));
    LocalMux I__607 (
            .O(N__4282),
            .I(N__4279));
    Span4Mux_h I__606 (
            .O(N__4279),
            .I(N__4276));
    Odrv4 I__605 (
            .O(N__4276),
            .I(n1167));
    InMux I__604 (
            .O(N__4273),
            .I(N__4265));
    InMux I__603 (
            .O(N__4272),
            .I(N__4265));
    InMux I__602 (
            .O(N__4271),
            .I(N__4258));
    CascadeMux I__601 (
            .O(N__4270),
            .I(N__4254));
    LocalMux I__600 (
            .O(N__4265),
            .I(N__4250));
    InMux I__599 (
            .O(N__4264),
            .I(N__4247));
    InMux I__598 (
            .O(N__4263),
            .I(N__4242));
    InMux I__597 (
            .O(N__4262),
            .I(N__4242));
    InMux I__596 (
            .O(N__4261),
            .I(N__4239));
    LocalMux I__595 (
            .O(N__4258),
            .I(N__4236));
    InMux I__594 (
            .O(N__4257),
            .I(N__4229));
    InMux I__593 (
            .O(N__4254),
            .I(N__4229));
    InMux I__592 (
            .O(N__4253),
            .I(N__4229));
    Span4Mux_v I__591 (
            .O(N__4250),
            .I(N__4226));
    LocalMux I__590 (
            .O(N__4247),
            .I(bit_cnt_0));
    LocalMux I__589 (
            .O(N__4242),
            .I(bit_cnt_0));
    LocalMux I__588 (
            .O(N__4239),
            .I(bit_cnt_0));
    Odrv4 I__587 (
            .O(N__4236),
            .I(bit_cnt_0));
    LocalMux I__586 (
            .O(N__4229),
            .I(bit_cnt_0));
    Odrv4 I__585 (
            .O(N__4226),
            .I(bit_cnt_0));
    InMux I__584 (
            .O(N__4213),
            .I(N__4207));
    InMux I__583 (
            .O(N__4212),
            .I(N__4201));
    InMux I__582 (
            .O(N__4211),
            .I(N__4201));
    InMux I__581 (
            .O(N__4210),
            .I(N__4198));
    LocalMux I__580 (
            .O(N__4207),
            .I(N__4195));
    InMux I__579 (
            .O(N__4206),
            .I(N__4192));
    LocalMux I__578 (
            .O(N__4201),
            .I(N__4189));
    LocalMux I__577 (
            .O(N__4198),
            .I(\uart_rx_inst.n677 ));
    Odrv4 I__576 (
            .O(N__4195),
            .I(\uart_rx_inst.n677 ));
    LocalMux I__575 (
            .O(N__4192),
            .I(\uart_rx_inst.n677 ));
    Odrv4 I__574 (
            .O(N__4189),
            .I(\uart_rx_inst.n677 ));
    CascadeMux I__573 (
            .O(N__4180),
            .I(N__4177));
    InMux I__572 (
            .O(N__4177),
            .I(N__4174));
    LocalMux I__571 (
            .O(N__4174),
            .I(N__4170));
    InMux I__570 (
            .O(N__4173),
            .I(N__4167));
    Odrv4 I__569 (
            .O(N__4170),
            .I(\uart_rx_inst.output_axis_tvalid_N_172 ));
    LocalMux I__568 (
            .O(N__4167),
            .I(\uart_rx_inst.output_axis_tvalid_N_172 ));
    InMux I__567 (
            .O(N__4162),
            .I(N__4156));
    InMux I__566 (
            .O(N__4161),
            .I(N__4149));
    InMux I__565 (
            .O(N__4160),
            .I(N__4149));
    InMux I__564 (
            .O(N__4159),
            .I(N__4149));
    LocalMux I__563 (
            .O(N__4156),
            .I(\uart_rx_inst.output_axis_tvalid_N_173 ));
    LocalMux I__562 (
            .O(N__4149),
            .I(\uart_rx_inst.output_axis_tvalid_N_173 ));
    CascadeMux I__561 (
            .O(N__4144),
            .I(n695_cascade_));
    InMux I__560 (
            .O(N__4141),
            .I(N__4138));
    LocalMux I__559 (
            .O(N__4138),
            .I(n695));
    InMux I__558 (
            .O(N__4135),
            .I(N__4131));
    InMux I__557 (
            .O(N__4134),
            .I(N__4128));
    LocalMux I__556 (
            .O(N__4131),
            .I(N__4120));
    LocalMux I__555 (
            .O(N__4128),
            .I(N__4120));
    InMux I__554 (
            .O(N__4127),
            .I(N__4117));
    InMux I__553 (
            .O(N__4126),
            .I(N__4114));
    InMux I__552 (
            .O(N__4125),
            .I(N__4111));
    Span4Mux_v I__551 (
            .O(N__4120),
            .I(N__4104));
    LocalMux I__550 (
            .O(N__4117),
            .I(N__4104));
    LocalMux I__549 (
            .O(N__4114),
            .I(N__4104));
    LocalMux I__548 (
            .O(N__4111),
            .I(output_axis_tvalid_N_175));
    Odrv4 I__547 (
            .O(N__4104),
            .I(output_axis_tvalid_N_175));
    InMux I__546 (
            .O(N__4099),
            .I(N__4095));
    InMux I__545 (
            .O(N__4098),
            .I(N__4092));
    LocalMux I__544 (
            .O(N__4095),
            .I(N__4086));
    LocalMux I__543 (
            .O(N__4092),
            .I(N__4086));
    InMux I__542 (
            .O(N__4091),
            .I(N__4083));
    Span12Mux_s4_v I__541 (
            .O(N__4086),
            .I(N__4080));
    LocalMux I__540 (
            .O(N__4083),
            .I(n680));
    Odrv12 I__539 (
            .O(N__4080),
            .I(n680));
    InMux I__538 (
            .O(N__4075),
            .I(N__4071));
    InMux I__537 (
            .O(N__4074),
            .I(N__4068));
    LocalMux I__536 (
            .O(N__4071),
            .I(N__4065));
    LocalMux I__535 (
            .O(N__4068),
            .I(N__4062));
    Odrv4 I__534 (
            .O(N__4065),
            .I(data_reg_0));
    Odrv4 I__533 (
            .O(N__4062),
            .I(data_reg_0));
    IoInMux I__532 (
            .O(N__4057),
            .I(N__4054));
    LocalMux I__531 (
            .O(N__4054),
            .I(N__4051));
    Span4Mux_s3_v I__530 (
            .O(N__4051),
            .I(N__4048));
    Odrv4 I__529 (
            .O(N__4048),
            .I(output_axis_tdata_c_0));
    InMux I__528 (
            .O(N__4045),
            .I(N__4042));
    LocalMux I__527 (
            .O(N__4042),
            .I(N__4039));
    Span4Mux_v I__526 (
            .O(N__4039),
            .I(N__4036));
    Odrv4 I__525 (
            .O(N__4036),
            .I(rxd_c));
    CascadeMux I__524 (
            .O(N__4033),
            .I(\uart_tx_inst.n910_cascade_ ));
    CascadeMux I__523 (
            .O(N__4030),
            .I(N__4024));
    InMux I__522 (
            .O(N__4029),
            .I(N__4019));
    InMux I__521 (
            .O(N__4028),
            .I(N__4019));
    InMux I__520 (
            .O(N__4027),
            .I(N__4016));
    InMux I__519 (
            .O(N__4024),
            .I(N__4013));
    LocalMux I__518 (
            .O(N__4019),
            .I(\uart_rx_inst.output_axis_tvalid_N_174 ));
    LocalMux I__517 (
            .O(N__4016),
            .I(\uart_rx_inst.output_axis_tvalid_N_174 ));
    LocalMux I__516 (
            .O(N__4013),
            .I(\uart_rx_inst.output_axis_tvalid_N_174 ));
    CascadeMux I__515 (
            .O(N__4006),
            .I(n1711_cascade_));
    CascadeMux I__514 (
            .O(N__4003),
            .I(n1220_cascade_));
    InMux I__513 (
            .O(N__4000),
            .I(N__3994));
    InMux I__512 (
            .O(N__3999),
            .I(N__3989));
    InMux I__511 (
            .O(N__3998),
            .I(N__3989));
    InMux I__510 (
            .O(N__3997),
            .I(N__3986));
    LocalMux I__509 (
            .O(N__3994),
            .I(\uart_rx_inst.bit_cnt_3 ));
    LocalMux I__508 (
            .O(N__3989),
            .I(\uart_rx_inst.bit_cnt_3 ));
    LocalMux I__507 (
            .O(N__3986),
            .I(\uart_rx_inst.bit_cnt_3 ));
    CascadeMux I__506 (
            .O(N__3979),
            .I(\uart_rx_inst.output_axis_tvalid_N_172_cascade_ ));
    CascadeMux I__505 (
            .O(N__3976),
            .I(\uart_rx_inst.n232_cascade_ ));
    InMux I__504 (
            .O(N__3973),
            .I(N__3969));
    InMux I__503 (
            .O(N__3972),
            .I(N__3966));
    LocalMux I__502 (
            .O(N__3969),
            .I(N__3961));
    LocalMux I__501 (
            .O(N__3966),
            .I(N__3961));
    Span4Mux_v I__500 (
            .O(N__3961),
            .I(N__3957));
    InMux I__499 (
            .O(N__3960),
            .I(N__3954));
    Odrv4 I__498 (
            .O(N__3957),
            .I(\uart_rx_inst.n1468 ));
    LocalMux I__497 (
            .O(N__3954),
            .I(\uart_rx_inst.n1468 ));
    InMux I__496 (
            .O(N__3949),
            .I(N__3946));
    LocalMux I__495 (
            .O(N__3946),
            .I(\uart_rx_inst.n1502 ));
    InMux I__494 (
            .O(N__3943),
            .I(N__3939));
    InMux I__493 (
            .O(N__3942),
            .I(N__3936));
    LocalMux I__492 (
            .O(N__3939),
            .I(\uart_rx_inst.n235 ));
    LocalMux I__491 (
            .O(N__3936),
            .I(\uart_rx_inst.n235 ));
    CascadeMux I__490 (
            .O(N__3931),
            .I(N__3927));
    InMux I__489 (
            .O(N__3930),
            .I(N__3920));
    InMux I__488 (
            .O(N__3927),
            .I(N__3917));
    InMux I__487 (
            .O(N__3926),
            .I(N__3912));
    InMux I__486 (
            .O(N__3925),
            .I(N__3912));
    InMux I__485 (
            .O(N__3924),
            .I(N__3909));
    InMux I__484 (
            .O(N__3923),
            .I(N__3906));
    LocalMux I__483 (
            .O(N__3920),
            .I(\uart_rx_inst.bit_cnt_1 ));
    LocalMux I__482 (
            .O(N__3917),
            .I(\uart_rx_inst.bit_cnt_1 ));
    LocalMux I__481 (
            .O(N__3912),
            .I(\uart_rx_inst.bit_cnt_1 ));
    LocalMux I__480 (
            .O(N__3909),
            .I(\uart_rx_inst.bit_cnt_1 ));
    LocalMux I__479 (
            .O(N__3906),
            .I(\uart_rx_inst.bit_cnt_1 ));
    InMux I__478 (
            .O(N__3895),
            .I(N__3888));
    InMux I__477 (
            .O(N__3894),
            .I(N__3885));
    InMux I__476 (
            .O(N__3893),
            .I(N__3880));
    InMux I__475 (
            .O(N__3892),
            .I(N__3880));
    InMux I__474 (
            .O(N__3891),
            .I(N__3877));
    LocalMux I__473 (
            .O(N__3888),
            .I(\uart_rx_inst.bit_cnt_2 ));
    LocalMux I__472 (
            .O(N__3885),
            .I(\uart_rx_inst.bit_cnt_2 ));
    LocalMux I__471 (
            .O(N__3880),
            .I(\uart_rx_inst.bit_cnt_2 ));
    LocalMux I__470 (
            .O(N__3877),
            .I(\uart_rx_inst.bit_cnt_2 ));
    CEMux I__469 (
            .O(N__3868),
            .I(N__3864));
    CEMux I__468 (
            .O(N__3867),
            .I(N__3861));
    LocalMux I__467 (
            .O(N__3864),
            .I(N__3858));
    LocalMux I__466 (
            .O(N__3861),
            .I(N__3855));
    Span4Mux_h I__465 (
            .O(N__3858),
            .I(N__3851));
    Span4Mux_h I__464 (
            .O(N__3855),
            .I(N__3848));
    InMux I__463 (
            .O(N__3854),
            .I(N__3845));
    Odrv4 I__462 (
            .O(N__3851),
            .I(n705));
    Odrv4 I__461 (
            .O(N__3848),
            .I(n705));
    LocalMux I__460 (
            .O(N__3845),
            .I(n705));
    CascadeMux I__459 (
            .O(N__3838),
            .I(\uart_rx_inst.n509_cascade_ ));
    InMux I__458 (
            .O(N__3835),
            .I(N__3832));
    LocalMux I__457 (
            .O(N__3832),
            .I(\uart_rx_inst.n31 ));
    InMux I__456 (
            .O(N__3829),
            .I(N__3826));
    LocalMux I__455 (
            .O(N__3826),
            .I(\uart_rx_inst.n33 ));
    CascadeMux I__454 (
            .O(N__3823),
            .I(N__3800));
    InMux I__453 (
            .O(N__3822),
            .I(N__3796));
    InMux I__452 (
            .O(N__3821),
            .I(N__3779));
    InMux I__451 (
            .O(N__3820),
            .I(N__3779));
    InMux I__450 (
            .O(N__3819),
            .I(N__3779));
    InMux I__449 (
            .O(N__3818),
            .I(N__3779));
    InMux I__448 (
            .O(N__3817),
            .I(N__3779));
    InMux I__447 (
            .O(N__3816),
            .I(N__3779));
    InMux I__446 (
            .O(N__3815),
            .I(N__3779));
    InMux I__445 (
            .O(N__3814),
            .I(N__3779));
    InMux I__444 (
            .O(N__3813),
            .I(N__3766));
    InMux I__443 (
            .O(N__3812),
            .I(N__3766));
    InMux I__442 (
            .O(N__3811),
            .I(N__3766));
    InMux I__441 (
            .O(N__3810),
            .I(N__3766));
    InMux I__440 (
            .O(N__3809),
            .I(N__3766));
    InMux I__439 (
            .O(N__3808),
            .I(N__3766));
    InMux I__438 (
            .O(N__3807),
            .I(N__3761));
    InMux I__437 (
            .O(N__3806),
            .I(N__3761));
    InMux I__436 (
            .O(N__3805),
            .I(N__3750));
    InMux I__435 (
            .O(N__3804),
            .I(N__3750));
    InMux I__434 (
            .O(N__3803),
            .I(N__3750));
    InMux I__433 (
            .O(N__3800),
            .I(N__3750));
    InMux I__432 (
            .O(N__3799),
            .I(N__3750));
    LocalMux I__431 (
            .O(N__3796),
            .I(\uart_rx_inst.n1479 ));
    LocalMux I__430 (
            .O(N__3779),
            .I(\uart_rx_inst.n1479 ));
    LocalMux I__429 (
            .O(N__3766),
            .I(\uart_rx_inst.n1479 ));
    LocalMux I__428 (
            .O(N__3761),
            .I(\uart_rx_inst.n1479 ));
    LocalMux I__427 (
            .O(N__3750),
            .I(\uart_rx_inst.n1479 ));
    CEMux I__426 (
            .O(N__3739),
            .I(N__3735));
    CEMux I__425 (
            .O(N__3738),
            .I(N__3730));
    LocalMux I__424 (
            .O(N__3735),
            .I(N__3727));
    CEMux I__423 (
            .O(N__3734),
            .I(N__3724));
    CEMux I__422 (
            .O(N__3733),
            .I(N__3721));
    LocalMux I__421 (
            .O(N__3730),
            .I(\uart_rx_inst.n1045 ));
    Odrv4 I__420 (
            .O(N__3727),
            .I(\uart_rx_inst.n1045 ));
    LocalMux I__419 (
            .O(N__3724),
            .I(\uart_rx_inst.n1045 ));
    LocalMux I__418 (
            .O(N__3721),
            .I(\uart_rx_inst.n1045 ));
    CascadeMux I__417 (
            .O(N__3712),
            .I(\uart_rx_inst.n30_cascade_ ));
    CascadeMux I__416 (
            .O(N__3709),
            .I(\uart_rx_inst.n32_cascade_ ));
    InMux I__415 (
            .O(N__3706),
            .I(N__3703));
    LocalMux I__414 (
            .O(N__3703),
            .I(\uart_rx_inst.n34 ));
    CascadeMux I__413 (
            .O(N__3700),
            .I(output_axis_tvalid_N_175_cascade_));
    CascadeMux I__412 (
            .O(N__3697),
            .I(N__3691));
    CascadeMux I__411 (
            .O(N__3696),
            .I(N__3686));
    CascadeMux I__410 (
            .O(N__3695),
            .I(N__3683));
    InMux I__409 (
            .O(N__3694),
            .I(N__3675));
    InMux I__408 (
            .O(N__3691),
            .I(N__3675));
    InMux I__407 (
            .O(N__3690),
            .I(N__3675));
    InMux I__406 (
            .O(N__3689),
            .I(N__3666));
    InMux I__405 (
            .O(N__3686),
            .I(N__3666));
    InMux I__404 (
            .O(N__3683),
            .I(N__3666));
    InMux I__403 (
            .O(N__3682),
            .I(N__3666));
    LocalMux I__402 (
            .O(N__3675),
            .I(bit_cnt_2));
    LocalMux I__401 (
            .O(N__3666),
            .I(bit_cnt_2));
    InMux I__400 (
            .O(N__3661),
            .I(N__3649));
    InMux I__399 (
            .O(N__3660),
            .I(N__3649));
    InMux I__398 (
            .O(N__3659),
            .I(N__3649));
    InMux I__397 (
            .O(N__3658),
            .I(N__3642));
    InMux I__396 (
            .O(N__3657),
            .I(N__3642));
    InMux I__395 (
            .O(N__3656),
            .I(N__3642));
    LocalMux I__394 (
            .O(N__3649),
            .I(\uart_tx_inst.bit_cnt_3 ));
    LocalMux I__393 (
            .O(N__3642),
            .I(\uart_tx_inst.bit_cnt_3 ));
    CascadeMux I__392 (
            .O(N__3637),
            .I(\uart_tx_inst.n1723_cascade_ ));
    SRMux I__391 (
            .O(N__3634),
            .I(N__3631));
    LocalMux I__390 (
            .O(N__3631),
            .I(N__3628));
    Odrv4 I__389 (
            .O(N__3628),
            .I(\uart_rx_inst.n681 ));
    InMux I__388 (
            .O(N__3625),
            .I(N__3622));
    LocalMux I__387 (
            .O(N__3622),
            .I(\uart_tx_inst.n13 ));
    InMux I__386 (
            .O(N__3619),
            .I(N__3616));
    LocalMux I__385 (
            .O(N__3616),
            .I(N__3613));
    Span4Mux_h I__384 (
            .O(N__3613),
            .I(N__3610));
    Odrv4 I__383 (
            .O(N__3610),
            .I(output_axis_tready_c));
    IoInMux I__382 (
            .O(N__3607),
            .I(N__3604));
    LocalMux I__381 (
            .O(N__3604),
            .I(N__3601));
    Span4Mux_s3_v I__380 (
            .O(N__3601),
            .I(N__3596));
    InMux I__379 (
            .O(N__3600),
            .I(N__3593));
    InMux I__378 (
            .O(N__3599),
            .I(N__3590));
    Odrv4 I__377 (
            .O(N__3596),
            .I(output_axis_tvalid_c));
    LocalMux I__376 (
            .O(N__3593),
            .I(output_axis_tvalid_c));
    LocalMux I__375 (
            .O(N__3590),
            .I(output_axis_tvalid_c));
    InMux I__374 (
            .O(N__3583),
            .I(N__3579));
    InMux I__373 (
            .O(N__3582),
            .I(N__3576));
    LocalMux I__372 (
            .O(N__3579),
            .I(N__3573));
    LocalMux I__371 (
            .O(N__3576),
            .I(n1471));
    Odrv4 I__370 (
            .O(N__3573),
            .I(n1471));
    CascadeMux I__369 (
            .O(N__3568),
            .I(\uart_tx_inst.n485_cascade_ ));
    CascadeMux I__368 (
            .O(N__3565),
            .I(\uart_tx_inst.n30_adj_196_cascade_ ));
    CascadeMux I__367 (
            .O(N__3562),
            .I(\uart_tx_inst.n34_cascade_ ));
    CascadeMux I__366 (
            .O(N__3559),
            .I(\uart_tx_inst.n189_cascade_ ));
    InMux I__365 (
            .O(N__3556),
            .I(N__3552));
    CascadeMux I__364 (
            .O(N__3555),
            .I(N__3545));
    LocalMux I__363 (
            .O(N__3552),
            .I(N__3542));
    InMux I__362 (
            .O(N__3551),
            .I(N__3539));
    InMux I__361 (
            .O(N__3550),
            .I(N__3536));
    InMux I__360 (
            .O(N__3549),
            .I(N__3533));
    InMux I__359 (
            .O(N__3548),
            .I(N__3528));
    InMux I__358 (
            .O(N__3545),
            .I(N__3528));
    Odrv4 I__357 (
            .O(N__3542),
            .I(\uart_tx_inst.bit_cnt_0 ));
    LocalMux I__356 (
            .O(N__3539),
            .I(\uart_tx_inst.bit_cnt_0 ));
    LocalMux I__355 (
            .O(N__3536),
            .I(\uart_tx_inst.bit_cnt_0 ));
    LocalMux I__354 (
            .O(N__3533),
            .I(\uart_tx_inst.bit_cnt_0 ));
    LocalMux I__353 (
            .O(N__3528),
            .I(\uart_tx_inst.bit_cnt_0 ));
    CascadeMux I__352 (
            .O(N__3517),
            .I(N__3514));
    InMux I__351 (
            .O(N__3514),
            .I(N__3511));
    LocalMux I__350 (
            .O(N__3511),
            .I(\uart_tx_inst.n7_adj_195 ));
    InMux I__349 (
            .O(N__3508),
            .I(N__3499));
    InMux I__348 (
            .O(N__3507),
            .I(N__3494));
    InMux I__347 (
            .O(N__3506),
            .I(N__3494));
    InMux I__346 (
            .O(N__3505),
            .I(N__3485));
    InMux I__345 (
            .O(N__3504),
            .I(N__3485));
    InMux I__344 (
            .O(N__3503),
            .I(N__3485));
    InMux I__343 (
            .O(N__3502),
            .I(N__3485));
    LocalMux I__342 (
            .O(N__3499),
            .I(\uart_tx_inst.bit_cnt_1 ));
    LocalMux I__341 (
            .O(N__3494),
            .I(\uart_tx_inst.bit_cnt_1 ));
    LocalMux I__340 (
            .O(N__3485),
            .I(\uart_tx_inst.bit_cnt_1 ));
    CascadeMux I__339 (
            .O(N__3478),
            .I(\uart_tx_inst.n15_cascade_ ));
    CascadeMux I__338 (
            .O(N__3475),
            .I(n1167_cascade_));
    InMux I__337 (
            .O(N__3472),
            .I(N__3469));
    LocalMux I__336 (
            .O(N__3469),
            .I(n1698));
    CascadeMux I__335 (
            .O(N__3466),
            .I(\uart_rx_inst.n677_cascade_ ));
    CascadeMux I__334 (
            .O(N__3463),
            .I(\uart_rx_inst.n607_cascade_ ));
    CascadeMux I__333 (
            .O(N__3460),
            .I(\uart_rx_inst.n603_cascade_ ));
    CEMux I__332 (
            .O(N__3457),
            .I(N__3454));
    LocalMux I__331 (
            .O(N__3454),
            .I(N__3451));
    Odrv12 I__330 (
            .O(N__3451),
            .I(\uart_rx_inst.n984 ));
    CascadeMux I__329 (
            .O(N__3448),
            .I(n705_cascade_));
    CascadeMux I__328 (
            .O(N__3445),
            .I(\uart_tx_inst.n7_cascade_ ));
    SRMux I__327 (
            .O(N__3442),
            .I(N__3439));
    LocalMux I__326 (
            .O(N__3439),
            .I(N__3436));
    Span4Mux_s0_v I__325 (
            .O(N__3436),
            .I(N__3432));
    InMux I__324 (
            .O(N__3435),
            .I(N__3429));
    Odrv4 I__323 (
            .O(N__3432),
            .I(n1165));
    LocalMux I__322 (
            .O(N__3429),
            .I(n1165));
    CascadeMux I__321 (
            .O(N__3424),
            .I(N__3421));
    InMux I__320 (
            .O(N__3421),
            .I(N__3418));
    LocalMux I__319 (
            .O(N__3418),
            .I(n4));
    InMux I__318 (
            .O(N__3415),
            .I(N__3412));
    LocalMux I__317 (
            .O(N__3412),
            .I(\uart_tx_inst.n613 ));
    CEMux I__316 (
            .O(N__3409),
            .I(N__3406));
    LocalMux I__315 (
            .O(N__3406),
            .I(N__3402));
    CEMux I__314 (
            .O(N__3405),
            .I(N__3399));
    Span4Mux_v I__313 (
            .O(N__3402),
            .I(N__3394));
    LocalMux I__312 (
            .O(N__3399),
            .I(N__3394));
    Span4Mux_s1_v I__311 (
            .O(N__3394),
            .I(N__3390));
    InMux I__310 (
            .O(N__3393),
            .I(N__3387));
    Odrv4 I__309 (
            .O(N__3390),
            .I(n707));
    LocalMux I__308 (
            .O(N__3387),
            .I(n707));
    IoInMux I__307 (
            .O(N__3382),
            .I(N__3379));
    LocalMux I__306 (
            .O(N__3379),
            .I(N__3376));
    IoSpan4Mux I__305 (
            .O(N__3376),
            .I(N__3373));
    Span4Mux_s0_v I__304 (
            .O(N__3373),
            .I(N__3370));
    Odrv4 I__303 (
            .O(N__3370),
            .I(rx_overrun_error_c));
    CEMux I__302 (
            .O(N__3367),
            .I(N__3364));
    LocalMux I__301 (
            .O(N__3364),
            .I(N__3361));
    Odrv4 I__300 (
            .O(N__3361),
            .I(\uart_tx_inst.n721 ));
    IoInMux I__299 (
            .O(N__3358),
            .I(N__3355));
    LocalMux I__298 (
            .O(N__3355),
            .I(N__3352));
    Span4Mux_s1_v I__297 (
            .O(N__3352),
            .I(N__3348));
    InMux I__296 (
            .O(N__3351),
            .I(N__3345));
    Odrv4 I__295 (
            .O(N__3348),
            .I(input_axis_tready_c));
    LocalMux I__294 (
            .O(N__3345),
            .I(input_axis_tready_c));
    CEMux I__293 (
            .O(N__3340),
            .I(N__3337));
    LocalMux I__292 (
            .O(N__3337),
            .I(N__3334));
    Span4Mux_h I__291 (
            .O(N__3334),
            .I(N__3331));
    Odrv4 I__290 (
            .O(N__3331),
            .I(\uart_tx_inst.n701 ));
    SRMux I__289 (
            .O(N__3328),
            .I(N__3325));
    LocalMux I__288 (
            .O(N__3325),
            .I(\uart_tx_inst.n535 ));
    IoInMux I__287 (
            .O(N__3322),
            .I(N__3319));
    LocalMux I__286 (
            .O(N__3319),
            .I(N__3316));
    Span12Mux_s5_v I__285 (
            .O(N__3316),
            .I(N__3313));
    Odrv12 I__284 (
            .O(N__3313),
            .I(rx_busy_c));
    CascadeMux I__283 (
            .O(N__3310),
            .I(n588_cascade_));
    CascadeMux I__282 (
            .O(N__3307),
            .I(n707_cascade_));
    IoInMux I__281 (
            .O(N__3304),
            .I(N__3301));
    LocalMux I__280 (
            .O(N__3301),
            .I(tx_busy_c));
    defparam IN_MUX_bfv_12_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_5_0_));
    defparam IN_MUX_bfv_12_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_6_0_ (
            .carryinitin(\uart_tx_inst.n1589 ),
            .carryinitout(bfn_12_6_0_));
    defparam IN_MUX_bfv_11_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_2_0_));
    defparam IN_MUX_bfv_11_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_3_0_ (
            .carryinitin(\uart_tx_inst.n1553 ),
            .carryinitout(bfn_11_3_0_));
    defparam IN_MUX_bfv_11_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_4_0_ (
            .carryinitin(\uart_tx_inst.n1561 ),
            .carryinitout(bfn_11_4_0_));
    defparam IN_MUX_bfv_9_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_5_0_));
    defparam IN_MUX_bfv_9_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_6_0_ (
            .carryinitin(\uart_rx_inst.n1571 ),
            .carryinitout(bfn_9_6_0_));
    defparam IN_MUX_bfv_9_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_7_0_ (
            .carryinitin(\uart_rx_inst.n1579 ),
            .carryinitout(bfn_9_7_0_));
    defparam IN_MUX_bfv_11_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_5_0_));
    defparam IN_MUX_bfv_11_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_6_0_ (
            .carryinitin(\uart_rx_inst.n1537 ),
            .carryinitout(bfn_11_6_0_));
    defparam IN_MUX_bfv_11_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_7_0_ (
            .carryinitin(\uart_rx_inst.n1545 ),
            .carryinitout(bfn_11_7_0_));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \uart_tx_inst.busy_reg_53_LC_5_1_0 .C_ON=1'b0;
    defparam \uart_tx_inst.busy_reg_53_LC_5_1_0 .SEQ_MODE=4'b1000;
    defparam \uart_tx_inst.busy_reg_53_LC_5_1_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_tx_inst.busy_reg_53_LC_5_1_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7660),
            .lcout(tx_busy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7365),
            .ce(N__3367),
            .sr(N__7188));
    defparam \uart_tx_inst.i1_2_lut_3_lut_LC_6_1_0 .C_ON=1'b0;
    defparam \uart_tx_inst.i1_2_lut_3_lut_LC_6_1_0 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.i1_2_lut_3_lut_LC_6_1_0 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \uart_tx_inst.i1_2_lut_3_lut_LC_6_1_0  (
            .in0(N__7185),
            .in1(N__7485),
            .in2(_gnd_net_),
            .in3(N__6708),
            .lcout(\uart_tx_inst.n701 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.i1_3_lut_adj_25_LC_6_1_1 .C_ON=1'b0;
    defparam \uart_tx_inst.i1_3_lut_adj_25_LC_6_1_1 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.i1_3_lut_adj_25_LC_6_1_1 .LUT_INIT=16'b1100110011011101;
    LogicCell40 \uart_tx_inst.i1_3_lut_adj_25_LC_6_1_1  (
            .in0(N__6709),
            .in1(N__7186),
            .in2(_gnd_net_),
            .in3(N__7486),
            .lcout(\uart_tx_inst.n721 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.i407_2_lut_LC_6_1_4 .C_ON=1'b0;
    defparam \uart_tx_inst.i407_2_lut_LC_6_1_4 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.i407_2_lut_LC_6_1_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \uart_tx_inst.i407_2_lut_LC_6_1_4  (
            .in0(N__7187),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6707),
            .lcout(\uart_tx_inst.n535 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.input_axis_tready_reg_49_LC_6_2_0 .C_ON=1'b0;
    defparam \uart_tx_inst.input_axis_tready_reg_49_LC_6_2_0 .SEQ_MODE=4'b1000;
    defparam \uart_tx_inst.input_axis_tready_reg_49_LC_6_2_0 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \uart_tx_inst.input_axis_tready_reg_49_LC_6_2_0  (
            .in0(N__7649),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3351),
            .lcout(input_axis_tready_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7366),
            .ce(N__3340),
            .sr(N__3328));
    defparam \uart_rx_inst.busy_reg_86_LC_6_6_6 .C_ON=1'b0;
    defparam \uart_rx_inst.busy_reg_86_LC_6_6_6 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.busy_reg_86_LC_6_6_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \uart_rx_inst.busy_reg_86_LC_6_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5291),
            .lcout(rx_busy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7354),
            .ce(N__3457),
            .sr(N__7237));
    defparam CONSTANT_ONE_LUT4_LC_6_7_2.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_6_7_2.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_6_7_2.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_6_7_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.bit_cnt__i1_LC_7_1_1 .C_ON=1'b0;
    defparam \uart_tx_inst.bit_cnt__i1_LC_7_1_1 .SEQ_MODE=4'b1000;
    defparam \uart_tx_inst.bit_cnt__i1_LC_7_1_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \uart_tx_inst.bit_cnt__i1_LC_7_1_1  (
            .in0(_gnd_net_),
            .in1(N__3556),
            .in2(_gnd_net_),
            .in3(N__3508),
            .lcout(\uart_tx_inst.bit_cnt_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7373),
            .ce(N__3405),
            .sr(N__3442));
    defparam \uart_tx_inst.i2_2_lut_4_lut_LC_7_2_0 .C_ON=1'b0;
    defparam \uart_tx_inst.i2_2_lut_4_lut_LC_7_2_0 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.i2_2_lut_4_lut_LC_7_2_0 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \uart_tx_inst.i2_2_lut_4_lut_LC_7_2_0  (
            .in0(N__3657),
            .in1(N__3503),
            .in2(N__3695),
            .in3(N__7430),
            .lcout(),
            .ltout(n588_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_LC_7_2_1.C_ON=1'b0;
    defparam i1_4_lut_LC_7_2_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_LC_7_2_1.LUT_INIT=16'b1010101010101110;
    LogicCell40 i1_4_lut_LC_7_2_1 (
            .in0(N__7161),
            .in1(N__3582),
            .in2(N__3310),
            .in3(N__6667),
            .lcout(n707),
            .ltout(n707_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.i1035_4_lut_LC_7_2_2 .C_ON=1'b0;
    defparam \uart_tx_inst.i1035_4_lut_LC_7_2_2 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.i1035_4_lut_LC_7_2_2 .LUT_INIT=16'b1111000011010000;
    LogicCell40 \uart_tx_inst.i1035_4_lut_LC_7_2_2  (
            .in0(N__7484),
            .in1(N__7162),
            .in2(N__3307),
            .in3(N__7431),
            .lcout(n1165),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.i1_2_lut_4_lut_adj_24_LC_7_2_3 .C_ON=1'b0;
    defparam \uart_tx_inst.i1_2_lut_4_lut_adj_24_LC_7_2_3 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.i1_2_lut_4_lut_adj_24_LC_7_2_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \uart_tx_inst.i1_2_lut_4_lut_adj_24_LC_7_2_3  (
            .in0(N__3502),
            .in1(N__3682),
            .in2(N__3555),
            .in3(N__3656),
            .lcout(\uart_tx_inst.n7 ),
            .ltout(\uart_tx_inst.n7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.i1343_2_lut_LC_7_2_4 .C_ON=1'b0;
    defparam \uart_tx_inst.i1343_2_lut_LC_7_2_4 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.i1343_2_lut_LC_7_2_4 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \uart_tx_inst.i1343_2_lut_LC_7_2_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3445),
            .in3(N__7645),
            .lcout(n1471),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.bit_cnt__i2_LC_7_2_5 .C_ON=1'b0;
    defparam \uart_tx_inst.bit_cnt__i2_LC_7_2_5 .SEQ_MODE=4'b1000;
    defparam \uart_tx_inst.bit_cnt__i2_LC_7_2_5 .LUT_INIT=16'b0000000011000110;
    LogicCell40 \uart_tx_inst.bit_cnt__i2_LC_7_2_5  (
            .in0(N__3393),
            .in1(N__3689),
            .in2(N__3424),
            .in3(N__3435),
            .lcout(bit_cnt_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7370),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.i1_3_lut_4_lut_LC_7_2_6 .C_ON=1'b0;
    defparam \uart_tx_inst.i1_3_lut_4_lut_LC_7_2_6 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.i1_3_lut_4_lut_LC_7_2_6 .LUT_INIT=16'b0101010101010110;
    LogicCell40 \uart_tx_inst.i1_3_lut_4_lut_LC_7_2_6  (
            .in0(N__3658),
            .in1(N__3505),
            .in2(N__3696),
            .in3(N__3548),
            .lcout(\uart_tx_inst.n613 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.i266_2_lut_LC_7_2_7 .C_ON=1'b0;
    defparam \uart_tx_inst.i266_2_lut_LC_7_2_7 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.i266_2_lut_LC_7_2_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \uart_tx_inst.i266_2_lut_LC_7_2_7  (
            .in0(N__3504),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3550),
            .lcout(n4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.bit_cnt__i3_LC_7_3_1 .C_ON=1'b0;
    defparam \uart_tx_inst.bit_cnt__i3_LC_7_3_1 .SEQ_MODE=4'b1000;
    defparam \uart_tx_inst.bit_cnt__i3_LC_7_3_1 .LUT_INIT=16'b0001000111110000;
    LogicCell40 \uart_tx_inst.bit_cnt__i3_LC_7_3_1  (
            .in0(N__7437),
            .in1(N__3415),
            .in2(N__7659),
            .in3(N__7519),
            .lcout(\uart_tx_inst.bit_cnt_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7367),
            .ce(N__3409),
            .sr(N__7231));
    defparam \uart_tx_inst.bit_cnt__i0_LC_7_3_3 .C_ON=1'b0;
    defparam \uart_tx_inst.bit_cnt__i0_LC_7_3_3 .SEQ_MODE=4'b1000;
    defparam \uart_tx_inst.bit_cnt__i0_LC_7_3_3 .LUT_INIT=16'b0011000001110100;
    LogicCell40 \uart_tx_inst.bit_cnt__i0_LC_7_3_3  (
            .in0(N__7436),
            .in1(N__7518),
            .in2(N__7658),
            .in3(N__3551),
            .lcout(\uart_tx_inst.bit_cnt_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7367),
            .ce(N__3409),
            .sr(N__7231));
    defparam \uart_rx_inst.overrun_error_reg_87_LC_7_4_0 .C_ON=1'b0;
    defparam \uart_rx_inst.overrun_error_reg_87_LC_7_4_0 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.overrun_error_reg_87_LC_7_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_rx_inst.overrun_error_reg_87_LC_7_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3600),
            .lcout(rx_overrun_error_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7362),
            .ce(),
            .sr(N__3634));
    defparam \uart_rx_inst.prescale_reg__i5_LC_7_5_1 .C_ON=1'b0;
    defparam \uart_rx_inst.prescale_reg__i5_LC_7_5_1 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.prescale_reg__i5_LC_7_5_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \uart_rx_inst.prescale_reg__i5_LC_7_5_1  (
            .in0(N__6181),
            .in1(N__3804),
            .in2(_gnd_net_),
            .in3(N__4384),
            .lcout(\uart_rx_inst.prescale_reg_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7359),
            .ce(N__3733),
            .sr(N__7239));
    defparam \uart_rx_inst.prescale_reg__i4_LC_7_5_2 .C_ON=1'b0;
    defparam \uart_rx_inst.prescale_reg__i4_LC_7_5_2 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.prescale_reg__i4_LC_7_5_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \uart_rx_inst.prescale_reg__i4_LC_7_5_2  (
            .in0(N__3803),
            .in1(N__5866),
            .in2(_gnd_net_),
            .in3(N__4423),
            .lcout(\uart_rx_inst.prescale_reg_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7359),
            .ce(N__3733),
            .sr(N__7239));
    defparam \uart_rx_inst.prescale_reg__i8_LC_7_5_3 .C_ON=1'b0;
    defparam \uart_rx_inst.prescale_reg__i8_LC_7_5_3 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.prescale_reg__i8_LC_7_5_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \uart_rx_inst.prescale_reg__i8_LC_7_5_3  (
            .in0(N__6142),
            .in1(N__3805),
            .in2(_gnd_net_),
            .in3(N__4774),
            .lcout(\uart_rx_inst.prescale_reg_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7359),
            .ce(N__3733),
            .sr(N__7239));
    defparam \uart_rx_inst.i1585_4_lut_LC_7_5_6 .C_ON=1'b0;
    defparam \uart_rx_inst.i1585_4_lut_LC_7_5_6 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i1585_4_lut_LC_7_5_6 .LUT_INIT=16'b1111110111011101;
    LogicCell40 \uart_rx_inst.i1585_4_lut_LC_7_5_6  (
            .in0(N__4596),
            .in1(N__7243),
            .in2(N__3823),
            .in3(N__3972),
            .lcout(\uart_rx_inst.n1648 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.i1011_2_lut_4_lut_LC_7_5_7 .C_ON=1'b0;
    defparam \uart_rx_inst.i1011_2_lut_4_lut_LC_7_5_7 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i1011_2_lut_4_lut_LC_7_5_7 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \uart_rx_inst.i1011_2_lut_4_lut_LC_7_5_7  (
            .in0(N__7242),
            .in1(N__3799),
            .in2(_gnd_net_),
            .in3(N__4595),
            .lcout(\uart_rx_inst.n1141 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.i1596_4_lut_4_lut_LC_7_6_3 .C_ON=1'b0;
    defparam \uart_rx_inst.i1596_4_lut_4_lut_LC_7_6_3 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i1596_4_lut_4_lut_LC_7_6_3 .LUT_INIT=16'b1111100011111111;
    LogicCell40 \uart_rx_inst.i1596_4_lut_4_lut_LC_7_6_3  (
            .in0(N__3973),
            .in1(N__3806),
            .in2(N__7263),
            .in3(N__4597),
            .lcout(\uart_rx_inst.n1045 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.i854_2_lut_LC_7_6_6 .C_ON=1'b0;
    defparam \uart_rx_inst.i854_2_lut_LC_7_6_6 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i854_2_lut_LC_7_6_6 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \uart_rx_inst.i854_2_lut_LC_7_6_6  (
            .in0(N__3807),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7236),
            .lcout(\uart_rx_inst.n984 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.prescale_reg__i2_LC_7_7_1 .C_ON=1'b0;
    defparam \uart_rx_inst.prescale_reg__i2_LC_7_7_1 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.prescale_reg__i2_LC_7_7_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \uart_rx_inst.prescale_reg__i2_LC_7_7_1  (
            .in0(N__5893),
            .in1(N__3822),
            .in2(_gnd_net_),
            .in3(N__4477),
            .lcout(\uart_rx_inst.prescale_reg_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7355),
            .ce(N__3734),
            .sr(N__7232));
    defparam \uart_rx_inst.i1568_2_lut_LC_7_7_4 .C_ON=1'b0;
    defparam \uart_rx_inst.i1568_2_lut_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i1568_2_lut_LC_7_7_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uart_rx_inst.i1568_2_lut_LC_7_7_4  (
            .in0(N__6904),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6287),
            .lcout(\uart_rx_inst.n1756 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.i1571_2_lut_LC_7_7_7 .C_ON=1'b0;
    defparam \uart_rx_inst.i1571_2_lut_LC_7_7_7 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i1571_2_lut_LC_7_7_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uart_rx_inst.i1571_2_lut_LC_7_7_7  (
            .in0(N__6288),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8002),
            .lcout(\uart_rx_inst.n1744 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_LC_7_8_0.C_ON=1'b0;
    defparam i1_3_lut_LC_7_8_0.SEQ_MODE=4'b0000;
    defparam i1_3_lut_LC_7_8_0.LUT_INIT=16'b1010101010111011;
    LogicCell40 i1_3_lut_LC_7_8_0 (
            .in0(N__7252),
            .in1(N__3472),
            .in2(_gnd_net_),
            .in3(N__4127),
            .lcout(n705),
            .ltout(n705_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.i1037_4_lut_LC_7_8_1 .C_ON=1'b0;
    defparam \uart_rx_inst.i1037_4_lut_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i1037_4_lut_LC_7_8_1 .LUT_INIT=16'b1011000011110000;
    LogicCell40 \uart_rx_inst.i1037_4_lut_LC_7_8_1  (
            .in0(N__7253),
            .in1(N__4027),
            .in2(N__3448),
            .in3(N__6311),
            .lcout(n1167),
            .ltout(n1167_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.bit_cnt__i0_LC_7_8_2 .C_ON=1'b0;
    defparam \uart_rx_inst.bit_cnt__i0_LC_7_8_2 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.bit_cnt__i0_LC_7_8_2 .LUT_INIT=16'b0000001100001100;
    LogicCell40 \uart_rx_inst.bit_cnt__i0_LC_7_8_2  (
            .in0(_gnd_net_),
            .in1(N__4257),
            .in2(N__3475),
            .in3(N__3854),
            .lcout(bit_cnt_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7352),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.i1_4_lut_4_lut_LC_7_8_3 .C_ON=1'b0;
    defparam \uart_rx_inst.i1_4_lut_4_lut_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i1_4_lut_4_lut_LC_7_8_3 .LUT_INIT=16'b0000001011001110;
    LogicCell40 \uart_rx_inst.i1_4_lut_4_lut_LC_7_8_3  (
            .in0(N__5293),
            .in1(N__4206),
            .in2(N__4270),
            .in3(N__3960),
            .lcout(n1698),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.i2_3_lut_adj_22_LC_7_8_5 .C_ON=1'b0;
    defparam \uart_rx_inst.i2_3_lut_adj_22_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i2_3_lut_adj_22_LC_7_8_5 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \uart_rx_inst.i2_3_lut_adj_22_LC_7_8_5  (
            .in0(N__4000),
            .in1(N__3894),
            .in2(_gnd_net_),
            .in3(N__3923),
            .lcout(\uart_rx_inst.n677 ),
            .ltout(\uart_rx_inst.n677_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.i1_2_lut_adj_23_LC_7_8_6 .C_ON=1'b0;
    defparam \uart_rx_inst.i1_2_lut_adj_23_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i1_2_lut_adj_23_LC_7_8_6 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \uart_rx_inst.i1_2_lut_adj_23_LC_7_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3466),
            .in3(N__4253),
            .lcout(\uart_rx_inst.output_axis_tvalid_N_174 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.i1_3_lut_4_lut_LC_7_9_0 .C_ON=1'b0;
    defparam \uart_rx_inst.i1_3_lut_4_lut_LC_7_9_0 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i1_3_lut_4_lut_LC_7_9_0 .LUT_INIT=16'b0101010101010110;
    LogicCell40 \uart_rx_inst.i1_3_lut_4_lut_LC_7_9_0  (
            .in0(N__3999),
            .in1(N__3893),
            .in2(N__3931),
            .in3(N__4263),
            .lcout(),
            .ltout(\uart_rx_inst.n607_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.bit_cnt__i3_LC_7_9_1 .C_ON=1'b0;
    defparam \uart_rx_inst.bit_cnt__i3_LC_7_9_1 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.bit_cnt__i3_LC_7_9_1 .LUT_INIT=16'b0000100001011101;
    LogicCell40 \uart_rx_inst.bit_cnt__i3_LC_7_9_1  (
            .in0(N__4029),
            .in1(N__6313),
            .in2(N__3463),
            .in3(N__5296),
            .lcout(\uart_rx_inst.bit_cnt_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7356),
            .ce(N__3867),
            .sr(N__7264));
    defparam \uart_rx_inst.i1_2_lut_LC_7_9_2 .C_ON=1'b0;
    defparam \uart_rx_inst.i1_2_lut_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i1_2_lut_LC_7_9_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uart_rx_inst.i1_2_lut_LC_7_9_2  (
            .in0(_gnd_net_),
            .in1(N__4262),
            .in2(_gnd_net_),
            .in3(N__3926),
            .lcout(),
            .ltout(\uart_rx_inst.n603_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.bit_cnt__i1_LC_7_9_3 .C_ON=1'b0;
    defparam \uart_rx_inst.bit_cnt__i1_LC_7_9_3 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.bit_cnt__i1_LC_7_9_3 .LUT_INIT=16'b0000100001011101;
    LogicCell40 \uart_rx_inst.bit_cnt__i1_LC_7_9_3  (
            .in0(N__4028),
            .in1(N__6312),
            .in2(N__3460),
            .in3(N__5295),
            .lcout(\uart_rx_inst.bit_cnt_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7356),
            .ce(N__3867),
            .sr(N__7264));
    defparam \uart_rx_inst.i209_2_lut_3_lut_LC_7_9_6 .C_ON=1'b0;
    defparam \uart_rx_inst.i209_2_lut_3_lut_LC_7_9_6 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i209_2_lut_3_lut_LC_7_9_6 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \uart_rx_inst.i209_2_lut_3_lut_LC_7_9_6  (
            .in0(N__3998),
            .in1(N__3892),
            .in2(_gnd_net_),
            .in3(N__3925),
            .lcout(\uart_rx_inst.output_axis_tvalid_N_173 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.i319_4_lut_LC_8_1_0 .C_ON=1'b0;
    defparam \uart_tx_inst.i319_4_lut_LC_8_1_0 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.i319_4_lut_LC_8_1_0 .LUT_INIT=16'b0000000010101110;
    LogicCell40 \uart_tx_inst.i319_4_lut_LC_8_1_0  (
            .in0(N__6554),
            .in1(N__3583),
            .in2(N__3517),
            .in3(N__6668),
            .lcout(\uart_tx_inst.n485 ),
            .ltout(\uart_tx_inst.n485_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.i787_3_lut_LC_8_1_1 .C_ON=1'b0;
    defparam \uart_tx_inst.i787_3_lut_LC_8_1_1 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.i787_3_lut_LC_8_1_1 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \uart_tx_inst.i787_3_lut_LC_8_1_1  (
            .in0(_gnd_net_),
            .in1(N__8803),
            .in2(N__3568),
            .in3(N__6052),
            .lcout(\uart_tx_inst.n915 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.i11_4_lut_LC_8_1_3 .C_ON=1'b0;
    defparam \uart_tx_inst.i11_4_lut_LC_8_1_3 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.i11_4_lut_LC_8_1_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \uart_tx_inst.i11_4_lut_LC_8_1_3  (
            .in0(N__5850),
            .in1(N__5754),
            .in2(N__5928),
            .in3(N__5587),
            .lcout(),
            .ltout(\uart_tx_inst.n30_adj_196_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.i15_4_lut_LC_8_1_4 .C_ON=1'b0;
    defparam \uart_tx_inst.i15_4_lut_LC_8_1_4 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.i15_4_lut_LC_8_1_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \uart_tx_inst.i15_4_lut_LC_8_1_4  (
            .in0(N__5724),
            .in1(N__5823),
            .in2(N__3565),
            .in3(N__6063),
            .lcout(),
            .ltout(\uart_tx_inst.n34_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.i18_4_lut_LC_8_1_5 .C_ON=1'b0;
    defparam \uart_tx_inst.i18_4_lut_LC_8_1_5 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.i18_4_lut_LC_8_1_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \uart_tx_inst.i18_4_lut_LC_8_1_5  (
            .in0(N__4300),
            .in1(N__6196),
            .in2(N__3562),
            .in3(N__5374),
            .lcout(input_axis_tready_N_72),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.i2_3_lut_LC_8_2_0 .C_ON=1'b0;
    defparam \uart_tx_inst.i2_3_lut_LC_8_2_0 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.i2_3_lut_LC_8_2_0 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \uart_tx_inst.i2_3_lut_LC_8_2_0  (
            .in0(N__7133),
            .in1(N__6569),
            .in2(_gnd_net_),
            .in3(N__6669),
            .lcout(\uart_tx_inst.n189 ),
            .ltout(\uart_tx_inst.n189_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.data_reg_i0_i8_LC_8_2_1 .C_ON=1'b0;
    defparam \uart_tx_inst.data_reg_i0_i8_LC_8_2_1 .SEQ_MODE=4'b1000;
    defparam \uart_tx_inst.data_reg_i0_i8_LC_8_2_1 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \uart_tx_inst.data_reg_i0_i8_LC_8_2_1  (
            .in0(N__7605),
            .in1(N__7563),
            .in2(N__3559),
            .in3(N__7483),
            .lcout(\uart_tx_inst.data_reg_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7375),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.i1_2_lut_4_lut_LC_8_2_2 .C_ON=1'b0;
    defparam \uart_tx_inst.i1_2_lut_4_lut_LC_8_2_2 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.i1_2_lut_4_lut_LC_8_2_2 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \uart_tx_inst.i1_2_lut_4_lut_LC_8_2_2  (
            .in0(N__3660),
            .in1(N__3549),
            .in2(N__3697),
            .in3(N__3507),
            .lcout(\uart_tx_inst.n7_adj_195 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.i1_4_lut_LC_8_2_3 .C_ON=1'b0;
    defparam \uart_tx_inst.i1_4_lut_LC_8_2_3 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.i1_4_lut_LC_8_2_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \uart_tx_inst.i1_4_lut_LC_8_2_3  (
            .in0(N__3506),
            .in1(N__3690),
            .in2(_gnd_net_),
            .in3(N__3659),
            .lcout(\uart_tx_inst.n15 ),
            .ltout(\uart_tx_inst.n15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.i146_3_lut_LC_8_2_4 .C_ON=1'b0;
    defparam \uart_tx_inst.i146_3_lut_LC_8_2_4 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.i146_3_lut_LC_8_2_4 .LUT_INIT=16'b0101111100001010;
    LogicCell40 \uart_tx_inst.i146_3_lut_LC_8_2_4  (
            .in0(N__7481),
            .in1(_gnd_net_),
            .in2(N__3478),
            .in3(N__7606),
            .lcout(\uart_tx_inst.n165 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.i1527_2_lut_LC_8_2_5 .C_ON=1'b0;
    defparam \uart_tx_inst.i1527_2_lut_LC_8_2_5 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.i1527_2_lut_LC_8_2_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \uart_tx_inst.i1527_2_lut_LC_8_2_5  (
            .in0(_gnd_net_),
            .in1(N__3694),
            .in2(_gnd_net_),
            .in3(N__3661),
            .lcout(),
            .ltout(\uart_tx_inst.n1723_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.i29_4_lut_LC_8_2_6 .C_ON=1'b0;
    defparam \uart_tx_inst.i29_4_lut_LC_8_2_6 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.i29_4_lut_LC_8_2_6 .LUT_INIT=16'b0100111011101110;
    LogicCell40 \uart_tx_inst.i29_4_lut_LC_8_2_6  (
            .in0(N__7482),
            .in1(N__7607),
            .in2(N__3637),
            .in3(N__7432),
            .lcout(\uart_tx_inst.n13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.i1587_2_lut_LC_8_3_0 .C_ON=1'b0;
    defparam \uart_rx_inst.i1587_2_lut_LC_8_3_0 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i1587_2_lut_LC_8_3_0 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \uart_rx_inst.i1587_2_lut_LC_8_3_0  (
            .in0(_gnd_net_),
            .in1(N__7176),
            .in2(_gnd_net_),
            .in3(N__4098),
            .lcout(\uart_rx_inst.n681 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.i1_3_lut_LC_8_3_6 .C_ON=1'b0;
    defparam \uart_tx_inst.i1_3_lut_LC_8_3_6 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.i1_3_lut_LC_8_3_6 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \uart_tx_inst.i1_3_lut_LC_8_3_6  (
            .in0(N__7177),
            .in1(N__3625),
            .in2(_gnd_net_),
            .in3(N__6721),
            .lcout(\uart_tx_inst.n719 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.output_axis_tvalid_reg_82_LC_8_4_3 .C_ON=1'b0;
    defparam \uart_rx_inst.output_axis_tvalid_reg_82_LC_8_4_3 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.output_axis_tvalid_reg_82_LC_8_4_3 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \uart_rx_inst.output_axis_tvalid_reg_82_LC_8_4_3  (
            .in0(N__3619),
            .in1(N__3599),
            .in2(_gnd_net_),
            .in3(N__4099),
            .lcout(output_axis_tvalid_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7368),
            .ce(),
            .sr(N__7163));
    defparam \uart_rx_inst.prescale_reg__i3_LC_8_5_0 .C_ON=1'b0;
    defparam \uart_rx_inst.prescale_reg__i3_LC_8_5_0 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.prescale_reg__i3_LC_8_5_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \uart_rx_inst.prescale_reg__i3_LC_8_5_0  (
            .in0(N__5878),
            .in1(N__3818),
            .in2(_gnd_net_),
            .in3(N__4450),
            .lcout(\uart_rx_inst.prescale_reg_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7363),
            .ce(N__3739),
            .sr(N__7241));
    defparam \uart_rx_inst.prescale_reg__i18_LC_8_5_1 .C_ON=1'b0;
    defparam \uart_rx_inst.prescale_reg__i18_LC_8_5_1 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.prescale_reg__i18_LC_8_5_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \uart_rx_inst.prescale_reg__i18_LC_8_5_1  (
            .in0(N__3817),
            .in1(N__6334),
            .in2(_gnd_net_),
            .in3(N__4834),
            .lcout(\uart_rx_inst.prescale_reg_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7363),
            .ce(N__3739),
            .sr(N__7241));
    defparam \uart_rx_inst.prescale_reg__i14_LC_8_5_2 .C_ON=1'b0;
    defparam \uart_rx_inst.prescale_reg__i14_LC_8_5_2 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.prescale_reg__i14_LC_8_5_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \uart_rx_inst.prescale_reg__i14_LC_8_5_2  (
            .in0(N__6397),
            .in1(N__3816),
            .in2(_gnd_net_),
            .in3(N__4606),
            .lcout(\uart_rx_inst.prescale_reg_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7363),
            .ce(N__3739),
            .sr(N__7241));
    defparam \uart_rx_inst.prescale_reg__i11_LC_8_5_3 .C_ON=1'b0;
    defparam \uart_rx_inst.prescale_reg__i11_LC_8_5_3 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.prescale_reg__i11_LC_8_5_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \uart_rx_inst.prescale_reg__i11_LC_8_5_3  (
            .in0(N__3815),
            .in1(N__6100),
            .in2(_gnd_net_),
            .in3(N__4678),
            .lcout(\uart_rx_inst.prescale_reg_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7363),
            .ce(N__3739),
            .sr(N__7241));
    defparam \uart_rx_inst.prescale_reg__i10_LC_8_5_4 .C_ON=1'b0;
    defparam \uart_rx_inst.prescale_reg__i10_LC_8_5_4 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.prescale_reg__i10_LC_8_5_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \uart_rx_inst.prescale_reg__i10_LC_8_5_4  (
            .in0(N__6115),
            .in1(N__3814),
            .in2(_gnd_net_),
            .in3(N__4702),
            .lcout(\uart_rx_inst.prescale_reg_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7363),
            .ce(N__3739),
            .sr(N__7241));
    defparam \uart_rx_inst.prescale_reg__i9_LC_8_5_5 .C_ON=1'b0;
    defparam \uart_rx_inst.prescale_reg__i9_LC_8_5_5 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.prescale_reg__i9_LC_8_5_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \uart_rx_inst.prescale_reg__i9_LC_8_5_5  (
            .in0(N__3821),
            .in1(N__6127),
            .in2(_gnd_net_),
            .in3(N__4738),
            .lcout(\uart_rx_inst.prescale_reg_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7363),
            .ce(N__3739),
            .sr(N__7241));
    defparam \uart_rx_inst.prescale_reg__i7_LC_8_5_6 .C_ON=1'b0;
    defparam \uart_rx_inst.prescale_reg__i7_LC_8_5_6 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.prescale_reg__i7_LC_8_5_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \uart_rx_inst.prescale_reg__i7_LC_8_5_6  (
            .in0(N__6154),
            .in1(N__3820),
            .in2(_gnd_net_),
            .in3(N__4336),
            .lcout(\uart_rx_inst.prescale_reg_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7363),
            .ce(N__3739),
            .sr(N__7241));
    defparam \uart_rx_inst.prescale_reg__i6_LC_8_5_7 .C_ON=1'b0;
    defparam \uart_rx_inst.prescale_reg__i6_LC_8_5_7 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.prescale_reg__i6_LC_8_5_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \uart_rx_inst.prescale_reg__i6_LC_8_5_7  (
            .in0(N__3819),
            .in1(_gnd_net_),
            .in2(N__6169),
            .in3(N__4357),
            .lcout(\uart_rx_inst.prescale_reg_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7363),
            .ce(N__3739),
            .sr(N__7241));
    defparam \uart_rx_inst.i1351_2_lut_3_lut_LC_8_6_0 .C_ON=1'b0;
    defparam \uart_rx_inst.i1351_2_lut_3_lut_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i1351_2_lut_3_lut_LC_8_6_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \uart_rx_inst.i1351_2_lut_3_lut_LC_8_6_0  (
            .in0(N__4273),
            .in1(N__4212),
            .in2(_gnd_net_),
            .in3(N__4125),
            .lcout(\uart_rx_inst.n1479 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.i11_4_lut_LC_8_6_2 .C_ON=1'b0;
    defparam \uart_rx_inst.i11_4_lut_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i11_4_lut_LC_8_6_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \uart_rx_inst.i11_4_lut_LC_8_6_2  (
            .in0(N__4848),
            .in1(N__4461),
            .in2(N__4717),
            .in3(N__4368),
            .lcout(),
            .ltout(\uart_rx_inst.n30_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.i15_4_lut_LC_8_6_3 .C_ON=1'b0;
    defparam \uart_rx_inst.i15_4_lut_LC_8_6_3 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i15_4_lut_LC_8_6_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \uart_rx_inst.i15_4_lut_LC_8_6_3  (
            .in0(N__4689),
            .in1(N__4347),
            .in2(N__3712),
            .in3(N__4617),
            .lcout(\uart_rx_inst.n34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.i13_4_lut_LC_8_6_4 .C_ON=1'b0;
    defparam \uart_rx_inst.i13_4_lut_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i13_4_lut_LC_8_6_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \uart_rx_inst.i13_4_lut_LC_8_6_4  (
            .in0(N__4575),
            .in1(N__4434),
            .in2(N__4791),
            .in3(N__4395),
            .lcout(),
            .ltout(\uart_rx_inst.n32_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.i18_4_lut_LC_8_6_5 .C_ON=1'b0;
    defparam \uart_rx_inst.i18_4_lut_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i18_4_lut_LC_8_6_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \uart_rx_inst.i18_4_lut_LC_8_6_5  (
            .in0(N__3829),
            .in1(N__3835),
            .in2(N__3709),
            .in3(N__3706),
            .lcout(output_axis_tvalid_N_175),
            .ltout(output_axis_tvalid_N_175_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.i362_3_lut_4_lut_LC_8_6_6 .C_ON=1'b0;
    defparam \uart_rx_inst.i362_3_lut_4_lut_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i362_3_lut_4_lut_LC_8_6_6 .LUT_INIT=16'b0000111100001110;
    LogicCell40 \uart_rx_inst.i362_3_lut_4_lut_LC_8_6_6  (
            .in0(N__4272),
            .in1(N__5292),
            .in2(N__3700),
            .in3(N__4211),
            .lcout(\uart_rx_inst.n509 ),
            .ltout(\uart_rx_inst.n509_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.i584_1_lut_LC_8_6_7 .C_ON=1'b0;
    defparam \uart_rx_inst.i584_1_lut_LC_8_6_7 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i584_1_lut_LC_8_6_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \uart_rx_inst.i584_1_lut_LC_8_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3838),
            .in3(_gnd_net_),
            .lcout(\uart_rx_inst.n712 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.i12_4_lut_LC_8_7_0 .C_ON=1'b0;
    defparam \uart_rx_inst.i12_4_lut_LC_8_7_0 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i12_4_lut_LC_8_7_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \uart_rx_inst.i12_4_lut_LC_8_7_0  (
            .in0(N__4962),
            .in1(N__5013),
            .in2(N__4993),
            .in3(N__4641),
            .lcout(\uart_rx_inst.n31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.prescale_reg__i13_LC_8_7_1 .C_ON=1'b0;
    defparam \uart_rx_inst.prescale_reg__i13_LC_8_7_1 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.prescale_reg__i13_LC_8_7_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \uart_rx_inst.prescale_reg__i13_LC_8_7_1  (
            .in0(N__6412),
            .in1(N__3810),
            .in2(_gnd_net_),
            .in3(N__4630),
            .lcout(\uart_rx_inst.prescale_reg_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7357),
            .ce(N__3738),
            .sr(N__7244));
    defparam \uart_rx_inst.prescale_reg__i15_LC_8_7_2 .C_ON=1'b0;
    defparam \uart_rx_inst.prescale_reg__i15_LC_8_7_2 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.prescale_reg__i15_LC_8_7_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \uart_rx_inst.prescale_reg__i15_LC_8_7_2  (
            .in0(N__3811),
            .in1(N__6382),
            .in2(_gnd_net_),
            .in3(N__5002),
            .lcout(\uart_rx_inst.prescale_reg_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7357),
            .ce(N__3738),
            .sr(N__7244));
    defparam \uart_rx_inst.prescale_reg__i17_LC_8_7_3 .C_ON=1'b0;
    defparam \uart_rx_inst.prescale_reg__i17_LC_8_7_3 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.prescale_reg__i17_LC_8_7_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \uart_rx_inst.prescale_reg__i17_LC_8_7_3  (
            .in0(N__6352),
            .in1(N__3813),
            .in2(_gnd_net_),
            .in3(N__4951),
            .lcout(\uart_rx_inst.prescale_reg_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7357),
            .ce(N__3738),
            .sr(N__7244));
    defparam \uart_rx_inst.prescale_reg__i16_LC_8_7_4 .C_ON=1'b0;
    defparam \uart_rx_inst.prescale_reg__i16_LC_8_7_4 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.prescale_reg__i16_LC_8_7_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \uart_rx_inst.prescale_reg__i16_LC_8_7_4  (
            .in0(N__3812),
            .in1(N__6367),
            .in2(_gnd_net_),
            .in3(N__4978),
            .lcout(\uart_rx_inst.prescale_reg_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7357),
            .ce(N__3738),
            .sr(N__7244));
    defparam \uart_rx_inst.prescale_reg__i1_LC_8_7_5 .C_ON=1'b0;
    defparam \uart_rx_inst.prescale_reg__i1_LC_8_7_5 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.prescale_reg__i1_LC_8_7_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \uart_rx_inst.prescale_reg__i1_LC_8_7_5  (
            .in0(_gnd_net_),
            .in1(N__3808),
            .in2(_gnd_net_),
            .in3(N__4510),
            .lcout(\uart_rx_inst.prescale_reg_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7357),
            .ce(N__3738),
            .sr(N__7244));
    defparam \uart_rx_inst.i14_4_lut_LC_8_7_6 .C_ON=1'b0;
    defparam \uart_rx_inst.i14_4_lut_LC_8_7_6 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i14_4_lut_LC_8_7_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \uart_rx_inst.i14_4_lut_LC_8_7_6  (
            .in0(N__4521),
            .in1(N__4488),
            .in2(N__4759),
            .in3(N__4668),
            .lcout(\uart_rx_inst.n33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.prescale_reg__i12_LC_8_7_7 .C_ON=1'b0;
    defparam \uart_rx_inst.prescale_reg__i12_LC_8_7_7 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.prescale_reg__i12_LC_8_7_7 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \uart_rx_inst.prescale_reg__i12_LC_8_7_7  (
            .in0(_gnd_net_),
            .in1(N__3809),
            .in2(N__4657),
            .in3(N__6085),
            .lcout(\uart_rx_inst.prescale_reg_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7357),
            .ce(N__3738),
            .sr(N__7244));
    defparam \uart_rx_inst.i1516_4_lut_LC_8_8_0 .C_ON=1'b0;
    defparam \uart_rx_inst.i1516_4_lut_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i1516_4_lut_LC_8_8_0 .LUT_INIT=16'b1111111101011100;
    LogicCell40 \uart_rx_inst.i1516_4_lut_LC_8_8_0  (
            .in0(N__3942),
            .in1(N__5271),
            .in2(N__4030),
            .in3(N__3949),
            .lcout(n1711),
            .ltout(n1711_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.i1384_3_lut_4_lut_LC_8_8_1 .C_ON=1'b0;
    defparam \uart_rx_inst.i1384_3_lut_4_lut_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i1384_3_lut_4_lut_LC_8_8_1 .LUT_INIT=16'b1111101011111000;
    LogicCell40 \uart_rx_inst.i1384_3_lut_4_lut_LC_8_8_1  (
            .in0(N__3943),
            .in1(N__4261),
            .in2(N__4006),
            .in3(N__4210),
            .lcout(n1220),
            .ltout(n1220_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.data_reg__i7_LC_8_8_2 .C_ON=1'b0;
    defparam \uart_rx_inst.data_reg__i7_LC_8_8_2 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.data_reg__i7_LC_8_8_2 .LUT_INIT=16'b1011000010000000;
    LogicCell40 \uart_rx_inst.data_reg__i7_LC_8_8_2  (
            .in0(N__5111),
            .in1(N__5355),
            .in2(N__4003),
            .in3(N__5272),
            .lcout(data_reg_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7353),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.i208_2_lut_3_lut_LC_8_8_3 .C_ON=1'b0;
    defparam \uart_rx_inst.i208_2_lut_3_lut_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i208_2_lut_3_lut_LC_8_8_3 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \uart_rx_inst.i208_2_lut_3_lut_LC_8_8_3  (
            .in0(N__3997),
            .in1(N__3891),
            .in2(_gnd_net_),
            .in3(N__3924),
            .lcout(\uart_rx_inst.output_axis_tvalid_N_172 ),
            .ltout(\uart_rx_inst.output_axis_tvalid_N_172_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.i149_3_lut_LC_8_8_4 .C_ON=1'b0;
    defparam \uart_rx_inst.i149_3_lut_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i149_3_lut_LC_8_8_4 .LUT_INIT=16'b0101000011111010;
    LogicCell40 \uart_rx_inst.i149_3_lut_LC_8_8_4  (
            .in0(N__4159),
            .in1(_gnd_net_),
            .in2(N__3979),
            .in3(N__5269),
            .lcout(\uart_rx_inst.n232 ),
            .ltout(\uart_rx_inst.n232_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.i1340_3_lut_LC_8_8_5 .C_ON=1'b0;
    defparam \uart_rx_inst.i1340_3_lut_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i1340_3_lut_LC_8_8_5 .LUT_INIT=16'b1111101011110000;
    LogicCell40 \uart_rx_inst.i1340_3_lut_LC_8_8_5  (
            .in0(N__5270),
            .in1(_gnd_net_),
            .in2(N__3976),
            .in3(N__4160),
            .lcout(\uart_rx_inst.n1468 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.i1374_2_lut_LC_8_8_6 .C_ON=1'b0;
    defparam \uart_rx_inst.i1374_2_lut_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i1374_2_lut_LC_8_8_6 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \uart_rx_inst.i1374_2_lut_LC_8_8_6  (
            .in0(N__7245),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4126),
            .lcout(\uart_rx_inst.n1502 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.i78_2_lut_LC_8_8_7 .C_ON=1'b0;
    defparam \uart_rx_inst.i78_2_lut_LC_8_8_7 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i78_2_lut_LC_8_8_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \uart_rx_inst.i78_2_lut_LC_8_8_7  (
            .in0(_gnd_net_),
            .in1(N__4173),
            .in2(_gnd_net_),
            .in3(N__4161),
            .lcout(\uart_rx_inst.n235 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.bit_cnt__i2_LC_8_9_0 .C_ON=1'b0;
    defparam \uart_rx_inst.bit_cnt__i2_LC_8_9_0 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.bit_cnt__i2_LC_8_9_0 .LUT_INIT=16'b1100110010011001;
    LogicCell40 \uart_rx_inst.bit_cnt__i2_LC_8_9_0  (
            .in0(N__4264),
            .in1(N__3895),
            .in2(_gnd_net_),
            .in3(N__3930),
            .lcout(\uart_rx_inst.bit_cnt_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7358),
            .ce(N__3868),
            .sr(N__4285));
    defparam \uart_rx_inst.i2_4_lut_LC_8_10_2 .C_ON=1'b0;
    defparam \uart_rx_inst.i2_4_lut_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i2_4_lut_LC_8_10_2 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \uart_rx_inst.i2_4_lut_LC_8_10_2  (
            .in0(N__4271),
            .in1(N__4213),
            .in2(N__4180),
            .in3(N__4162),
            .lcout(n695),
            .ltout(n695_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.i1589_2_lut_3_lut_LC_8_10_3 .C_ON=1'b0;
    defparam \uart_tx_inst.i1589_2_lut_3_lut_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.i1589_2_lut_3_lut_LC_8_10_3 .LUT_INIT=16'b1111111110101111;
    LogicCell40 \uart_tx_inst.i1589_2_lut_3_lut_LC_8_10_3  (
            .in0(N__7238),
            .in1(_gnd_net_),
            .in2(N__4144),
            .in3(N__4135),
            .lcout(n697),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.data_reg__i0_LC_8_10_6 .C_ON=1'b0;
    defparam \uart_rx_inst.data_reg__i0_LC_8_10_6 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.data_reg__i0_LC_8_10_6 .LUT_INIT=16'b1011100000000000;
    LogicCell40 \uart_rx_inst.data_reg__i0_LC_8_10_6  (
            .in0(N__4074),
            .in1(N__5365),
            .in2(N__5494),
            .in3(N__5326),
            .lcout(data_reg_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7360),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.i2_3_lut_LC_8_11_6 .C_ON=1'b0;
    defparam \uart_rx_inst.i2_3_lut_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i2_3_lut_LC_8_11_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \uart_rx_inst.i2_3_lut_LC_8_11_6  (
            .in0(N__4141),
            .in1(N__5282),
            .in2(_gnd_net_),
            .in3(N__4134),
            .lcout(n680),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_LC_8_12_4.C_ON=1'b0;
    defparam i1_2_lut_LC_8_12_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_LC_8_12_4.LUT_INIT=16'b1111111110101010;
    LogicCell40 i1_2_lut_LC_8_12_4 (
            .in0(N__7255),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4091),
            .lcout(n703),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.output_axis_tdata_reg__i1_LC_8_13_3 .C_ON=1'b0;
    defparam \uart_rx_inst.output_axis_tdata_reg__i1_LC_8_13_3 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.output_axis_tdata_reg__i1_LC_8_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_rx_inst.output_axis_tdata_reg__i1_LC_8_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4075),
            .lcout(output_axis_tdata_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7371),
            .ce(N__5418),
            .sr(N__7266));
    defparam \uart_rx_inst.rxd_reg_83_LC_8_14_4 .C_ON=1'b0;
    defparam \uart_rx_inst.rxd_reg_83_LC_8_14_4 .SEQ_MODE=4'b1001;
    defparam \uart_rx_inst.rxd_reg_83_LC_8_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_rx_inst.rxd_reg_83_LC_8_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4045),
            .lcout(rxd_reg),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7374),
            .ce(),
            .sr(N__7267));
    defparam \uart_tx_inst.i782_3_lut_LC_9_1_0 .C_ON=1'b0;
    defparam \uart_tx_inst.i782_3_lut_LC_9_1_0 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.i782_3_lut_LC_9_1_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \uart_tx_inst.i782_3_lut_LC_9_1_0  (
            .in0(N__7714),
            .in1(N__5647),
            .in2(_gnd_net_),
            .in3(N__6775),
            .lcout(),
            .ltout(\uart_tx_inst.n910_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.prescale_reg__i13_LC_9_1_1 .C_ON=1'b0;
    defparam \uart_tx_inst.prescale_reg__i13_LC_9_1_1 .SEQ_MODE=4'b1000;
    defparam \uart_tx_inst.prescale_reg__i13_LC_9_1_1 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \uart_tx_inst.prescale_reg__i13_LC_9_1_1  (
            .in0(N__6566),
            .in1(N__7784),
            .in2(N__4033),
            .in3(N__6690),
            .lcout(\uart_tx_inst.prescale_reg_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7379),
            .ce(N__6476),
            .sr(N__7072));
    defparam \uart_tx_inst.i792_3_lut_LC_9_1_2 .C_ON=1'b0;
    defparam \uart_tx_inst.i792_3_lut_LC_9_1_2 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.i792_3_lut_LC_9_1_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \uart_tx_inst.i792_3_lut_LC_9_1_2  (
            .in0(N__8701),
            .in1(N__6016),
            .in2(_gnd_net_),
            .in3(N__6776),
            .lcout(),
            .ltout(\uart_tx_inst.n920_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.prescale_reg__i15_LC_9_1_3 .C_ON=1'b0;
    defparam \uart_tx_inst.prescale_reg__i15_LC_9_1_3 .SEQ_MODE=4'b1000;
    defparam \uart_tx_inst.prescale_reg__i15_LC_9_1_3 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \uart_tx_inst.prescale_reg__i15_LC_9_1_3  (
            .in0(N__6567),
            .in1(N__8775),
            .in2(N__4306),
            .in3(N__6691),
            .lcout(\uart_tx_inst.prescale_reg_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7379),
            .ce(N__6476),
            .sr(N__7072));
    defparam \uart_tx_inst.i802_3_lut_LC_9_1_4 .C_ON=1'b0;
    defparam \uart_tx_inst.i802_3_lut_LC_9_1_4 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.i802_3_lut_LC_9_1_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \uart_tx_inst.i802_3_lut_LC_9_1_4  (
            .in0(N__8491),
            .in1(N__5944),
            .in2(_gnd_net_),
            .in3(N__6777),
            .lcout(),
            .ltout(\uart_tx_inst.n930_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.prescale_reg__i17_LC_9_1_5 .C_ON=1'b0;
    defparam \uart_tx_inst.prescale_reg__i17_LC_9_1_5 .SEQ_MODE=4'b1000;
    defparam \uart_tx_inst.prescale_reg__i17_LC_9_1_5 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \uart_tx_inst.prescale_reg__i17_LC_9_1_5  (
            .in0(N__6568),
            .in1(N__8571),
            .in2(N__4303),
            .in3(N__6692),
            .lcout(\uart_tx_inst.prescale_reg_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7379),
            .ce(N__6476),
            .sr(N__7072));
    defparam \uart_tx_inst.i12_4_lut_LC_9_1_6 .C_ON=1'b0;
    defparam \uart_tx_inst.i12_4_lut_LC_9_1_6 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.i12_4_lut_LC_9_1_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \uart_tx_inst.i12_4_lut_LC_9_1_6  (
            .in0(N__5955),
            .in1(N__6027),
            .in2(N__6000),
            .in3(N__5658),
            .lcout(\uart_tx_inst.n31_adj_199 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.i2_3_lut_4_lut_LC_9_1_7 .C_ON=1'b0;
    defparam \uart_tx_inst.i2_3_lut_4_lut_LC_9_1_7 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.i2_3_lut_4_lut_LC_9_1_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \uart_tx_inst.i2_3_lut_4_lut_LC_9_1_7  (
            .in0(N__6774),
            .in1(N__7073),
            .in2(N__6592),
            .in3(N__6689),
            .lcout(\uart_tx_inst.n873 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.prescale_reg__i14_LC_9_2_0 .C_ON=1'b0;
    defparam \uart_tx_inst.prescale_reg__i14_LC_9_2_0 .SEQ_MODE=4'b1000;
    defparam \uart_tx_inst.prescale_reg__i14_LC_9_2_0 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \uart_tx_inst.prescale_reg__i14_LC_9_2_0  (
            .in0(N__6570),
            .in1(N__4294),
            .in2(N__8872),
            .in3(N__6697),
            .lcout(\uart_tx_inst.prescale_reg_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7378),
            .ce(N__6464),
            .sr(N__7175));
    defparam \uart_tx_inst.i747_3_lut_LC_9_2_1 .C_ON=1'b0;
    defparam \uart_tx_inst.i747_3_lut_LC_9_2_1 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.i747_3_lut_LC_9_2_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \uart_tx_inst.i747_3_lut_LC_9_2_1  (
            .in0(N__8107),
            .in1(N__5836),
            .in2(_gnd_net_),
            .in3(N__6804),
            .lcout(),
            .ltout(\uart_tx_inst.n875_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.prescale_reg__i6_LC_9_2_2 .C_ON=1'b0;
    defparam \uart_tx_inst.prescale_reg__i6_LC_9_2_2 .SEQ_MODE=4'b1000;
    defparam \uart_tx_inst.prescale_reg__i6_LC_9_2_2 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \uart_tx_inst.prescale_reg__i6_LC_9_2_2  (
            .in0(N__8871),
            .in1(N__6574),
            .in2(N__4288),
            .in3(N__6698),
            .lcout(\uart_tx_inst.prescale_reg_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7378),
            .ce(N__6464),
            .sr(N__7175));
    defparam \uart_tx_inst.i752_3_lut_LC_9_2_3 .C_ON=1'b0;
    defparam \uart_tx_inst.i752_3_lut_LC_9_2_3 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.i752_3_lut_LC_9_2_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \uart_tx_inst.i752_3_lut_LC_9_2_3  (
            .in0(N__8080),
            .in1(N__5809),
            .in2(_gnd_net_),
            .in3(N__6805),
            .lcout(),
            .ltout(\uart_tx_inst.n880_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.prescale_reg__i7_LC_9_2_4 .C_ON=1'b0;
    defparam \uart_tx_inst.prescale_reg__i7_LC_9_2_4 .SEQ_MODE=4'b1000;
    defparam \uart_tx_inst.prescale_reg__i7_LC_9_2_4 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \uart_tx_inst.prescale_reg__i7_LC_9_2_4  (
            .in0(N__8776),
            .in1(N__6575),
            .in2(N__4327),
            .in3(N__6699),
            .lcout(\uart_tx_inst.prescale_reg_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7378),
            .ce(N__6464),
            .sr(N__7175));
    defparam \uart_tx_inst.i767_3_lut_LC_9_2_5 .C_ON=1'b0;
    defparam \uart_tx_inst.i767_3_lut_LC_9_2_5 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.i767_3_lut_LC_9_2_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \uart_tx_inst.i767_3_lut_LC_9_2_5  (
            .in0(N__5743),
            .in1(N__7998),
            .in2(_gnd_net_),
            .in3(N__6806),
            .lcout(),
            .ltout(\uart_tx_inst.n895_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.prescale_reg__i10_LC_9_2_6 .C_ON=1'b0;
    defparam \uart_tx_inst.prescale_reg__i10_LC_9_2_6 .SEQ_MODE=4'b1000;
    defparam \uart_tx_inst.prescale_reg__i10_LC_9_2_6 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \uart_tx_inst.prescale_reg__i10_LC_9_2_6  (
            .in0(N__8462),
            .in1(N__6573),
            .in2(N__4324),
            .in3(N__6696),
            .lcout(\uart_tx_inst.prescale_reg_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7378),
            .ce(N__6464),
            .sr(N__7175));
    defparam \uart_tx_inst.prescale_reg__i16_LC_9_3_2 .C_ON=1'b0;
    defparam \uart_tx_inst.prescale_reg__i16_LC_9_3_2 .SEQ_MODE=4'b1000;
    defparam \uart_tx_inst.prescale_reg__i16_LC_9_3_2 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \uart_tx_inst.prescale_reg__i16_LC_9_3_2  (
            .in0(N__6571),
            .in1(N__4318),
            .in2(N__8674),
            .in3(N__6723),
            .lcout(\uart_tx_inst.prescale_reg_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7377),
            .ce(N__6465),
            .sr(N__7132));
    defparam \uart_tx_inst.prescale_reg__i18_LC_9_3_4 .C_ON=1'b0;
    defparam \uart_tx_inst.prescale_reg__i18_LC_9_3_4 .SEQ_MODE=4'b1000;
    defparam \uart_tx_inst.prescale_reg__i18_LC_9_3_4 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \uart_tx_inst.prescale_reg__i18_LC_9_3_4  (
            .in0(N__6572),
            .in1(N__4312),
            .in2(N__8464),
            .in3(N__6724),
            .lcout(\uart_tx_inst.prescale_reg_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7377),
            .ce(N__6465),
            .sr(N__7132));
    defparam \uart_tx_inst.i772_3_lut_LC_9_3_5 .C_ON=1'b0;
    defparam \uart_tx_inst.i772_3_lut_LC_9_3_5 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.i772_3_lut_LC_9_3_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \uart_tx_inst.i772_3_lut_LC_9_3_5  (
            .in0(N__7909),
            .in1(N__5707),
            .in2(_gnd_net_),
            .in3(N__6835),
            .lcout(),
            .ltout(\uart_tx_inst.n900_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.prescale_reg__i11_LC_9_3_6 .C_ON=1'b0;
    defparam \uart_tx_inst.prescale_reg__i11_LC_9_3_6 .SEQ_MODE=4'b1000;
    defparam \uart_tx_inst.prescale_reg__i11_LC_9_3_6 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \uart_tx_inst.prescale_reg__i11_LC_9_3_6  (
            .in0(N__7969),
            .in1(N__6576),
            .in2(N__4321),
            .in3(N__6722),
            .lcout(\uart_tx_inst.prescale_reg_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7377),
            .ce(N__6465),
            .sr(N__7132));
    defparam \uart_tx_inst.i797_3_lut_LC_9_4_1 .C_ON=1'b0;
    defparam \uart_tx_inst.i797_3_lut_LC_9_4_1 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.i797_3_lut_LC_9_4_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \uart_tx_inst.i797_3_lut_LC_9_4_1  (
            .in0(N__8596),
            .in1(N__5977),
            .in2(_gnd_net_),
            .in3(N__6834),
            .lcout(\uart_tx_inst.n925 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.i807_3_lut_LC_9_4_4 .C_ON=1'b0;
    defparam \uart_tx_inst.i807_3_lut_LC_9_4_4 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.i807_3_lut_LC_9_4_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uart_tx_inst.i807_3_lut_LC_9_4_4  (
            .in0(N__6833),
            .in1(N__8131),
            .in2(_gnd_net_),
            .in3(N__5902),
            .lcout(\uart_tx_inst.n935 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.prescale_reg__i0_LC_9_5_0 .C_ON=1'b1;
    defparam \uart_rx_inst.prescale_reg__i0_LC_9_5_0 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.prescale_reg__i0_LC_9_5_0 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \uart_rx_inst.prescale_reg__i0_LC_9_5_0  (
            .in0(N__6322),
            .in1(N__4594),
            .in2(N__4576),
            .in3(N__4558),
            .lcout(\uart_rx_inst.prescale_reg_0 ),
            .ltout(),
            .carryin(bfn_9_5_0_),
            .carryout(\uart_rx_inst.n1564 ),
            .clk(N__7369),
            .ce(N__4555),
            .sr(N__4543));
    defparam \uart_rx_inst.sub_10_add_2_3_lut_LC_9_5_1 .C_ON=1'b1;
    defparam \uart_rx_inst.sub_10_add_2_3_lut_LC_9_5_1 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.sub_10_add_2_3_lut_LC_9_5_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \uart_rx_inst.sub_10_add_2_3_lut_LC_9_5_1  (
            .in0(N__6320),
            .in1(N__4528),
            .in2(N__4934),
            .in3(N__4501),
            .lcout(\uart_rx_inst.n819 ),
            .ltout(),
            .carryin(\uart_rx_inst.n1564 ),
            .carryout(\uart_rx_inst.n1565 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.sub_10_add_2_4_lut_LC_9_5_2 .C_ON=1'b1;
    defparam \uart_rx_inst.sub_10_add_2_4_lut_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.sub_10_add_2_4_lut_LC_9_5_2 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \uart_rx_inst.sub_10_add_2_4_lut_LC_9_5_2  (
            .in0(N__6321),
            .in1(N__4901),
            .in2(N__4498),
            .in3(N__4465),
            .lcout(\uart_rx_inst.n814 ),
            .ltout(),
            .carryin(\uart_rx_inst.n1565 ),
            .carryout(\uart_rx_inst.n1566 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.sub_10_add_2_5_lut_LC_9_5_3 .C_ON=1'b1;
    defparam \uart_rx_inst.sub_10_add_2_5_lut_LC_9_5_3 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.sub_10_add_2_5_lut_LC_9_5_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \uart_rx_inst.sub_10_add_2_5_lut_LC_9_5_3  (
            .in0(N__5050),
            .in1(N__4462),
            .in2(N__4935),
            .in3(N__4444),
            .lcout(\uart_rx_inst.n809 ),
            .ltout(),
            .carryin(\uart_rx_inst.n1566 ),
            .carryout(\uart_rx_inst.n1567 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.sub_10_add_2_6_lut_LC_9_5_4 .C_ON=1'b1;
    defparam \uart_rx_inst.sub_10_add_2_6_lut_LC_9_5_4 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.sub_10_add_2_6_lut_LC_9_5_4 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \uart_rx_inst.sub_10_add_2_6_lut_LC_9_5_4  (
            .in0(N__5026),
            .in1(N__4905),
            .in2(N__4441),
            .in3(N__4414),
            .lcout(\uart_rx_inst.n804 ),
            .ltout(),
            .carryin(\uart_rx_inst.n1567 ),
            .carryout(\uart_rx_inst.n1568 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.sub_10_add_2_7_lut_LC_9_5_5 .C_ON=1'b1;
    defparam \uart_rx_inst.sub_10_add_2_7_lut_LC_9_5_5 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.sub_10_add_2_7_lut_LC_9_5_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \uart_rx_inst.sub_10_add_2_7_lut_LC_9_5_5  (
            .in0(N__4411),
            .in1(N__4399),
            .in2(N__4936),
            .in3(N__4375),
            .lcout(\uart_rx_inst.n799 ),
            .ltout(),
            .carryin(\uart_rx_inst.n1568 ),
            .carryout(\uart_rx_inst.n1569 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.sub_10_add_2_8_lut_LC_9_5_6 .C_ON=1'b1;
    defparam \uart_rx_inst.sub_10_add_2_8_lut_LC_9_5_6 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.sub_10_add_2_8_lut_LC_9_5_6 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \uart_rx_inst.sub_10_add_2_8_lut_LC_9_5_6  (
            .in0(N__5077),
            .in1(N__4909),
            .in2(N__4372),
            .in3(N__4351),
            .lcout(\uart_rx_inst.n794 ),
            .ltout(),
            .carryin(\uart_rx_inst.n1569 ),
            .carryout(\uart_rx_inst.n1570 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.sub_10_add_2_9_lut_LC_9_5_7 .C_ON=1'b1;
    defparam \uart_rx_inst.sub_10_add_2_9_lut_LC_9_5_7 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.sub_10_add_2_9_lut_LC_9_5_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \uart_rx_inst.sub_10_add_2_9_lut_LC_9_5_7  (
            .in0(N__5035),
            .in1(N__4348),
            .in2(N__4937),
            .in3(N__4330),
            .lcout(\uart_rx_inst.n789 ),
            .ltout(),
            .carryin(\uart_rx_inst.n1570 ),
            .carryout(\uart_rx_inst.n1571 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.sub_10_add_2_10_lut_LC_9_6_0 .C_ON=1'b1;
    defparam \uart_rx_inst.sub_10_add_2_10_lut_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.sub_10_add_2_10_lut_LC_9_6_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \uart_rx_inst.sub_10_add_2_10_lut_LC_9_6_0  (
            .in0(N__4813),
            .in1(N__4795),
            .in2(N__4938),
            .in3(N__4762),
            .lcout(\uart_rx_inst.n784 ),
            .ltout(),
            .carryin(bfn_9_6_0_),
            .carryout(\uart_rx_inst.n1572 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.sub_10_add_2_11_lut_LC_9_6_1 .C_ON=1'b1;
    defparam \uart_rx_inst.sub_10_add_2_11_lut_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.sub_10_add_2_11_lut_LC_9_6_1 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \uart_rx_inst.sub_10_add_2_11_lut_LC_9_6_1  (
            .in0(N__4825),
            .in1(N__4916),
            .in2(N__4758),
            .in3(N__4732),
            .lcout(\uart_rx_inst.n779 ),
            .ltout(),
            .carryin(\uart_rx_inst.n1572 ),
            .carryout(\uart_rx_inst.n1573 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.sub_10_add_2_12_lut_LC_9_6_2 .C_ON=1'b1;
    defparam \uart_rx_inst.sub_10_add_2_12_lut_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.sub_10_add_2_12_lut_LC_9_6_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \uart_rx_inst.sub_10_add_2_12_lut_LC_9_6_2  (
            .in0(N__4729),
            .in1(N__4716),
            .in2(N__4939),
            .in3(N__4696),
            .lcout(\uart_rx_inst.n774 ),
            .ltout(),
            .carryin(\uart_rx_inst.n1573 ),
            .carryout(\uart_rx_inst.n1574 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.sub_10_add_2_13_lut_LC_9_6_3 .C_ON=1'b1;
    defparam \uart_rx_inst.sub_10_add_2_13_lut_LC_9_6_3 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.sub_10_add_2_13_lut_LC_9_6_3 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \uart_rx_inst.sub_10_add_2_13_lut_LC_9_6_3  (
            .in0(N__4801),
            .in1(N__4920),
            .in2(N__4693),
            .in3(N__4672),
            .lcout(\uart_rx_inst.n769 ),
            .ltout(),
            .carryin(\uart_rx_inst.n1574 ),
            .carryout(\uart_rx_inst.n1575 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.sub_10_add_2_14_lut_LC_9_6_4 .C_ON=1'b1;
    defparam \uart_rx_inst.sub_10_add_2_14_lut_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.sub_10_add_2_14_lut_LC_9_6_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \uart_rx_inst.sub_10_add_2_14_lut_LC_9_6_4  (
            .in0(N__6220),
            .in1(N__4669),
            .in2(N__4940),
            .in3(N__4648),
            .lcout(\uart_rx_inst.n764 ),
            .ltout(),
            .carryin(\uart_rx_inst.n1575 ),
            .carryout(\uart_rx_inst.n1576 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.sub_10_add_2_15_lut_LC_9_6_5 .C_ON=1'b1;
    defparam \uart_rx_inst.sub_10_add_2_15_lut_LC_9_6_5 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.sub_10_add_2_15_lut_LC_9_6_5 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \uart_rx_inst.sub_10_add_2_15_lut_LC_9_6_5  (
            .in0(N__4807),
            .in1(N__4924),
            .in2(N__4645),
            .in3(N__4624),
            .lcout(\uart_rx_inst.n759 ),
            .ltout(),
            .carryin(\uart_rx_inst.n1576 ),
            .carryout(\uart_rx_inst.n1577 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.sub_10_add_2_16_lut_LC_9_6_6 .C_ON=1'b1;
    defparam \uart_rx_inst.sub_10_add_2_16_lut_LC_9_6_6 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.sub_10_add_2_16_lut_LC_9_6_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \uart_rx_inst.sub_10_add_2_16_lut_LC_9_6_6  (
            .in0(N__5086),
            .in1(N__4621),
            .in2(N__4941),
            .in3(N__4600),
            .lcout(\uart_rx_inst.n754 ),
            .ltout(),
            .carryin(\uart_rx_inst.n1577 ),
            .carryout(\uart_rx_inst.n1578 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.sub_10_add_2_17_lut_LC_9_6_7 .C_ON=1'b1;
    defparam \uart_rx_inst.sub_10_add_2_17_lut_LC_9_6_7 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.sub_10_add_2_17_lut_LC_9_6_7 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \uart_rx_inst.sub_10_add_2_17_lut_LC_9_6_7  (
            .in0(N__4819),
            .in1(N__4928),
            .in2(N__5017),
            .in3(N__4996),
            .lcout(\uart_rx_inst.n749 ),
            .ltout(),
            .carryin(\uart_rx_inst.n1578 ),
            .carryout(\uart_rx_inst.n1579 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.sub_10_add_2_18_lut_LC_9_7_0 .C_ON=1'b1;
    defparam \uart_rx_inst.sub_10_add_2_18_lut_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.sub_10_add_2_18_lut_LC_9_7_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \uart_rx_inst.sub_10_add_2_18_lut_LC_9_7_0  (
            .in0(N__5041),
            .in1(N__4992),
            .in2(N__4942),
            .in3(N__4972),
            .lcout(\uart_rx_inst.n744 ),
            .ltout(),
            .carryin(bfn_9_7_0_),
            .carryout(\uart_rx_inst.n1580 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.sub_10_add_2_19_lut_LC_9_7_1 .C_ON=1'b1;
    defparam \uart_rx_inst.sub_10_add_2_19_lut_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.sub_10_add_2_19_lut_LC_9_7_1 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \uart_rx_inst.sub_10_add_2_19_lut_LC_9_7_1  (
            .in0(N__5059),
            .in1(N__4932),
            .in2(N__4969),
            .in3(N__4945),
            .lcout(\uart_rx_inst.n739 ),
            .ltout(),
            .carryin(\uart_rx_inst.n1580 ),
            .carryout(\uart_rx_inst.n1581 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.sub_10_add_2_20_lut_LC_9_7_2 .C_ON=1'b0;
    defparam \uart_rx_inst.sub_10_add_2_20_lut_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.sub_10_add_2_20_lut_LC_9_7_2 .LUT_INIT=16'b1101100001110010;
    LogicCell40 \uart_rx_inst.sub_10_add_2_20_lut_LC_9_7_2  (
            .in0(N__4933),
            .in1(N__4852),
            .in2(N__5068),
            .in3(N__4837),
            .lcout(\uart_rx_inst.n729 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.i1578_2_lut_LC_9_7_3 .C_ON=1'b0;
    defparam \uart_rx_inst.i1578_2_lut_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i1578_2_lut_LC_9_7_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uart_rx_inst.i1578_2_lut_LC_9_7_3  (
            .in0(N__6302),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8028),
            .lcout(\uart_rx_inst.n1743 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.i1569_2_lut_LC_9_7_4 .C_ON=1'b0;
    defparam \uart_rx_inst.i1569_2_lut_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i1569_2_lut_LC_9_7_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uart_rx_inst.i1569_2_lut_LC_9_7_4  (
            .in0(N__8697),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6303),
            .lcout(\uart_rx_inst.n1740 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.i1577_2_lut_LC_9_7_5 .C_ON=1'b0;
    defparam \uart_rx_inst.i1577_2_lut_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i1577_2_lut_LC_9_7_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uart_rx_inst.i1577_2_lut_LC_9_7_5  (
            .in0(N__6300),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8056),
            .lcout(\uart_rx_inst.n1741 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.i1574_2_lut_LC_9_7_6 .C_ON=1'b0;
    defparam \uart_rx_inst.i1574_2_lut_LC_9_7_6 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i1574_2_lut_LC_9_7_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uart_rx_inst.i1574_2_lut_LC_9_7_6  (
            .in0(N__7707),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6304),
            .lcout(\uart_rx_inst.n1747 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.i1572_2_lut_LC_9_7_7 .C_ON=1'b0;
    defparam \uart_rx_inst.i1572_2_lut_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i1572_2_lut_LC_9_7_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uart_rx_inst.i1572_2_lut_LC_9_7_7  (
            .in0(N__6301),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7905),
            .lcout(\uart_rx_inst.n1745 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.i1563_2_lut_LC_9_8_0 .C_ON=1'b0;
    defparam \uart_rx_inst.i1563_2_lut_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i1563_2_lut_LC_9_8_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uart_rx_inst.i1563_2_lut_LC_9_8_0  (
            .in0(N__8799),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6296),
            .lcout(\uart_rx_inst.n1750 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.i1580_2_lut_LC_9_8_1 .C_ON=1'b0;
    defparam \uart_rx_inst.i1580_2_lut_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i1580_2_lut_LC_9_8_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uart_rx_inst.i1580_2_lut_LC_9_8_1  (
            .in0(N__6295),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8106),
            .lcout(\uart_rx_inst.n1755 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.i1565_2_lut_LC_9_8_2 .C_ON=1'b0;
    defparam \uart_rx_inst.i1565_2_lut_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i1565_2_lut_LC_9_8_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_rx_inst.i1565_2_lut_LC_9_8_2  (
            .in0(_gnd_net_),
            .in1(N__8130),
            .in2(_gnd_net_),
            .in3(N__6298),
            .lcout(\uart_rx_inst.n1754 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.i1576_2_lut_LC_9_8_3 .C_ON=1'b0;
    defparam \uart_rx_inst.i1576_2_lut_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i1576_2_lut_LC_9_8_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uart_rx_inst.i1576_2_lut_LC_9_8_3  (
            .in0(N__6294),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8487),
            .lcout(\uart_rx_inst.n1751 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.i1566_2_lut_LC_9_8_4 .C_ON=1'b0;
    defparam \uart_rx_inst.i1566_2_lut_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i1566_2_lut_LC_9_8_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_rx_inst.i1566_2_lut_LC_9_8_4  (
            .in0(_gnd_net_),
            .in1(N__6961),
            .in2(_gnd_net_),
            .in3(N__6297),
            .lcout(\uart_rx_inst.n1758 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.i1570_2_lut_LC_9_8_5 .C_ON=1'b0;
    defparam \uart_rx_inst.i1570_2_lut_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i1570_2_lut_LC_9_8_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uart_rx_inst.i1570_2_lut_LC_9_8_5  (
            .in0(N__6299),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8595),
            .lcout(\uart_rx_inst.n1742 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.i1581_2_lut_LC_9_8_6 .C_ON=1'b0;
    defparam \uart_rx_inst.i1581_2_lut_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i1581_2_lut_LC_9_8_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_rx_inst.i1581_2_lut_LC_9_8_6  (
            .in0(_gnd_net_),
            .in1(N__8079),
            .in2(_gnd_net_),
            .in3(N__6293),
            .lcout(\uart_rx_inst.n1739 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.i1567_2_lut_LC_9_8_7 .C_ON=1'b0;
    defparam \uart_rx_inst.i1567_2_lut_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i1567_2_lut_LC_9_8_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uart_rx_inst.i1567_2_lut_LC_9_8_7  (
            .in0(N__6292),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6934),
            .lcout(\uart_rx_inst.n1757 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.data_reg__i2_LC_9_9_0 .C_ON=1'b0;
    defparam \uart_rx_inst.data_reg__i2_LC_9_9_0 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.data_reg__i2_LC_9_9_0 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \uart_rx_inst.data_reg__i2_LC_9_9_0  (
            .in0(N__5321),
            .in1(N__5453),
            .in2(N__5163),
            .in3(N__5362),
            .lcout(data_reg_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7361),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.data_reg__i5_LC_9_9_1 .C_ON=1'b0;
    defparam \uart_rx_inst.data_reg__i5_LC_9_9_1 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.data_reg__i5_LC_9_9_1 .LUT_INIT=16'b1011100000000000;
    LogicCell40 \uart_rx_inst.data_reg__i5_LC_9_9_1  (
            .in0(N__5519),
            .in1(N__5361),
            .in2(N__5193),
            .in3(N__5324),
            .lcout(data_reg_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7361),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.data_reg__i3_LC_9_9_2 .C_ON=1'b0;
    defparam \uart_rx_inst.data_reg__i3_LC_9_9_2 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.data_reg__i3_LC_9_9_2 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \uart_rx_inst.data_reg__i3_LC_9_9_2  (
            .in0(N__5322),
            .in1(N__5553),
            .in2(N__5455),
            .in3(N__5363),
            .lcout(data_reg_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7361),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.data_reg__i1_LC_9_9_5 .C_ON=1'b0;
    defparam \uart_rx_inst.data_reg__i1_LC_9_9_5 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.data_reg__i1_LC_9_9_5 .LUT_INIT=16'b1011100000000000;
    LogicCell40 \uart_rx_inst.data_reg__i1_LC_9_9_5  (
            .in0(N__5483),
            .in1(N__5359),
            .in2(N__5164),
            .in3(N__5320),
            .lcout(data_reg_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7361),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.data_reg__i6_LC_9_9_6 .C_ON=1'b0;
    defparam \uart_rx_inst.data_reg__i6_LC_9_9_6 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.data_reg__i6_LC_9_9_6 .LUT_INIT=16'b1000100010100000;
    LogicCell40 \uart_rx_inst.data_reg__i6_LC_9_9_6  (
            .in0(N__5325),
            .in1(N__5186),
            .in2(N__5118),
            .in3(N__5364),
            .lcout(data_reg_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7361),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.data_reg__i4_LC_9_9_7 .C_ON=1'b0;
    defparam \uart_rx_inst.data_reg__i4_LC_9_9_7 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.data_reg__i4_LC_9_9_7 .LUT_INIT=16'b1011100000000000;
    LogicCell40 \uart_rx_inst.data_reg__i4_LC_9_9_7  (
            .in0(N__5552),
            .in1(N__5360),
            .in2(N__5526),
            .in3(N__5323),
            .lcout(data_reg_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7361),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.frame_error_reg_88_LC_9_10_3 .C_ON=1'b0;
    defparam \uart_rx_inst.frame_error_reg_88_LC_9_10_3 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.frame_error_reg_88_LC_9_10_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \uart_rx_inst.frame_error_reg_88_LC_9_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5294),
            .lcout(rx_frame_error_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7364),
            .ce(),
            .sr(N__5206));
    defparam \uart_rx_inst.output_axis_tdata_reg__i7_LC_9_12_1 .C_ON=1'b0;
    defparam \uart_rx_inst.output_axis_tdata_reg__i7_LC_9_12_1 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.output_axis_tdata_reg__i7_LC_9_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_rx_inst.output_axis_tdata_reg__i7_LC_9_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5194),
            .lcout(output_axis_tdata_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7372),
            .ce(N__5408),
            .sr(N__7254));
    defparam \uart_rx_inst.output_axis_tdata_reg__i3_LC_9_12_2 .C_ON=1'b0;
    defparam \uart_rx_inst.output_axis_tdata_reg__i3_LC_9_12_2 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.output_axis_tdata_reg__i3_LC_9_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_rx_inst.output_axis_tdata_reg__i3_LC_9_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5162),
            .lcout(output_axis_tdata_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7372),
            .ce(N__5408),
            .sr(N__7254));
    defparam \uart_rx_inst.output_axis_tdata_reg__i8_LC_9_12_3 .C_ON=1'b0;
    defparam \uart_rx_inst.output_axis_tdata_reg__i8_LC_9_12_3 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.output_axis_tdata_reg__i8_LC_9_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_rx_inst.output_axis_tdata_reg__i8_LC_9_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5122),
            .lcout(output_axis_tdata_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7372),
            .ce(N__5408),
            .sr(N__7254));
    defparam \uart_rx_inst.output_axis_tdata_reg__i5_LC_9_12_4 .C_ON=1'b0;
    defparam \uart_rx_inst.output_axis_tdata_reg__i5_LC_9_12_4 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.output_axis_tdata_reg__i5_LC_9_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_rx_inst.output_axis_tdata_reg__i5_LC_9_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5557),
            .lcout(output_axis_tdata_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7372),
            .ce(N__5408),
            .sr(N__7254));
    defparam \uart_rx_inst.output_axis_tdata_reg__i6_LC_9_12_5 .C_ON=1'b0;
    defparam \uart_rx_inst.output_axis_tdata_reg__i6_LC_9_12_5 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.output_axis_tdata_reg__i6_LC_9_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_rx_inst.output_axis_tdata_reg__i6_LC_9_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5527),
            .lcout(output_axis_tdata_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7372),
            .ce(N__5408),
            .sr(N__7254));
    defparam \uart_rx_inst.output_axis_tdata_reg__i2_LC_9_13_3 .C_ON=1'b0;
    defparam \uart_rx_inst.output_axis_tdata_reg__i2_LC_9_13_3 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.output_axis_tdata_reg__i2_LC_9_13_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart_rx_inst.output_axis_tdata_reg__i2_LC_9_13_3  (
            .in0(N__5493),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(output_axis_tdata_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7376),
            .ce(N__5419),
            .sr(N__7265));
    defparam \uart_rx_inst.output_axis_tdata_reg__i4_LC_9_13_7 .C_ON=1'b0;
    defparam \uart_rx_inst.output_axis_tdata_reg__i4_LC_9_13_7 .SEQ_MODE=4'b1000;
    defparam \uart_rx_inst.output_axis_tdata_reg__i4_LC_9_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_rx_inst.output_axis_tdata_reg__i4_LC_9_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5454),
            .lcout(output_axis_tdata_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7376),
            .ce(N__5419),
            .sr(N__7265));
    defparam \uart_tx_inst.i777_3_lut_LC_11_1_0 .C_ON=1'b0;
    defparam \uart_tx_inst.i777_3_lut_LC_11_1_0 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.i777_3_lut_LC_11_1_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uart_tx_inst.i777_3_lut_LC_11_1_0  (
            .in0(N__6809),
            .in1(N__7813),
            .in2(_gnd_net_),
            .in3(N__5680),
            .lcout(),
            .ltout(\uart_tx_inst.n905_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.prescale_reg__i12_LC_11_1_1 .C_ON=1'b0;
    defparam \uart_tx_inst.prescale_reg__i12_LC_11_1_1 .SEQ_MODE=4'b1000;
    defparam \uart_tx_inst.prescale_reg__i12_LC_11_1_1 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \uart_tx_inst.prescale_reg__i12_LC_11_1_1  (
            .in0(N__6594),
            .in1(N__7883),
            .in2(N__5380),
            .in3(N__6711),
            .lcout(\uart_tx_inst.prescale_reg_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7382),
            .ce(N__6477),
            .sr(N__7181));
    defparam \uart_tx_inst.i762_3_lut_LC_11_1_2 .C_ON=1'b0;
    defparam \uart_tx_inst.i762_3_lut_LC_11_1_2 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.i762_3_lut_LC_11_1_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uart_tx_inst.i762_3_lut_LC_11_1_2  (
            .in0(N__6808),
            .in1(N__8029),
            .in2(_gnd_net_),
            .in3(N__5773),
            .lcout(),
            .ltout(\uart_tx_inst.n890_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.prescale_reg__i9_LC_11_1_3 .C_ON=1'b0;
    defparam \uart_tx_inst.prescale_reg__i9_LC_11_1_3 .SEQ_MODE=4'b1000;
    defparam \uart_tx_inst.prescale_reg__i9_LC_11_1_3 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \uart_tx_inst.prescale_reg__i9_LC_11_1_3  (
            .in0(N__6595),
            .in1(N__8570),
            .in2(N__5377),
            .in3(N__6713),
            .lcout(\uart_tx_inst.prescale_reg_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7382),
            .ce(N__6477),
            .sr(N__7181));
    defparam \uart_tx_inst.i14_4_lut_LC_11_1_4 .C_ON=1'b0;
    defparam \uart_tx_inst.i14_4_lut_LC_11_1_4 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.i14_4_lut_LC_11_1_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \uart_tx_inst.i14_4_lut_LC_11_1_4  (
            .in0(N__5625),
            .in1(N__5610),
            .in2(N__5790),
            .in3(N__5691),
            .lcout(\uart_tx_inst.n33_adj_198 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.i732_3_lut_LC_11_1_5 .C_ON=1'b0;
    defparam \uart_tx_inst.i732_3_lut_LC_11_1_5 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.i732_3_lut_LC_11_1_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \uart_tx_inst.i732_3_lut_LC_11_1_5  (
            .in0(N__5572),
            .in1(N__6960),
            .in2(_gnd_net_),
            .in3(N__6810),
            .lcout(),
            .ltout(\uart_tx_inst.n860_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.prescale_reg__i3_LC_11_1_6 .C_ON=1'b0;
    defparam \uart_tx_inst.prescale_reg__i3_LC_11_1_6 .SEQ_MODE=4'b1000;
    defparam \uart_tx_inst.prescale_reg__i3_LC_11_1_6 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \uart_tx_inst.prescale_reg__i3_LC_11_1_6  (
            .in0(N__6712),
            .in1(N__7970),
            .in2(N__5632),
            .in3(N__6596),
            .lcout(\uart_tx_inst.prescale_reg_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7382),
            .ce(N__6477),
            .sr(N__7181));
    defparam \uart_tx_inst.i1524_3_lut_4_lut_LC_11_1_7 .C_ON=1'b0;
    defparam \uart_tx_inst.i1524_3_lut_4_lut_LC_11_1_7 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.i1524_3_lut_4_lut_LC_11_1_7 .LUT_INIT=16'b1111000011110100;
    LogicCell40 \uart_tx_inst.i1524_3_lut_4_lut_LC_11_1_7  (
            .in0(N__6593),
            .in1(N__6807),
            .in2(N__7240),
            .in3(N__6710),
            .lcout(\uart_tx_inst.n1170 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.prescale_reg__i0_LC_11_2_0 .C_ON=1'b1;
    defparam \uart_tx_inst.prescale_reg__i0_LC_11_2_0 .SEQ_MODE=4'b1000;
    defparam \uart_tx_inst.prescale_reg__i0_LC_11_2_0 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \uart_tx_inst.prescale_reg__i0_LC_11_2_0  (
            .in0(N__6837),
            .in1(N__6208),
            .in2(_gnd_net_),
            .in3(N__5629),
            .lcout(\uart_tx_inst.prescale_reg_0 ),
            .ltout(),
            .carryin(bfn_11_2_0_),
            .carryout(\uart_tx_inst.n1546 ),
            .clk(N__7380),
            .ce(N__6481),
            .sr(N__5596));
    defparam \uart_tx_inst.prescale_reg__i1_LC_11_2_1 .C_ON=1'b1;
    defparam \uart_tx_inst.prescale_reg__i1_LC_11_2_1 .SEQ_MODE=4'b1000;
    defparam \uart_tx_inst.prescale_reg__i1_LC_11_2_1 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \uart_tx_inst.prescale_reg__i1_LC_11_2_1  (
            .in0(N__6836),
            .in1(N__5626),
            .in2(N__8380),
            .in3(N__5614),
            .lcout(\uart_tx_inst.prescale_reg_1 ),
            .ltout(),
            .carryin(\uart_tx_inst.n1546 ),
            .carryout(\uart_tx_inst.n1547 ),
            .clk(N__7380),
            .ce(N__6481),
            .sr(N__5596));
    defparam \uart_tx_inst.prescale_reg__i2_LC_11_2_2 .C_ON=1'b1;
    defparam \uart_tx_inst.prescale_reg__i2_LC_11_2_2 .SEQ_MODE=4'b1000;
    defparam \uart_tx_inst.prescale_reg__i2_LC_11_2_2 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \uart_tx_inst.prescale_reg__i2_LC_11_2_2  (
            .in0(N__6838),
            .in1(N__5611),
            .in2(N__8374),
            .in3(N__5599),
            .lcout(\uart_tx_inst.prescale_reg_2 ),
            .ltout(),
            .carryin(\uart_tx_inst.n1547 ),
            .carryout(\uart_tx_inst.n1548 ),
            .clk(N__7380),
            .ce(N__6481),
            .sr(N__5596));
    defparam \uart_tx_inst.sub_5_add_2_5_lut_LC_11_2_3 .C_ON=1'b1;
    defparam \uart_tx_inst.sub_5_add_2_5_lut_LC_11_2_3 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.sub_5_add_2_5_lut_LC_11_2_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_tx_inst.sub_5_add_2_5_lut_LC_11_2_3  (
            .in0(_gnd_net_),
            .in1(N__5586),
            .in2(N__8381),
            .in3(N__5566),
            .lcout(\uart_tx_inst.n33 ),
            .ltout(),
            .carryin(\uart_tx_inst.n1548 ),
            .carryout(\uart_tx_inst.n1549 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.sub_5_add_2_6_lut_LC_11_2_4 .C_ON=1'b1;
    defparam \uart_tx_inst.sub_5_add_2_6_lut_LC_11_2_4 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.sub_5_add_2_6_lut_LC_11_2_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_tx_inst.sub_5_add_2_6_lut_LC_11_2_4  (
            .in0(_gnd_net_),
            .in1(N__8366),
            .in2(N__6877),
            .in3(N__5563),
            .lcout(\uart_tx_inst.n32 ),
            .ltout(),
            .carryin(\uart_tx_inst.n1549 ),
            .carryout(\uart_tx_inst.n1550 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.sub_5_add_2_7_lut_LC_11_2_5 .C_ON=1'b1;
    defparam \uart_tx_inst.sub_5_add_2_7_lut_LC_11_2_5 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.sub_5_add_2_7_lut_LC_11_2_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_tx_inst.sub_5_add_2_7_lut_LC_11_2_5  (
            .in0(_gnd_net_),
            .in1(N__6850),
            .in2(N__8382),
            .in3(N__5560),
            .lcout(\uart_tx_inst.n31 ),
            .ltout(),
            .carryin(\uart_tx_inst.n1550 ),
            .carryout(\uart_tx_inst.n1551 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.sub_5_add_2_8_lut_LC_11_2_6 .C_ON=1'b1;
    defparam \uart_tx_inst.sub_5_add_2_8_lut_LC_11_2_6 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.sub_5_add_2_8_lut_LC_11_2_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_tx_inst.sub_5_add_2_8_lut_LC_11_2_6  (
            .in0(_gnd_net_),
            .in1(N__8370),
            .in2(N__5854),
            .in3(N__5827),
            .lcout(\uart_tx_inst.n30 ),
            .ltout(),
            .carryin(\uart_tx_inst.n1551 ),
            .carryout(\uart_tx_inst.n1552 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.sub_5_add_2_9_lut_LC_11_2_7 .C_ON=1'b1;
    defparam \uart_tx_inst.sub_5_add_2_9_lut_LC_11_2_7 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.sub_5_add_2_9_lut_LC_11_2_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_tx_inst.sub_5_add_2_9_lut_LC_11_2_7  (
            .in0(_gnd_net_),
            .in1(N__5824),
            .in2(N__8383),
            .in3(N__5800),
            .lcout(\uart_tx_inst.n29 ),
            .ltout(),
            .carryin(\uart_tx_inst.n1552 ),
            .carryout(\uart_tx_inst.n1553 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.sub_5_add_2_10_lut_LC_11_3_0 .C_ON=1'b1;
    defparam \uart_tx_inst.sub_5_add_2_10_lut_LC_11_3_0 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.sub_5_add_2_10_lut_LC_11_3_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_tx_inst.sub_5_add_2_10_lut_LC_11_3_0  (
            .in0(_gnd_net_),
            .in1(N__6499),
            .in2(N__8376),
            .in3(N__5797),
            .lcout(\uart_tx_inst.n28 ),
            .ltout(),
            .carryin(bfn_11_3_0_),
            .carryout(\uart_tx_inst.n1554 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.sub_5_add_2_11_lut_LC_11_3_1 .C_ON=1'b1;
    defparam \uart_tx_inst.sub_5_add_2_11_lut_LC_11_3_1 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.sub_5_add_2_11_lut_LC_11_3_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_tx_inst.sub_5_add_2_11_lut_LC_11_3_1  (
            .in0(_gnd_net_),
            .in1(N__8347),
            .in2(N__5794),
            .in3(N__5764),
            .lcout(\uart_tx_inst.n27 ),
            .ltout(),
            .carryin(\uart_tx_inst.n1554 ),
            .carryout(\uart_tx_inst.n1555 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.sub_5_add_2_12_lut_LC_11_3_2 .C_ON=1'b1;
    defparam \uart_tx_inst.sub_5_add_2_12_lut_LC_11_3_2 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.sub_5_add_2_12_lut_LC_11_3_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_tx_inst.sub_5_add_2_12_lut_LC_11_3_2  (
            .in0(_gnd_net_),
            .in1(N__5761),
            .in2(N__8377),
            .in3(N__5731),
            .lcout(\uart_tx_inst.n26 ),
            .ltout(),
            .carryin(\uart_tx_inst.n1555 ),
            .carryout(\uart_tx_inst.n1556 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.sub_5_add_2_13_lut_LC_11_3_3 .C_ON=1'b1;
    defparam \uart_tx_inst.sub_5_add_2_13_lut_LC_11_3_3 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.sub_5_add_2_13_lut_LC_11_3_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_tx_inst.sub_5_add_2_13_lut_LC_11_3_3  (
            .in0(_gnd_net_),
            .in1(N__8351),
            .in2(N__5728),
            .in3(N__5698),
            .lcout(\uart_tx_inst.n25 ),
            .ltout(),
            .carryin(\uart_tx_inst.n1556 ),
            .carryout(\uart_tx_inst.n1557 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.sub_5_add_2_14_lut_LC_11_3_4 .C_ON=1'b1;
    defparam \uart_tx_inst.sub_5_add_2_14_lut_LC_11_3_4 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.sub_5_add_2_14_lut_LC_11_3_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_tx_inst.sub_5_add_2_14_lut_LC_11_3_4  (
            .in0(_gnd_net_),
            .in1(N__5695),
            .in2(N__8378),
            .in3(N__5671),
            .lcout(\uart_tx_inst.n24 ),
            .ltout(),
            .carryin(\uart_tx_inst.n1557 ),
            .carryout(\uart_tx_inst.n1558 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.sub_5_add_2_15_lut_LC_11_3_5 .C_ON=1'b1;
    defparam \uart_tx_inst.sub_5_add_2_15_lut_LC_11_3_5 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.sub_5_add_2_15_lut_LC_11_3_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_tx_inst.sub_5_add_2_15_lut_LC_11_3_5  (
            .in0(_gnd_net_),
            .in1(N__8355),
            .in2(N__5668),
            .in3(N__5635),
            .lcout(\uart_tx_inst.n23 ),
            .ltout(),
            .carryin(\uart_tx_inst.n1558 ),
            .carryout(\uart_tx_inst.n1559 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.sub_5_add_2_16_lut_LC_11_3_6 .C_ON=1'b1;
    defparam \uart_tx_inst.sub_5_add_2_16_lut_LC_11_3_6 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.sub_5_add_2_16_lut_LC_11_3_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_tx_inst.sub_5_add_2_16_lut_LC_11_3_6  (
            .in0(_gnd_net_),
            .in1(N__6070),
            .in2(N__8379),
            .in3(N__6040),
            .lcout(\uart_tx_inst.n22 ),
            .ltout(),
            .carryin(\uart_tx_inst.n1559 ),
            .carryout(\uart_tx_inst.n1560 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.sub_5_add_2_17_lut_LC_11_3_7 .C_ON=1'b1;
    defparam \uart_tx_inst.sub_5_add_2_17_lut_LC_11_3_7 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.sub_5_add_2_17_lut_LC_11_3_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_tx_inst.sub_5_add_2_17_lut_LC_11_3_7  (
            .in0(_gnd_net_),
            .in1(N__8359),
            .in2(N__6037),
            .in3(N__6004),
            .lcout(\uart_tx_inst.n21 ),
            .ltout(),
            .carryin(\uart_tx_inst.n1560 ),
            .carryout(\uart_tx_inst.n1561 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.sub_5_add_2_18_lut_LC_11_4_0 .C_ON=1'b1;
    defparam \uart_tx_inst.sub_5_add_2_18_lut_LC_11_4_0 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.sub_5_add_2_18_lut_LC_11_4_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_tx_inst.sub_5_add_2_18_lut_LC_11_4_0  (
            .in0(_gnd_net_),
            .in1(N__6001),
            .in2(N__8375),
            .in3(N__5968),
            .lcout(\uart_tx_inst.n20 ),
            .ltout(),
            .carryin(bfn_11_4_0_),
            .carryout(\uart_tx_inst.n1562 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.sub_5_add_2_19_lut_LC_11_4_1 .C_ON=1'b1;
    defparam \uart_tx_inst.sub_5_add_2_19_lut_LC_11_4_1 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.sub_5_add_2_19_lut_LC_11_4_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_tx_inst.sub_5_add_2_19_lut_LC_11_4_1  (
            .in0(_gnd_net_),
            .in1(N__8342),
            .in2(N__5965),
            .in3(N__5932),
            .lcout(\uart_tx_inst.n19 ),
            .ltout(),
            .carryin(\uart_tx_inst.n1562 ),
            .carryout(\uart_tx_inst.n1563 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.sub_5_add_2_20_lut_LC_11_4_2 .C_ON=1'b0;
    defparam \uart_tx_inst.sub_5_add_2_20_lut_LC_11_4_2 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.sub_5_add_2_20_lut_LC_11_4_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_tx_inst.sub_5_add_2_20_lut_LC_11_4_2  (
            .in0(N__8343),
            .in1(N__5929),
            .in2(_gnd_net_),
            .in3(N__5905),
            .lcout(\uart_tx_inst.n18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.add_144_2_lut_LC_11_5_0 .C_ON=1'b1;
    defparam \uart_rx_inst.add_144_2_lut_LC_11_5_0 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.add_144_2_lut_LC_11_5_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_rx_inst.add_144_2_lut_LC_11_5_0  (
            .in0(_gnd_net_),
            .in1(N__7959),
            .in2(_gnd_net_),
            .in3(N__5881),
            .lcout(\uart_rx_inst.n328 ),
            .ltout(),
            .carryin(bfn_11_5_0_),
            .carryout(\uart_rx_inst.n1530 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.add_144_3_lut_LC_11_5_1 .C_ON=1'b1;
    defparam \uart_rx_inst.add_144_3_lut_LC_11_5_1 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.add_144_3_lut_LC_11_5_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_rx_inst.add_144_3_lut_LC_11_5_1  (
            .in0(_gnd_net_),
            .in1(N__8241),
            .in2(N__7881),
            .in3(N__5869),
            .lcout(\uart_rx_inst.n327 ),
            .ltout(),
            .carryin(\uart_rx_inst.n1530 ),
            .carryout(\uart_rx_inst.n1531 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.add_144_4_lut_LC_11_5_2 .C_ON=1'b1;
    defparam \uart_rx_inst.add_144_4_lut_LC_11_5_2 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.add_144_4_lut_LC_11_5_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_rx_inst.add_144_4_lut_LC_11_5_2  (
            .in0(_gnd_net_),
            .in1(N__8245),
            .in2(N__7785),
            .in3(N__5857),
            .lcout(\uart_rx_inst.n326 ),
            .ltout(),
            .carryin(\uart_rx_inst.n1531 ),
            .carryout(\uart_rx_inst.n1532 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.add_144_5_lut_LC_11_5_3 .C_ON=1'b1;
    defparam \uart_rx_inst.add_144_5_lut_LC_11_5_3 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.add_144_5_lut_LC_11_5_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_rx_inst.add_144_5_lut_LC_11_5_3  (
            .in0(_gnd_net_),
            .in1(N__8242),
            .in2(N__8858),
            .in3(N__6172),
            .lcout(\uart_rx_inst.n325 ),
            .ltout(),
            .carryin(\uart_rx_inst.n1532 ),
            .carryout(\uart_rx_inst.n1533 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.add_144_6_lut_LC_11_5_4 .C_ON=1'b1;
    defparam \uart_rx_inst.add_144_6_lut_LC_11_5_4 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.add_144_6_lut_LC_11_5_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_rx_inst.add_144_6_lut_LC_11_5_4  (
            .in0(_gnd_net_),
            .in1(N__8246),
            .in2(N__8770),
            .in3(N__6157),
            .lcout(\uart_rx_inst.n324 ),
            .ltout(),
            .carryin(\uart_rx_inst.n1533 ),
            .carryout(\uart_rx_inst.n1534 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.add_144_7_lut_LC_11_5_5 .C_ON=1'b1;
    defparam \uart_rx_inst.add_144_7_lut_LC_11_5_5 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.add_144_7_lut_LC_11_5_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_rx_inst.add_144_7_lut_LC_11_5_5  (
            .in0(_gnd_net_),
            .in1(N__8243),
            .in2(N__8669),
            .in3(N__6145),
            .lcout(\uart_rx_inst.n323 ),
            .ltout(),
            .carryin(\uart_rx_inst.n1534 ),
            .carryout(\uart_rx_inst.n1535 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.add_144_8_lut_LC_11_5_6 .C_ON=1'b1;
    defparam \uart_rx_inst.add_144_8_lut_LC_11_5_6 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.add_144_8_lut_LC_11_5_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_rx_inst.add_144_8_lut_LC_11_5_6  (
            .in0(_gnd_net_),
            .in1(N__8247),
            .in2(N__8566),
            .in3(N__6130),
            .lcout(\uart_rx_inst.n322 ),
            .ltout(),
            .carryin(\uart_rx_inst.n1535 ),
            .carryout(\uart_rx_inst.n1536 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.add_144_9_lut_LC_11_5_7 .C_ON=1'b1;
    defparam \uart_rx_inst.add_144_9_lut_LC_11_5_7 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.add_144_9_lut_LC_11_5_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_rx_inst.add_144_9_lut_LC_11_5_7  (
            .in0(_gnd_net_),
            .in1(N__8244),
            .in2(N__8463),
            .in3(N__6118),
            .lcout(\uart_rx_inst.n321 ),
            .ltout(),
            .carryin(\uart_rx_inst.n1536 ),
            .carryout(\uart_rx_inst.n1537 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.add_144_10_lut_LC_11_6_0 .C_ON=1'b1;
    defparam \uart_rx_inst.add_144_10_lut_LC_11_6_0 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.add_144_10_lut_LC_11_6_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_rx_inst.add_144_10_lut_LC_11_6_0  (
            .in0(_gnd_net_),
            .in1(N__8262),
            .in2(N__7972),
            .in3(N__6103),
            .lcout(\uart_rx_inst.n320 ),
            .ltout(),
            .carryin(bfn_11_6_0_),
            .carryout(\uart_rx_inst.n1538 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.add_144_11_lut_LC_11_6_1 .C_ON=1'b1;
    defparam \uart_rx_inst.add_144_11_lut_LC_11_6_1 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.add_144_11_lut_LC_11_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_rx_inst.add_144_11_lut_LC_11_6_1  (
            .in0(_gnd_net_),
            .in1(N__8328),
            .in2(N__7882),
            .in3(N__6088),
            .lcout(\uart_rx_inst.n319 ),
            .ltout(),
            .carryin(\uart_rx_inst.n1538 ),
            .carryout(\uart_rx_inst.n1539 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.add_144_12_lut_LC_11_6_2 .C_ON=1'b1;
    defparam \uart_rx_inst.add_144_12_lut_LC_11_6_2 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.add_144_12_lut_LC_11_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_rx_inst.add_144_12_lut_LC_11_6_2  (
            .in0(_gnd_net_),
            .in1(N__8263),
            .in2(N__7787),
            .in3(N__6073),
            .lcout(\uart_rx_inst.n318 ),
            .ltout(),
            .carryin(\uart_rx_inst.n1539 ),
            .carryout(\uart_rx_inst.n1540 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.add_144_13_lut_LC_11_6_3 .C_ON=1'b1;
    defparam \uart_rx_inst.add_144_13_lut_LC_11_6_3 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.add_144_13_lut_LC_11_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_rx_inst.add_144_13_lut_LC_11_6_3  (
            .in0(_gnd_net_),
            .in1(N__8329),
            .in2(N__8848),
            .in3(N__6400),
            .lcout(\uart_rx_inst.n317 ),
            .ltout(),
            .carryin(\uart_rx_inst.n1540 ),
            .carryout(\uart_rx_inst.n1541 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.add_144_14_lut_LC_11_6_4 .C_ON=1'b1;
    defparam \uart_rx_inst.add_144_14_lut_LC_11_6_4 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.add_144_14_lut_LC_11_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_rx_inst.add_144_14_lut_LC_11_6_4  (
            .in0(_gnd_net_),
            .in1(N__8264),
            .in2(N__8757),
            .in3(N__6385),
            .lcout(\uart_rx_inst.n316 ),
            .ltout(),
            .carryin(\uart_rx_inst.n1541 ),
            .carryout(\uart_rx_inst.n1542 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.add_144_15_lut_LC_11_6_5 .C_ON=1'b1;
    defparam \uart_rx_inst.add_144_15_lut_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.add_144_15_lut_LC_11_6_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_rx_inst.add_144_15_lut_LC_11_6_5  (
            .in0(_gnd_net_),
            .in1(N__8330),
            .in2(N__8663),
            .in3(N__6370),
            .lcout(\uart_rx_inst.n315 ),
            .ltout(),
            .carryin(\uart_rx_inst.n1542 ),
            .carryout(\uart_rx_inst.n1543 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.add_144_16_lut_LC_11_6_6 .C_ON=1'b1;
    defparam \uart_rx_inst.add_144_16_lut_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.add_144_16_lut_LC_11_6_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_rx_inst.add_144_16_lut_LC_11_6_6  (
            .in0(_gnd_net_),
            .in1(N__8265),
            .in2(N__8564),
            .in3(N__6355),
            .lcout(\uart_rx_inst.n314 ),
            .ltout(),
            .carryin(\uart_rx_inst.n1543 ),
            .carryout(\uart_rx_inst.n1544 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.add_144_17_lut_LC_11_6_7 .C_ON=1'b1;
    defparam \uart_rx_inst.add_144_17_lut_LC_11_6_7 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.add_144_17_lut_LC_11_6_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_rx_inst.add_144_17_lut_LC_11_6_7  (
            .in0(_gnd_net_),
            .in1(N__8331),
            .in2(N__8453),
            .in3(N__6340),
            .lcout(\uart_rx_inst.n313 ),
            .ltout(),
            .carryin(\uart_rx_inst.n1544 ),
            .carryout(\uart_rx_inst.n1545 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.add_144_18_lut_LC_11_7_0 .C_ON=1'b0;
    defparam \uart_rx_inst.add_144_18_lut_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.add_144_18_lut_LC_11_7_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_rx_inst.add_144_18_lut_LC_11_7_0  (
            .in0(_gnd_net_),
            .in1(N__8169),
            .in2(_gnd_net_),
            .in3(N__6337),
            .lcout(\uart_rx_inst.n312 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx_inst.i1573_2_lut_LC_11_8_1 .C_ON=1'b0;
    defparam \uart_rx_inst.i1573_2_lut_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \uart_rx_inst.i1573_2_lut_LC_11_8_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_rx_inst.i1573_2_lut_LC_11_8_1  (
            .in0(_gnd_net_),
            .in1(N__7809),
            .in2(_gnd_net_),
            .in3(N__6314),
            .lcout(\uart_rx_inst.n1746 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.i13_4_lut_LC_12_1_0 .C_ON=1'b0;
    defparam \uart_tx_inst.i13_4_lut_LC_12_1_0 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.i13_4_lut_LC_12_1_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \uart_tx_inst.i13_4_lut_LC_12_1_0  (
            .in0(N__6873),
            .in1(N__6207),
            .in2(N__6498),
            .in3(N__6849),
            .lcout(\uart_tx_inst.n32_adj_197 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.i737_3_lut_LC_12_1_1 .C_ON=1'b0;
    defparam \uart_tx_inst.i737_3_lut_LC_12_1_1 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.i737_3_lut_LC_12_1_1 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \uart_tx_inst.i737_3_lut_LC_12_1_1  (
            .in0(_gnd_net_),
            .in1(N__6187),
            .in2(N__6832),
            .in3(N__6930),
            .lcout(),
            .ltout(\uart_tx_inst.n865_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.prescale_reg__i4_LC_12_1_2 .C_ON=1'b0;
    defparam \uart_tx_inst.prescale_reg__i4_LC_12_1_2 .SEQ_MODE=4'b1000;
    defparam \uart_tx_inst.prescale_reg__i4_LC_12_1_2 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \uart_tx_inst.prescale_reg__i4_LC_12_1_2  (
            .in0(N__7877),
            .in1(N__6597),
            .in2(N__6880),
            .in3(N__6725),
            .lcout(\uart_tx_inst.prescale_reg_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7384),
            .ce(N__6475),
            .sr(N__7227));
    defparam \uart_tx_inst.i742_3_lut_LC_12_1_4 .C_ON=1'b0;
    defparam \uart_tx_inst.i742_3_lut_LC_12_1_4 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.i742_3_lut_LC_12_1_4 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \uart_tx_inst.i742_3_lut_LC_12_1_4  (
            .in0(_gnd_net_),
            .in1(N__6811),
            .in2(N__6862),
            .in3(N__6897),
            .lcout(),
            .ltout(\uart_tx_inst.n870_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.prescale_reg__i5_LC_12_1_5 .C_ON=1'b0;
    defparam \uart_tx_inst.prescale_reg__i5_LC_12_1_5 .SEQ_MODE=4'b1000;
    defparam \uart_tx_inst.prescale_reg__i5_LC_12_1_5 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \uart_tx_inst.prescale_reg__i5_LC_12_1_5  (
            .in0(N__6726),
            .in1(N__7788),
            .in2(N__6853),
            .in3(N__6603),
            .lcout(\uart_tx_inst.prescale_reg_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7384),
            .ce(N__6475),
            .sr(N__7227));
    defparam \uart_tx_inst.i757_3_lut_LC_12_1_6 .C_ON=1'b0;
    defparam \uart_tx_inst.i757_3_lut_LC_12_1_6 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.i757_3_lut_LC_12_1_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \uart_tx_inst.i757_3_lut_LC_12_1_6  (
            .in0(N__8055),
            .in1(N__6812),
            .in2(_gnd_net_),
            .in3(N__6736),
            .lcout(),
            .ltout(\uart_tx_inst.n885_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.prescale_reg__i8_LC_12_1_7 .C_ON=1'b0;
    defparam \uart_tx_inst.prescale_reg__i8_LC_12_1_7 .SEQ_MODE=4'b1000;
    defparam \uart_tx_inst.prescale_reg__i8_LC_12_1_7 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \uart_tx_inst.prescale_reg__i8_LC_12_1_7  (
            .in0(N__6727),
            .in1(N__8667),
            .in2(N__6607),
            .in3(N__6604),
            .lcout(\uart_tx_inst.prescale_reg_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7384),
            .ce(N__6475),
            .sr(N__7227));
    defparam \uart_tx_inst.data_reg_i0_i0_LC_12_2_0 .C_ON=1'b0;
    defparam \uart_tx_inst.data_reg_i0_i0_LC_12_2_0 .SEQ_MODE=4'b1000;
    defparam \uart_tx_inst.data_reg_i0_i0_LC_12_2_0 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \uart_tx_inst.data_reg_i0_i0_LC_12_2_0  (
            .in0(N__7650),
            .in1(N__6424),
            .in2(N__7939),
            .in3(N__7520),
            .lcout(\uart_tx_inst.data_reg_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7383),
            .ce(N__7546),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.data_reg_i0_i1_LC_12_2_1 .C_ON=1'b0;
    defparam \uart_tx_inst.data_reg_i0_i1_LC_12_2_1 .SEQ_MODE=4'b1000;
    defparam \uart_tx_inst.data_reg_i0_i1_LC_12_2_1 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \uart_tx_inst.data_reg_i0_i1_LC_12_2_1  (
            .in0(N__7521),
            .in1(N__7651),
            .in2(N__7884),
            .in3(N__6418),
            .lcout(\uart_tx_inst.data_reg_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7383),
            .ce(N__7546),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.data_reg_i0_i2_LC_12_2_2 .C_ON=1'b0;
    defparam \uart_tx_inst.data_reg_i0_i2_LC_12_2_2 .SEQ_MODE=4'b1000;
    defparam \uart_tx_inst.data_reg_i0_i2_LC_12_2_2 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \uart_tx_inst.data_reg_i0_i2_LC_12_2_2  (
            .in0(N__7652),
            .in1(N__7687),
            .in2(N__7789),
            .in3(N__7522),
            .lcout(\uart_tx_inst.data_reg_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7383),
            .ce(N__7546),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.data_reg_i0_i3_LC_12_2_3 .C_ON=1'b0;
    defparam \uart_tx_inst.data_reg_i0_i3_LC_12_2_3 .SEQ_MODE=4'b1000;
    defparam \uart_tx_inst.data_reg_i0_i3_LC_12_2_3 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \uart_tx_inst.data_reg_i0_i3_LC_12_2_3  (
            .in0(N__7523),
            .in1(N__7653),
            .in2(N__8867),
            .in3(N__7681),
            .lcout(\uart_tx_inst.data_reg_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7383),
            .ce(N__7546),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.data_reg_i0_i4_LC_12_2_4 .C_ON=1'b0;
    defparam \uart_tx_inst.data_reg_i0_i4_LC_12_2_4 .SEQ_MODE=4'b1000;
    defparam \uart_tx_inst.data_reg_i0_i4_LC_12_2_4 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_tx_inst.data_reg_i0_i4_LC_12_2_4  (
            .in0(N__7654),
            .in1(N__8771),
            .in2(N__7675),
            .in3(N__7524),
            .lcout(\uart_tx_inst.data_reg_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7383),
            .ce(N__7546),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.data_reg_i0_i5_LC_12_2_5 .C_ON=1'b0;
    defparam \uart_tx_inst.data_reg_i0_i5_LC_12_2_5 .SEQ_MODE=4'b1000;
    defparam \uart_tx_inst.data_reg_i0_i5_LC_12_2_5 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \uart_tx_inst.data_reg_i0_i5_LC_12_2_5  (
            .in0(N__7525),
            .in1(N__7655),
            .in2(N__8673),
            .in3(N__7666),
            .lcout(\uart_tx_inst.data_reg_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7383),
            .ce(N__7546),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.data_reg_i0_i6_LC_12_2_6 .C_ON=1'b0;
    defparam \uart_tx_inst.data_reg_i0_i6_LC_12_2_6 .SEQ_MODE=4'b1000;
    defparam \uart_tx_inst.data_reg_i0_i6_LC_12_2_6 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \uart_tx_inst.data_reg_i0_i6_LC_12_2_6  (
            .in0(N__7656),
            .in1(N__7552),
            .in2(N__8572),
            .in3(N__7526),
            .lcout(\uart_tx_inst.data_reg_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7383),
            .ce(N__7546),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.data_reg_i0_i7_LC_12_2_7 .C_ON=1'b0;
    defparam \uart_tx_inst.data_reg_i0_i7_LC_12_2_7 .SEQ_MODE=4'b1000;
    defparam \uart_tx_inst.data_reg_i0_i7_LC_12_2_7 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \uart_tx_inst.data_reg_i0_i7_LC_12_2_7  (
            .in0(N__7527),
            .in1(N__7657),
            .in2(N__8458),
            .in3(N__7570),
            .lcout(\uart_tx_inst.data_reg_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7383),
            .ce(N__7546),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.txd_reg_50_LC_12_3_0 .C_ON=1'b0;
    defparam \uart_tx_inst.txd_reg_50_LC_12_3_0 .SEQ_MODE=4'b1001;
    defparam \uart_tx_inst.txd_reg_50_LC_12_3_0 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \uart_tx_inst.txd_reg_50_LC_12_3_0  (
            .in0(N__7534),
            .in1(N__7528),
            .in2(_gnd_net_),
            .in3(N__7441),
            .lcout(txd_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7381),
            .ce(N__7279),
            .sr(N__7262));
    defparam \uart_tx_inst.sub_8_add_2_2_lut_LC_12_5_0 .C_ON=1'b1;
    defparam \uart_tx_inst.sub_8_add_2_2_lut_LC_12_5_0 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.sub_8_add_2_2_lut_LC_12_5_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_tx_inst.sub_8_add_2_2_lut_LC_12_5_0  (
            .in0(_gnd_net_),
            .in1(N__7958),
            .in2(_gnd_net_),
            .in3(N__6937),
            .lcout(n108),
            .ltout(),
            .carryin(bfn_12_5_0_),
            .carryout(\uart_tx_inst.n1582 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.sub_8_add_2_3_lut_LC_12_5_1 .C_ON=1'b1;
    defparam \uart_tx_inst.sub_8_add_2_3_lut_LC_12_5_1 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.sub_8_add_2_3_lut_LC_12_5_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_tx_inst.sub_8_add_2_3_lut_LC_12_5_1  (
            .in0(_gnd_net_),
            .in1(N__8255),
            .in2(N__7846),
            .in3(N__6907),
            .lcout(n107),
            .ltout(),
            .carryin(\uart_tx_inst.n1582 ),
            .carryout(\uart_tx_inst.n1583 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.sub_8_add_2_4_lut_LC_12_5_2 .C_ON=1'b1;
    defparam \uart_tx_inst.sub_8_add_2_4_lut_LC_12_5_2 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.sub_8_add_2_4_lut_LC_12_5_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_tx_inst.sub_8_add_2_4_lut_LC_12_5_2  (
            .in0(_gnd_net_),
            .in1(N__8259),
            .in2(N__7750),
            .in3(N__8110),
            .lcout(n106),
            .ltout(),
            .carryin(\uart_tx_inst.n1583 ),
            .carryout(\uart_tx_inst.n1584 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.sub_8_add_2_5_lut_LC_12_5_3 .C_ON=1'b1;
    defparam \uart_tx_inst.sub_8_add_2_5_lut_LC_12_5_3 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.sub_8_add_2_5_lut_LC_12_5_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_tx_inst.sub_8_add_2_5_lut_LC_12_5_3  (
            .in0(_gnd_net_),
            .in1(N__8256),
            .in2(N__8847),
            .in3(N__8083),
            .lcout(n105),
            .ltout(),
            .carryin(\uart_tx_inst.n1584 ),
            .carryout(\uart_tx_inst.n1585 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.sub_8_add_2_6_lut_LC_12_5_4 .C_ON=1'b1;
    defparam \uart_tx_inst.sub_8_add_2_6_lut_LC_12_5_4 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.sub_8_add_2_6_lut_LC_12_5_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_tx_inst.sub_8_add_2_6_lut_LC_12_5_4  (
            .in0(_gnd_net_),
            .in1(N__8260),
            .in2(N__8753),
            .in3(N__8059),
            .lcout(n104),
            .ltout(),
            .carryin(\uart_tx_inst.n1585 ),
            .carryout(\uart_tx_inst.n1586 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.sub_8_add_2_7_lut_LC_12_5_5 .C_ON=1'b1;
    defparam \uart_tx_inst.sub_8_add_2_7_lut_LC_12_5_5 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.sub_8_add_2_7_lut_LC_12_5_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_tx_inst.sub_8_add_2_7_lut_LC_12_5_5  (
            .in0(_gnd_net_),
            .in1(N__8257),
            .in2(N__8668),
            .in3(N__8032),
            .lcout(n103),
            .ltout(),
            .carryin(\uart_tx_inst.n1586 ),
            .carryout(\uart_tx_inst.n1587 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.sub_8_add_2_8_lut_LC_12_5_6 .C_ON=1'b1;
    defparam \uart_tx_inst.sub_8_add_2_8_lut_LC_12_5_6 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.sub_8_add_2_8_lut_LC_12_5_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_tx_inst.sub_8_add_2_8_lut_LC_12_5_6  (
            .in0(_gnd_net_),
            .in1(N__8261),
            .in2(N__8565),
            .in3(N__8005),
            .lcout(n102),
            .ltout(),
            .carryin(\uart_tx_inst.n1587 ),
            .carryout(\uart_tx_inst.n1588 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.sub_8_add_2_9_lut_LC_12_5_7 .C_ON=1'b1;
    defparam \uart_tx_inst.sub_8_add_2_9_lut_LC_12_5_7 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.sub_8_add_2_9_lut_LC_12_5_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_tx_inst.sub_8_add_2_9_lut_LC_12_5_7  (
            .in0(_gnd_net_),
            .in1(N__8258),
            .in2(N__8454),
            .in3(N__7975),
            .lcout(n101),
            .ltout(),
            .carryin(\uart_tx_inst.n1588 ),
            .carryout(\uart_tx_inst.n1589 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.sub_8_add_2_10_lut_LC_12_6_0 .C_ON=1'b1;
    defparam \uart_tx_inst.sub_8_add_2_10_lut_LC_12_6_0 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.sub_8_add_2_10_lut_LC_12_6_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_tx_inst.sub_8_add_2_10_lut_LC_12_6_0  (
            .in0(_gnd_net_),
            .in1(N__8332),
            .in2(N__7971),
            .in3(N__7888),
            .lcout(n100),
            .ltout(),
            .carryin(bfn_12_6_0_),
            .carryout(\uart_tx_inst.n1590 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.sub_8_add_2_11_lut_LC_12_6_1 .C_ON=1'b1;
    defparam \uart_tx_inst.sub_8_add_2_11_lut_LC_12_6_1 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.sub_8_add_2_11_lut_LC_12_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_tx_inst.sub_8_add_2_11_lut_LC_12_6_1  (
            .in0(_gnd_net_),
            .in1(N__8266),
            .in2(N__7885),
            .in3(N__7792),
            .lcout(n99),
            .ltout(),
            .carryin(\uart_tx_inst.n1590 ),
            .carryout(\uart_tx_inst.n1591 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.sub_8_add_2_12_lut_LC_12_6_2 .C_ON=1'b1;
    defparam \uart_tx_inst.sub_8_add_2_12_lut_LC_12_6_2 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.sub_8_add_2_12_lut_LC_12_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_tx_inst.sub_8_add_2_12_lut_LC_12_6_2  (
            .in0(_gnd_net_),
            .in1(N__8333),
            .in2(N__7786),
            .in3(N__7690),
            .lcout(n98),
            .ltout(),
            .carryin(\uart_tx_inst.n1591 ),
            .carryout(\uart_tx_inst.n1592 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.sub_8_add_2_13_lut_LC_12_6_3 .C_ON=1'b1;
    defparam \uart_tx_inst.sub_8_add_2_13_lut_LC_12_6_3 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.sub_8_add_2_13_lut_LC_12_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_tx_inst.sub_8_add_2_13_lut_LC_12_6_3  (
            .in0(_gnd_net_),
            .in1(N__8267),
            .in2(N__8835),
            .in3(N__8779),
            .lcout(n97),
            .ltout(),
            .carryin(\uart_tx_inst.n1592 ),
            .carryout(\uart_tx_inst.n1593 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.sub_8_add_2_14_lut_LC_12_6_4 .C_ON=1'b1;
    defparam \uart_tx_inst.sub_8_add_2_14_lut_LC_12_6_4 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.sub_8_add_2_14_lut_LC_12_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_tx_inst.sub_8_add_2_14_lut_LC_12_6_4  (
            .in0(_gnd_net_),
            .in1(N__8334),
            .in2(N__8741),
            .in3(N__8677),
            .lcout(n96),
            .ltout(),
            .carryin(\uart_tx_inst.n1593 ),
            .carryout(\uart_tx_inst.n1594 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.sub_8_add_2_15_lut_LC_12_6_5 .C_ON=1'b1;
    defparam \uart_tx_inst.sub_8_add_2_15_lut_LC_12_6_5 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.sub_8_add_2_15_lut_LC_12_6_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_tx_inst.sub_8_add_2_15_lut_LC_12_6_5  (
            .in0(_gnd_net_),
            .in1(N__8268),
            .in2(N__8626),
            .in3(N__8575),
            .lcout(n95),
            .ltout(),
            .carryin(\uart_tx_inst.n1594 ),
            .carryout(\uart_tx_inst.n1595 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.sub_8_add_2_16_lut_LC_12_6_6 .C_ON=1'b1;
    defparam \uart_tx_inst.sub_8_add_2_16_lut_LC_12_6_6 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.sub_8_add_2_16_lut_LC_12_6_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_tx_inst.sub_8_add_2_16_lut_LC_12_6_6  (
            .in0(_gnd_net_),
            .in1(N__8335),
            .in2(N__8528),
            .in3(N__8467),
            .lcout(n94),
            .ltout(),
            .carryin(\uart_tx_inst.n1595 ),
            .carryout(\uart_tx_inst.n1596 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx_inst.sub_8_add_2_17_lut_LC_12_6_7 .C_ON=1'b0;
    defparam \uart_tx_inst.sub_8_add_2_17_lut_LC_12_6_7 .SEQ_MODE=4'b0000;
    defparam \uart_tx_inst.sub_8_add_2_17_lut_LC_12_6_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_tx_inst.sub_8_add_2_17_lut_LC_12_6_7  (
            .in0(N__8434),
            .in1(N__8269),
            .in2(_gnd_net_),
            .in3(N__8134),
            .lcout(n93),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // uart
