// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 12 2017 08:25:46

// File Generated:     Jan 24 2019 13:59:16

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "big_counter" view "INTERFACE"

module big_counter (
    rco,
    en_in,
    clk);

    output [199:0] rco;
    input en_in;
    input clk;

    wire N__95452;
    wire N__95451;
    wire N__95450;
    wire N__95441;
    wire N__95440;
    wire N__95439;
    wire N__95432;
    wire N__95431;
    wire N__95430;
    wire N__95423;
    wire N__95422;
    wire N__95421;
    wire N__95414;
    wire N__95413;
    wire N__95412;
    wire N__95405;
    wire N__95404;
    wire N__95403;
    wire N__95396;
    wire N__95395;
    wire N__95394;
    wire N__95387;
    wire N__95386;
    wire N__95385;
    wire N__95378;
    wire N__95377;
    wire N__95376;
    wire N__95369;
    wire N__95368;
    wire N__95367;
    wire N__95360;
    wire N__95359;
    wire N__95358;
    wire N__95351;
    wire N__95350;
    wire N__95349;
    wire N__95342;
    wire N__95341;
    wire N__95340;
    wire N__95333;
    wire N__95332;
    wire N__95331;
    wire N__95324;
    wire N__95323;
    wire N__95322;
    wire N__95315;
    wire N__95314;
    wire N__95313;
    wire N__95306;
    wire N__95305;
    wire N__95304;
    wire N__95297;
    wire N__95296;
    wire N__95295;
    wire N__95288;
    wire N__95287;
    wire N__95286;
    wire N__95279;
    wire N__95278;
    wire N__95277;
    wire N__95270;
    wire N__95269;
    wire N__95268;
    wire N__95261;
    wire N__95260;
    wire N__95259;
    wire N__95252;
    wire N__95251;
    wire N__95250;
    wire N__95243;
    wire N__95242;
    wire N__95241;
    wire N__95234;
    wire N__95233;
    wire N__95232;
    wire N__95225;
    wire N__95224;
    wire N__95223;
    wire N__95216;
    wire N__95215;
    wire N__95214;
    wire N__95207;
    wire N__95206;
    wire N__95205;
    wire N__95198;
    wire N__95197;
    wire N__95196;
    wire N__95189;
    wire N__95188;
    wire N__95187;
    wire N__95180;
    wire N__95179;
    wire N__95178;
    wire N__95171;
    wire N__95170;
    wire N__95169;
    wire N__95162;
    wire N__95161;
    wire N__95160;
    wire N__95153;
    wire N__95152;
    wire N__95151;
    wire N__95144;
    wire N__95143;
    wire N__95142;
    wire N__95135;
    wire N__95134;
    wire N__95133;
    wire N__95126;
    wire N__95125;
    wire N__95124;
    wire N__95117;
    wire N__95116;
    wire N__95115;
    wire N__95108;
    wire N__95107;
    wire N__95106;
    wire N__95099;
    wire N__95098;
    wire N__95097;
    wire N__95090;
    wire N__95089;
    wire N__95088;
    wire N__95081;
    wire N__95080;
    wire N__95079;
    wire N__95072;
    wire N__95071;
    wire N__95070;
    wire N__95063;
    wire N__95062;
    wire N__95061;
    wire N__95054;
    wire N__95053;
    wire N__95052;
    wire N__95045;
    wire N__95044;
    wire N__95043;
    wire N__95036;
    wire N__95035;
    wire N__95034;
    wire N__95027;
    wire N__95026;
    wire N__95025;
    wire N__95018;
    wire N__95017;
    wire N__95016;
    wire N__95009;
    wire N__95008;
    wire N__95007;
    wire N__95000;
    wire N__94999;
    wire N__94998;
    wire N__94991;
    wire N__94990;
    wire N__94989;
    wire N__94982;
    wire N__94981;
    wire N__94980;
    wire N__94973;
    wire N__94972;
    wire N__94971;
    wire N__94964;
    wire N__94963;
    wire N__94962;
    wire N__94955;
    wire N__94954;
    wire N__94953;
    wire N__94946;
    wire N__94945;
    wire N__94944;
    wire N__94937;
    wire N__94936;
    wire N__94935;
    wire N__94928;
    wire N__94927;
    wire N__94926;
    wire N__94919;
    wire N__94918;
    wire N__94917;
    wire N__94910;
    wire N__94909;
    wire N__94908;
    wire N__94901;
    wire N__94900;
    wire N__94899;
    wire N__94892;
    wire N__94891;
    wire N__94890;
    wire N__94883;
    wire N__94882;
    wire N__94881;
    wire N__94874;
    wire N__94873;
    wire N__94872;
    wire N__94865;
    wire N__94864;
    wire N__94863;
    wire N__94856;
    wire N__94855;
    wire N__94854;
    wire N__94847;
    wire N__94846;
    wire N__94845;
    wire N__94838;
    wire N__94837;
    wire N__94836;
    wire N__94829;
    wire N__94828;
    wire N__94827;
    wire N__94820;
    wire N__94819;
    wire N__94818;
    wire N__94811;
    wire N__94810;
    wire N__94809;
    wire N__94802;
    wire N__94801;
    wire N__94800;
    wire N__94793;
    wire N__94792;
    wire N__94791;
    wire N__94784;
    wire N__94783;
    wire N__94782;
    wire N__94775;
    wire N__94774;
    wire N__94773;
    wire N__94766;
    wire N__94765;
    wire N__94764;
    wire N__94757;
    wire N__94756;
    wire N__94755;
    wire N__94748;
    wire N__94747;
    wire N__94746;
    wire N__94739;
    wire N__94738;
    wire N__94737;
    wire N__94730;
    wire N__94729;
    wire N__94728;
    wire N__94721;
    wire N__94720;
    wire N__94719;
    wire N__94712;
    wire N__94711;
    wire N__94710;
    wire N__94703;
    wire N__94702;
    wire N__94701;
    wire N__94694;
    wire N__94693;
    wire N__94692;
    wire N__94685;
    wire N__94684;
    wire N__94683;
    wire N__94676;
    wire N__94675;
    wire N__94674;
    wire N__94667;
    wire N__94666;
    wire N__94665;
    wire N__94658;
    wire N__94657;
    wire N__94656;
    wire N__94649;
    wire N__94648;
    wire N__94647;
    wire N__94640;
    wire N__94639;
    wire N__94638;
    wire N__94631;
    wire N__94630;
    wire N__94629;
    wire N__94622;
    wire N__94621;
    wire N__94620;
    wire N__94613;
    wire N__94612;
    wire N__94611;
    wire N__94604;
    wire N__94603;
    wire N__94602;
    wire N__94595;
    wire N__94594;
    wire N__94593;
    wire N__94586;
    wire N__94585;
    wire N__94584;
    wire N__94577;
    wire N__94576;
    wire N__94575;
    wire N__94568;
    wire N__94567;
    wire N__94566;
    wire N__94559;
    wire N__94558;
    wire N__94557;
    wire N__94550;
    wire N__94549;
    wire N__94548;
    wire N__94541;
    wire N__94540;
    wire N__94539;
    wire N__94532;
    wire N__94531;
    wire N__94530;
    wire N__94523;
    wire N__94522;
    wire N__94521;
    wire N__94514;
    wire N__94513;
    wire N__94512;
    wire N__94505;
    wire N__94504;
    wire N__94503;
    wire N__94496;
    wire N__94495;
    wire N__94494;
    wire N__94487;
    wire N__94486;
    wire N__94485;
    wire N__94478;
    wire N__94477;
    wire N__94476;
    wire N__94469;
    wire N__94468;
    wire N__94467;
    wire N__94460;
    wire N__94459;
    wire N__94458;
    wire N__94451;
    wire N__94450;
    wire N__94449;
    wire N__94442;
    wire N__94441;
    wire N__94440;
    wire N__94433;
    wire N__94432;
    wire N__94431;
    wire N__94424;
    wire N__94423;
    wire N__94422;
    wire N__94415;
    wire N__94414;
    wire N__94413;
    wire N__94406;
    wire N__94405;
    wire N__94404;
    wire N__94397;
    wire N__94396;
    wire N__94395;
    wire N__94388;
    wire N__94387;
    wire N__94386;
    wire N__94379;
    wire N__94378;
    wire N__94377;
    wire N__94370;
    wire N__94369;
    wire N__94368;
    wire N__94361;
    wire N__94360;
    wire N__94359;
    wire N__94352;
    wire N__94351;
    wire N__94350;
    wire N__94343;
    wire N__94342;
    wire N__94341;
    wire N__94334;
    wire N__94333;
    wire N__94332;
    wire N__94325;
    wire N__94324;
    wire N__94323;
    wire N__94316;
    wire N__94315;
    wire N__94314;
    wire N__94307;
    wire N__94306;
    wire N__94305;
    wire N__94298;
    wire N__94297;
    wire N__94296;
    wire N__94289;
    wire N__94288;
    wire N__94287;
    wire N__94280;
    wire N__94279;
    wire N__94278;
    wire N__94271;
    wire N__94270;
    wire N__94269;
    wire N__94262;
    wire N__94261;
    wire N__94260;
    wire N__94253;
    wire N__94252;
    wire N__94251;
    wire N__94244;
    wire N__94243;
    wire N__94242;
    wire N__94235;
    wire N__94234;
    wire N__94233;
    wire N__94226;
    wire N__94225;
    wire N__94224;
    wire N__94217;
    wire N__94216;
    wire N__94215;
    wire N__94208;
    wire N__94207;
    wire N__94206;
    wire N__94199;
    wire N__94198;
    wire N__94197;
    wire N__94190;
    wire N__94189;
    wire N__94188;
    wire N__94181;
    wire N__94180;
    wire N__94179;
    wire N__94172;
    wire N__94171;
    wire N__94170;
    wire N__94163;
    wire N__94162;
    wire N__94161;
    wire N__94154;
    wire N__94153;
    wire N__94152;
    wire N__94145;
    wire N__94144;
    wire N__94143;
    wire N__94136;
    wire N__94135;
    wire N__94134;
    wire N__94127;
    wire N__94126;
    wire N__94125;
    wire N__94118;
    wire N__94117;
    wire N__94116;
    wire N__94109;
    wire N__94108;
    wire N__94107;
    wire N__94100;
    wire N__94099;
    wire N__94098;
    wire N__94091;
    wire N__94090;
    wire N__94089;
    wire N__94082;
    wire N__94081;
    wire N__94080;
    wire N__94073;
    wire N__94072;
    wire N__94071;
    wire N__94064;
    wire N__94063;
    wire N__94062;
    wire N__94055;
    wire N__94054;
    wire N__94053;
    wire N__94046;
    wire N__94045;
    wire N__94044;
    wire N__94037;
    wire N__94036;
    wire N__94035;
    wire N__94028;
    wire N__94027;
    wire N__94026;
    wire N__94019;
    wire N__94018;
    wire N__94017;
    wire N__94010;
    wire N__94009;
    wire N__94008;
    wire N__94001;
    wire N__94000;
    wire N__93999;
    wire N__93992;
    wire N__93991;
    wire N__93990;
    wire N__93983;
    wire N__93982;
    wire N__93981;
    wire N__93974;
    wire N__93973;
    wire N__93972;
    wire N__93965;
    wire N__93964;
    wire N__93963;
    wire N__93956;
    wire N__93955;
    wire N__93954;
    wire N__93947;
    wire N__93946;
    wire N__93945;
    wire N__93938;
    wire N__93937;
    wire N__93936;
    wire N__93929;
    wire N__93928;
    wire N__93927;
    wire N__93920;
    wire N__93919;
    wire N__93918;
    wire N__93911;
    wire N__93910;
    wire N__93909;
    wire N__93902;
    wire N__93901;
    wire N__93900;
    wire N__93893;
    wire N__93892;
    wire N__93891;
    wire N__93884;
    wire N__93883;
    wire N__93882;
    wire N__93875;
    wire N__93874;
    wire N__93873;
    wire N__93866;
    wire N__93865;
    wire N__93864;
    wire N__93857;
    wire N__93856;
    wire N__93855;
    wire N__93848;
    wire N__93847;
    wire N__93846;
    wire N__93839;
    wire N__93838;
    wire N__93837;
    wire N__93830;
    wire N__93829;
    wire N__93828;
    wire N__93821;
    wire N__93820;
    wire N__93819;
    wire N__93812;
    wire N__93811;
    wire N__93810;
    wire N__93803;
    wire N__93802;
    wire N__93801;
    wire N__93794;
    wire N__93793;
    wire N__93792;
    wire N__93785;
    wire N__93784;
    wire N__93783;
    wire N__93776;
    wire N__93775;
    wire N__93774;
    wire N__93767;
    wire N__93766;
    wire N__93765;
    wire N__93758;
    wire N__93757;
    wire N__93756;
    wire N__93749;
    wire N__93748;
    wire N__93747;
    wire N__93740;
    wire N__93739;
    wire N__93738;
    wire N__93731;
    wire N__93730;
    wire N__93729;
    wire N__93722;
    wire N__93721;
    wire N__93720;
    wire N__93713;
    wire N__93712;
    wire N__93711;
    wire N__93704;
    wire N__93703;
    wire N__93702;
    wire N__93695;
    wire N__93694;
    wire N__93693;
    wire N__93686;
    wire N__93685;
    wire N__93684;
    wire N__93677;
    wire N__93676;
    wire N__93675;
    wire N__93668;
    wire N__93667;
    wire N__93666;
    wire N__93659;
    wire N__93658;
    wire N__93657;
    wire N__93650;
    wire N__93649;
    wire N__93648;
    wire N__93641;
    wire N__93640;
    wire N__93639;
    wire N__93622;
    wire N__93619;
    wire N__93616;
    wire N__93615;
    wire N__93612;
    wire N__93609;
    wire N__93604;
    wire N__93603;
    wire N__93600;
    wire N__93597;
    wire N__93596;
    wire N__93595;
    wire N__93594;
    wire N__93593;
    wire N__93588;
    wire N__93587;
    wire N__93584;
    wire N__93577;
    wire N__93576;
    wire N__93573;
    wire N__93570;
    wire N__93567;
    wire N__93566;
    wire N__93565;
    wire N__93564;
    wire N__93561;
    wire N__93558;
    wire N__93557;
    wire N__93556;
    wire N__93555;
    wire N__93554;
    wire N__93553;
    wire N__93552;
    wire N__93549;
    wire N__93544;
    wire N__93541;
    wire N__93538;
    wire N__93535;
    wire N__93532;
    wire N__93521;
    wire N__93516;
    wire N__93499;
    wire N__93496;
    wire N__93495;
    wire N__93492;
    wire N__93491;
    wire N__93488;
    wire N__93485;
    wire N__93482;
    wire N__93479;
    wire N__93478;
    wire N__93477;
    wire N__93474;
    wire N__93471;
    wire N__93468;
    wire N__93465;
    wire N__93462;
    wire N__93451;
    wire N__93448;
    wire N__93445;
    wire N__93442;
    wire N__93439;
    wire N__93436;
    wire N__93433;
    wire N__93430;
    wire N__93427;
    wire N__93426;
    wire N__93425;
    wire N__93424;
    wire N__93423;
    wire N__93422;
    wire N__93421;
    wire N__93420;
    wire N__93419;
    wire N__93418;
    wire N__93417;
    wire N__93416;
    wire N__93415;
    wire N__93414;
    wire N__93413;
    wire N__93412;
    wire N__93411;
    wire N__93410;
    wire N__93409;
    wire N__93408;
    wire N__93407;
    wire N__93406;
    wire N__93405;
    wire N__93404;
    wire N__93403;
    wire N__93402;
    wire N__93401;
    wire N__93400;
    wire N__93399;
    wire N__93398;
    wire N__93397;
    wire N__93396;
    wire N__93395;
    wire N__93394;
    wire N__93393;
    wire N__93392;
    wire N__93391;
    wire N__93390;
    wire N__93389;
    wire N__93388;
    wire N__93387;
    wire N__93386;
    wire N__93385;
    wire N__93384;
    wire N__93383;
    wire N__93382;
    wire N__93381;
    wire N__93380;
    wire N__93379;
    wire N__93378;
    wire N__93377;
    wire N__93376;
    wire N__93375;
    wire N__93374;
    wire N__93373;
    wire N__93372;
    wire N__93371;
    wire N__93370;
    wire N__93369;
    wire N__93368;
    wire N__93367;
    wire N__93366;
    wire N__93365;
    wire N__93364;
    wire N__93363;
    wire N__93362;
    wire N__93361;
    wire N__93360;
    wire N__93359;
    wire N__93358;
    wire N__93357;
    wire N__93356;
    wire N__93355;
    wire N__93354;
    wire N__93353;
    wire N__93352;
    wire N__93351;
    wire N__93350;
    wire N__93349;
    wire N__93348;
    wire N__93347;
    wire N__93346;
    wire N__93345;
    wire N__93344;
    wire N__93343;
    wire N__93342;
    wire N__93341;
    wire N__93340;
    wire N__93339;
    wire N__93338;
    wire N__93337;
    wire N__93336;
    wire N__93335;
    wire N__93334;
    wire N__93333;
    wire N__93332;
    wire N__93331;
    wire N__93330;
    wire N__93329;
    wire N__93328;
    wire N__93327;
    wire N__93326;
    wire N__93325;
    wire N__93324;
    wire N__93323;
    wire N__93322;
    wire N__93321;
    wire N__93320;
    wire N__93319;
    wire N__93318;
    wire N__93317;
    wire N__93316;
    wire N__93315;
    wire N__93314;
    wire N__93313;
    wire N__93312;
    wire N__93311;
    wire N__93310;
    wire N__93309;
    wire N__93308;
    wire N__93307;
    wire N__93306;
    wire N__93305;
    wire N__93304;
    wire N__93303;
    wire N__93302;
    wire N__93301;
    wire N__93300;
    wire N__93299;
    wire N__93298;
    wire N__93297;
    wire N__93296;
    wire N__93295;
    wire N__93294;
    wire N__93293;
    wire N__93292;
    wire N__93291;
    wire N__93290;
    wire N__93289;
    wire N__93288;
    wire N__93287;
    wire N__93286;
    wire N__93285;
    wire N__93284;
    wire N__93283;
    wire N__93282;
    wire N__93281;
    wire N__93280;
    wire N__93279;
    wire N__93278;
    wire N__93277;
    wire N__93276;
    wire N__93275;
    wire N__93274;
    wire N__93273;
    wire N__93272;
    wire N__93271;
    wire N__93270;
    wire N__93269;
    wire N__93268;
    wire N__93267;
    wire N__93266;
    wire N__93265;
    wire N__93264;
    wire N__93263;
    wire N__93262;
    wire N__93261;
    wire N__93260;
    wire N__93259;
    wire N__93258;
    wire N__93257;
    wire N__93256;
    wire N__93255;
    wire N__93254;
    wire N__93253;
    wire N__93252;
    wire N__93251;
    wire N__93250;
    wire N__93249;
    wire N__93248;
    wire N__93247;
    wire N__93246;
    wire N__93245;
    wire N__93244;
    wire N__93243;
    wire N__93242;
    wire N__93241;
    wire N__93240;
    wire N__93239;
    wire N__93238;
    wire N__93237;
    wire N__93236;
    wire N__93235;
    wire N__93234;
    wire N__93233;
    wire N__93232;
    wire N__93231;
    wire N__93230;
    wire N__93229;
    wire N__93228;
    wire N__93227;
    wire N__93226;
    wire N__93225;
    wire N__93224;
    wire N__93223;
    wire N__93222;
    wire N__93221;
    wire N__93220;
    wire N__93219;
    wire N__93218;
    wire N__93217;
    wire N__93216;
    wire N__93215;
    wire N__93214;
    wire N__93213;
    wire N__93212;
    wire N__93211;
    wire N__93210;
    wire N__93209;
    wire N__93208;
    wire N__93207;
    wire N__93206;
    wire N__93205;
    wire N__93204;
    wire N__93203;
    wire N__93202;
    wire N__93201;
    wire N__93200;
    wire N__93199;
    wire N__93198;
    wire N__93197;
    wire N__93196;
    wire N__93195;
    wire N__93194;
    wire N__93193;
    wire N__93192;
    wire N__93191;
    wire N__93190;
    wire N__93189;
    wire N__93188;
    wire N__93187;
    wire N__93186;
    wire N__93185;
    wire N__93184;
    wire N__93183;
    wire N__93182;
    wire N__93181;
    wire N__93180;
    wire N__93179;
    wire N__93178;
    wire N__93177;
    wire N__93176;
    wire N__93175;
    wire N__93174;
    wire N__93173;
    wire N__93172;
    wire N__93171;
    wire N__93170;
    wire N__93169;
    wire N__93168;
    wire N__93167;
    wire N__93166;
    wire N__93165;
    wire N__93164;
    wire N__93163;
    wire N__93162;
    wire N__93161;
    wire N__93160;
    wire N__93159;
    wire N__93158;
    wire N__93157;
    wire N__93156;
    wire N__93155;
    wire N__93154;
    wire N__93153;
    wire N__93152;
    wire N__93151;
    wire N__93150;
    wire N__93149;
    wire N__93148;
    wire N__93147;
    wire N__93146;
    wire N__93145;
    wire N__93144;
    wire N__93143;
    wire N__93142;
    wire N__93141;
    wire N__93140;
    wire N__93139;
    wire N__93138;
    wire N__93137;
    wire N__93136;
    wire N__93135;
    wire N__93134;
    wire N__93133;
    wire N__93132;
    wire N__93131;
    wire N__93130;
    wire N__93129;
    wire N__93128;
    wire N__93127;
    wire N__93126;
    wire N__93125;
    wire N__93124;
    wire N__93123;
    wire N__93122;
    wire N__93121;
    wire N__93120;
    wire N__93119;
    wire N__93118;
    wire N__93117;
    wire N__93116;
    wire N__93115;
    wire N__93114;
    wire N__93113;
    wire N__93112;
    wire N__93111;
    wire N__93110;
    wire N__93109;
    wire N__93108;
    wire N__93107;
    wire N__93106;
    wire N__93105;
    wire N__93104;
    wire N__93103;
    wire N__93102;
    wire N__93101;
    wire N__93100;
    wire N__93099;
    wire N__93098;
    wire N__93097;
    wire N__93096;
    wire N__93095;
    wire N__93094;
    wire N__93093;
    wire N__93092;
    wire N__93091;
    wire N__93090;
    wire N__93089;
    wire N__93088;
    wire N__93087;
    wire N__93086;
    wire N__93085;
    wire N__93084;
    wire N__93083;
    wire N__93082;
    wire N__93081;
    wire N__93080;
    wire N__93079;
    wire N__93078;
    wire N__93077;
    wire N__93076;
    wire N__93075;
    wire N__93074;
    wire N__93073;
    wire N__93072;
    wire N__93071;
    wire N__93070;
    wire N__93069;
    wire N__93068;
    wire N__93067;
    wire N__93066;
    wire N__93065;
    wire N__93064;
    wire N__93063;
    wire N__93062;
    wire N__93061;
    wire N__93060;
    wire N__93059;
    wire N__93058;
    wire N__93057;
    wire N__93056;
    wire N__93055;
    wire N__93054;
    wire N__93053;
    wire N__93052;
    wire N__93051;
    wire N__93050;
    wire N__93049;
    wire N__93048;
    wire N__93047;
    wire N__93046;
    wire N__93045;
    wire N__93044;
    wire N__93043;
    wire N__93042;
    wire N__93041;
    wire N__93040;
    wire N__93039;
    wire N__93038;
    wire N__93037;
    wire N__93036;
    wire N__93035;
    wire N__93034;
    wire N__93033;
    wire N__93032;
    wire N__93031;
    wire N__93030;
    wire N__93029;
    wire N__93028;
    wire N__93027;
    wire N__93026;
    wire N__93025;
    wire N__93024;
    wire N__93023;
    wire N__93022;
    wire N__93021;
    wire N__93020;
    wire N__93019;
    wire N__93018;
    wire N__93017;
    wire N__93016;
    wire N__93015;
    wire N__93014;
    wire N__93013;
    wire N__93012;
    wire N__93011;
    wire N__93010;
    wire N__93009;
    wire N__93008;
    wire N__93007;
    wire N__93006;
    wire N__93005;
    wire N__93004;
    wire N__93003;
    wire N__93002;
    wire N__93001;
    wire N__93000;
    wire N__92999;
    wire N__92998;
    wire N__92997;
    wire N__92996;
    wire N__92995;
    wire N__92994;
    wire N__92993;
    wire N__92992;
    wire N__92991;
    wire N__92990;
    wire N__92989;
    wire N__92988;
    wire N__92987;
    wire N__92986;
    wire N__92985;
    wire N__92984;
    wire N__92983;
    wire N__92982;
    wire N__92981;
    wire N__92980;
    wire N__92979;
    wire N__92978;
    wire N__92977;
    wire N__92976;
    wire N__92975;
    wire N__92974;
    wire N__92973;
    wire N__92972;
    wire N__92971;
    wire N__92970;
    wire N__92969;
    wire N__92968;
    wire N__92967;
    wire N__92966;
    wire N__92965;
    wire N__92964;
    wire N__92963;
    wire N__92962;
    wire N__92961;
    wire N__92960;
    wire N__92959;
    wire N__92958;
    wire N__92957;
    wire N__92956;
    wire N__92955;
    wire N__92954;
    wire N__92953;
    wire N__92952;
    wire N__92951;
    wire N__92950;
    wire N__92949;
    wire N__92948;
    wire N__92947;
    wire N__92946;
    wire N__92945;
    wire N__92944;
    wire N__92943;
    wire N__92942;
    wire N__92941;
    wire N__92940;
    wire N__92939;
    wire N__92938;
    wire N__92937;
    wire N__92936;
    wire N__92935;
    wire N__92934;
    wire N__92933;
    wire N__92932;
    wire N__92931;
    wire N__92930;
    wire N__92929;
    wire N__92928;
    wire N__92927;
    wire N__92926;
    wire N__92925;
    wire N__92924;
    wire N__92923;
    wire N__92922;
    wire N__92921;
    wire N__92920;
    wire N__92919;
    wire N__92918;
    wire N__92917;
    wire N__92916;
    wire N__92915;
    wire N__92914;
    wire N__92913;
    wire N__92912;
    wire N__92911;
    wire N__92910;
    wire N__92909;
    wire N__92908;
    wire N__92907;
    wire N__91864;
    wire N__91861;
    wire N__91858;
    wire N__91857;
    wire N__91856;
    wire N__91855;
    wire N__91852;
    wire N__91849;
    wire N__91846;
    wire N__91843;
    wire N__91838;
    wire N__91835;
    wire N__91832;
    wire N__91825;
    wire N__91822;
    wire N__91821;
    wire N__91818;
    wire N__91815;
    wire N__91814;
    wire N__91811;
    wire N__91808;
    wire N__91807;
    wire N__91804;
    wire N__91799;
    wire N__91798;
    wire N__91795;
    wire N__91792;
    wire N__91789;
    wire N__91786;
    wire N__91777;
    wire N__91774;
    wire N__91771;
    wire N__91768;
    wire N__91767;
    wire N__91764;
    wire N__91763;
    wire N__91762;
    wire N__91761;
    wire N__91758;
    wire N__91755;
    wire N__91752;
    wire N__91749;
    wire N__91746;
    wire N__91743;
    wire N__91742;
    wire N__91737;
    wire N__91736;
    wire N__91733;
    wire N__91728;
    wire N__91725;
    wire N__91722;
    wire N__91719;
    wire N__91716;
    wire N__91713;
    wire N__91710;
    wire N__91699;
    wire N__91698;
    wire N__91695;
    wire N__91692;
    wire N__91691;
    wire N__91690;
    wire N__91689;
    wire N__91688;
    wire N__91683;
    wire N__91682;
    wire N__91679;
    wire N__91676;
    wire N__91673;
    wire N__91670;
    wire N__91667;
    wire N__91664;
    wire N__91661;
    wire N__91658;
    wire N__91653;
    wire N__91648;
    wire N__91647;
    wire N__91646;
    wire N__91643;
    wire N__91638;
    wire N__91635;
    wire N__91630;
    wire N__91621;
    wire N__91618;
    wire N__91615;
    wire N__91612;
    wire N__91609;
    wire N__91608;
    wire N__91607;
    wire N__91606;
    wire N__91603;
    wire N__91600;
    wire N__91597;
    wire N__91594;
    wire N__91589;
    wire N__91582;
    wire N__91579;
    wire N__91576;
    wire N__91573;
    wire N__91570;
    wire N__91567;
    wire N__91566;
    wire N__91565;
    wire N__91562;
    wire N__91559;
    wire N__91556;
    wire N__91553;
    wire N__91550;
    wire N__91547;
    wire N__91540;
    wire N__91539;
    wire N__91538;
    wire N__91537;
    wire N__91534;
    wire N__91533;
    wire N__91532;
    wire N__91531;
    wire N__91530;
    wire N__91529;
    wire N__91528;
    wire N__91527;
    wire N__91526;
    wire N__91525;
    wire N__91522;
    wire N__91517;
    wire N__91516;
    wire N__91513;
    wire N__91512;
    wire N__91511;
    wire N__91506;
    wire N__91497;
    wire N__91494;
    wire N__91493;
    wire N__91488;
    wire N__91483;
    wire N__91480;
    wire N__91479;
    wire N__91478;
    wire N__91475;
    wire N__91470;
    wire N__91465;
    wire N__91462;
    wire N__91459;
    wire N__91458;
    wire N__91457;
    wire N__91454;
    wire N__91451;
    wire N__91448;
    wire N__91443;
    wire N__91438;
    wire N__91435;
    wire N__91430;
    wire N__91425;
    wire N__91422;
    wire N__91415;
    wire N__91412;
    wire N__91399;
    wire N__91396;
    wire N__91393;
    wire N__91390;
    wire N__91387;
    wire N__91384;
    wire N__91381;
    wire N__91378;
    wire N__91375;
    wire N__91374;
    wire N__91371;
    wire N__91368;
    wire N__91365;
    wire N__91362;
    wire N__91359;
    wire N__91356;
    wire N__91351;
    wire N__91348;
    wire N__91345;
    wire N__91342;
    wire N__91339;
    wire N__91336;
    wire N__91335;
    wire N__91334;
    wire N__91329;
    wire N__91326;
    wire N__91325;
    wire N__91322;
    wire N__91319;
    wire N__91316;
    wire N__91313;
    wire N__91310;
    wire N__91307;
    wire N__91306;
    wire N__91303;
    wire N__91300;
    wire N__91297;
    wire N__91294;
    wire N__91291;
    wire N__91284;
    wire N__91279;
    wire N__91276;
    wire N__91273;
    wire N__91270;
    wire N__91269;
    wire N__91268;
    wire N__91267;
    wire N__91266;
    wire N__91263;
    wire N__91260;
    wire N__91257;
    wire N__91256;
    wire N__91251;
    wire N__91250;
    wire N__91249;
    wire N__91248;
    wire N__91247;
    wire N__91246;
    wire N__91245;
    wire N__91242;
    wire N__91239;
    wire N__91236;
    wire N__91233;
    wire N__91230;
    wire N__91221;
    wire N__91218;
    wire N__91215;
    wire N__91214;
    wire N__91213;
    wire N__91210;
    wire N__91205;
    wire N__91200;
    wire N__91195;
    wire N__91192;
    wire N__91187;
    wire N__91174;
    wire N__91171;
    wire N__91168;
    wire N__91165;
    wire N__91162;
    wire N__91159;
    wire N__91156;
    wire N__91155;
    wire N__91152;
    wire N__91149;
    wire N__91146;
    wire N__91143;
    wire N__91140;
    wire N__91137;
    wire N__91134;
    wire N__91131;
    wire N__91126;
    wire N__91123;
    wire N__91120;
    wire N__91117;
    wire N__91114;
    wire N__91113;
    wire N__91112;
    wire N__91111;
    wire N__91110;
    wire N__91107;
    wire N__91104;
    wire N__91101;
    wire N__91096;
    wire N__91093;
    wire N__91090;
    wire N__91087;
    wire N__91084;
    wire N__91083;
    wire N__91082;
    wire N__91077;
    wire N__91074;
    wire N__91071;
    wire N__91066;
    wire N__91061;
    wire N__91058;
    wire N__91055;
    wire N__91048;
    wire N__91045;
    wire N__91042;
    wire N__91039;
    wire N__91036;
    wire N__91033;
    wire N__91030;
    wire N__91027;
    wire N__91024;
    wire N__91021;
    wire N__91018;
    wire N__91015;
    wire N__91012;
    wire N__91009;
    wire N__91006;
    wire N__91003;
    wire N__91000;
    wire N__90997;
    wire N__90996;
    wire N__90993;
    wire N__90990;
    wire N__90987;
    wire N__90984;
    wire N__90981;
    wire N__90976;
    wire N__90973;
    wire N__90970;
    wire N__90967;
    wire N__90964;
    wire N__90961;
    wire N__90958;
    wire N__90955;
    wire N__90952;
    wire N__90949;
    wire N__90946;
    wire N__90943;
    wire N__90942;
    wire N__90939;
    wire N__90938;
    wire N__90935;
    wire N__90932;
    wire N__90929;
    wire N__90926;
    wire N__90923;
    wire N__90920;
    wire N__90919;
    wire N__90918;
    wire N__90915;
    wire N__90910;
    wire N__90907;
    wire N__90904;
    wire N__90901;
    wire N__90898;
    wire N__90895;
    wire N__90892;
    wire N__90883;
    wire N__90882;
    wire N__90879;
    wire N__90876;
    wire N__90875;
    wire N__90870;
    wire N__90869;
    wire N__90866;
    wire N__90863;
    wire N__90860;
    wire N__90857;
    wire N__90854;
    wire N__90847;
    wire N__90846;
    wire N__90843;
    wire N__90840;
    wire N__90839;
    wire N__90838;
    wire N__90835;
    wire N__90834;
    wire N__90831;
    wire N__90828;
    wire N__90827;
    wire N__90824;
    wire N__90821;
    wire N__90818;
    wire N__90813;
    wire N__90808;
    wire N__90799;
    wire N__90796;
    wire N__90793;
    wire N__90790;
    wire N__90787;
    wire N__90786;
    wire N__90785;
    wire N__90782;
    wire N__90779;
    wire N__90776;
    wire N__90775;
    wire N__90770;
    wire N__90767;
    wire N__90766;
    wire N__90763;
    wire N__90758;
    wire N__90755;
    wire N__90752;
    wire N__90749;
    wire N__90746;
    wire N__90739;
    wire N__90738;
    wire N__90735;
    wire N__90734;
    wire N__90733;
    wire N__90730;
    wire N__90729;
    wire N__90728;
    wire N__90727;
    wire N__90724;
    wire N__90721;
    wire N__90718;
    wire N__90715;
    wire N__90714;
    wire N__90713;
    wire N__90710;
    wire N__90707;
    wire N__90704;
    wire N__90697;
    wire N__90696;
    wire N__90695;
    wire N__90694;
    wire N__90693;
    wire N__90690;
    wire N__90685;
    wire N__90680;
    wire N__90677;
    wire N__90674;
    wire N__90667;
    wire N__90664;
    wire N__90659;
    wire N__90656;
    wire N__90653;
    wire N__90646;
    wire N__90643;
    wire N__90640;
    wire N__90631;
    wire N__90628;
    wire N__90625;
    wire N__90622;
    wire N__90619;
    wire N__90616;
    wire N__90613;
    wire N__90610;
    wire N__90607;
    wire N__90604;
    wire N__90601;
    wire N__90598;
    wire N__90595;
    wire N__90592;
    wire N__90589;
    wire N__90586;
    wire N__90585;
    wire N__90584;
    wire N__90581;
    wire N__90580;
    wire N__90579;
    wire N__90572;
    wire N__90571;
    wire N__90570;
    wire N__90569;
    wire N__90566;
    wire N__90565;
    wire N__90564;
    wire N__90563;
    wire N__90562;
    wire N__90561;
    wire N__90560;
    wire N__90559;
    wire N__90558;
    wire N__90557;
    wire N__90556;
    wire N__90555;
    wire N__90554;
    wire N__90553;
    wire N__90552;
    wire N__90551;
    wire N__90550;
    wire N__90547;
    wire N__90546;
    wire N__90543;
    wire N__90534;
    wire N__90533;
    wire N__90532;
    wire N__90531;
    wire N__90530;
    wire N__90523;
    wire N__90520;
    wire N__90519;
    wire N__90518;
    wire N__90517;
    wire N__90514;
    wire N__90513;
    wire N__90510;
    wire N__90501;
    wire N__90498;
    wire N__90495;
    wire N__90494;
    wire N__90493;
    wire N__90492;
    wire N__90489;
    wire N__90488;
    wire N__90487;
    wire N__90486;
    wire N__90485;
    wire N__90484;
    wire N__90483;
    wire N__90482;
    wire N__90479;
    wire N__90476;
    wire N__90475;
    wire N__90474;
    wire N__90473;
    wire N__90472;
    wire N__90471;
    wire N__90468;
    wire N__90465;
    wire N__90464;
    wire N__90463;
    wire N__90462;
    wire N__90461;
    wire N__90460;
    wire N__90459;
    wire N__90458;
    wire N__90455;
    wire N__90454;
    wire N__90453;
    wire N__90452;
    wire N__90451;
    wire N__90450;
    wire N__90449;
    wire N__90444;
    wire N__90443;
    wire N__90440;
    wire N__90439;
    wire N__90436;
    wire N__90435;
    wire N__90434;
    wire N__90433;
    wire N__90432;
    wire N__90431;
    wire N__90430;
    wire N__90429;
    wire N__90428;
    wire N__90427;
    wire N__90426;
    wire N__90425;
    wire N__90424;
    wire N__90423;
    wire N__90422;
    wire N__90421;
    wire N__90420;
    wire N__90417;
    wire N__90414;
    wire N__90413;
    wire N__90410;
    wire N__90407;
    wire N__90406;
    wire N__90405;
    wire N__90404;
    wire N__90403;
    wire N__90400;
    wire N__90399;
    wire N__90396;
    wire N__90395;
    wire N__90392;
    wire N__90391;
    wire N__90390;
    wire N__90389;
    wire N__90386;
    wire N__90381;
    wire N__90378;
    wire N__90371;
    wire N__90370;
    wire N__90367;
    wire N__90364;
    wire N__90357;
    wire N__90354;
    wire N__90351;
    wire N__90350;
    wire N__90349;
    wire N__90346;
    wire N__90345;
    wire N__90344;
    wire N__90341;
    wire N__90338;
    wire N__90335;
    wire N__90330;
    wire N__90329;
    wire N__90328;
    wire N__90325;
    wire N__90322;
    wire N__90321;
    wire N__90320;
    wire N__90319;
    wire N__90318;
    wire N__90313;
    wire N__90310;
    wire N__90309;
    wire N__90308;
    wire N__90307;
    wire N__90304;
    wire N__90301;
    wire N__90298;
    wire N__90293;
    wire N__90292;
    wire N__90289;
    wire N__90286;
    wire N__90285;
    wire N__90282;
    wire N__90279;
    wire N__90278;
    wire N__90273;
    wire N__90266;
    wire N__90265;
    wire N__90264;
    wire N__90263;
    wire N__90260;
    wire N__90257;
    wire N__90248;
    wire N__90245;
    wire N__90244;
    wire N__90243;
    wire N__90242;
    wire N__90239;
    wire N__90238;
    wire N__90237;
    wire N__90236;
    wire N__90235;
    wire N__90234;
    wire N__90231;
    wire N__90230;
    wire N__90229;
    wire N__90228;
    wire N__90227;
    wire N__90226;
    wire N__90225;
    wire N__90224;
    wire N__90221;
    wire N__90218;
    wire N__90213;
    wire N__90212;
    wire N__90211;
    wire N__90210;
    wire N__90207;
    wire N__90204;
    wire N__90201;
    wire N__90198;
    wire N__90195;
    wire N__90190;
    wire N__90187;
    wire N__90186;
    wire N__90185;
    wire N__90184;
    wire N__90183;
    wire N__90180;
    wire N__90175;
    wire N__90172;
    wire N__90167;
    wire N__90164;
    wire N__90163;
    wire N__90158;
    wire N__90153;
    wire N__90150;
    wire N__90147;
    wire N__90142;
    wire N__90141;
    wire N__90134;
    wire N__90133;
    wire N__90130;
    wire N__90123;
    wire N__90120;
    wire N__90117;
    wire N__90114;
    wire N__90109;
    wire N__90106;
    wire N__90101;
    wire N__90092;
    wire N__90085;
    wire N__90078;
    wire N__90077;
    wire N__90076;
    wire N__90075;
    wire N__90072;
    wire N__90071;
    wire N__90068;
    wire N__90065;
    wire N__90062;
    wire N__90059;
    wire N__90054;
    wire N__90051;
    wire N__90048;
    wire N__90045;
    wire N__90044;
    wire N__90043;
    wire N__90042;
    wire N__90041;
    wire N__90040;
    wire N__90033;
    wire N__90030;
    wire N__90027;
    wire N__90026;
    wire N__90025;
    wire N__90024;
    wire N__90023;
    wire N__90022;
    wire N__90017;
    wire N__90014;
    wire N__90013;
    wire N__90010;
    wire N__90007;
    wire N__90004;
    wire N__90001;
    wire N__89998;
    wire N__89993;
    wire N__89990;
    wire N__89987;
    wire N__89982;
    wire N__89979;
    wire N__89978;
    wire N__89975;
    wire N__89974;
    wire N__89973;
    wire N__89972;
    wire N__89969;
    wire N__89968;
    wire N__89967;
    wire N__89964;
    wire N__89959;
    wire N__89952;
    wire N__89951;
    wire N__89950;
    wire N__89947;
    wire N__89946;
    wire N__89945;
    wire N__89944;
    wire N__89943;
    wire N__89940;
    wire N__89935;
    wire N__89932;
    wire N__89931;
    wire N__89930;
    wire N__89927;
    wire N__89922;
    wire N__89917;
    wire N__89916;
    wire N__89911;
    wire N__89908;
    wire N__89903;
    wire N__89902;
    wire N__89897;
    wire N__89892;
    wire N__89887;
    wire N__89884;
    wire N__89881;
    wire N__89876;
    wire N__89873;
    wire N__89866;
    wire N__89863;
    wire N__89858;
    wire N__89853;
    wire N__89850;
    wire N__89845;
    wire N__89842;
    wire N__89839;
    wire N__89836;
    wire N__89831;
    wire N__89826;
    wire N__89823;
    wire N__89820;
    wire N__89809;
    wire N__89806;
    wire N__89803;
    wire N__89800;
    wire N__89799;
    wire N__89798;
    wire N__89795;
    wire N__89794;
    wire N__89793;
    wire N__89792;
    wire N__89789;
    wire N__89788;
    wire N__89787;
    wire N__89786;
    wire N__89777;
    wire N__89774;
    wire N__89769;
    wire N__89766;
    wire N__89765;
    wire N__89762;
    wire N__89761;
    wire N__89760;
    wire N__89759;
    wire N__89756;
    wire N__89753;
    wire N__89748;
    wire N__89743;
    wire N__89740;
    wire N__89729;
    wire N__89726;
    wire N__89723;
    wire N__89720;
    wire N__89717;
    wire N__89704;
    wire N__89701;
    wire N__89696;
    wire N__89687;
    wire N__89684;
    wire N__89681;
    wire N__89674;
    wire N__89671;
    wire N__89668;
    wire N__89663;
    wire N__89660;
    wire N__89659;
    wire N__89658;
    wire N__89655;
    wire N__89648;
    wire N__89645;
    wire N__89642;
    wire N__89635;
    wire N__89628;
    wire N__89625;
    wire N__89622;
    wire N__89619;
    wire N__89618;
    wire N__89617;
    wire N__89616;
    wire N__89615;
    wire N__89614;
    wire N__89613;
    wire N__89610;
    wire N__89607;
    wire N__89600;
    wire N__89593;
    wire N__89590;
    wire N__89587;
    wire N__89582;
    wire N__89579;
    wire N__89574;
    wire N__89571;
    wire N__89568;
    wire N__89565;
    wire N__89562;
    wire N__89559;
    wire N__89552;
    wire N__89549;
    wire N__89546;
    wire N__89539;
    wire N__89536;
    wire N__89531;
    wire N__89526;
    wire N__89525;
    wire N__89524;
    wire N__89519;
    wire N__89516;
    wire N__89509;
    wire N__89506;
    wire N__89503;
    wire N__89500;
    wire N__89497;
    wire N__89494;
    wire N__89491;
    wire N__89486;
    wire N__89483;
    wire N__89480;
    wire N__89465;
    wire N__89460;
    wire N__89459;
    wire N__89458;
    wire N__89455;
    wire N__89450;
    wire N__89447;
    wire N__89444;
    wire N__89437;
    wire N__89430;
    wire N__89421;
    wire N__89418;
    wire N__89411;
    wire N__89408;
    wire N__89405;
    wire N__89402;
    wire N__89395;
    wire N__89390;
    wire N__89385;
    wire N__89378;
    wire N__89373;
    wire N__89360;
    wire N__89347;
    wire N__89344;
    wire N__89341;
    wire N__89338;
    wire N__89335;
    wire N__89332;
    wire N__89331;
    wire N__89328;
    wire N__89325;
    wire N__89320;
    wire N__89317;
    wire N__89304;
    wire N__89301;
    wire N__89298;
    wire N__89293;
    wire N__89286;
    wire N__89283;
    wire N__89276;
    wire N__89255;
    wire N__89244;
    wire N__89241;
    wire N__89234;
    wire N__89229;
    wire N__89214;
    wire N__89211;
    wire N__89200;
    wire N__89197;
    wire N__89194;
    wire N__89191;
    wire N__89188;
    wire N__89185;
    wire N__89182;
    wire N__89181;
    wire N__89180;
    wire N__89179;
    wire N__89178;
    wire N__89171;
    wire N__89170;
    wire N__89165;
    wire N__89162;
    wire N__89159;
    wire N__89156;
    wire N__89153;
    wire N__89146;
    wire N__89143;
    wire N__89140;
    wire N__89137;
    wire N__89134;
    wire N__89131;
    wire N__89128;
    wire N__89125;
    wire N__89122;
    wire N__89119;
    wire N__89116;
    wire N__89113;
    wire N__89110;
    wire N__89107;
    wire N__89106;
    wire N__89105;
    wire N__89104;
    wire N__89101;
    wire N__89098;
    wire N__89095;
    wire N__89092;
    wire N__89085;
    wire N__89082;
    wire N__89079;
    wire N__89076;
    wire N__89073;
    wire N__89068;
    wire N__89065;
    wire N__89062;
    wire N__89059;
    wire N__89056;
    wire N__89053;
    wire N__89050;
    wire N__89047;
    wire N__89044;
    wire N__89041;
    wire N__89038;
    wire N__89035;
    wire N__89032;
    wire N__89029;
    wire N__89026;
    wire N__89023;
    wire N__89020;
    wire N__89017;
    wire N__89014;
    wire N__89011;
    wire N__89008;
    wire N__89005;
    wire N__89004;
    wire N__89001;
    wire N__88998;
    wire N__88993;
    wire N__88990;
    wire N__88987;
    wire N__88984;
    wire N__88981;
    wire N__88978;
    wire N__88975;
    wire N__88972;
    wire N__88969;
    wire N__88966;
    wire N__88963;
    wire N__88960;
    wire N__88957;
    wire N__88954;
    wire N__88951;
    wire N__88948;
    wire N__88945;
    wire N__88942;
    wire N__88939;
    wire N__88938;
    wire N__88935;
    wire N__88932;
    wire N__88929;
    wire N__88924;
    wire N__88921;
    wire N__88918;
    wire N__88915;
    wire N__88912;
    wire N__88911;
    wire N__88908;
    wire N__88905;
    wire N__88900;
    wire N__88897;
    wire N__88894;
    wire N__88891;
    wire N__88888;
    wire N__88885;
    wire N__88882;
    wire N__88881;
    wire N__88878;
    wire N__88875;
    wire N__88870;
    wire N__88867;
    wire N__88864;
    wire N__88861;
    wire N__88858;
    wire N__88855;
    wire N__88852;
    wire N__88849;
    wire N__88846;
    wire N__88843;
    wire N__88840;
    wire N__88837;
    wire N__88834;
    wire N__88833;
    wire N__88832;
    wire N__88829;
    wire N__88826;
    wire N__88825;
    wire N__88822;
    wire N__88817;
    wire N__88814;
    wire N__88811;
    wire N__88808;
    wire N__88805;
    wire N__88802;
    wire N__88799;
    wire N__88792;
    wire N__88789;
    wire N__88786;
    wire N__88783;
    wire N__88780;
    wire N__88777;
    wire N__88774;
    wire N__88771;
    wire N__88768;
    wire N__88765;
    wire N__88762;
    wire N__88759;
    wire N__88756;
    wire N__88753;
    wire N__88750;
    wire N__88747;
    wire N__88744;
    wire N__88741;
    wire N__88738;
    wire N__88735;
    wire N__88732;
    wire N__88729;
    wire N__88726;
    wire N__88723;
    wire N__88720;
    wire N__88717;
    wire N__88714;
    wire N__88711;
    wire N__88708;
    wire N__88705;
    wire N__88702;
    wire N__88701;
    wire N__88700;
    wire N__88697;
    wire N__88694;
    wire N__88691;
    wire N__88688;
    wire N__88685;
    wire N__88682;
    wire N__88679;
    wire N__88676;
    wire N__88673;
    wire N__88666;
    wire N__88663;
    wire N__88660;
    wire N__88657;
    wire N__88654;
    wire N__88651;
    wire N__88648;
    wire N__88645;
    wire N__88642;
    wire N__88639;
    wire N__88636;
    wire N__88633;
    wire N__88630;
    wire N__88627;
    wire N__88624;
    wire N__88621;
    wire N__88618;
    wire N__88615;
    wire N__88612;
    wire N__88611;
    wire N__88610;
    wire N__88609;
    wire N__88606;
    wire N__88605;
    wire N__88602;
    wire N__88597;
    wire N__88594;
    wire N__88591;
    wire N__88586;
    wire N__88585;
    wire N__88584;
    wire N__88581;
    wire N__88578;
    wire N__88575;
    wire N__88570;
    wire N__88561;
    wire N__88558;
    wire N__88555;
    wire N__88552;
    wire N__88549;
    wire N__88546;
    wire N__88545;
    wire N__88544;
    wire N__88543;
    wire N__88542;
    wire N__88541;
    wire N__88538;
    wire N__88535;
    wire N__88534;
    wire N__88533;
    wire N__88524;
    wire N__88523;
    wire N__88518;
    wire N__88513;
    wire N__88510;
    wire N__88509;
    wire N__88508;
    wire N__88505;
    wire N__88500;
    wire N__88497;
    wire N__88492;
    wire N__88489;
    wire N__88486;
    wire N__88481;
    wire N__88478;
    wire N__88475;
    wire N__88472;
    wire N__88465;
    wire N__88464;
    wire N__88461;
    wire N__88460;
    wire N__88457;
    wire N__88454;
    wire N__88451;
    wire N__88448;
    wire N__88447;
    wire N__88444;
    wire N__88439;
    wire N__88438;
    wire N__88435;
    wire N__88432;
    wire N__88429;
    wire N__88424;
    wire N__88417;
    wire N__88414;
    wire N__88411;
    wire N__88408;
    wire N__88405;
    wire N__88404;
    wire N__88403;
    wire N__88398;
    wire N__88395;
    wire N__88394;
    wire N__88391;
    wire N__88390;
    wire N__88387;
    wire N__88384;
    wire N__88381;
    wire N__88378;
    wire N__88373;
    wire N__88366;
    wire N__88363;
    wire N__88360;
    wire N__88357;
    wire N__88354;
    wire N__88351;
    wire N__88348;
    wire N__88345;
    wire N__88342;
    wire N__88339;
    wire N__88336;
    wire N__88333;
    wire N__88330;
    wire N__88329;
    wire N__88326;
    wire N__88325;
    wire N__88324;
    wire N__88321;
    wire N__88320;
    wire N__88317;
    wire N__88310;
    wire N__88307;
    wire N__88304;
    wire N__88301;
    wire N__88298;
    wire N__88291;
    wire N__88288;
    wire N__88285;
    wire N__88282;
    wire N__88279;
    wire N__88278;
    wire N__88275;
    wire N__88272;
    wire N__88269;
    wire N__88266;
    wire N__88261;
    wire N__88258;
    wire N__88255;
    wire N__88252;
    wire N__88249;
    wire N__88246;
    wire N__88243;
    wire N__88240;
    wire N__88237;
    wire N__88234;
    wire N__88231;
    wire N__88228;
    wire N__88225;
    wire N__88222;
    wire N__88219;
    wire N__88216;
    wire N__88213;
    wire N__88210;
    wire N__88207;
    wire N__88204;
    wire N__88203;
    wire N__88200;
    wire N__88197;
    wire N__88194;
    wire N__88191;
    wire N__88186;
    wire N__88183;
    wire N__88180;
    wire N__88177;
    wire N__88174;
    wire N__88171;
    wire N__88168;
    wire N__88165;
    wire N__88162;
    wire N__88159;
    wire N__88156;
    wire N__88153;
    wire N__88150;
    wire N__88147;
    wire N__88144;
    wire N__88141;
    wire N__88138;
    wire N__88135;
    wire N__88132;
    wire N__88129;
    wire N__88128;
    wire N__88125;
    wire N__88122;
    wire N__88117;
    wire N__88114;
    wire N__88113;
    wire N__88112;
    wire N__88109;
    wire N__88106;
    wire N__88103;
    wire N__88102;
    wire N__88101;
    wire N__88098;
    wire N__88097;
    wire N__88092;
    wire N__88087;
    wire N__88084;
    wire N__88081;
    wire N__88076;
    wire N__88069;
    wire N__88066;
    wire N__88063;
    wire N__88060;
    wire N__88057;
    wire N__88054;
    wire N__88051;
    wire N__88048;
    wire N__88045;
    wire N__88042;
    wire N__88039;
    wire N__88036;
    wire N__88033;
    wire N__88030;
    wire N__88027;
    wire N__88024;
    wire N__88021;
    wire N__88018;
    wire N__88015;
    wire N__88012;
    wire N__88011;
    wire N__88010;
    wire N__88009;
    wire N__88006;
    wire N__88005;
    wire N__88004;
    wire N__87997;
    wire N__87996;
    wire N__87993;
    wire N__87992;
    wire N__87989;
    wire N__87988;
    wire N__87985;
    wire N__87984;
    wire N__87981;
    wire N__87978;
    wire N__87975;
    wire N__87972;
    wire N__87967;
    wire N__87964;
    wire N__87961;
    wire N__87960;
    wire N__87957;
    wire N__87954;
    wire N__87947;
    wire N__87944;
    wire N__87941;
    wire N__87938;
    wire N__87933;
    wire N__87930;
    wire N__87925;
    wire N__87916;
    wire N__87913;
    wire N__87910;
    wire N__87909;
    wire N__87908;
    wire N__87907;
    wire N__87906;
    wire N__87905;
    wire N__87904;
    wire N__87901;
    wire N__87900;
    wire N__87887;
    wire N__87884;
    wire N__87881;
    wire N__87880;
    wire N__87879;
    wire N__87876;
    wire N__87875;
    wire N__87874;
    wire N__87873;
    wire N__87870;
    wire N__87869;
    wire N__87866;
    wire N__87861;
    wire N__87858;
    wire N__87851;
    wire N__87848;
    wire N__87845;
    wire N__87844;
    wire N__87843;
    wire N__87842;
    wire N__87839;
    wire N__87836;
    wire N__87833;
    wire N__87830;
    wire N__87827;
    wire N__87818;
    wire N__87815;
    wire N__87812;
    wire N__87807;
    wire N__87796;
    wire N__87795;
    wire N__87792;
    wire N__87789;
    wire N__87786;
    wire N__87785;
    wire N__87782;
    wire N__87779;
    wire N__87776;
    wire N__87773;
    wire N__87768;
    wire N__87763;
    wire N__87762;
    wire N__87761;
    wire N__87758;
    wire N__87753;
    wire N__87750;
    wire N__87749;
    wire N__87746;
    wire N__87743;
    wire N__87742;
    wire N__87739;
    wire N__87734;
    wire N__87731;
    wire N__87724;
    wire N__87721;
    wire N__87720;
    wire N__87719;
    wire N__87718;
    wire N__87717;
    wire N__87716;
    wire N__87713;
    wire N__87712;
    wire N__87709;
    wire N__87708;
    wire N__87699;
    wire N__87698;
    wire N__87695;
    wire N__87692;
    wire N__87691;
    wire N__87688;
    wire N__87685;
    wire N__87682;
    wire N__87679;
    wire N__87676;
    wire N__87671;
    wire N__87670;
    wire N__87669;
    wire N__87666;
    wire N__87663;
    wire N__87662;
    wire N__87657;
    wire N__87654;
    wire N__87651;
    wire N__87648;
    wire N__87645;
    wire N__87642;
    wire N__87639;
    wire N__87636;
    wire N__87635;
    wire N__87634;
    wire N__87633;
    wire N__87630;
    wire N__87627;
    wire N__87624;
    wire N__87619;
    wire N__87614;
    wire N__87605;
    wire N__87602;
    wire N__87595;
    wire N__87586;
    wire N__87583;
    wire N__87580;
    wire N__87577;
    wire N__87574;
    wire N__87571;
    wire N__87568;
    wire N__87565;
    wire N__87562;
    wire N__87559;
    wire N__87556;
    wire N__87553;
    wire N__87550;
    wire N__87547;
    wire N__87544;
    wire N__87541;
    wire N__87538;
    wire N__87535;
    wire N__87532;
    wire N__87529;
    wire N__87526;
    wire N__87523;
    wire N__87520;
    wire N__87517;
    wire N__87514;
    wire N__87511;
    wire N__87508;
    wire N__87505;
    wire N__87502;
    wire N__87499;
    wire N__87496;
    wire N__87495;
    wire N__87494;
    wire N__87491;
    wire N__87488;
    wire N__87485;
    wire N__87480;
    wire N__87475;
    wire N__87472;
    wire N__87469;
    wire N__87466;
    wire N__87463;
    wire N__87462;
    wire N__87461;
    wire N__87458;
    wire N__87453;
    wire N__87450;
    wire N__87447;
    wire N__87442;
    wire N__87439;
    wire N__87436;
    wire N__87433;
    wire N__87430;
    wire N__87429;
    wire N__87426;
    wire N__87425;
    wire N__87420;
    wire N__87419;
    wire N__87416;
    wire N__87415;
    wire N__87414;
    wire N__87411;
    wire N__87406;
    wire N__87401;
    wire N__87398;
    wire N__87395;
    wire N__87388;
    wire N__87385;
    wire N__87382;
    wire N__87379;
    wire N__87376;
    wire N__87373;
    wire N__87370;
    wire N__87367;
    wire N__87364;
    wire N__87363;
    wire N__87360;
    wire N__87357;
    wire N__87354;
    wire N__87351;
    wire N__87348;
    wire N__87347;
    wire N__87344;
    wire N__87341;
    wire N__87338;
    wire N__87335;
    wire N__87330;
    wire N__87325;
    wire N__87324;
    wire N__87323;
    wire N__87320;
    wire N__87319;
    wire N__87318;
    wire N__87313;
    wire N__87310;
    wire N__87305;
    wire N__87302;
    wire N__87299;
    wire N__87298;
    wire N__87295;
    wire N__87292;
    wire N__87289;
    wire N__87286;
    wire N__87283;
    wire N__87280;
    wire N__87277;
    wire N__87268;
    wire N__87265;
    wire N__87262;
    wire N__87259;
    wire N__87256;
    wire N__87255;
    wire N__87252;
    wire N__87249;
    wire N__87246;
    wire N__87243;
    wire N__87242;
    wire N__87239;
    wire N__87236;
    wire N__87233;
    wire N__87226;
    wire N__87223;
    wire N__87220;
    wire N__87217;
    wire N__87214;
    wire N__87211;
    wire N__87208;
    wire N__87205;
    wire N__87202;
    wire N__87199;
    wire N__87196;
    wire N__87193;
    wire N__87190;
    wire N__87187;
    wire N__87186;
    wire N__87183;
    wire N__87180;
    wire N__87177;
    wire N__87174;
    wire N__87171;
    wire N__87170;
    wire N__87167;
    wire N__87164;
    wire N__87161;
    wire N__87154;
    wire N__87151;
    wire N__87148;
    wire N__87145;
    wire N__87142;
    wire N__87139;
    wire N__87136;
    wire N__87135;
    wire N__87132;
    wire N__87131;
    wire N__87128;
    wire N__87125;
    wire N__87122;
    wire N__87121;
    wire N__87120;
    wire N__87117;
    wire N__87112;
    wire N__87109;
    wire N__87106;
    wire N__87103;
    wire N__87100;
    wire N__87097;
    wire N__87094;
    wire N__87085;
    wire N__87082;
    wire N__87079;
    wire N__87076;
    wire N__87073;
    wire N__87070;
    wire N__87067;
    wire N__87064;
    wire N__87061;
    wire N__87058;
    wire N__87055;
    wire N__87052;
    wire N__87049;
    wire N__87046;
    wire N__87043;
    wire N__87040;
    wire N__87037;
    wire N__87034;
    wire N__87031;
    wire N__87028;
    wire N__87025;
    wire N__87022;
    wire N__87019;
    wire N__87016;
    wire N__87013;
    wire N__87010;
    wire N__87007;
    wire N__87004;
    wire N__87003;
    wire N__87002;
    wire N__86999;
    wire N__86996;
    wire N__86993;
    wire N__86986;
    wire N__86983;
    wire N__86980;
    wire N__86977;
    wire N__86974;
    wire N__86971;
    wire N__86968;
    wire N__86965;
    wire N__86962;
    wire N__86959;
    wire N__86956;
    wire N__86953;
    wire N__86950;
    wire N__86947;
    wire N__86944;
    wire N__86941;
    wire N__86938;
    wire N__86935;
    wire N__86934;
    wire N__86931;
    wire N__86928;
    wire N__86927;
    wire N__86926;
    wire N__86925;
    wire N__86920;
    wire N__86917;
    wire N__86914;
    wire N__86911;
    wire N__86908;
    wire N__86901;
    wire N__86896;
    wire N__86893;
    wire N__86892;
    wire N__86891;
    wire N__86888;
    wire N__86885;
    wire N__86882;
    wire N__86879;
    wire N__86876;
    wire N__86869;
    wire N__86868;
    wire N__86865;
    wire N__86862;
    wire N__86861;
    wire N__86860;
    wire N__86857;
    wire N__86856;
    wire N__86853;
    wire N__86848;
    wire N__86845;
    wire N__86842;
    wire N__86839;
    wire N__86834;
    wire N__86829;
    wire N__86824;
    wire N__86821;
    wire N__86818;
    wire N__86817;
    wire N__86816;
    wire N__86815;
    wire N__86812;
    wire N__86811;
    wire N__86810;
    wire N__86809;
    wire N__86806;
    wire N__86805;
    wire N__86804;
    wire N__86801;
    wire N__86800;
    wire N__86797;
    wire N__86794;
    wire N__86791;
    wire N__86786;
    wire N__86783;
    wire N__86778;
    wire N__86775;
    wire N__86772;
    wire N__86769;
    wire N__86766;
    wire N__86763;
    wire N__86760;
    wire N__86755;
    wire N__86754;
    wire N__86751;
    wire N__86742;
    wire N__86737;
    wire N__86734;
    wire N__86731;
    wire N__86728;
    wire N__86719;
    wire N__86718;
    wire N__86715;
    wire N__86714;
    wire N__86711;
    wire N__86708;
    wire N__86705;
    wire N__86698;
    wire N__86697;
    wire N__86696;
    wire N__86695;
    wire N__86694;
    wire N__86689;
    wire N__86686;
    wire N__86683;
    wire N__86680;
    wire N__86677;
    wire N__86672;
    wire N__86665;
    wire N__86664;
    wire N__86661;
    wire N__86660;
    wire N__86657;
    wire N__86656;
    wire N__86655;
    wire N__86654;
    wire N__86651;
    wire N__86648;
    wire N__86645;
    wire N__86640;
    wire N__86637;
    wire N__86626;
    wire N__86623;
    wire N__86620;
    wire N__86617;
    wire N__86614;
    wire N__86611;
    wire N__86608;
    wire N__86605;
    wire N__86602;
    wire N__86599;
    wire N__86596;
    wire N__86593;
    wire N__86590;
    wire N__86589;
    wire N__86586;
    wire N__86583;
    wire N__86580;
    wire N__86577;
    wire N__86572;
    wire N__86569;
    wire N__86566;
    wire N__86563;
    wire N__86560;
    wire N__86557;
    wire N__86554;
    wire N__86551;
    wire N__86548;
    wire N__86545;
    wire N__86542;
    wire N__86539;
    wire N__86536;
    wire N__86533;
    wire N__86530;
    wire N__86527;
    wire N__86524;
    wire N__86521;
    wire N__86518;
    wire N__86515;
    wire N__86512;
    wire N__86509;
    wire N__86506;
    wire N__86503;
    wire N__86500;
    wire N__86497;
    wire N__86494;
    wire N__86491;
    wire N__86488;
    wire N__86485;
    wire N__86482;
    wire N__86479;
    wire N__86476;
    wire N__86475;
    wire N__86474;
    wire N__86471;
    wire N__86470;
    wire N__86465;
    wire N__86462;
    wire N__86459;
    wire N__86452;
    wire N__86449;
    wire N__86446;
    wire N__86443;
    wire N__86440;
    wire N__86437;
    wire N__86434;
    wire N__86431;
    wire N__86428;
    wire N__86427;
    wire N__86426;
    wire N__86423;
    wire N__86420;
    wire N__86417;
    wire N__86414;
    wire N__86411;
    wire N__86408;
    wire N__86403;
    wire N__86400;
    wire N__86395;
    wire N__86392;
    wire N__86389;
    wire N__86386;
    wire N__86383;
    wire N__86380;
    wire N__86377;
    wire N__86374;
    wire N__86371;
    wire N__86368;
    wire N__86365;
    wire N__86362;
    wire N__86359;
    wire N__86356;
    wire N__86353;
    wire N__86350;
    wire N__86349;
    wire N__86348;
    wire N__86347;
    wire N__86344;
    wire N__86339;
    wire N__86338;
    wire N__86335;
    wire N__86334;
    wire N__86331;
    wire N__86328;
    wire N__86325;
    wire N__86322;
    wire N__86319;
    wire N__86314;
    wire N__86311;
    wire N__86302;
    wire N__86299;
    wire N__86296;
    wire N__86293;
    wire N__86290;
    wire N__86287;
    wire N__86284;
    wire N__86283;
    wire N__86280;
    wire N__86277;
    wire N__86272;
    wire N__86269;
    wire N__86266;
    wire N__86263;
    wire N__86260;
    wire N__86257;
    wire N__86254;
    wire N__86251;
    wire N__86248;
    wire N__86245;
    wire N__86242;
    wire N__86239;
    wire N__86236;
    wire N__86233;
    wire N__86230;
    wire N__86227;
    wire N__86224;
    wire N__86221;
    wire N__86218;
    wire N__86215;
    wire N__86212;
    wire N__86209;
    wire N__86206;
    wire N__86203;
    wire N__86200;
    wire N__86197;
    wire N__86194;
    wire N__86191;
    wire N__86188;
    wire N__86185;
    wire N__86182;
    wire N__86179;
    wire N__86176;
    wire N__86173;
    wire N__86170;
    wire N__86169;
    wire N__86166;
    wire N__86163;
    wire N__86162;
    wire N__86159;
    wire N__86156;
    wire N__86153;
    wire N__86150;
    wire N__86147;
    wire N__86140;
    wire N__86137;
    wire N__86136;
    wire N__86135;
    wire N__86132;
    wire N__86129;
    wire N__86126;
    wire N__86123;
    wire N__86120;
    wire N__86117;
    wire N__86112;
    wire N__86107;
    wire N__86104;
    wire N__86103;
    wire N__86100;
    wire N__86097;
    wire N__86096;
    wire N__86095;
    wire N__86094;
    wire N__86091;
    wire N__86088;
    wire N__86085;
    wire N__86080;
    wire N__86077;
    wire N__86074;
    wire N__86065;
    wire N__86062;
    wire N__86061;
    wire N__86058;
    wire N__86055;
    wire N__86050;
    wire N__86047;
    wire N__86044;
    wire N__86041;
    wire N__86040;
    wire N__86039;
    wire N__86038;
    wire N__86037;
    wire N__86036;
    wire N__86035;
    wire N__86034;
    wire N__86031;
    wire N__86018;
    wire N__86015;
    wire N__86010;
    wire N__86009;
    wire N__86006;
    wire N__86003;
    wire N__86000;
    wire N__85993;
    wire N__85992;
    wire N__85991;
    wire N__85990;
    wire N__85989;
    wire N__85986;
    wire N__85985;
    wire N__85984;
    wire N__85975;
    wire N__85972;
    wire N__85971;
    wire N__85970;
    wire N__85969;
    wire N__85968;
    wire N__85965;
    wire N__85964;
    wire N__85961;
    wire N__85958;
    wire N__85955;
    wire N__85952;
    wire N__85949;
    wire N__85948;
    wire N__85945;
    wire N__85942;
    wire N__85941;
    wire N__85936;
    wire N__85933;
    wire N__85932;
    wire N__85931;
    wire N__85930;
    wire N__85927;
    wire N__85922;
    wire N__85917;
    wire N__85914;
    wire N__85909;
    wire N__85904;
    wire N__85901;
    wire N__85900;
    wire N__85899;
    wire N__85896;
    wire N__85895;
    wire N__85892;
    wire N__85889;
    wire N__85886;
    wire N__85883;
    wire N__85878;
    wire N__85875;
    wire N__85862;
    wire N__85849;
    wire N__85846;
    wire N__85843;
    wire N__85840;
    wire N__85837;
    wire N__85834;
    wire N__85831;
    wire N__85828;
    wire N__85825;
    wire N__85822;
    wire N__85819;
    wire N__85816;
    wire N__85813;
    wire N__85810;
    wire N__85807;
    wire N__85804;
    wire N__85803;
    wire N__85800;
    wire N__85797;
    wire N__85796;
    wire N__85791;
    wire N__85788;
    wire N__85783;
    wire N__85780;
    wire N__85777;
    wire N__85776;
    wire N__85773;
    wire N__85770;
    wire N__85767;
    wire N__85762;
    wire N__85759;
    wire N__85756;
    wire N__85753;
    wire N__85750;
    wire N__85747;
    wire N__85744;
    wire N__85741;
    wire N__85738;
    wire N__85735;
    wire N__85732;
    wire N__85729;
    wire N__85726;
    wire N__85723;
    wire N__85720;
    wire N__85717;
    wire N__85714;
    wire N__85711;
    wire N__85708;
    wire N__85705;
    wire N__85702;
    wire N__85699;
    wire N__85696;
    wire N__85693;
    wire N__85690;
    wire N__85687;
    wire N__85684;
    wire N__85681;
    wire N__85678;
    wire N__85675;
    wire N__85672;
    wire N__85669;
    wire N__85666;
    wire N__85663;
    wire N__85660;
    wire N__85657;
    wire N__85654;
    wire N__85651;
    wire N__85648;
    wire N__85645;
    wire N__85644;
    wire N__85641;
    wire N__85638;
    wire N__85635;
    wire N__85632;
    wire N__85627;
    wire N__85624;
    wire N__85621;
    wire N__85618;
    wire N__85615;
    wire N__85612;
    wire N__85609;
    wire N__85606;
    wire N__85603;
    wire N__85600;
    wire N__85597;
    wire N__85594;
    wire N__85591;
    wire N__85588;
    wire N__85585;
    wire N__85582;
    wire N__85579;
    wire N__85576;
    wire N__85575;
    wire N__85574;
    wire N__85569;
    wire N__85566;
    wire N__85563;
    wire N__85560;
    wire N__85557;
    wire N__85556;
    wire N__85555;
    wire N__85552;
    wire N__85549;
    wire N__85546;
    wire N__85543;
    wire N__85540;
    wire N__85537;
    wire N__85528;
    wire N__85525;
    wire N__85522;
    wire N__85519;
    wire N__85516;
    wire N__85513;
    wire N__85510;
    wire N__85509;
    wire N__85506;
    wire N__85503;
    wire N__85498;
    wire N__85495;
    wire N__85492;
    wire N__85489;
    wire N__85486;
    wire N__85483;
    wire N__85480;
    wire N__85477;
    wire N__85474;
    wire N__85471;
    wire N__85468;
    wire N__85465;
    wire N__85462;
    wire N__85459;
    wire N__85456;
    wire N__85453;
    wire N__85450;
    wire N__85447;
    wire N__85444;
    wire N__85441;
    wire N__85438;
    wire N__85435;
    wire N__85432;
    wire N__85429;
    wire N__85426;
    wire N__85423;
    wire N__85422;
    wire N__85421;
    wire N__85418;
    wire N__85415;
    wire N__85412;
    wire N__85407;
    wire N__85404;
    wire N__85401;
    wire N__85398;
    wire N__85395;
    wire N__85390;
    wire N__85387;
    wire N__85384;
    wire N__85381;
    wire N__85378;
    wire N__85375;
    wire N__85372;
    wire N__85369;
    wire N__85366;
    wire N__85363;
    wire N__85360;
    wire N__85357;
    wire N__85354;
    wire N__85351;
    wire N__85348;
    wire N__85345;
    wire N__85342;
    wire N__85339;
    wire N__85336;
    wire N__85333;
    wire N__85330;
    wire N__85327;
    wire N__85324;
    wire N__85321;
    wire N__85318;
    wire N__85315;
    wire N__85312;
    wire N__85309;
    wire N__85306;
    wire N__85303;
    wire N__85300;
    wire N__85297;
    wire N__85296;
    wire N__85293;
    wire N__85290;
    wire N__85285;
    wire N__85282;
    wire N__85279;
    wire N__85276;
    wire N__85273;
    wire N__85270;
    wire N__85267;
    wire N__85266;
    wire N__85265;
    wire N__85262;
    wire N__85261;
    wire N__85258;
    wire N__85255;
    wire N__85250;
    wire N__85247;
    wire N__85244;
    wire N__85241;
    wire N__85238;
    wire N__85231;
    wire N__85230;
    wire N__85229;
    wire N__85228;
    wire N__85227;
    wire N__85226;
    wire N__85225;
    wire N__85224;
    wire N__85221;
    wire N__85218;
    wire N__85217;
    wire N__85216;
    wire N__85215;
    wire N__85204;
    wire N__85201;
    wire N__85198;
    wire N__85197;
    wire N__85196;
    wire N__85195;
    wire N__85194;
    wire N__85191;
    wire N__85186;
    wire N__85183;
    wire N__85180;
    wire N__85179;
    wire N__85178;
    wire N__85177;
    wire N__85176;
    wire N__85173;
    wire N__85172;
    wire N__85169;
    wire N__85166;
    wire N__85161;
    wire N__85160;
    wire N__85157;
    wire N__85152;
    wire N__85149;
    wire N__85146;
    wire N__85143;
    wire N__85136;
    wire N__85133;
    wire N__85130;
    wire N__85129;
    wire N__85126;
    wire N__85123;
    wire N__85120;
    wire N__85117;
    wire N__85116;
    wire N__85113;
    wire N__85110;
    wire N__85105;
    wire N__85100;
    wire N__85097;
    wire N__85094;
    wire N__85091;
    wire N__85090;
    wire N__85087;
    wire N__85084;
    wire N__85081;
    wire N__85078;
    wire N__85075;
    wire N__85066;
    wire N__85063;
    wire N__85058;
    wire N__85055;
    wire N__85052;
    wire N__85049;
    wire N__85044;
    wire N__85033;
    wire N__85024;
    wire N__85021;
    wire N__85020;
    wire N__85019;
    wire N__85018;
    wire N__85009;
    wire N__85008;
    wire N__85005;
    wire N__85004;
    wire N__85003;
    wire N__85000;
    wire N__84999;
    wire N__84998;
    wire N__84997;
    wire N__84994;
    wire N__84991;
    wire N__84988;
    wire N__84985;
    wire N__84982;
    wire N__84979;
    wire N__84976;
    wire N__84971;
    wire N__84968;
    wire N__84965;
    wire N__84962;
    wire N__84957;
    wire N__84952;
    wire N__84951;
    wire N__84948;
    wire N__84945;
    wire N__84942;
    wire N__84939;
    wire N__84936;
    wire N__84925;
    wire N__84924;
    wire N__84923;
    wire N__84922;
    wire N__84921;
    wire N__84912;
    wire N__84909;
    wire N__84906;
    wire N__84905;
    wire N__84904;
    wire N__84903;
    wire N__84902;
    wire N__84899;
    wire N__84896;
    wire N__84895;
    wire N__84890;
    wire N__84887;
    wire N__84884;
    wire N__84881;
    wire N__84878;
    wire N__84875;
    wire N__84870;
    wire N__84867;
    wire N__84866;
    wire N__84865;
    wire N__84864;
    wire N__84861;
    wire N__84856;
    wire N__84851;
    wire N__84844;
    wire N__84835;
    wire N__84834;
    wire N__84833;
    wire N__84832;
    wire N__84829;
    wire N__84828;
    wire N__84825;
    wire N__84822;
    wire N__84819;
    wire N__84816;
    wire N__84809;
    wire N__84802;
    wire N__84799;
    wire N__84796;
    wire N__84793;
    wire N__84790;
    wire N__84787;
    wire N__84784;
    wire N__84781;
    wire N__84778;
    wire N__84775;
    wire N__84772;
    wire N__84769;
    wire N__84766;
    wire N__84763;
    wire N__84760;
    wire N__84757;
    wire N__84754;
    wire N__84751;
    wire N__84748;
    wire N__84745;
    wire N__84742;
    wire N__84739;
    wire N__84736;
    wire N__84733;
    wire N__84730;
    wire N__84729;
    wire N__84726;
    wire N__84723;
    wire N__84718;
    wire N__84715;
    wire N__84712;
    wire N__84709;
    wire N__84706;
    wire N__84703;
    wire N__84700;
    wire N__84697;
    wire N__84694;
    wire N__84691;
    wire N__84688;
    wire N__84685;
    wire N__84682;
    wire N__84679;
    wire N__84678;
    wire N__84675;
    wire N__84674;
    wire N__84671;
    wire N__84668;
    wire N__84665;
    wire N__84658;
    wire N__84655;
    wire N__84652;
    wire N__84649;
    wire N__84646;
    wire N__84643;
    wire N__84640;
    wire N__84637;
    wire N__84634;
    wire N__84631;
    wire N__84628;
    wire N__84625;
    wire N__84622;
    wire N__84619;
    wire N__84616;
    wire N__84613;
    wire N__84612;
    wire N__84609;
    wire N__84606;
    wire N__84605;
    wire N__84602;
    wire N__84599;
    wire N__84596;
    wire N__84593;
    wire N__84590;
    wire N__84587;
    wire N__84580;
    wire N__84577;
    wire N__84576;
    wire N__84573;
    wire N__84572;
    wire N__84569;
    wire N__84566;
    wire N__84563;
    wire N__84556;
    wire N__84553;
    wire N__84550;
    wire N__84547;
    wire N__84544;
    wire N__84541;
    wire N__84538;
    wire N__84535;
    wire N__84532;
    wire N__84529;
    wire N__84526;
    wire N__84523;
    wire N__84520;
    wire N__84517;
    wire N__84514;
    wire N__84511;
    wire N__84508;
    wire N__84507;
    wire N__84506;
    wire N__84505;
    wire N__84504;
    wire N__84501;
    wire N__84500;
    wire N__84497;
    wire N__84490;
    wire N__84487;
    wire N__84484;
    wire N__84475;
    wire N__84472;
    wire N__84469;
    wire N__84466;
    wire N__84463;
    wire N__84460;
    wire N__84457;
    wire N__84454;
    wire N__84451;
    wire N__84448;
    wire N__84445;
    wire N__84442;
    wire N__84439;
    wire N__84436;
    wire N__84433;
    wire N__84430;
    wire N__84427;
    wire N__84424;
    wire N__84421;
    wire N__84418;
    wire N__84415;
    wire N__84412;
    wire N__84409;
    wire N__84406;
    wire N__84403;
    wire N__84400;
    wire N__84397;
    wire N__84394;
    wire N__84391;
    wire N__84388;
    wire N__84385;
    wire N__84382;
    wire N__84379;
    wire N__84376;
    wire N__84373;
    wire N__84370;
    wire N__84367;
    wire N__84364;
    wire N__84361;
    wire N__84358;
    wire N__84355;
    wire N__84352;
    wire N__84349;
    wire N__84346;
    wire N__84343;
    wire N__84340;
    wire N__84337;
    wire N__84334;
    wire N__84331;
    wire N__84328;
    wire N__84325;
    wire N__84322;
    wire N__84319;
    wire N__84316;
    wire N__84313;
    wire N__84310;
    wire N__84307;
    wire N__84304;
    wire N__84301;
    wire N__84298;
    wire N__84295;
    wire N__84292;
    wire N__84289;
    wire N__84288;
    wire N__84285;
    wire N__84282;
    wire N__84279;
    wire N__84274;
    wire N__84273;
    wire N__84272;
    wire N__84271;
    wire N__84268;
    wire N__84265;
    wire N__84260;
    wire N__84255;
    wire N__84250;
    wire N__84247;
    wire N__84244;
    wire N__84241;
    wire N__84240;
    wire N__84237;
    wire N__84236;
    wire N__84235;
    wire N__84234;
    wire N__84231;
    wire N__84230;
    wire N__84227;
    wire N__84224;
    wire N__84221;
    wire N__84220;
    wire N__84213;
    wire N__84212;
    wire N__84211;
    wire N__84206;
    wire N__84203;
    wire N__84200;
    wire N__84197;
    wire N__84192;
    wire N__84187;
    wire N__84184;
    wire N__84181;
    wire N__84176;
    wire N__84173;
    wire N__84168;
    wire N__84163;
    wire N__84160;
    wire N__84159;
    wire N__84156;
    wire N__84155;
    wire N__84154;
    wire N__84151;
    wire N__84146;
    wire N__84143;
    wire N__84140;
    wire N__84137;
    wire N__84134;
    wire N__84131;
    wire N__84128;
    wire N__84125;
    wire N__84120;
    wire N__84117;
    wire N__84112;
    wire N__84109;
    wire N__84106;
    wire N__84103;
    wire N__84100;
    wire N__84097;
    wire N__84094;
    wire N__84091;
    wire N__84088;
    wire N__84085;
    wire N__84082;
    wire N__84079;
    wire N__84076;
    wire N__84073;
    wire N__84070;
    wire N__84067;
    wire N__84064;
    wire N__84061;
    wire N__84058;
    wire N__84055;
    wire N__84052;
    wire N__84049;
    wire N__84046;
    wire N__84043;
    wire N__84040;
    wire N__84037;
    wire N__84034;
    wire N__84031;
    wire N__84028;
    wire N__84025;
    wire N__84022;
    wire N__84019;
    wire N__84016;
    wire N__84013;
    wire N__84012;
    wire N__84011;
    wire N__84010;
    wire N__84007;
    wire N__84004;
    wire N__84001;
    wire N__83998;
    wire N__83995;
    wire N__83992;
    wire N__83983;
    wire N__83980;
    wire N__83977;
    wire N__83974;
    wire N__83971;
    wire N__83970;
    wire N__83969;
    wire N__83966;
    wire N__83965;
    wire N__83964;
    wire N__83959;
    wire N__83956;
    wire N__83953;
    wire N__83950;
    wire N__83949;
    wire N__83946;
    wire N__83943;
    wire N__83940;
    wire N__83937;
    wire N__83934;
    wire N__83931;
    wire N__83926;
    wire N__83923;
    wire N__83914;
    wire N__83911;
    wire N__83910;
    wire N__83907;
    wire N__83904;
    wire N__83901;
    wire N__83896;
    wire N__83893;
    wire N__83892;
    wire N__83889;
    wire N__83888;
    wire N__83885;
    wire N__83884;
    wire N__83883;
    wire N__83880;
    wire N__83877;
    wire N__83872;
    wire N__83869;
    wire N__83866;
    wire N__83861;
    wire N__83856;
    wire N__83853;
    wire N__83848;
    wire N__83845;
    wire N__83842;
    wire N__83841;
    wire N__83840;
    wire N__83839;
    wire N__83838;
    wire N__83837;
    wire N__83834;
    wire N__83829;
    wire N__83826;
    wire N__83823;
    wire N__83820;
    wire N__83817;
    wire N__83814;
    wire N__83803;
    wire N__83802;
    wire N__83797;
    wire N__83796;
    wire N__83795;
    wire N__83794;
    wire N__83793;
    wire N__83792;
    wire N__83791;
    wire N__83790;
    wire N__83787;
    wire N__83784;
    wire N__83779;
    wire N__83776;
    wire N__83773;
    wire N__83770;
    wire N__83767;
    wire N__83764;
    wire N__83761;
    wire N__83758;
    wire N__83755;
    wire N__83750;
    wire N__83747;
    wire N__83742;
    wire N__83739;
    wire N__83736;
    wire N__83733;
    wire N__83722;
    wire N__83721;
    wire N__83720;
    wire N__83719;
    wire N__83718;
    wire N__83713;
    wire N__83708;
    wire N__83705;
    wire N__83700;
    wire N__83699;
    wire N__83696;
    wire N__83693;
    wire N__83690;
    wire N__83685;
    wire N__83680;
    wire N__83677;
    wire N__83674;
    wire N__83671;
    wire N__83668;
    wire N__83665;
    wire N__83662;
    wire N__83661;
    wire N__83658;
    wire N__83657;
    wire N__83652;
    wire N__83651;
    wire N__83648;
    wire N__83645;
    wire N__83642;
    wire N__83639;
    wire N__83636;
    wire N__83629;
    wire N__83626;
    wire N__83623;
    wire N__83620;
    wire N__83617;
    wire N__83616;
    wire N__83613;
    wire N__83610;
    wire N__83609;
    wire N__83606;
    wire N__83603;
    wire N__83600;
    wire N__83597;
    wire N__83594;
    wire N__83591;
    wire N__83584;
    wire N__83583;
    wire N__83582;
    wire N__83579;
    wire N__83578;
    wire N__83573;
    wire N__83568;
    wire N__83563;
    wire N__83560;
    wire N__83559;
    wire N__83554;
    wire N__83551;
    wire N__83548;
    wire N__83545;
    wire N__83542;
    wire N__83539;
    wire N__83536;
    wire N__83533;
    wire N__83530;
    wire N__83527;
    wire N__83526;
    wire N__83523;
    wire N__83520;
    wire N__83515;
    wire N__83512;
    wire N__83509;
    wire N__83506;
    wire N__83503;
    wire N__83500;
    wire N__83499;
    wire N__83496;
    wire N__83493;
    wire N__83488;
    wire N__83485;
    wire N__83484;
    wire N__83481;
    wire N__83478;
    wire N__83473;
    wire N__83470;
    wire N__83469;
    wire N__83468;
    wire N__83465;
    wire N__83462;
    wire N__83459;
    wire N__83452;
    wire N__83449;
    wire N__83446;
    wire N__83445;
    wire N__83442;
    wire N__83437;
    wire N__83434;
    wire N__83433;
    wire N__83430;
    wire N__83427;
    wire N__83424;
    wire N__83419;
    wire N__83416;
    wire N__83413;
    wire N__83410;
    wire N__83407;
    wire N__83404;
    wire N__83401;
    wire N__83398;
    wire N__83395;
    wire N__83392;
    wire N__83389;
    wire N__83386;
    wire N__83383;
    wire N__83380;
    wire N__83377;
    wire N__83374;
    wire N__83371;
    wire N__83368;
    wire N__83365;
    wire N__83362;
    wire N__83359;
    wire N__83356;
    wire N__83353;
    wire N__83350;
    wire N__83349;
    wire N__83348;
    wire N__83343;
    wire N__83340;
    wire N__83339;
    wire N__83338;
    wire N__83335;
    wire N__83332;
    wire N__83329;
    wire N__83326;
    wire N__83323;
    wire N__83320;
    wire N__83313;
    wire N__83310;
    wire N__83305;
    wire N__83302;
    wire N__83299;
    wire N__83296;
    wire N__83293;
    wire N__83290;
    wire N__83287;
    wire N__83284;
    wire N__83281;
    wire N__83278;
    wire N__83275;
    wire N__83272;
    wire N__83269;
    wire N__83266;
    wire N__83263;
    wire N__83260;
    wire N__83257;
    wire N__83254;
    wire N__83251;
    wire N__83248;
    wire N__83245;
    wire N__83242;
    wire N__83239;
    wire N__83236;
    wire N__83233;
    wire N__83230;
    wire N__83227;
    wire N__83224;
    wire N__83221;
    wire N__83218;
    wire N__83215;
    wire N__83212;
    wire N__83209;
    wire N__83206;
    wire N__83203;
    wire N__83200;
    wire N__83197;
    wire N__83194;
    wire N__83191;
    wire N__83188;
    wire N__83185;
    wire N__83182;
    wire N__83179;
    wire N__83176;
    wire N__83173;
    wire N__83170;
    wire N__83167;
    wire N__83164;
    wire N__83161;
    wire N__83158;
    wire N__83155;
    wire N__83152;
    wire N__83149;
    wire N__83146;
    wire N__83143;
    wire N__83140;
    wire N__83137;
    wire N__83134;
    wire N__83131;
    wire N__83128;
    wire N__83125;
    wire N__83122;
    wire N__83119;
    wire N__83116;
    wire N__83113;
    wire N__83110;
    wire N__83107;
    wire N__83104;
    wire N__83101;
    wire N__83098;
    wire N__83095;
    wire N__83092;
    wire N__83089;
    wire N__83086;
    wire N__83083;
    wire N__83080;
    wire N__83077;
    wire N__83074;
    wire N__83071;
    wire N__83068;
    wire N__83065;
    wire N__83062;
    wire N__83059;
    wire N__83056;
    wire N__83053;
    wire N__83050;
    wire N__83047;
    wire N__83044;
    wire N__83041;
    wire N__83038;
    wire N__83035;
    wire N__83032;
    wire N__83029;
    wire N__83026;
    wire N__83023;
    wire N__83020;
    wire N__83017;
    wire N__83014;
    wire N__83011;
    wire N__83008;
    wire N__83005;
    wire N__83002;
    wire N__82999;
    wire N__82996;
    wire N__82993;
    wire N__82990;
    wire N__82987;
    wire N__82984;
    wire N__82981;
    wire N__82978;
    wire N__82975;
    wire N__82972;
    wire N__82969;
    wire N__82966;
    wire N__82963;
    wire N__82960;
    wire N__82957;
    wire N__82954;
    wire N__82951;
    wire N__82948;
    wire N__82945;
    wire N__82942;
    wire N__82939;
    wire N__82936;
    wire N__82933;
    wire N__82930;
    wire N__82927;
    wire N__82924;
    wire N__82921;
    wire N__82918;
    wire N__82915;
    wire N__82912;
    wire N__82909;
    wire N__82906;
    wire N__82903;
    wire N__82900;
    wire N__82897;
    wire N__82894;
    wire N__82891;
    wire N__82888;
    wire N__82885;
    wire N__82882;
    wire N__82879;
    wire N__82876;
    wire N__82873;
    wire N__82870;
    wire N__82867;
    wire N__82864;
    wire N__82861;
    wire N__82858;
    wire N__82855;
    wire N__82852;
    wire N__82849;
    wire N__82846;
    wire N__82845;
    wire N__82842;
    wire N__82839;
    wire N__82836;
    wire N__82833;
    wire N__82830;
    wire N__82825;
    wire N__82822;
    wire N__82819;
    wire N__82816;
    wire N__82813;
    wire N__82810;
    wire N__82807;
    wire N__82804;
    wire N__82801;
    wire N__82798;
    wire N__82797;
    wire N__82796;
    wire N__82793;
    wire N__82790;
    wire N__82787;
    wire N__82782;
    wire N__82779;
    wire N__82776;
    wire N__82771;
    wire N__82768;
    wire N__82765;
    wire N__82762;
    wire N__82759;
    wire N__82756;
    wire N__82753;
    wire N__82752;
    wire N__82751;
    wire N__82750;
    wire N__82743;
    wire N__82742;
    wire N__82739;
    wire N__82736;
    wire N__82731;
    wire N__82730;
    wire N__82725;
    wire N__82722;
    wire N__82719;
    wire N__82714;
    wire N__82711;
    wire N__82708;
    wire N__82705;
    wire N__82702;
    wire N__82699;
    wire N__82696;
    wire N__82693;
    wire N__82690;
    wire N__82689;
    wire N__82686;
    wire N__82683;
    wire N__82680;
    wire N__82677;
    wire N__82674;
    wire N__82671;
    wire N__82666;
    wire N__82663;
    wire N__82660;
    wire N__82657;
    wire N__82654;
    wire N__82651;
    wire N__82648;
    wire N__82645;
    wire N__82642;
    wire N__82639;
    wire N__82636;
    wire N__82633;
    wire N__82630;
    wire N__82627;
    wire N__82624;
    wire N__82621;
    wire N__82618;
    wire N__82615;
    wire N__82612;
    wire N__82609;
    wire N__82606;
    wire N__82603;
    wire N__82600;
    wire N__82599;
    wire N__82598;
    wire N__82595;
    wire N__82592;
    wire N__82589;
    wire N__82582;
    wire N__82579;
    wire N__82576;
    wire N__82573;
    wire N__82570;
    wire N__82567;
    wire N__82564;
    wire N__82561;
    wire N__82558;
    wire N__82555;
    wire N__82552;
    wire N__82549;
    wire N__82546;
    wire N__82545;
    wire N__82544;
    wire N__82541;
    wire N__82538;
    wire N__82535;
    wire N__82528;
    wire N__82525;
    wire N__82522;
    wire N__82519;
    wire N__82516;
    wire N__82513;
    wire N__82510;
    wire N__82507;
    wire N__82504;
    wire N__82501;
    wire N__82498;
    wire N__82495;
    wire N__82492;
    wire N__82489;
    wire N__82486;
    wire N__82483;
    wire N__82480;
    wire N__82479;
    wire N__82476;
    wire N__82473;
    wire N__82468;
    wire N__82465;
    wire N__82462;
    wire N__82459;
    wire N__82456;
    wire N__82453;
    wire N__82450;
    wire N__82447;
    wire N__82444;
    wire N__82441;
    wire N__82438;
    wire N__82435;
    wire N__82432;
    wire N__82429;
    wire N__82428;
    wire N__82427;
    wire N__82426;
    wire N__82425;
    wire N__82422;
    wire N__82419;
    wire N__82416;
    wire N__82415;
    wire N__82412;
    wire N__82409;
    wire N__82404;
    wire N__82401;
    wire N__82396;
    wire N__82393;
    wire N__82390;
    wire N__82387;
    wire N__82382;
    wire N__82379;
    wire N__82376;
    wire N__82373;
    wire N__82366;
    wire N__82363;
    wire N__82362;
    wire N__82359;
    wire N__82356;
    wire N__82353;
    wire N__82350;
    wire N__82345;
    wire N__82342;
    wire N__82341;
    wire N__82340;
    wire N__82339;
    wire N__82336;
    wire N__82335;
    wire N__82334;
    wire N__82331;
    wire N__82328;
    wire N__82327;
    wire N__82324;
    wire N__82321;
    wire N__82316;
    wire N__82313;
    wire N__82312;
    wire N__82309;
    wire N__82306;
    wire N__82303;
    wire N__82296;
    wire N__82295;
    wire N__82294;
    wire N__82293;
    wire N__82292;
    wire N__82289;
    wire N__82288;
    wire N__82285;
    wire N__82282;
    wire N__82279;
    wire N__82276;
    wire N__82267;
    wire N__82264;
    wire N__82261;
    wire N__82256;
    wire N__82253;
    wire N__82250;
    wire N__82245;
    wire N__82242;
    wire N__82237;
    wire N__82234;
    wire N__82231;
    wire N__82222;
    wire N__82221;
    wire N__82220;
    wire N__82217;
    wire N__82216;
    wire N__82213;
    wire N__82212;
    wire N__82209;
    wire N__82206;
    wire N__82203;
    wire N__82202;
    wire N__82199;
    wire N__82198;
    wire N__82195;
    wire N__82194;
    wire N__82191;
    wire N__82186;
    wire N__82185;
    wire N__82182;
    wire N__82179;
    wire N__82176;
    wire N__82175;
    wire N__82170;
    wire N__82167;
    wire N__82164;
    wire N__82161;
    wire N__82160;
    wire N__82157;
    wire N__82152;
    wire N__82149;
    wire N__82148;
    wire N__82147;
    wire N__82146;
    wire N__82145;
    wire N__82142;
    wire N__82139;
    wire N__82134;
    wire N__82131;
    wire N__82128;
    wire N__82125;
    wire N__82122;
    wire N__82113;
    wire N__82110;
    wire N__82105;
    wire N__82102;
    wire N__82099;
    wire N__82096;
    wire N__82091;
    wire N__82086;
    wire N__82083;
    wire N__82080;
    wire N__82069;
    wire N__82066;
    wire N__82063;
    wire N__82060;
    wire N__82057;
    wire N__82054;
    wire N__82051;
    wire N__82048;
    wire N__82045;
    wire N__82042;
    wire N__82039;
    wire N__82036;
    wire N__82033;
    wire N__82030;
    wire N__82027;
    wire N__82024;
    wire N__82023;
    wire N__82020;
    wire N__82017;
    wire N__82016;
    wire N__82013;
    wire N__82010;
    wire N__82007;
    wire N__82000;
    wire N__81997;
    wire N__81994;
    wire N__81991;
    wire N__81988;
    wire N__81985;
    wire N__81982;
    wire N__81979;
    wire N__81976;
    wire N__81973;
    wire N__81970;
    wire N__81967;
    wire N__81964;
    wire N__81961;
    wire N__81958;
    wire N__81955;
    wire N__81952;
    wire N__81949;
    wire N__81946;
    wire N__81943;
    wire N__81940;
    wire N__81937;
    wire N__81934;
    wire N__81931;
    wire N__81928;
    wire N__81925;
    wire N__81922;
    wire N__81919;
    wire N__81916;
    wire N__81913;
    wire N__81910;
    wire N__81907;
    wire N__81904;
    wire N__81903;
    wire N__81902;
    wire N__81899;
    wire N__81896;
    wire N__81893;
    wire N__81890;
    wire N__81887;
    wire N__81882;
    wire N__81877;
    wire N__81874;
    wire N__81871;
    wire N__81868;
    wire N__81865;
    wire N__81862;
    wire N__81859;
    wire N__81856;
    wire N__81853;
    wire N__81850;
    wire N__81847;
    wire N__81844;
    wire N__81841;
    wire N__81838;
    wire N__81835;
    wire N__81832;
    wire N__81829;
    wire N__81826;
    wire N__81823;
    wire N__81822;
    wire N__81819;
    wire N__81816;
    wire N__81811;
    wire N__81808;
    wire N__81805;
    wire N__81804;
    wire N__81801;
    wire N__81798;
    wire N__81797;
    wire N__81794;
    wire N__81791;
    wire N__81788;
    wire N__81783;
    wire N__81780;
    wire N__81775;
    wire N__81772;
    wire N__81769;
    wire N__81766;
    wire N__81763;
    wire N__81760;
    wire N__81757;
    wire N__81754;
    wire N__81751;
    wire N__81748;
    wire N__81745;
    wire N__81742;
    wire N__81739;
    wire N__81736;
    wire N__81733;
    wire N__81730;
    wire N__81727;
    wire N__81724;
    wire N__81721;
    wire N__81718;
    wire N__81717;
    wire N__81714;
    wire N__81711;
    wire N__81708;
    wire N__81703;
    wire N__81700;
    wire N__81697;
    wire N__81694;
    wire N__81691;
    wire N__81688;
    wire N__81685;
    wire N__81682;
    wire N__81681;
    wire N__81678;
    wire N__81675;
    wire N__81670;
    wire N__81667;
    wire N__81664;
    wire N__81661;
    wire N__81658;
    wire N__81655;
    wire N__81652;
    wire N__81649;
    wire N__81646;
    wire N__81643;
    wire N__81640;
    wire N__81637;
    wire N__81634;
    wire N__81631;
    wire N__81628;
    wire N__81625;
    wire N__81622;
    wire N__81619;
    wire N__81616;
    wire N__81613;
    wire N__81610;
    wire N__81607;
    wire N__81604;
    wire N__81601;
    wire N__81598;
    wire N__81595;
    wire N__81592;
    wire N__81589;
    wire N__81588;
    wire N__81587;
    wire N__81586;
    wire N__81583;
    wire N__81580;
    wire N__81577;
    wire N__81574;
    wire N__81571;
    wire N__81568;
    wire N__81565;
    wire N__81558;
    wire N__81553;
    wire N__81552;
    wire N__81551;
    wire N__81550;
    wire N__81549;
    wire N__81544;
    wire N__81541;
    wire N__81540;
    wire N__81539;
    wire N__81536;
    wire N__81533;
    wire N__81532;
    wire N__81527;
    wire N__81526;
    wire N__81523;
    wire N__81520;
    wire N__81515;
    wire N__81512;
    wire N__81509;
    wire N__81506;
    wire N__81499;
    wire N__81490;
    wire N__81489;
    wire N__81486;
    wire N__81483;
    wire N__81480;
    wire N__81479;
    wire N__81478;
    wire N__81475;
    wire N__81472;
    wire N__81469;
    wire N__81466;
    wire N__81463;
    wire N__81460;
    wire N__81455;
    wire N__81452;
    wire N__81445;
    wire N__81444;
    wire N__81443;
    wire N__81442;
    wire N__81441;
    wire N__81440;
    wire N__81437;
    wire N__81432;
    wire N__81429;
    wire N__81424;
    wire N__81423;
    wire N__81418;
    wire N__81415;
    wire N__81414;
    wire N__81411;
    wire N__81408;
    wire N__81403;
    wire N__81400;
    wire N__81397;
    wire N__81394;
    wire N__81391;
    wire N__81382;
    wire N__81379;
    wire N__81376;
    wire N__81373;
    wire N__81370;
    wire N__81367;
    wire N__81364;
    wire N__81363;
    wire N__81360;
    wire N__81357;
    wire N__81354;
    wire N__81351;
    wire N__81346;
    wire N__81343;
    wire N__81340;
    wire N__81337;
    wire N__81334;
    wire N__81333;
    wire N__81332;
    wire N__81331;
    wire N__81328;
    wire N__81327;
    wire N__81324;
    wire N__81323;
    wire N__81322;
    wire N__81319;
    wire N__81316;
    wire N__81313;
    wire N__81310;
    wire N__81307;
    wire N__81304;
    wire N__81301;
    wire N__81298;
    wire N__81295;
    wire N__81290;
    wire N__81289;
    wire N__81288;
    wire N__81285;
    wire N__81282;
    wire N__81279;
    wire N__81272;
    wire N__81269;
    wire N__81266;
    wire N__81261;
    wire N__81250;
    wire N__81247;
    wire N__81246;
    wire N__81243;
    wire N__81240;
    wire N__81237;
    wire N__81234;
    wire N__81229;
    wire N__81226;
    wire N__81223;
    wire N__81220;
    wire N__81217;
    wire N__81214;
    wire N__81211;
    wire N__81208;
    wire N__81205;
    wire N__81202;
    wire N__81199;
    wire N__81196;
    wire N__81193;
    wire N__81190;
    wire N__81187;
    wire N__81184;
    wire N__81181;
    wire N__81178;
    wire N__81175;
    wire N__81172;
    wire N__81169;
    wire N__81166;
    wire N__81163;
    wire N__81160;
    wire N__81157;
    wire N__81154;
    wire N__81151;
    wire N__81148;
    wire N__81145;
    wire N__81142;
    wire N__81139;
    wire N__81138;
    wire N__81137;
    wire N__81134;
    wire N__81133;
    wire N__81132;
    wire N__81129;
    wire N__81126;
    wire N__81125;
    wire N__81124;
    wire N__81117;
    wire N__81112;
    wire N__81107;
    wire N__81104;
    wire N__81101;
    wire N__81094;
    wire N__81093;
    wire N__81092;
    wire N__81087;
    wire N__81084;
    wire N__81083;
    wire N__81082;
    wire N__81079;
    wire N__81076;
    wire N__81073;
    wire N__81070;
    wire N__81065;
    wire N__81058;
    wire N__81057;
    wire N__81056;
    wire N__81055;
    wire N__81054;
    wire N__81051;
    wire N__81048;
    wire N__81045;
    wire N__81038;
    wire N__81033;
    wire N__81032;
    wire N__81029;
    wire N__81028;
    wire N__81025;
    wire N__81022;
    wire N__81019;
    wire N__81016;
    wire N__81013;
    wire N__81010;
    wire N__81007;
    wire N__80998;
    wire N__80995;
    wire N__80994;
    wire N__80991;
    wire N__80990;
    wire N__80987;
    wire N__80984;
    wire N__80981;
    wire N__80974;
    wire N__80971;
    wire N__80968;
    wire N__80965;
    wire N__80962;
    wire N__80959;
    wire N__80956;
    wire N__80953;
    wire N__80950;
    wire N__80947;
    wire N__80944;
    wire N__80941;
    wire N__80938;
    wire N__80935;
    wire N__80932;
    wire N__80929;
    wire N__80926;
    wire N__80923;
    wire N__80920;
    wire N__80917;
    wire N__80914;
    wire N__80911;
    wire N__80908;
    wire N__80905;
    wire N__80902;
    wire N__80899;
    wire N__80896;
    wire N__80893;
    wire N__80890;
    wire N__80887;
    wire N__80884;
    wire N__80881;
    wire N__80878;
    wire N__80875;
    wire N__80872;
    wire N__80869;
    wire N__80868;
    wire N__80865;
    wire N__80864;
    wire N__80861;
    wire N__80858;
    wire N__80855;
    wire N__80852;
    wire N__80845;
    wire N__80842;
    wire N__80841;
    wire N__80838;
    wire N__80835;
    wire N__80832;
    wire N__80829;
    wire N__80824;
    wire N__80823;
    wire N__80822;
    wire N__80821;
    wire N__80814;
    wire N__80811;
    wire N__80808;
    wire N__80803;
    wire N__80800;
    wire N__80799;
    wire N__80796;
    wire N__80793;
    wire N__80790;
    wire N__80785;
    wire N__80782;
    wire N__80779;
    wire N__80776;
    wire N__80775;
    wire N__80774;
    wire N__80771;
    wire N__80768;
    wire N__80765;
    wire N__80760;
    wire N__80757;
    wire N__80754;
    wire N__80749;
    wire N__80746;
    wire N__80743;
    wire N__80740;
    wire N__80737;
    wire N__80734;
    wire N__80731;
    wire N__80728;
    wire N__80725;
    wire N__80722;
    wire N__80719;
    wire N__80716;
    wire N__80713;
    wire N__80710;
    wire N__80707;
    wire N__80704;
    wire N__80701;
    wire N__80698;
    wire N__80695;
    wire N__80692;
    wire N__80689;
    wire N__80686;
    wire N__80683;
    wire N__80680;
    wire N__80677;
    wire N__80674;
    wire N__80673;
    wire N__80672;
    wire N__80669;
    wire N__80666;
    wire N__80663;
    wire N__80658;
    wire N__80655;
    wire N__80652;
    wire N__80647;
    wire N__80644;
    wire N__80641;
    wire N__80638;
    wire N__80635;
    wire N__80632;
    wire N__80629;
    wire N__80626;
    wire N__80623;
    wire N__80620;
    wire N__80617;
    wire N__80614;
    wire N__80611;
    wire N__80608;
    wire N__80605;
    wire N__80602;
    wire N__80599;
    wire N__80596;
    wire N__80593;
    wire N__80590;
    wire N__80587;
    wire N__80584;
    wire N__80583;
    wire N__80580;
    wire N__80579;
    wire N__80576;
    wire N__80573;
    wire N__80570;
    wire N__80567;
    wire N__80564;
    wire N__80561;
    wire N__80558;
    wire N__80553;
    wire N__80548;
    wire N__80545;
    wire N__80544;
    wire N__80543;
    wire N__80540;
    wire N__80539;
    wire N__80538;
    wire N__80535;
    wire N__80532;
    wire N__80529;
    wire N__80526;
    wire N__80523;
    wire N__80522;
    wire N__80517;
    wire N__80514;
    wire N__80511;
    wire N__80508;
    wire N__80505;
    wire N__80502;
    wire N__80497;
    wire N__80494;
    wire N__80491;
    wire N__80488;
    wire N__80485;
    wire N__80476;
    wire N__80475;
    wire N__80474;
    wire N__80471;
    wire N__80468;
    wire N__80465;
    wire N__80462;
    wire N__80459;
    wire N__80456;
    wire N__80455;
    wire N__80452;
    wire N__80451;
    wire N__80450;
    wire N__80449;
    wire N__80446;
    wire N__80443;
    wire N__80440;
    wire N__80437;
    wire N__80430;
    wire N__80419;
    wire N__80416;
    wire N__80415;
    wire N__80412;
    wire N__80409;
    wire N__80406;
    wire N__80405;
    wire N__80402;
    wire N__80401;
    wire N__80400;
    wire N__80397;
    wire N__80394;
    wire N__80391;
    wire N__80386;
    wire N__80377;
    wire N__80374;
    wire N__80371;
    wire N__80368;
    wire N__80365;
    wire N__80362;
    wire N__80359;
    wire N__80356;
    wire N__80355;
    wire N__80354;
    wire N__80351;
    wire N__80346;
    wire N__80345;
    wire N__80342;
    wire N__80339;
    wire N__80336;
    wire N__80335;
    wire N__80334;
    wire N__80329;
    wire N__80326;
    wire N__80321;
    wire N__80314;
    wire N__80311;
    wire N__80308;
    wire N__80305;
    wire N__80302;
    wire N__80299;
    wire N__80296;
    wire N__80293;
    wire N__80290;
    wire N__80287;
    wire N__80284;
    wire N__80281;
    wire N__80278;
    wire N__80275;
    wire N__80272;
    wire N__80269;
    wire N__80266;
    wire N__80263;
    wire N__80260;
    wire N__80257;
    wire N__80254;
    wire N__80251;
    wire N__80248;
    wire N__80245;
    wire N__80242;
    wire N__80239;
    wire N__80236;
    wire N__80233;
    wire N__80230;
    wire N__80227;
    wire N__80224;
    wire N__80221;
    wire N__80218;
    wire N__80215;
    wire N__80212;
    wire N__80209;
    wire N__80206;
    wire N__80203;
    wire N__80200;
    wire N__80197;
    wire N__80194;
    wire N__80191;
    wire N__80188;
    wire N__80185;
    wire N__80182;
    wire N__80179;
    wire N__80176;
    wire N__80173;
    wire N__80170;
    wire N__80167;
    wire N__80164;
    wire N__80161;
    wire N__80158;
    wire N__80155;
    wire N__80152;
    wire N__80149;
    wire N__80146;
    wire N__80143;
    wire N__80140;
    wire N__80137;
    wire N__80134;
    wire N__80131;
    wire N__80128;
    wire N__80125;
    wire N__80122;
    wire N__80119;
    wire N__80116;
    wire N__80113;
    wire N__80110;
    wire N__80107;
    wire N__80104;
    wire N__80101;
    wire N__80098;
    wire N__80095;
    wire N__80092;
    wire N__80089;
    wire N__80086;
    wire N__80083;
    wire N__80080;
    wire N__80077;
    wire N__80074;
    wire N__80071;
    wire N__80068;
    wire N__80065;
    wire N__80062;
    wire N__80059;
    wire N__80056;
    wire N__80053;
    wire N__80050;
    wire N__80047;
    wire N__80044;
    wire N__80041;
    wire N__80038;
    wire N__80035;
    wire N__80032;
    wire N__80029;
    wire N__80026;
    wire N__80023;
    wire N__80020;
    wire N__80017;
    wire N__80014;
    wire N__80011;
    wire N__80010;
    wire N__80007;
    wire N__80004;
    wire N__79999;
    wire N__79996;
    wire N__79993;
    wire N__79990;
    wire N__79987;
    wire N__79984;
    wire N__79981;
    wire N__79978;
    wire N__79975;
    wire N__79972;
    wire N__79969;
    wire N__79966;
    wire N__79963;
    wire N__79960;
    wire N__79957;
    wire N__79954;
    wire N__79951;
    wire N__79948;
    wire N__79945;
    wire N__79942;
    wire N__79939;
    wire N__79936;
    wire N__79933;
    wire N__79930;
    wire N__79929;
    wire N__79926;
    wire N__79923;
    wire N__79920;
    wire N__79917;
    wire N__79916;
    wire N__79913;
    wire N__79910;
    wire N__79907;
    wire N__79900;
    wire N__79897;
    wire N__79894;
    wire N__79893;
    wire N__79890;
    wire N__79887;
    wire N__79882;
    wire N__79879;
    wire N__79876;
    wire N__79873;
    wire N__79870;
    wire N__79867;
    wire N__79864;
    wire N__79861;
    wire N__79858;
    wire N__79855;
    wire N__79852;
    wire N__79849;
    wire N__79846;
    wire N__79843;
    wire N__79840;
    wire N__79837;
    wire N__79834;
    wire N__79831;
    wire N__79830;
    wire N__79827;
    wire N__79824;
    wire N__79823;
    wire N__79820;
    wire N__79817;
    wire N__79814;
    wire N__79811;
    wire N__79808;
    wire N__79805;
    wire N__79798;
    wire N__79795;
    wire N__79792;
    wire N__79789;
    wire N__79786;
    wire N__79785;
    wire N__79782;
    wire N__79779;
    wire N__79774;
    wire N__79771;
    wire N__79768;
    wire N__79765;
    wire N__79762;
    wire N__79761;
    wire N__79758;
    wire N__79755;
    wire N__79754;
    wire N__79751;
    wire N__79748;
    wire N__79745;
    wire N__79744;
    wire N__79741;
    wire N__79738;
    wire N__79735;
    wire N__79732;
    wire N__79729;
    wire N__79726;
    wire N__79723;
    wire N__79714;
    wire N__79711;
    wire N__79708;
    wire N__79705;
    wire N__79702;
    wire N__79699;
    wire N__79696;
    wire N__79693;
    wire N__79690;
    wire N__79689;
    wire N__79688;
    wire N__79685;
    wire N__79682;
    wire N__79679;
    wire N__79678;
    wire N__79677;
    wire N__79676;
    wire N__79675;
    wire N__79674;
    wire N__79673;
    wire N__79670;
    wire N__79667;
    wire N__79658;
    wire N__79651;
    wire N__79642;
    wire N__79639;
    wire N__79638;
    wire N__79635;
    wire N__79632;
    wire N__79629;
    wire N__79626;
    wire N__79623;
    wire N__79620;
    wire N__79617;
    wire N__79614;
    wire N__79609;
    wire N__79606;
    wire N__79603;
    wire N__79600;
    wire N__79597;
    wire N__79596;
    wire N__79595;
    wire N__79592;
    wire N__79587;
    wire N__79586;
    wire N__79585;
    wire N__79584;
    wire N__79579;
    wire N__79572;
    wire N__79567;
    wire N__79564;
    wire N__79563;
    wire N__79560;
    wire N__79557;
    wire N__79556;
    wire N__79555;
    wire N__79552;
    wire N__79551;
    wire N__79550;
    wire N__79549;
    wire N__79548;
    wire N__79547;
    wire N__79546;
    wire N__79545;
    wire N__79544;
    wire N__79543;
    wire N__79542;
    wire N__79541;
    wire N__79538;
    wire N__79533;
    wire N__79532;
    wire N__79531;
    wire N__79530;
    wire N__79529;
    wire N__79528;
    wire N__79527;
    wire N__79526;
    wire N__79525;
    wire N__79522;
    wire N__79519;
    wire N__79512;
    wire N__79511;
    wire N__79510;
    wire N__79499;
    wire N__79498;
    wire N__79497;
    wire N__79496;
    wire N__79493;
    wire N__79490;
    wire N__79487;
    wire N__79484;
    wire N__79483;
    wire N__79482;
    wire N__79479;
    wire N__79476;
    wire N__79467;
    wire N__79466;
    wire N__79465;
    wire N__79464;
    wire N__79459;
    wire N__79456;
    wire N__79455;
    wire N__79452;
    wire N__79449;
    wire N__79446;
    wire N__79443;
    wire N__79440;
    wire N__79437;
    wire N__79432;
    wire N__79427;
    wire N__79422;
    wire N__79417;
    wire N__79416;
    wire N__79415;
    wire N__79412;
    wire N__79409;
    wire N__79406;
    wire N__79399;
    wire N__79398;
    wire N__79397;
    wire N__79396;
    wire N__79393;
    wire N__79392;
    wire N__79391;
    wire N__79390;
    wire N__79389;
    wire N__79386;
    wire N__79383;
    wire N__79380;
    wire N__79375;
    wire N__79366;
    wire N__79359;
    wire N__79356;
    wire N__79353;
    wire N__79348;
    wire N__79343;
    wire N__79336;
    wire N__79335;
    wire N__79334;
    wire N__79331;
    wire N__79328;
    wire N__79325;
    wire N__79322;
    wire N__79321;
    wire N__79320;
    wire N__79317;
    wire N__79314;
    wire N__79311;
    wire N__79300;
    wire N__79291;
    wire N__79286;
    wire N__79277;
    wire N__79272;
    wire N__79269;
    wire N__79252;
    wire N__79249;
    wire N__79248;
    wire N__79245;
    wire N__79242;
    wire N__79239;
    wire N__79236;
    wire N__79233;
    wire N__79230;
    wire N__79227;
    wire N__79224;
    wire N__79221;
    wire N__79218;
    wire N__79213;
    wire N__79210;
    wire N__79207;
    wire N__79204;
    wire N__79201;
    wire N__79198;
    wire N__79195;
    wire N__79192;
    wire N__79191;
    wire N__79188;
    wire N__79185;
    wire N__79184;
    wire N__79181;
    wire N__79178;
    wire N__79175;
    wire N__79172;
    wire N__79167;
    wire N__79162;
    wire N__79159;
    wire N__79156;
    wire N__79153;
    wire N__79150;
    wire N__79147;
    wire N__79144;
    wire N__79141;
    wire N__79138;
    wire N__79135;
    wire N__79132;
    wire N__79129;
    wire N__79126;
    wire N__79123;
    wire N__79120;
    wire N__79117;
    wire N__79114;
    wire N__79111;
    wire N__79108;
    wire N__79105;
    wire N__79102;
    wire N__79101;
    wire N__79098;
    wire N__79095;
    wire N__79092;
    wire N__79089;
    wire N__79086;
    wire N__79081;
    wire N__79080;
    wire N__79079;
    wire N__79076;
    wire N__79075;
    wire N__79072;
    wire N__79069;
    wire N__79066;
    wire N__79063;
    wire N__79060;
    wire N__79057;
    wire N__79054;
    wire N__79051;
    wire N__79048;
    wire N__79045;
    wire N__79036;
    wire N__79033;
    wire N__79030;
    wire N__79027;
    wire N__79024;
    wire N__79021;
    wire N__79018;
    wire N__79015;
    wire N__79012;
    wire N__79009;
    wire N__79006;
    wire N__79003;
    wire N__79002;
    wire N__78999;
    wire N__78996;
    wire N__78993;
    wire N__78988;
    wire N__78985;
    wire N__78982;
    wire N__78979;
    wire N__78976;
    wire N__78973;
    wire N__78970;
    wire N__78969;
    wire N__78966;
    wire N__78963;
    wire N__78958;
    wire N__78955;
    wire N__78952;
    wire N__78949;
    wire N__78946;
    wire N__78943;
    wire N__78940;
    wire N__78937;
    wire N__78934;
    wire N__78931;
    wire N__78928;
    wire N__78925;
    wire N__78922;
    wire N__78919;
    wire N__78916;
    wire N__78913;
    wire N__78910;
    wire N__78907;
    wire N__78904;
    wire N__78901;
    wire N__78898;
    wire N__78895;
    wire N__78892;
    wire N__78889;
    wire N__78886;
    wire N__78883;
    wire N__78880;
    wire N__78877;
    wire N__78874;
    wire N__78871;
    wire N__78868;
    wire N__78865;
    wire N__78862;
    wire N__78859;
    wire N__78856;
    wire N__78853;
    wire N__78850;
    wire N__78847;
    wire N__78844;
    wire N__78841;
    wire N__78838;
    wire N__78835;
    wire N__78832;
    wire N__78829;
    wire N__78828;
    wire N__78825;
    wire N__78822;
    wire N__78819;
    wire N__78816;
    wire N__78813;
    wire N__78810;
    wire N__78805;
    wire N__78802;
    wire N__78799;
    wire N__78798;
    wire N__78797;
    wire N__78794;
    wire N__78793;
    wire N__78790;
    wire N__78787;
    wire N__78786;
    wire N__78783;
    wire N__78780;
    wire N__78779;
    wire N__78778;
    wire N__78775;
    wire N__78772;
    wire N__78769;
    wire N__78764;
    wire N__78759;
    wire N__78754;
    wire N__78745;
    wire N__78742;
    wire N__78739;
    wire N__78736;
    wire N__78733;
    wire N__78730;
    wire N__78727;
    wire N__78724;
    wire N__78721;
    wire N__78718;
    wire N__78715;
    wire N__78712;
    wire N__78709;
    wire N__78706;
    wire N__78703;
    wire N__78700;
    wire N__78697;
    wire N__78694;
    wire N__78691;
    wire N__78688;
    wire N__78687;
    wire N__78684;
    wire N__78681;
    wire N__78676;
    wire N__78673;
    wire N__78670;
    wire N__78667;
    wire N__78664;
    wire N__78661;
    wire N__78658;
    wire N__78655;
    wire N__78652;
    wire N__78649;
    wire N__78646;
    wire N__78643;
    wire N__78640;
    wire N__78637;
    wire N__78634;
    wire N__78631;
    wire N__78628;
    wire N__78625;
    wire N__78622;
    wire N__78619;
    wire N__78616;
    wire N__78613;
    wire N__78610;
    wire N__78607;
    wire N__78604;
    wire N__78601;
    wire N__78598;
    wire N__78595;
    wire N__78592;
    wire N__78589;
    wire N__78586;
    wire N__78583;
    wire N__78580;
    wire N__78577;
    wire N__78574;
    wire N__78571;
    wire N__78568;
    wire N__78565;
    wire N__78562;
    wire N__78559;
    wire N__78556;
    wire N__78553;
    wire N__78550;
    wire N__78547;
    wire N__78544;
    wire N__78541;
    wire N__78538;
    wire N__78535;
    wire N__78532;
    wire N__78531;
    wire N__78528;
    wire N__78525;
    wire N__78520;
    wire N__78519;
    wire N__78516;
    wire N__78513;
    wire N__78510;
    wire N__78509;
    wire N__78508;
    wire N__78505;
    wire N__78502;
    wire N__78497;
    wire N__78492;
    wire N__78489;
    wire N__78486;
    wire N__78483;
    wire N__78478;
    wire N__78475;
    wire N__78474;
    wire N__78473;
    wire N__78472;
    wire N__78469;
    wire N__78466;
    wire N__78463;
    wire N__78460;
    wire N__78457;
    wire N__78454;
    wire N__78451;
    wire N__78448;
    wire N__78447;
    wire N__78446;
    wire N__78443;
    wire N__78440;
    wire N__78437;
    wire N__78434;
    wire N__78431;
    wire N__78428;
    wire N__78415;
    wire N__78412;
    wire N__78409;
    wire N__78406;
    wire N__78403;
    wire N__78400;
    wire N__78397;
    wire N__78394;
    wire N__78391;
    wire N__78388;
    wire N__78385;
    wire N__78382;
    wire N__78379;
    wire N__78376;
    wire N__78373;
    wire N__78370;
    wire N__78367;
    wire N__78364;
    wire N__78361;
    wire N__78358;
    wire N__78355;
    wire N__78352;
    wire N__78351;
    wire N__78350;
    wire N__78347;
    wire N__78344;
    wire N__78339;
    wire N__78334;
    wire N__78331;
    wire N__78328;
    wire N__78325;
    wire N__78322;
    wire N__78319;
    wire N__78316;
    wire N__78313;
    wire N__78310;
    wire N__78307;
    wire N__78304;
    wire N__78301;
    wire N__78298;
    wire N__78295;
    wire N__78292;
    wire N__78289;
    wire N__78286;
    wire N__78283;
    wire N__78280;
    wire N__78277;
    wire N__78274;
    wire N__78271;
    wire N__78268;
    wire N__78265;
    wire N__78262;
    wire N__78259;
    wire N__78256;
    wire N__78253;
    wire N__78250;
    wire N__78247;
    wire N__78244;
    wire N__78241;
    wire N__78238;
    wire N__78235;
    wire N__78232;
    wire N__78229;
    wire N__78226;
    wire N__78223;
    wire N__78220;
    wire N__78217;
    wire N__78214;
    wire N__78211;
    wire N__78210;
    wire N__78207;
    wire N__78204;
    wire N__78199;
    wire N__78196;
    wire N__78193;
    wire N__78190;
    wire N__78187;
    wire N__78184;
    wire N__78181;
    wire N__78178;
    wire N__78175;
    wire N__78172;
    wire N__78169;
    wire N__78166;
    wire N__78163;
    wire N__78162;
    wire N__78161;
    wire N__78160;
    wire N__78159;
    wire N__78156;
    wire N__78153;
    wire N__78148;
    wire N__78145;
    wire N__78138;
    wire N__78133;
    wire N__78132;
    wire N__78131;
    wire N__78126;
    wire N__78123;
    wire N__78120;
    wire N__78115;
    wire N__78112;
    wire N__78109;
    wire N__78106;
    wire N__78103;
    wire N__78102;
    wire N__78099;
    wire N__78096;
    wire N__78093;
    wire N__78090;
    wire N__78085;
    wire N__78082;
    wire N__78079;
    wire N__78076;
    wire N__78073;
    wire N__78070;
    wire N__78067;
    wire N__78064;
    wire N__78061;
    wire N__78060;
    wire N__78057;
    wire N__78054;
    wire N__78051;
    wire N__78048;
    wire N__78045;
    wire N__78042;
    wire N__78039;
    wire N__78034;
    wire N__78031;
    wire N__78028;
    wire N__78025;
    wire N__78022;
    wire N__78019;
    wire N__78016;
    wire N__78013;
    wire N__78010;
    wire N__78007;
    wire N__78004;
    wire N__78001;
    wire N__77998;
    wire N__77995;
    wire N__77992;
    wire N__77989;
    wire N__77986;
    wire N__77983;
    wire N__77980;
    wire N__77977;
    wire N__77974;
    wire N__77971;
    wire N__77968;
    wire N__77965;
    wire N__77962;
    wire N__77959;
    wire N__77956;
    wire N__77955;
    wire N__77952;
    wire N__77949;
    wire N__77944;
    wire N__77941;
    wire N__77938;
    wire N__77935;
    wire N__77932;
    wire N__77929;
    wire N__77926;
    wire N__77923;
    wire N__77920;
    wire N__77917;
    wire N__77914;
    wire N__77911;
    wire N__77908;
    wire N__77907;
    wire N__77904;
    wire N__77903;
    wire N__77902;
    wire N__77899;
    wire N__77898;
    wire N__77895;
    wire N__77892;
    wire N__77887;
    wire N__77884;
    wire N__77881;
    wire N__77876;
    wire N__77873;
    wire N__77872;
    wire N__77871;
    wire N__77868;
    wire N__77865;
    wire N__77862;
    wire N__77859;
    wire N__77856;
    wire N__77853;
    wire N__77850;
    wire N__77847;
    wire N__77844;
    wire N__77833;
    wire N__77830;
    wire N__77827;
    wire N__77826;
    wire N__77825;
    wire N__77824;
    wire N__77823;
    wire N__77822;
    wire N__77821;
    wire N__77820;
    wire N__77817;
    wire N__77816;
    wire N__77815;
    wire N__77812;
    wire N__77809;
    wire N__77806;
    wire N__77805;
    wire N__77804;
    wire N__77801;
    wire N__77796;
    wire N__77793;
    wire N__77790;
    wire N__77785;
    wire N__77782;
    wire N__77775;
    wire N__77774;
    wire N__77771;
    wire N__77768;
    wire N__77765;
    wire N__77764;
    wire N__77757;
    wire N__77752;
    wire N__77749;
    wire N__77746;
    wire N__77743;
    wire N__77740;
    wire N__77737;
    wire N__77734;
    wire N__77729;
    wire N__77720;
    wire N__77717;
    wire N__77710;
    wire N__77707;
    wire N__77706;
    wire N__77703;
    wire N__77702;
    wire N__77699;
    wire N__77696;
    wire N__77693;
    wire N__77690;
    wire N__77687;
    wire N__77684;
    wire N__77681;
    wire N__77674;
    wire N__77671;
    wire N__77670;
    wire N__77667;
    wire N__77664;
    wire N__77661;
    wire N__77656;
    wire N__77653;
    wire N__77652;
    wire N__77651;
    wire N__77648;
    wire N__77645;
    wire N__77642;
    wire N__77639;
    wire N__77636;
    wire N__77633;
    wire N__77632;
    wire N__77629;
    wire N__77624;
    wire N__77621;
    wire N__77616;
    wire N__77611;
    wire N__77608;
    wire N__77607;
    wire N__77606;
    wire N__77605;
    wire N__77604;
    wire N__77601;
    wire N__77598;
    wire N__77591;
    wire N__77588;
    wire N__77585;
    wire N__77582;
    wire N__77581;
    wire N__77578;
    wire N__77575;
    wire N__77572;
    wire N__77569;
    wire N__77564;
    wire N__77557;
    wire N__77556;
    wire N__77553;
    wire N__77552;
    wire N__77551;
    wire N__77548;
    wire N__77547;
    wire N__77544;
    wire N__77541;
    wire N__77534;
    wire N__77533;
    wire N__77530;
    wire N__77529;
    wire N__77526;
    wire N__77523;
    wire N__77520;
    wire N__77519;
    wire N__77516;
    wire N__77513;
    wire N__77510;
    wire N__77505;
    wire N__77502;
    wire N__77491;
    wire N__77488;
    wire N__77485;
    wire N__77482;
    wire N__77479;
    wire N__77476;
    wire N__77473;
    wire N__77470;
    wire N__77467;
    wire N__77464;
    wire N__77461;
    wire N__77458;
    wire N__77455;
    wire N__77452;
    wire N__77449;
    wire N__77446;
    wire N__77443;
    wire N__77440;
    wire N__77437;
    wire N__77434;
    wire N__77431;
    wire N__77430;
    wire N__77427;
    wire N__77424;
    wire N__77421;
    wire N__77420;
    wire N__77417;
    wire N__77414;
    wire N__77411;
    wire N__77408;
    wire N__77405;
    wire N__77398;
    wire N__77395;
    wire N__77392;
    wire N__77391;
    wire N__77388;
    wire N__77385;
    wire N__77382;
    wire N__77377;
    wire N__77376;
    wire N__77373;
    wire N__77370;
    wire N__77369;
    wire N__77366;
    wire N__77363;
    wire N__77360;
    wire N__77357;
    wire N__77354;
    wire N__77351;
    wire N__77350;
    wire N__77347;
    wire N__77344;
    wire N__77341;
    wire N__77338;
    wire N__77335;
    wire N__77332;
    wire N__77323;
    wire N__77320;
    wire N__77317;
    wire N__77314;
    wire N__77311;
    wire N__77308;
    wire N__77305;
    wire N__77304;
    wire N__77301;
    wire N__77300;
    wire N__77297;
    wire N__77294;
    wire N__77291;
    wire N__77284;
    wire N__77281;
    wire N__77280;
    wire N__77279;
    wire N__77278;
    wire N__77277;
    wire N__77274;
    wire N__77271;
    wire N__77268;
    wire N__77265;
    wire N__77262;
    wire N__77255;
    wire N__77248;
    wire N__77245;
    wire N__77242;
    wire N__77239;
    wire N__77236;
    wire N__77233;
    wire N__77230;
    wire N__77227;
    wire N__77224;
    wire N__77221;
    wire N__77218;
    wire N__77215;
    wire N__77212;
    wire N__77209;
    wire N__77206;
    wire N__77203;
    wire N__77200;
    wire N__77197;
    wire N__77194;
    wire N__77191;
    wire N__77188;
    wire N__77185;
    wire N__77182;
    wire N__77179;
    wire N__77176;
    wire N__77173;
    wire N__77170;
    wire N__77167;
    wire N__77164;
    wire N__77161;
    wire N__77158;
    wire N__77155;
    wire N__77152;
    wire N__77149;
    wire N__77146;
    wire N__77143;
    wire N__77140;
    wire N__77137;
    wire N__77134;
    wire N__77131;
    wire N__77128;
    wire N__77125;
    wire N__77122;
    wire N__77119;
    wire N__77116;
    wire N__77113;
    wire N__77110;
    wire N__77107;
    wire N__77104;
    wire N__77101;
    wire N__77098;
    wire N__77095;
    wire N__77092;
    wire N__77089;
    wire N__77086;
    wire N__77083;
    wire N__77082;
    wire N__77079;
    wire N__77076;
    wire N__77073;
    wire N__77070;
    wire N__77069;
    wire N__77064;
    wire N__77061;
    wire N__77058;
    wire N__77055;
    wire N__77052;
    wire N__77049;
    wire N__77048;
    wire N__77047;
    wire N__77046;
    wire N__77041;
    wire N__77034;
    wire N__77031;
    wire N__77028;
    wire N__77023;
    wire N__77020;
    wire N__77017;
    wire N__77014;
    wire N__77013;
    wire N__77010;
    wire N__77007;
    wire N__77006;
    wire N__77005;
    wire N__77004;
    wire N__77001;
    wire N__76998;
    wire N__76993;
    wire N__76990;
    wire N__76981;
    wire N__76978;
    wire N__76975;
    wire N__76972;
    wire N__76969;
    wire N__76966;
    wire N__76963;
    wire N__76960;
    wire N__76957;
    wire N__76954;
    wire N__76951;
    wire N__76948;
    wire N__76945;
    wire N__76942;
    wire N__76941;
    wire N__76940;
    wire N__76939;
    wire N__76930;
    wire N__76929;
    wire N__76928;
    wire N__76925;
    wire N__76922;
    wire N__76919;
    wire N__76912;
    wire N__76911;
    wire N__76908;
    wire N__76907;
    wire N__76906;
    wire N__76903;
    wire N__76900;
    wire N__76897;
    wire N__76894;
    wire N__76893;
    wire N__76890;
    wire N__76887;
    wire N__76884;
    wire N__76881;
    wire N__76878;
    wire N__76875;
    wire N__76864;
    wire N__76861;
    wire N__76858;
    wire N__76857;
    wire N__76856;
    wire N__76855;
    wire N__76854;
    wire N__76851;
    wire N__76848;
    wire N__76843;
    wire N__76842;
    wire N__76841;
    wire N__76838;
    wire N__76833;
    wire N__76832;
    wire N__76829;
    wire N__76824;
    wire N__76821;
    wire N__76818;
    wire N__76815;
    wire N__76810;
    wire N__76807;
    wire N__76798;
    wire N__76797;
    wire N__76796;
    wire N__76795;
    wire N__76792;
    wire N__76789;
    wire N__76784;
    wire N__76781;
    wire N__76774;
    wire N__76771;
    wire N__76768;
    wire N__76765;
    wire N__76762;
    wire N__76759;
    wire N__76756;
    wire N__76753;
    wire N__76750;
    wire N__76747;
    wire N__76744;
    wire N__76741;
    wire N__76738;
    wire N__76735;
    wire N__76732;
    wire N__76729;
    wire N__76726;
    wire N__76725;
    wire N__76722;
    wire N__76719;
    wire N__76716;
    wire N__76713;
    wire N__76708;
    wire N__76705;
    wire N__76702;
    wire N__76699;
    wire N__76696;
    wire N__76693;
    wire N__76690;
    wire N__76689;
    wire N__76686;
    wire N__76683;
    wire N__76678;
    wire N__76675;
    wire N__76672;
    wire N__76669;
    wire N__76666;
    wire N__76663;
    wire N__76660;
    wire N__76657;
    wire N__76654;
    wire N__76651;
    wire N__76648;
    wire N__76645;
    wire N__76642;
    wire N__76639;
    wire N__76636;
    wire N__76633;
    wire N__76630;
    wire N__76627;
    wire N__76624;
    wire N__76621;
    wire N__76618;
    wire N__76617;
    wire N__76614;
    wire N__76613;
    wire N__76612;
    wire N__76609;
    wire N__76608;
    wire N__76605;
    wire N__76602;
    wire N__76601;
    wire N__76598;
    wire N__76595;
    wire N__76594;
    wire N__76593;
    wire N__76592;
    wire N__76589;
    wire N__76584;
    wire N__76581;
    wire N__76578;
    wire N__76575;
    wire N__76568;
    wire N__76565;
    wire N__76560;
    wire N__76549;
    wire N__76548;
    wire N__76547;
    wire N__76546;
    wire N__76543;
    wire N__76538;
    wire N__76533;
    wire N__76532;
    wire N__76527;
    wire N__76526;
    wire N__76523;
    wire N__76520;
    wire N__76517;
    wire N__76510;
    wire N__76507;
    wire N__76504;
    wire N__76501;
    wire N__76498;
    wire N__76495;
    wire N__76492;
    wire N__76489;
    wire N__76486;
    wire N__76483;
    wire N__76482;
    wire N__76479;
    wire N__76476;
    wire N__76475;
    wire N__76474;
    wire N__76469;
    wire N__76466;
    wire N__76463;
    wire N__76458;
    wire N__76455;
    wire N__76450;
    wire N__76449;
    wire N__76446;
    wire N__76443;
    wire N__76442;
    wire N__76441;
    wire N__76438;
    wire N__76435;
    wire N__76432;
    wire N__76429;
    wire N__76426;
    wire N__76417;
    wire N__76414;
    wire N__76411;
    wire N__76408;
    wire N__76405;
    wire N__76402;
    wire N__76399;
    wire N__76396;
    wire N__76393;
    wire N__76390;
    wire N__76387;
    wire N__76384;
    wire N__76381;
    wire N__76378;
    wire N__76375;
    wire N__76372;
    wire N__76369;
    wire N__76366;
    wire N__76363;
    wire N__76360;
    wire N__76357;
    wire N__76354;
    wire N__76351;
    wire N__76348;
    wire N__76347;
    wire N__76346;
    wire N__76343;
    wire N__76340;
    wire N__76337;
    wire N__76334;
    wire N__76327;
    wire N__76324;
    wire N__76321;
    wire N__76320;
    wire N__76317;
    wire N__76314;
    wire N__76309;
    wire N__76306;
    wire N__76303;
    wire N__76300;
    wire N__76297;
    wire N__76294;
    wire N__76291;
    wire N__76288;
    wire N__76285;
    wire N__76282;
    wire N__76279;
    wire N__76276;
    wire N__76273;
    wire N__76270;
    wire N__76267;
    wire N__76264;
    wire N__76261;
    wire N__76258;
    wire N__76255;
    wire N__76254;
    wire N__76251;
    wire N__76248;
    wire N__76243;
    wire N__76240;
    wire N__76237;
    wire N__76234;
    wire N__76231;
    wire N__76228;
    wire N__76225;
    wire N__76224;
    wire N__76221;
    wire N__76218;
    wire N__76213;
    wire N__76210;
    wire N__76209;
    wire N__76206;
    wire N__76203;
    wire N__76202;
    wire N__76201;
    wire N__76196;
    wire N__76191;
    wire N__76190;
    wire N__76189;
    wire N__76184;
    wire N__76181;
    wire N__76178;
    wire N__76175;
    wire N__76168;
    wire N__76165;
    wire N__76162;
    wire N__76159;
    wire N__76156;
    wire N__76153;
    wire N__76150;
    wire N__76147;
    wire N__76144;
    wire N__76141;
    wire N__76138;
    wire N__76135;
    wire N__76132;
    wire N__76129;
    wire N__76126;
    wire N__76123;
    wire N__76120;
    wire N__76117;
    wire N__76114;
    wire N__76111;
    wire N__76108;
    wire N__76105;
    wire N__76102;
    wire N__76101;
    wire N__76098;
    wire N__76095;
    wire N__76092;
    wire N__76087;
    wire N__76084;
    wire N__76081;
    wire N__76078;
    wire N__76075;
    wire N__76072;
    wire N__76069;
    wire N__76066;
    wire N__76063;
    wire N__76060;
    wire N__76057;
    wire N__76054;
    wire N__76051;
    wire N__76050;
    wire N__76049;
    wire N__76048;
    wire N__76047;
    wire N__76044;
    wire N__76035;
    wire N__76032;
    wire N__76029;
    wire N__76024;
    wire N__76023;
    wire N__76022;
    wire N__76019;
    wire N__76016;
    wire N__76015;
    wire N__76014;
    wire N__76011;
    wire N__76010;
    wire N__76005;
    wire N__75996;
    wire N__75991;
    wire N__75990;
    wire N__75987;
    wire N__75984;
    wire N__75981;
    wire N__75976;
    wire N__75973;
    wire N__75970;
    wire N__75969;
    wire N__75966;
    wire N__75965;
    wire N__75962;
    wire N__75959;
    wire N__75956;
    wire N__75953;
    wire N__75952;
    wire N__75949;
    wire N__75946;
    wire N__75943;
    wire N__75940;
    wire N__75939;
    wire N__75938;
    wire N__75937;
    wire N__75936;
    wire N__75935;
    wire N__75932;
    wire N__75929;
    wire N__75924;
    wire N__75913;
    wire N__75904;
    wire N__75901;
    wire N__75900;
    wire N__75897;
    wire N__75894;
    wire N__75891;
    wire N__75886;
    wire N__75885;
    wire N__75882;
    wire N__75877;
    wire N__75876;
    wire N__75875;
    wire N__75872;
    wire N__75869;
    wire N__75866;
    wire N__75863;
    wire N__75860;
    wire N__75853;
    wire N__75850;
    wire N__75847;
    wire N__75844;
    wire N__75841;
    wire N__75838;
    wire N__75837;
    wire N__75834;
    wire N__75831;
    wire N__75830;
    wire N__75829;
    wire N__75824;
    wire N__75819;
    wire N__75816;
    wire N__75813;
    wire N__75810;
    wire N__75807;
    wire N__75802;
    wire N__75799;
    wire N__75796;
    wire N__75793;
    wire N__75790;
    wire N__75787;
    wire N__75784;
    wire N__75781;
    wire N__75778;
    wire N__75775;
    wire N__75772;
    wire N__75769;
    wire N__75766;
    wire N__75763;
    wire N__75760;
    wire N__75757;
    wire N__75754;
    wire N__75751;
    wire N__75748;
    wire N__75745;
    wire N__75742;
    wire N__75739;
    wire N__75736;
    wire N__75733;
    wire N__75730;
    wire N__75727;
    wire N__75724;
    wire N__75721;
    wire N__75718;
    wire N__75715;
    wire N__75712;
    wire N__75709;
    wire N__75706;
    wire N__75703;
    wire N__75700;
    wire N__75697;
    wire N__75694;
    wire N__75691;
    wire N__75688;
    wire N__75685;
    wire N__75682;
    wire N__75679;
    wire N__75676;
    wire N__75673;
    wire N__75670;
    wire N__75667;
    wire N__75664;
    wire N__75661;
    wire N__75658;
    wire N__75655;
    wire N__75652;
    wire N__75649;
    wire N__75646;
    wire N__75643;
    wire N__75640;
    wire N__75637;
    wire N__75634;
    wire N__75631;
    wire N__75628;
    wire N__75625;
    wire N__75622;
    wire N__75619;
    wire N__75616;
    wire N__75613;
    wire N__75610;
    wire N__75607;
    wire N__75604;
    wire N__75601;
    wire N__75598;
    wire N__75595;
    wire N__75592;
    wire N__75589;
    wire N__75586;
    wire N__75583;
    wire N__75580;
    wire N__75577;
    wire N__75574;
    wire N__75571;
    wire N__75568;
    wire N__75567;
    wire N__75564;
    wire N__75561;
    wire N__75558;
    wire N__75555;
    wire N__75550;
    wire N__75547;
    wire N__75544;
    wire N__75541;
    wire N__75538;
    wire N__75535;
    wire N__75532;
    wire N__75529;
    wire N__75526;
    wire N__75523;
    wire N__75520;
    wire N__75517;
    wire N__75514;
    wire N__75511;
    wire N__75508;
    wire N__75505;
    wire N__75502;
    wire N__75499;
    wire N__75496;
    wire N__75493;
    wire N__75490;
    wire N__75487;
    wire N__75484;
    wire N__75481;
    wire N__75478;
    wire N__75475;
    wire N__75472;
    wire N__75469;
    wire N__75466;
    wire N__75463;
    wire N__75460;
    wire N__75457;
    wire N__75454;
    wire N__75451;
    wire N__75448;
    wire N__75445;
    wire N__75442;
    wire N__75439;
    wire N__75436;
    wire N__75433;
    wire N__75430;
    wire N__75427;
    wire N__75424;
    wire N__75421;
    wire N__75418;
    wire N__75415;
    wire N__75412;
    wire N__75409;
    wire N__75406;
    wire N__75403;
    wire N__75400;
    wire N__75397;
    wire N__75394;
    wire N__75391;
    wire N__75388;
    wire N__75385;
    wire N__75382;
    wire N__75379;
    wire N__75376;
    wire N__75373;
    wire N__75370;
    wire N__75367;
    wire N__75364;
    wire N__75361;
    wire N__75358;
    wire N__75355;
    wire N__75352;
    wire N__75349;
    wire N__75346;
    wire N__75343;
    wire N__75340;
    wire N__75337;
    wire N__75334;
    wire N__75333;
    wire N__75332;
    wire N__75331;
    wire N__75330;
    wire N__75325;
    wire N__75318;
    wire N__75315;
    wire N__75312;
    wire N__75307;
    wire N__75304;
    wire N__75301;
    wire N__75298;
    wire N__75295;
    wire N__75292;
    wire N__75289;
    wire N__75286;
    wire N__75283;
    wire N__75280;
    wire N__75277;
    wire N__75274;
    wire N__75271;
    wire N__75268;
    wire N__75265;
    wire N__75262;
    wire N__75259;
    wire N__75256;
    wire N__75253;
    wire N__75250;
    wire N__75247;
    wire N__75244;
    wire N__75241;
    wire N__75238;
    wire N__75235;
    wire N__75232;
    wire N__75229;
    wire N__75226;
    wire N__75223;
    wire N__75220;
    wire N__75217;
    wire N__75214;
    wire N__75211;
    wire N__75208;
    wire N__75205;
    wire N__75202;
    wire N__75199;
    wire N__75196;
    wire N__75193;
    wire N__75190;
    wire N__75187;
    wire N__75184;
    wire N__75181;
    wire N__75178;
    wire N__75177;
    wire N__75176;
    wire N__75175;
    wire N__75172;
    wire N__75165;
    wire N__75160;
    wire N__75157;
    wire N__75154;
    wire N__75151;
    wire N__75148;
    wire N__75147;
    wire N__75146;
    wire N__75145;
    wire N__75138;
    wire N__75137;
    wire N__75136;
    wire N__75135;
    wire N__75132;
    wire N__75129;
    wire N__75124;
    wire N__75121;
    wire N__75118;
    wire N__75115;
    wire N__75112;
    wire N__75109;
    wire N__75106;
    wire N__75097;
    wire N__75094;
    wire N__75091;
    wire N__75090;
    wire N__75089;
    wire N__75082;
    wire N__75081;
    wire N__75080;
    wire N__75079;
    wire N__75078;
    wire N__75077;
    wire N__75074;
    wire N__75071;
    wire N__75066;
    wire N__75063;
    wire N__75060;
    wire N__75057;
    wire N__75054;
    wire N__75053;
    wire N__75050;
    wire N__75047;
    wire N__75044;
    wire N__75039;
    wire N__75036;
    wire N__75035;
    wire N__75032;
    wire N__75029;
    wire N__75026;
    wire N__75021;
    wire N__75018;
    wire N__75011;
    wire N__75008;
    wire N__75001;
    wire N__74998;
    wire N__74995;
    wire N__74992;
    wire N__74989;
    wire N__74986;
    wire N__74983;
    wire N__74980;
    wire N__74977;
    wire N__74974;
    wire N__74971;
    wire N__74968;
    wire N__74965;
    wire N__74962;
    wire N__74959;
    wire N__74956;
    wire N__74953;
    wire N__74950;
    wire N__74947;
    wire N__74944;
    wire N__74941;
    wire N__74938;
    wire N__74935;
    wire N__74932;
    wire N__74929;
    wire N__74926;
    wire N__74923;
    wire N__74920;
    wire N__74917;
    wire N__74914;
    wire N__74911;
    wire N__74908;
    wire N__74905;
    wire N__74902;
    wire N__74901;
    wire N__74898;
    wire N__74895;
    wire N__74894;
    wire N__74889;
    wire N__74886;
    wire N__74881;
    wire N__74878;
    wire N__74875;
    wire N__74874;
    wire N__74873;
    wire N__74870;
    wire N__74867;
    wire N__74864;
    wire N__74861;
    wire N__74854;
    wire N__74851;
    wire N__74848;
    wire N__74845;
    wire N__74842;
    wire N__74839;
    wire N__74836;
    wire N__74833;
    wire N__74830;
    wire N__74827;
    wire N__74824;
    wire N__74821;
    wire N__74818;
    wire N__74815;
    wire N__74812;
    wire N__74809;
    wire N__74806;
    wire N__74803;
    wire N__74800;
    wire N__74797;
    wire N__74794;
    wire N__74791;
    wire N__74788;
    wire N__74785;
    wire N__74782;
    wire N__74779;
    wire N__74776;
    wire N__74773;
    wire N__74770;
    wire N__74767;
    wire N__74764;
    wire N__74763;
    wire N__74760;
    wire N__74757;
    wire N__74756;
    wire N__74755;
    wire N__74754;
    wire N__74749;
    wire N__74742;
    wire N__74741;
    wire N__74740;
    wire N__74739;
    wire N__74736;
    wire N__74733;
    wire N__74730;
    wire N__74725;
    wire N__74716;
    wire N__74715;
    wire N__74714;
    wire N__74711;
    wire N__74710;
    wire N__74709;
    wire N__74706;
    wire N__74705;
    wire N__74704;
    wire N__74701;
    wire N__74700;
    wire N__74697;
    wire N__74692;
    wire N__74689;
    wire N__74684;
    wire N__74681;
    wire N__74678;
    wire N__74673;
    wire N__74670;
    wire N__74667;
    wire N__74664;
    wire N__74661;
    wire N__74656;
    wire N__74653;
    wire N__74648;
    wire N__74645;
    wire N__74638;
    wire N__74637;
    wire N__74636;
    wire N__74629;
    wire N__74628;
    wire N__74627;
    wire N__74626;
    wire N__74623;
    wire N__74620;
    wire N__74617;
    wire N__74614;
    wire N__74609;
    wire N__74602;
    wire N__74599;
    wire N__74596;
    wire N__74593;
    wire N__74590;
    wire N__74587;
    wire N__74584;
    wire N__74581;
    wire N__74578;
    wire N__74575;
    wire N__74572;
    wire N__74569;
    wire N__74566;
    wire N__74563;
    wire N__74560;
    wire N__74557;
    wire N__74554;
    wire N__74551;
    wire N__74548;
    wire N__74545;
    wire N__74542;
    wire N__74539;
    wire N__74536;
    wire N__74533;
    wire N__74530;
    wire N__74527;
    wire N__74524;
    wire N__74521;
    wire N__74518;
    wire N__74515;
    wire N__74512;
    wire N__74509;
    wire N__74506;
    wire N__74503;
    wire N__74500;
    wire N__74499;
    wire N__74498;
    wire N__74497;
    wire N__74496;
    wire N__74491;
    wire N__74484;
    wire N__74481;
    wire N__74480;
    wire N__74479;
    wire N__74476;
    wire N__74473;
    wire N__74470;
    wire N__74469;
    wire N__74466;
    wire N__74463;
    wire N__74460;
    wire N__74455;
    wire N__74452;
    wire N__74447;
    wire N__74444;
    wire N__74441;
    wire N__74434;
    wire N__74431;
    wire N__74428;
    wire N__74427;
    wire N__74426;
    wire N__74423;
    wire N__74420;
    wire N__74417;
    wire N__74412;
    wire N__74409;
    wire N__74408;
    wire N__74403;
    wire N__74400;
    wire N__74399;
    wire N__74396;
    wire N__74393;
    wire N__74390;
    wire N__74383;
    wire N__74382;
    wire N__74381;
    wire N__74378;
    wire N__74373;
    wire N__74370;
    wire N__74369;
    wire N__74366;
    wire N__74363;
    wire N__74360;
    wire N__74357;
    wire N__74350;
    wire N__74347;
    wire N__74344;
    wire N__74341;
    wire N__74338;
    wire N__74335;
    wire N__74332;
    wire N__74329;
    wire N__74326;
    wire N__74323;
    wire N__74320;
    wire N__74317;
    wire N__74314;
    wire N__74311;
    wire N__74308;
    wire N__74305;
    wire N__74302;
    wire N__74299;
    wire N__74296;
    wire N__74293;
    wire N__74290;
    wire N__74287;
    wire N__74284;
    wire N__74281;
    wire N__74278;
    wire N__74275;
    wire N__74272;
    wire N__74269;
    wire N__74266;
    wire N__74263;
    wire N__74260;
    wire N__74259;
    wire N__74258;
    wire N__74255;
    wire N__74252;
    wire N__74251;
    wire N__74248;
    wire N__74245;
    wire N__74242;
    wire N__74237;
    wire N__74234;
    wire N__74231;
    wire N__74228;
    wire N__74223;
    wire N__74218;
    wire N__74217;
    wire N__74216;
    wire N__74215;
    wire N__74212;
    wire N__74209;
    wire N__74204;
    wire N__74201;
    wire N__74194;
    wire N__74191;
    wire N__74188;
    wire N__74185;
    wire N__74182;
    wire N__74179;
    wire N__74176;
    wire N__74173;
    wire N__74170;
    wire N__74167;
    wire N__74164;
    wire N__74161;
    wire N__74158;
    wire N__74155;
    wire N__74152;
    wire N__74149;
    wire N__74146;
    wire N__74143;
    wire N__74140;
    wire N__74137;
    wire N__74134;
    wire N__74131;
    wire N__74128;
    wire N__74125;
    wire N__74124;
    wire N__74121;
    wire N__74118;
    wire N__74113;
    wire N__74110;
    wire N__74107;
    wire N__74104;
    wire N__74101;
    wire N__74098;
    wire N__74095;
    wire N__74092;
    wire N__74089;
    wire N__74086;
    wire N__74083;
    wire N__74080;
    wire N__74077;
    wire N__74074;
    wire N__74071;
    wire N__74068;
    wire N__74065;
    wire N__74062;
    wire N__74059;
    wire N__74056;
    wire N__74055;
    wire N__74052;
    wire N__74049;
    wire N__74044;
    wire N__74041;
    wire N__74038;
    wire N__74037;
    wire N__74034;
    wire N__74031;
    wire N__74026;
    wire N__74023;
    wire N__74020;
    wire N__74017;
    wire N__74014;
    wire N__74011;
    wire N__74008;
    wire N__74005;
    wire N__74002;
    wire N__73999;
    wire N__73996;
    wire N__73993;
    wire N__73990;
    wire N__73987;
    wire N__73984;
    wire N__73981;
    wire N__73978;
    wire N__73977;
    wire N__73974;
    wire N__73971;
    wire N__73966;
    wire N__73963;
    wire N__73960;
    wire N__73957;
    wire N__73954;
    wire N__73951;
    wire N__73948;
    wire N__73945;
    wire N__73942;
    wire N__73939;
    wire N__73936;
    wire N__73935;
    wire N__73934;
    wire N__73931;
    wire N__73928;
    wire N__73925;
    wire N__73920;
    wire N__73917;
    wire N__73914;
    wire N__73909;
    wire N__73906;
    wire N__73903;
    wire N__73902;
    wire N__73901;
    wire N__73900;
    wire N__73895;
    wire N__73892;
    wire N__73889;
    wire N__73886;
    wire N__73883;
    wire N__73880;
    wire N__73877;
    wire N__73874;
    wire N__73871;
    wire N__73864;
    wire N__73863;
    wire N__73858;
    wire N__73857;
    wire N__73854;
    wire N__73851;
    wire N__73846;
    wire N__73845;
    wire N__73842;
    wire N__73839;
    wire N__73834;
    wire N__73833;
    wire N__73832;
    wire N__73829;
    wire N__73828;
    wire N__73823;
    wire N__73822;
    wire N__73819;
    wire N__73816;
    wire N__73813;
    wire N__73810;
    wire N__73805;
    wire N__73800;
    wire N__73797;
    wire N__73792;
    wire N__73789;
    wire N__73786;
    wire N__73783;
    wire N__73780;
    wire N__73777;
    wire N__73774;
    wire N__73771;
    wire N__73768;
    wire N__73765;
    wire N__73762;
    wire N__73759;
    wire N__73756;
    wire N__73753;
    wire N__73750;
    wire N__73747;
    wire N__73744;
    wire N__73741;
    wire N__73738;
    wire N__73735;
    wire N__73732;
    wire N__73729;
    wire N__73726;
    wire N__73723;
    wire N__73720;
    wire N__73717;
    wire N__73714;
    wire N__73711;
    wire N__73708;
    wire N__73705;
    wire N__73702;
    wire N__73699;
    wire N__73698;
    wire N__73695;
    wire N__73692;
    wire N__73687;
    wire N__73684;
    wire N__73681;
    wire N__73678;
    wire N__73675;
    wire N__73672;
    wire N__73669;
    wire N__73666;
    wire N__73663;
    wire N__73660;
    wire N__73657;
    wire N__73654;
    wire N__73651;
    wire N__73648;
    wire N__73645;
    wire N__73642;
    wire N__73639;
    wire N__73636;
    wire N__73633;
    wire N__73630;
    wire N__73627;
    wire N__73624;
    wire N__73621;
    wire N__73618;
    wire N__73615;
    wire N__73612;
    wire N__73609;
    wire N__73606;
    wire N__73603;
    wire N__73600;
    wire N__73597;
    wire N__73594;
    wire N__73591;
    wire N__73588;
    wire N__73585;
    wire N__73582;
    wire N__73579;
    wire N__73576;
    wire N__73573;
    wire N__73570;
    wire N__73567;
    wire N__73564;
    wire N__73563;
    wire N__73560;
    wire N__73557;
    wire N__73554;
    wire N__73551;
    wire N__73546;
    wire N__73543;
    wire N__73540;
    wire N__73537;
    wire N__73534;
    wire N__73531;
    wire N__73528;
    wire N__73525;
    wire N__73522;
    wire N__73519;
    wire N__73516;
    wire N__73515;
    wire N__73512;
    wire N__73509;
    wire N__73504;
    wire N__73501;
    wire N__73498;
    wire N__73495;
    wire N__73492;
    wire N__73489;
    wire N__73486;
    wire N__73485;
    wire N__73482;
    wire N__73479;
    wire N__73474;
    wire N__73471;
    wire N__73468;
    wire N__73465;
    wire N__73462;
    wire N__73459;
    wire N__73456;
    wire N__73453;
    wire N__73450;
    wire N__73447;
    wire N__73444;
    wire N__73441;
    wire N__73438;
    wire N__73435;
    wire N__73434;
    wire N__73433;
    wire N__73430;
    wire N__73425;
    wire N__73420;
    wire N__73417;
    wire N__73416;
    wire N__73413;
    wire N__73410;
    wire N__73405;
    wire N__73402;
    wire N__73399;
    wire N__73396;
    wire N__73393;
    wire N__73390;
    wire N__73387;
    wire N__73384;
    wire N__73381;
    wire N__73380;
    wire N__73379;
    wire N__73376;
    wire N__73373;
    wire N__73370;
    wire N__73367;
    wire N__73362;
    wire N__73359;
    wire N__73356;
    wire N__73351;
    wire N__73348;
    wire N__73345;
    wire N__73342;
    wire N__73339;
    wire N__73336;
    wire N__73333;
    wire N__73330;
    wire N__73327;
    wire N__73324;
    wire N__73321;
    wire N__73318;
    wire N__73315;
    wire N__73312;
    wire N__73309;
    wire N__73306;
    wire N__73303;
    wire N__73300;
    wire N__73297;
    wire N__73294;
    wire N__73291;
    wire N__73290;
    wire N__73287;
    wire N__73284;
    wire N__73279;
    wire N__73278;
    wire N__73275;
    wire N__73272;
    wire N__73271;
    wire N__73268;
    wire N__73265;
    wire N__73262;
    wire N__73261;
    wire N__73256;
    wire N__73253;
    wire N__73250;
    wire N__73247;
    wire N__73240;
    wire N__73239;
    wire N__73238;
    wire N__73233;
    wire N__73232;
    wire N__73231;
    wire N__73230;
    wire N__73227;
    wire N__73224;
    wire N__73217;
    wire N__73214;
    wire N__73211;
    wire N__73206;
    wire N__73201;
    wire N__73198;
    wire N__73195;
    wire N__73192;
    wire N__73189;
    wire N__73186;
    wire N__73183;
    wire N__73180;
    wire N__73177;
    wire N__73174;
    wire N__73171;
    wire N__73168;
    wire N__73165;
    wire N__73162;
    wire N__73159;
    wire N__73156;
    wire N__73153;
    wire N__73150;
    wire N__73147;
    wire N__73144;
    wire N__73141;
    wire N__73138;
    wire N__73135;
    wire N__73132;
    wire N__73129;
    wire N__73126;
    wire N__73123;
    wire N__73120;
    wire N__73117;
    wire N__73114;
    wire N__73111;
    wire N__73108;
    wire N__73105;
    wire N__73102;
    wire N__73101;
    wire N__73098;
    wire N__73095;
    wire N__73090;
    wire N__73089;
    wire N__73086;
    wire N__73083;
    wire N__73078;
    wire N__73075;
    wire N__73072;
    wire N__73069;
    wire N__73068;
    wire N__73065;
    wire N__73062;
    wire N__73059;
    wire N__73056;
    wire N__73053;
    wire N__73050;
    wire N__73045;
    wire N__73042;
    wire N__73041;
    wire N__73038;
    wire N__73035;
    wire N__73030;
    wire N__73027;
    wire N__73024;
    wire N__73021;
    wire N__73018;
    wire N__73015;
    wire N__73012;
    wire N__73009;
    wire N__73008;
    wire N__73005;
    wire N__73002;
    wire N__72999;
    wire N__72996;
    wire N__72993;
    wire N__72990;
    wire N__72985;
    wire N__72982;
    wire N__72981;
    wire N__72978;
    wire N__72975;
    wire N__72970;
    wire N__72967;
    wire N__72964;
    wire N__72961;
    wire N__72958;
    wire N__72955;
    wire N__72952;
    wire N__72949;
    wire N__72946;
    wire N__72943;
    wire N__72940;
    wire N__72937;
    wire N__72934;
    wire N__72931;
    wire N__72928;
    wire N__72925;
    wire N__72922;
    wire N__72919;
    wire N__72916;
    wire N__72913;
    wire N__72910;
    wire N__72907;
    wire N__72904;
    wire N__72901;
    wire N__72898;
    wire N__72895;
    wire N__72892;
    wire N__72889;
    wire N__72886;
    wire N__72883;
    wire N__72882;
    wire N__72881;
    wire N__72878;
    wire N__72877;
    wire N__72874;
    wire N__72873;
    wire N__72868;
    wire N__72865;
    wire N__72862;
    wire N__72859;
    wire N__72856;
    wire N__72853;
    wire N__72846;
    wire N__72841;
    wire N__72838;
    wire N__72835;
    wire N__72832;
    wire N__72829;
    wire N__72826;
    wire N__72823;
    wire N__72820;
    wire N__72819;
    wire N__72816;
    wire N__72813;
    wire N__72810;
    wire N__72807;
    wire N__72804;
    wire N__72801;
    wire N__72796;
    wire N__72793;
    wire N__72790;
    wire N__72789;
    wire N__72788;
    wire N__72787;
    wire N__72784;
    wire N__72777;
    wire N__72776;
    wire N__72773;
    wire N__72770;
    wire N__72767;
    wire N__72766;
    wire N__72765;
    wire N__72764;
    wire N__72763;
    wire N__72758;
    wire N__72755;
    wire N__72750;
    wire N__72745;
    wire N__72736;
    wire N__72733;
    wire N__72730;
    wire N__72727;
    wire N__72724;
    wire N__72723;
    wire N__72718;
    wire N__72717;
    wire N__72714;
    wire N__72713;
    wire N__72712;
    wire N__72709;
    wire N__72706;
    wire N__72703;
    wire N__72700;
    wire N__72697;
    wire N__72688;
    wire N__72685;
    wire N__72682;
    wire N__72679;
    wire N__72676;
    wire N__72673;
    wire N__72670;
    wire N__72667;
    wire N__72664;
    wire N__72661;
    wire N__72658;
    wire N__72655;
    wire N__72654;
    wire N__72651;
    wire N__72650;
    wire N__72647;
    wire N__72646;
    wire N__72643;
    wire N__72640;
    wire N__72637;
    wire N__72634;
    wire N__72631;
    wire N__72628;
    wire N__72623;
    wire N__72620;
    wire N__72617;
    wire N__72614;
    wire N__72607;
    wire N__72604;
    wire N__72601;
    wire N__72598;
    wire N__72595;
    wire N__72592;
    wire N__72589;
    wire N__72586;
    wire N__72583;
    wire N__72580;
    wire N__72577;
    wire N__72574;
    wire N__72571;
    wire N__72568;
    wire N__72565;
    wire N__72562;
    wire N__72559;
    wire N__72556;
    wire N__72553;
    wire N__72550;
    wire N__72549;
    wire N__72546;
    wire N__72543;
    wire N__72538;
    wire N__72535;
    wire N__72532;
    wire N__72529;
    wire N__72526;
    wire N__72523;
    wire N__72520;
    wire N__72517;
    wire N__72514;
    wire N__72511;
    wire N__72508;
    wire N__72505;
    wire N__72504;
    wire N__72501;
    wire N__72498;
    wire N__72497;
    wire N__72494;
    wire N__72491;
    wire N__72488;
    wire N__72483;
    wire N__72480;
    wire N__72475;
    wire N__72472;
    wire N__72469;
    wire N__72466;
    wire N__72463;
    wire N__72460;
    wire N__72457;
    wire N__72454;
    wire N__72451;
    wire N__72448;
    wire N__72445;
    wire N__72442;
    wire N__72439;
    wire N__72436;
    wire N__72433;
    wire N__72430;
    wire N__72427;
    wire N__72424;
    wire N__72421;
    wire N__72418;
    wire N__72415;
    wire N__72412;
    wire N__72409;
    wire N__72406;
    wire N__72405;
    wire N__72402;
    wire N__72399;
    wire N__72396;
    wire N__72393;
    wire N__72388;
    wire N__72385;
    wire N__72384;
    wire N__72383;
    wire N__72380;
    wire N__72377;
    wire N__72376;
    wire N__72373;
    wire N__72370;
    wire N__72367;
    wire N__72362;
    wire N__72359;
    wire N__72352;
    wire N__72349;
    wire N__72346;
    wire N__72343;
    wire N__72340;
    wire N__72337;
    wire N__72334;
    wire N__72331;
    wire N__72328;
    wire N__72325;
    wire N__72322;
    wire N__72319;
    wire N__72316;
    wire N__72313;
    wire N__72310;
    wire N__72307;
    wire N__72304;
    wire N__72301;
    wire N__72298;
    wire N__72295;
    wire N__72292;
    wire N__72289;
    wire N__72286;
    wire N__72283;
    wire N__72280;
    wire N__72277;
    wire N__72274;
    wire N__72271;
    wire N__72268;
    wire N__72265;
    wire N__72262;
    wire N__72261;
    wire N__72258;
    wire N__72255;
    wire N__72254;
    wire N__72249;
    wire N__72246;
    wire N__72241;
    wire N__72238;
    wire N__72235;
    wire N__72234;
    wire N__72231;
    wire N__72228;
    wire N__72225;
    wire N__72222;
    wire N__72217;
    wire N__72216;
    wire N__72213;
    wire N__72210;
    wire N__72205;
    wire N__72204;
    wire N__72201;
    wire N__72200;
    wire N__72197;
    wire N__72194;
    wire N__72191;
    wire N__72188;
    wire N__72185;
    wire N__72182;
    wire N__72179;
    wire N__72172;
    wire N__72169;
    wire N__72166;
    wire N__72163;
    wire N__72160;
    wire N__72157;
    wire N__72154;
    wire N__72151;
    wire N__72148;
    wire N__72145;
    wire N__72142;
    wire N__72139;
    wire N__72136;
    wire N__72133;
    wire N__72130;
    wire N__72127;
    wire N__72124;
    wire N__72121;
    wire N__72118;
    wire N__72115;
    wire N__72112;
    wire N__72111;
    wire N__72110;
    wire N__72107;
    wire N__72104;
    wire N__72101;
    wire N__72098;
    wire N__72097;
    wire N__72096;
    wire N__72093;
    wire N__72090;
    wire N__72087;
    wire N__72084;
    wire N__72081;
    wire N__72078;
    wire N__72075;
    wire N__72072;
    wire N__72069;
    wire N__72066;
    wire N__72063;
    wire N__72060;
    wire N__72055;
    wire N__72052;
    wire N__72049;
    wire N__72044;
    wire N__72041;
    wire N__72034;
    wire N__72033;
    wire N__72030;
    wire N__72029;
    wire N__72028;
    wire N__72025;
    wire N__72022;
    wire N__72019;
    wire N__72016;
    wire N__72013;
    wire N__72010;
    wire N__72007;
    wire N__72004;
    wire N__72001;
    wire N__71998;
    wire N__71995;
    wire N__71990;
    wire N__71983;
    wire N__71980;
    wire N__71977;
    wire N__71976;
    wire N__71973;
    wire N__71970;
    wire N__71967;
    wire N__71964;
    wire N__71961;
    wire N__71956;
    wire N__71955;
    wire N__71952;
    wire N__71949;
    wire N__71946;
    wire N__71943;
    wire N__71938;
    wire N__71935;
    wire N__71932;
    wire N__71929;
    wire N__71926;
    wire N__71923;
    wire N__71920;
    wire N__71917;
    wire N__71914;
    wire N__71911;
    wire N__71908;
    wire N__71905;
    wire N__71902;
    wire N__71899;
    wire N__71896;
    wire N__71893;
    wire N__71890;
    wire N__71887;
    wire N__71884;
    wire N__71881;
    wire N__71878;
    wire N__71875;
    wire N__71872;
    wire N__71869;
    wire N__71866;
    wire N__71865;
    wire N__71864;
    wire N__71861;
    wire N__71858;
    wire N__71855;
    wire N__71852;
    wire N__71849;
    wire N__71846;
    wire N__71839;
    wire N__71836;
    wire N__71833;
    wire N__71830;
    wire N__71827;
    wire N__71824;
    wire N__71821;
    wire N__71818;
    wire N__71815;
    wire N__71812;
    wire N__71809;
    wire N__71806;
    wire N__71803;
    wire N__71800;
    wire N__71797;
    wire N__71794;
    wire N__71791;
    wire N__71788;
    wire N__71785;
    wire N__71782;
    wire N__71779;
    wire N__71776;
    wire N__71773;
    wire N__71770;
    wire N__71767;
    wire N__71764;
    wire N__71761;
    wire N__71758;
    wire N__71755;
    wire N__71752;
    wire N__71749;
    wire N__71746;
    wire N__71743;
    wire N__71740;
    wire N__71737;
    wire N__71734;
    wire N__71731;
    wire N__71728;
    wire N__71725;
    wire N__71722;
    wire N__71719;
    wire N__71716;
    wire N__71713;
    wire N__71710;
    wire N__71707;
    wire N__71704;
    wire N__71701;
    wire N__71698;
    wire N__71695;
    wire N__71692;
    wire N__71689;
    wire N__71686;
    wire N__71683;
    wire N__71680;
    wire N__71677;
    wire N__71674;
    wire N__71671;
    wire N__71668;
    wire N__71665;
    wire N__71662;
    wire N__71659;
    wire N__71656;
    wire N__71653;
    wire N__71650;
    wire N__71649;
    wire N__71646;
    wire N__71643;
    wire N__71638;
    wire N__71635;
    wire N__71634;
    wire N__71631;
    wire N__71628;
    wire N__71623;
    wire N__71620;
    wire N__71617;
    wire N__71614;
    wire N__71611;
    wire N__71608;
    wire N__71605;
    wire N__71602;
    wire N__71599;
    wire N__71596;
    wire N__71593;
    wire N__71590;
    wire N__71587;
    wire N__71584;
    wire N__71581;
    wire N__71578;
    wire N__71575;
    wire N__71572;
    wire N__71569;
    wire N__71566;
    wire N__71563;
    wire N__71560;
    wire N__71557;
    wire N__71554;
    wire N__71551;
    wire N__71548;
    wire N__71545;
    wire N__71544;
    wire N__71543;
    wire N__71542;
    wire N__71541;
    wire N__71536;
    wire N__71533;
    wire N__71528;
    wire N__71527;
    wire N__71526;
    wire N__71523;
    wire N__71518;
    wire N__71513;
    wire N__71510;
    wire N__71503;
    wire N__71502;
    wire N__71501;
    wire N__71500;
    wire N__71499;
    wire N__71496;
    wire N__71493;
    wire N__71492;
    wire N__71489;
    wire N__71486;
    wire N__71483;
    wire N__71480;
    wire N__71475;
    wire N__71470;
    wire N__71467;
    wire N__71464;
    wire N__71463;
    wire N__71460;
    wire N__71455;
    wire N__71452;
    wire N__71449;
    wire N__71446;
    wire N__71443;
    wire N__71440;
    wire N__71431;
    wire N__71430;
    wire N__71427;
    wire N__71426;
    wire N__71423;
    wire N__71422;
    wire N__71421;
    wire N__71418;
    wire N__71415;
    wire N__71410;
    wire N__71407;
    wire N__71400;
    wire N__71395;
    wire N__71392;
    wire N__71389;
    wire N__71386;
    wire N__71383;
    wire N__71380;
    wire N__71377;
    wire N__71374;
    wire N__71371;
    wire N__71368;
    wire N__71365;
    wire N__71362;
    wire N__71359;
    wire N__71356;
    wire N__71353;
    wire N__71350;
    wire N__71347;
    wire N__71344;
    wire N__71341;
    wire N__71338;
    wire N__71335;
    wire N__71332;
    wire N__71329;
    wire N__71326;
    wire N__71323;
    wire N__71320;
    wire N__71317;
    wire N__71314;
    wire N__71311;
    wire N__71308;
    wire N__71305;
    wire N__71302;
    wire N__71299;
    wire N__71296;
    wire N__71293;
    wire N__71290;
    wire N__71287;
    wire N__71284;
    wire N__71281;
    wire N__71278;
    wire N__71275;
    wire N__71272;
    wire N__71269;
    wire N__71266;
    wire N__71263;
    wire N__71260;
    wire N__71257;
    wire N__71254;
    wire N__71251;
    wire N__71248;
    wire N__71245;
    wire N__71242;
    wire N__71239;
    wire N__71236;
    wire N__71233;
    wire N__71230;
    wire N__71227;
    wire N__71224;
    wire N__71221;
    wire N__71218;
    wire N__71215;
    wire N__71212;
    wire N__71211;
    wire N__71208;
    wire N__71205;
    wire N__71200;
    wire N__71197;
    wire N__71194;
    wire N__71191;
    wire N__71188;
    wire N__71185;
    wire N__71182;
    wire N__71179;
    wire N__71176;
    wire N__71173;
    wire N__71170;
    wire N__71167;
    wire N__71164;
    wire N__71161;
    wire N__71158;
    wire N__71155;
    wire N__71152;
    wire N__71149;
    wire N__71146;
    wire N__71143;
    wire N__71140;
    wire N__71137;
    wire N__71134;
    wire N__71131;
    wire N__71128;
    wire N__71125;
    wire N__71122;
    wire N__71119;
    wire N__71116;
    wire N__71113;
    wire N__71110;
    wire N__71107;
    wire N__71104;
    wire N__71101;
    wire N__71098;
    wire N__71095;
    wire N__71092;
    wire N__71089;
    wire N__71086;
    wire N__71083;
    wire N__71080;
    wire N__71077;
    wire N__71074;
    wire N__71071;
    wire N__71068;
    wire N__71065;
    wire N__71062;
    wire N__71059;
    wire N__71056;
    wire N__71053;
    wire N__71050;
    wire N__71047;
    wire N__71044;
    wire N__71041;
    wire N__71038;
    wire N__71035;
    wire N__71032;
    wire N__71029;
    wire N__71026;
    wire N__71023;
    wire N__71020;
    wire N__71017;
    wire N__71014;
    wire N__71011;
    wire N__71008;
    wire N__71005;
    wire N__71002;
    wire N__70999;
    wire N__70996;
    wire N__70993;
    wire N__70990;
    wire N__70987;
    wire N__70984;
    wire N__70981;
    wire N__70978;
    wire N__70975;
    wire N__70972;
    wire N__70969;
    wire N__70966;
    wire N__70963;
    wire N__70960;
    wire N__70957;
    wire N__70954;
    wire N__70951;
    wire N__70948;
    wire N__70945;
    wire N__70944;
    wire N__70941;
    wire N__70938;
    wire N__70933;
    wire N__70930;
    wire N__70927;
    wire N__70924;
    wire N__70921;
    wire N__70918;
    wire N__70915;
    wire N__70912;
    wire N__70909;
    wire N__70906;
    wire N__70903;
    wire N__70900;
    wire N__70897;
    wire N__70894;
    wire N__70891;
    wire N__70888;
    wire N__70885;
    wire N__70882;
    wire N__70879;
    wire N__70876;
    wire N__70873;
    wire N__70872;
    wire N__70869;
    wire N__70866;
    wire N__70863;
    wire N__70860;
    wire N__70855;
    wire N__70852;
    wire N__70849;
    wire N__70848;
    wire N__70847;
    wire N__70844;
    wire N__70843;
    wire N__70838;
    wire N__70835;
    wire N__70832;
    wire N__70829;
    wire N__70826;
    wire N__70819;
    wire N__70816;
    wire N__70813;
    wire N__70810;
    wire N__70807;
    wire N__70804;
    wire N__70801;
    wire N__70798;
    wire N__70795;
    wire N__70792;
    wire N__70789;
    wire N__70786;
    wire N__70783;
    wire N__70780;
    wire N__70777;
    wire N__70774;
    wire N__70771;
    wire N__70768;
    wire N__70765;
    wire N__70762;
    wire N__70759;
    wire N__70758;
    wire N__70757;
    wire N__70754;
    wire N__70751;
    wire N__70748;
    wire N__70743;
    wire N__70740;
    wire N__70737;
    wire N__70734;
    wire N__70729;
    wire N__70726;
    wire N__70723;
    wire N__70720;
    wire N__70719;
    wire N__70718;
    wire N__70717;
    wire N__70716;
    wire N__70713;
    wire N__70710;
    wire N__70707;
    wire N__70702;
    wire N__70697;
    wire N__70694;
    wire N__70693;
    wire N__70692;
    wire N__70691;
    wire N__70690;
    wire N__70683;
    wire N__70674;
    wire N__70669;
    wire N__70666;
    wire N__70663;
    wire N__70660;
    wire N__70657;
    wire N__70654;
    wire N__70651;
    wire N__70648;
    wire N__70645;
    wire N__70642;
    wire N__70639;
    wire N__70636;
    wire N__70633;
    wire N__70630;
    wire N__70629;
    wire N__70626;
    wire N__70623;
    wire N__70620;
    wire N__70615;
    wire N__70612;
    wire N__70609;
    wire N__70606;
    wire N__70603;
    wire N__70600;
    wire N__70597;
    wire N__70594;
    wire N__70591;
    wire N__70588;
    wire N__70585;
    wire N__70582;
    wire N__70579;
    wire N__70576;
    wire N__70575;
    wire N__70572;
    wire N__70571;
    wire N__70568;
    wire N__70565;
    wire N__70562;
    wire N__70559;
    wire N__70554;
    wire N__70549;
    wire N__70546;
    wire N__70543;
    wire N__70540;
    wire N__70537;
    wire N__70534;
    wire N__70531;
    wire N__70528;
    wire N__70525;
    wire N__70522;
    wire N__70519;
    wire N__70516;
    wire N__70513;
    wire N__70510;
    wire N__70507;
    wire N__70504;
    wire N__70501;
    wire N__70498;
    wire N__70495;
    wire N__70492;
    wire N__70489;
    wire N__70486;
    wire N__70483;
    wire N__70480;
    wire N__70477;
    wire N__70474;
    wire N__70471;
    wire N__70468;
    wire N__70465;
    wire N__70462;
    wire N__70459;
    wire N__70456;
    wire N__70453;
    wire N__70452;
    wire N__70449;
    wire N__70446;
    wire N__70443;
    wire N__70440;
    wire N__70437;
    wire N__70434;
    wire N__70429;
    wire N__70426;
    wire N__70423;
    wire N__70420;
    wire N__70417;
    wire N__70416;
    wire N__70415;
    wire N__70412;
    wire N__70407;
    wire N__70404;
    wire N__70399;
    wire N__70396;
    wire N__70393;
    wire N__70390;
    wire N__70387;
    wire N__70384;
    wire N__70381;
    wire N__70378;
    wire N__70375;
    wire N__70372;
    wire N__70369;
    wire N__70366;
    wire N__70363;
    wire N__70360;
    wire N__70357;
    wire N__70354;
    wire N__70351;
    wire N__70348;
    wire N__70345;
    wire N__70342;
    wire N__70339;
    wire N__70336;
    wire N__70333;
    wire N__70330;
    wire N__70327;
    wire N__70324;
    wire N__70321;
    wire N__70318;
    wire N__70315;
    wire N__70312;
    wire N__70309;
    wire N__70306;
    wire N__70303;
    wire N__70300;
    wire N__70297;
    wire N__70294;
    wire N__70291;
    wire N__70288;
    wire N__70285;
    wire N__70282;
    wire N__70279;
    wire N__70276;
    wire N__70273;
    wire N__70270;
    wire N__70267;
    wire N__70264;
    wire N__70261;
    wire N__70258;
    wire N__70255;
    wire N__70252;
    wire N__70249;
    wire N__70246;
    wire N__70243;
    wire N__70240;
    wire N__70237;
    wire N__70234;
    wire N__70231;
    wire N__70228;
    wire N__70225;
    wire N__70222;
    wire N__70219;
    wire N__70216;
    wire N__70213;
    wire N__70210;
    wire N__70207;
    wire N__70204;
    wire N__70201;
    wire N__70198;
    wire N__70195;
    wire N__70192;
    wire N__70189;
    wire N__70186;
    wire N__70183;
    wire N__70180;
    wire N__70177;
    wire N__70174;
    wire N__70171;
    wire N__70168;
    wire N__70165;
    wire N__70162;
    wire N__70159;
    wire N__70156;
    wire N__70153;
    wire N__70150;
    wire N__70149;
    wire N__70146;
    wire N__70143;
    wire N__70140;
    wire N__70137;
    wire N__70134;
    wire N__70131;
    wire N__70126;
    wire N__70123;
    wire N__70120;
    wire N__70117;
    wire N__70114;
    wire N__70111;
    wire N__70108;
    wire N__70107;
    wire N__70104;
    wire N__70101;
    wire N__70096;
    wire N__70093;
    wire N__70090;
    wire N__70087;
    wire N__70084;
    wire N__70081;
    wire N__70078;
    wire N__70075;
    wire N__70072;
    wire N__70069;
    wire N__70066;
    wire N__70065;
    wire N__70064;
    wire N__70061;
    wire N__70056;
    wire N__70051;
    wire N__70048;
    wire N__70045;
    wire N__70044;
    wire N__70041;
    wire N__70038;
    wire N__70035;
    wire N__70032;
    wire N__70029;
    wire N__70026;
    wire N__70021;
    wire N__70018;
    wire N__70015;
    wire N__70012;
    wire N__70009;
    wire N__70006;
    wire N__70003;
    wire N__70000;
    wire N__69997;
    wire N__69994;
    wire N__69991;
    wire N__69988;
    wire N__69985;
    wire N__69982;
    wire N__69979;
    wire N__69976;
    wire N__69973;
    wire N__69970;
    wire N__69967;
    wire N__69964;
    wire N__69961;
    wire N__69958;
    wire N__69955;
    wire N__69952;
    wire N__69949;
    wire N__69946;
    wire N__69943;
    wire N__69940;
    wire N__69937;
    wire N__69934;
    wire N__69931;
    wire N__69928;
    wire N__69925;
    wire N__69922;
    wire N__69919;
    wire N__69916;
    wire N__69913;
    wire N__69910;
    wire N__69907;
    wire N__69904;
    wire N__69901;
    wire N__69898;
    wire N__69895;
    wire N__69892;
    wire N__69889;
    wire N__69888;
    wire N__69885;
    wire N__69882;
    wire N__69879;
    wire N__69876;
    wire N__69873;
    wire N__69870;
    wire N__69865;
    wire N__69862;
    wire N__69861;
    wire N__69860;
    wire N__69857;
    wire N__69852;
    wire N__69849;
    wire N__69846;
    wire N__69843;
    wire N__69842;
    wire N__69839;
    wire N__69836;
    wire N__69833;
    wire N__69826;
    wire N__69823;
    wire N__69820;
    wire N__69817;
    wire N__69814;
    wire N__69811;
    wire N__69808;
    wire N__69805;
    wire N__69802;
    wire N__69799;
    wire N__69796;
    wire N__69793;
    wire N__69790;
    wire N__69787;
    wire N__69784;
    wire N__69781;
    wire N__69780;
    wire N__69777;
    wire N__69774;
    wire N__69773;
    wire N__69768;
    wire N__69765;
    wire N__69762;
    wire N__69759;
    wire N__69754;
    wire N__69751;
    wire N__69748;
    wire N__69745;
    wire N__69742;
    wire N__69739;
    wire N__69736;
    wire N__69733;
    wire N__69730;
    wire N__69727;
    wire N__69724;
    wire N__69721;
    wire N__69718;
    wire N__69715;
    wire N__69712;
    wire N__69709;
    wire N__69706;
    wire N__69703;
    wire N__69700;
    wire N__69697;
    wire N__69694;
    wire N__69691;
    wire N__69688;
    wire N__69685;
    wire N__69682;
    wire N__69679;
    wire N__69676;
    wire N__69673;
    wire N__69672;
    wire N__69671;
    wire N__69664;
    wire N__69661;
    wire N__69658;
    wire N__69655;
    wire N__69652;
    wire N__69649;
    wire N__69646;
    wire N__69643;
    wire N__69640;
    wire N__69637;
    wire N__69634;
    wire N__69631;
    wire N__69628;
    wire N__69625;
    wire N__69622;
    wire N__69619;
    wire N__69616;
    wire N__69613;
    wire N__69610;
    wire N__69607;
    wire N__69604;
    wire N__69601;
    wire N__69598;
    wire N__69595;
    wire N__69592;
    wire N__69589;
    wire N__69586;
    wire N__69583;
    wire N__69580;
    wire N__69577;
    wire N__69574;
    wire N__69571;
    wire N__69568;
    wire N__69565;
    wire N__69562;
    wire N__69559;
    wire N__69556;
    wire N__69553;
    wire N__69552;
    wire N__69549;
    wire N__69548;
    wire N__69545;
    wire N__69542;
    wire N__69539;
    wire N__69536;
    wire N__69533;
    wire N__69530;
    wire N__69527;
    wire N__69520;
    wire N__69519;
    wire N__69516;
    wire N__69513;
    wire N__69510;
    wire N__69505;
    wire N__69502;
    wire N__69499;
    wire N__69496;
    wire N__69495;
    wire N__69490;
    wire N__69487;
    wire N__69484;
    wire N__69481;
    wire N__69478;
    wire N__69475;
    wire N__69472;
    wire N__69469;
    wire N__69466;
    wire N__69463;
    wire N__69460;
    wire N__69457;
    wire N__69454;
    wire N__69451;
    wire N__69450;
    wire N__69449;
    wire N__69448;
    wire N__69447;
    wire N__69446;
    wire N__69441;
    wire N__69438;
    wire N__69435;
    wire N__69430;
    wire N__69425;
    wire N__69418;
    wire N__69417;
    wire N__69414;
    wire N__69411;
    wire N__69408;
    wire N__69403;
    wire N__69400;
    wire N__69397;
    wire N__69394;
    wire N__69391;
    wire N__69388;
    wire N__69385;
    wire N__69382;
    wire N__69381;
    wire N__69378;
    wire N__69375;
    wire N__69370;
    wire N__69369;
    wire N__69366;
    wire N__69363;
    wire N__69358;
    wire N__69355;
    wire N__69352;
    wire N__69349;
    wire N__69346;
    wire N__69343;
    wire N__69340;
    wire N__69337;
    wire N__69334;
    wire N__69331;
    wire N__69328;
    wire N__69325;
    wire N__69322;
    wire N__69319;
    wire N__69316;
    wire N__69313;
    wire N__69310;
    wire N__69307;
    wire N__69304;
    wire N__69301;
    wire N__69298;
    wire N__69295;
    wire N__69294;
    wire N__69291;
    wire N__69288;
    wire N__69285;
    wire N__69282;
    wire N__69277;
    wire N__69276;
    wire N__69273;
    wire N__69272;
    wire N__69269;
    wire N__69266;
    wire N__69263;
    wire N__69260;
    wire N__69257;
    wire N__69254;
    wire N__69251;
    wire N__69248;
    wire N__69243;
    wire N__69238;
    wire N__69235;
    wire N__69232;
    wire N__69231;
    wire N__69228;
    wire N__69227;
    wire N__69224;
    wire N__69221;
    wire N__69218;
    wire N__69215;
    wire N__69212;
    wire N__69209;
    wire N__69206;
    wire N__69201;
    wire N__69196;
    wire N__69193;
    wire N__69192;
    wire N__69189;
    wire N__69188;
    wire N__69185;
    wire N__69182;
    wire N__69179;
    wire N__69178;
    wire N__69175;
    wire N__69172;
    wire N__69169;
    wire N__69166;
    wire N__69163;
    wire N__69160;
    wire N__69157;
    wire N__69154;
    wire N__69151;
    wire N__69148;
    wire N__69143;
    wire N__69140;
    wire N__69133;
    wire N__69130;
    wire N__69127;
    wire N__69124;
    wire N__69121;
    wire N__69120;
    wire N__69119;
    wire N__69116;
    wire N__69111;
    wire N__69110;
    wire N__69109;
    wire N__69106;
    wire N__69103;
    wire N__69102;
    wire N__69099;
    wire N__69096;
    wire N__69095;
    wire N__69092;
    wire N__69089;
    wire N__69080;
    wire N__69073;
    wire N__69072;
    wire N__69069;
    wire N__69066;
    wire N__69061;
    wire N__69058;
    wire N__69055;
    wire N__69052;
    wire N__69049;
    wire N__69046;
    wire N__69043;
    wire N__69040;
    wire N__69037;
    wire N__69034;
    wire N__69031;
    wire N__69028;
    wire N__69025;
    wire N__69022;
    wire N__69019;
    wire N__69016;
    wire N__69013;
    wire N__69010;
    wire N__69007;
    wire N__69004;
    wire N__69001;
    wire N__68998;
    wire N__68997;
    wire N__68994;
    wire N__68991;
    wire N__68990;
    wire N__68987;
    wire N__68984;
    wire N__68981;
    wire N__68976;
    wire N__68973;
    wire N__68970;
    wire N__68967;
    wire N__68962;
    wire N__68959;
    wire N__68956;
    wire N__68953;
    wire N__68950;
    wire N__68947;
    wire N__68944;
    wire N__68941;
    wire N__68938;
    wire N__68935;
    wire N__68932;
    wire N__68929;
    wire N__68926;
    wire N__68923;
    wire N__68920;
    wire N__68917;
    wire N__68914;
    wire N__68911;
    wire N__68908;
    wire N__68907;
    wire N__68904;
    wire N__68901;
    wire N__68898;
    wire N__68895;
    wire N__68890;
    wire N__68887;
    wire N__68884;
    wire N__68881;
    wire N__68878;
    wire N__68875;
    wire N__68872;
    wire N__68869;
    wire N__68866;
    wire N__68863;
    wire N__68860;
    wire N__68857;
    wire N__68854;
    wire N__68851;
    wire N__68848;
    wire N__68845;
    wire N__68842;
    wire N__68839;
    wire N__68836;
    wire N__68833;
    wire N__68830;
    wire N__68827;
    wire N__68824;
    wire N__68821;
    wire N__68818;
    wire N__68815;
    wire N__68812;
    wire N__68809;
    wire N__68806;
    wire N__68803;
    wire N__68800;
    wire N__68797;
    wire N__68794;
    wire N__68791;
    wire N__68788;
    wire N__68785;
    wire N__68782;
    wire N__68779;
    wire N__68776;
    wire N__68773;
    wire N__68770;
    wire N__68767;
    wire N__68764;
    wire N__68761;
    wire N__68758;
    wire N__68755;
    wire N__68752;
    wire N__68749;
    wire N__68746;
    wire N__68743;
    wire N__68740;
    wire N__68737;
    wire N__68734;
    wire N__68731;
    wire N__68728;
    wire N__68725;
    wire N__68722;
    wire N__68719;
    wire N__68716;
    wire N__68713;
    wire N__68710;
    wire N__68707;
    wire N__68704;
    wire N__68701;
    wire N__68698;
    wire N__68695;
    wire N__68692;
    wire N__68689;
    wire N__68686;
    wire N__68683;
    wire N__68682;
    wire N__68681;
    wire N__68680;
    wire N__68677;
    wire N__68672;
    wire N__68671;
    wire N__68668;
    wire N__68665;
    wire N__68662;
    wire N__68659;
    wire N__68656;
    wire N__68655;
    wire N__68648;
    wire N__68647;
    wire N__68644;
    wire N__68641;
    wire N__68638;
    wire N__68635;
    wire N__68626;
    wire N__68623;
    wire N__68620;
    wire N__68617;
    wire N__68614;
    wire N__68611;
    wire N__68610;
    wire N__68609;
    wire N__68608;
    wire N__68605;
    wire N__68602;
    wire N__68597;
    wire N__68594;
    wire N__68591;
    wire N__68588;
    wire N__68585;
    wire N__68582;
    wire N__68579;
    wire N__68572;
    wire N__68569;
    wire N__68566;
    wire N__68563;
    wire N__68560;
    wire N__68559;
    wire N__68554;
    wire N__68551;
    wire N__68550;
    wire N__68549;
    wire N__68546;
    wire N__68543;
    wire N__68540;
    wire N__68533;
    wire N__68530;
    wire N__68529;
    wire N__68526;
    wire N__68523;
    wire N__68522;
    wire N__68521;
    wire N__68520;
    wire N__68519;
    wire N__68518;
    wire N__68517;
    wire N__68516;
    wire N__68515;
    wire N__68510;
    wire N__68509;
    wire N__68506;
    wire N__68505;
    wire N__68502;
    wire N__68497;
    wire N__68488;
    wire N__68485;
    wire N__68482;
    wire N__68481;
    wire N__68480;
    wire N__68479;
    wire N__68478;
    wire N__68477;
    wire N__68474;
    wire N__68471;
    wire N__68464;
    wire N__68461;
    wire N__68452;
    wire N__68447;
    wire N__68440;
    wire N__68431;
    wire N__68428;
    wire N__68425;
    wire N__68422;
    wire N__68419;
    wire N__68418;
    wire N__68415;
    wire N__68412;
    wire N__68411;
    wire N__68408;
    wire N__68405;
    wire N__68402;
    wire N__68397;
    wire N__68392;
    wire N__68389;
    wire N__68386;
    wire N__68383;
    wire N__68380;
    wire N__68377;
    wire N__68374;
    wire N__68371;
    wire N__68368;
    wire N__68365;
    wire N__68362;
    wire N__68359;
    wire N__68356;
    wire N__68353;
    wire N__68350;
    wire N__68347;
    wire N__68344;
    wire N__68341;
    wire N__68338;
    wire N__68335;
    wire N__68332;
    wire N__68329;
    wire N__68326;
    wire N__68323;
    wire N__68320;
    wire N__68317;
    wire N__68314;
    wire N__68311;
    wire N__68308;
    wire N__68305;
    wire N__68302;
    wire N__68301;
    wire N__68298;
    wire N__68295;
    wire N__68294;
    wire N__68289;
    wire N__68286;
    wire N__68285;
    wire N__68280;
    wire N__68277;
    wire N__68274;
    wire N__68271;
    wire N__68268;
    wire N__68263;
    wire N__68260;
    wire N__68257;
    wire N__68254;
    wire N__68251;
    wire N__68248;
    wire N__68245;
    wire N__68242;
    wire N__68239;
    wire N__68236;
    wire N__68233;
    wire N__68230;
    wire N__68227;
    wire N__68224;
    wire N__68221;
    wire N__68218;
    wire N__68215;
    wire N__68214;
    wire N__68211;
    wire N__68208;
    wire N__68205;
    wire N__68202;
    wire N__68197;
    wire N__68194;
    wire N__68191;
    wire N__68188;
    wire N__68185;
    wire N__68182;
    wire N__68179;
    wire N__68176;
    wire N__68173;
    wire N__68170;
    wire N__68167;
    wire N__68164;
    wire N__68161;
    wire N__68158;
    wire N__68155;
    wire N__68152;
    wire N__68149;
    wire N__68146;
    wire N__68143;
    wire N__68140;
    wire N__68137;
    wire N__68134;
    wire N__68131;
    wire N__68128;
    wire N__68125;
    wire N__68124;
    wire N__68121;
    wire N__68118;
    wire N__68115;
    wire N__68114;
    wire N__68111;
    wire N__68108;
    wire N__68105;
    wire N__68098;
    wire N__68095;
    wire N__68092;
    wire N__68089;
    wire N__68086;
    wire N__68083;
    wire N__68082;
    wire N__68079;
    wire N__68076;
    wire N__68073;
    wire N__68068;
    wire N__68065;
    wire N__68062;
    wire N__68059;
    wire N__68056;
    wire N__68053;
    wire N__68050;
    wire N__68047;
    wire N__68044;
    wire N__68041;
    wire N__68038;
    wire N__68035;
    wire N__68032;
    wire N__68029;
    wire N__68026;
    wire N__68023;
    wire N__68020;
    wire N__68017;
    wire N__68014;
    wire N__68011;
    wire N__68008;
    wire N__68005;
    wire N__68002;
    wire N__67999;
    wire N__67996;
    wire N__67993;
    wire N__67990;
    wire N__67987;
    wire N__67984;
    wire N__67981;
    wire N__67978;
    wire N__67975;
    wire N__67972;
    wire N__67969;
    wire N__67966;
    wire N__67963;
    wire N__67960;
    wire N__67957;
    wire N__67954;
    wire N__67951;
    wire N__67948;
    wire N__67945;
    wire N__67942;
    wire N__67939;
    wire N__67936;
    wire N__67933;
    wire N__67930;
    wire N__67927;
    wire N__67924;
    wire N__67921;
    wire N__67918;
    wire N__67915;
    wire N__67912;
    wire N__67909;
    wire N__67906;
    wire N__67903;
    wire N__67900;
    wire N__67897;
    wire N__67894;
    wire N__67891;
    wire N__67888;
    wire N__67885;
    wire N__67882;
    wire N__67879;
    wire N__67876;
    wire N__67873;
    wire N__67870;
    wire N__67867;
    wire N__67864;
    wire N__67861;
    wire N__67858;
    wire N__67855;
    wire N__67852;
    wire N__67849;
    wire N__67846;
    wire N__67843;
    wire N__67840;
    wire N__67837;
    wire N__67834;
    wire N__67831;
    wire N__67828;
    wire N__67825;
    wire N__67822;
    wire N__67819;
    wire N__67816;
    wire N__67813;
    wire N__67810;
    wire N__67807;
    wire N__67804;
    wire N__67801;
    wire N__67798;
    wire N__67795;
    wire N__67792;
    wire N__67789;
    wire N__67786;
    wire N__67783;
    wire N__67780;
    wire N__67777;
    wire N__67774;
    wire N__67771;
    wire N__67768;
    wire N__67765;
    wire N__67762;
    wire N__67761;
    wire N__67758;
    wire N__67755;
    wire N__67752;
    wire N__67749;
    wire N__67744;
    wire N__67741;
    wire N__67738;
    wire N__67735;
    wire N__67732;
    wire N__67729;
    wire N__67726;
    wire N__67723;
    wire N__67720;
    wire N__67717;
    wire N__67716;
    wire N__67713;
    wire N__67710;
    wire N__67705;
    wire N__67704;
    wire N__67699;
    wire N__67696;
    wire N__67693;
    wire N__67690;
    wire N__67687;
    wire N__67684;
    wire N__67681;
    wire N__67678;
    wire N__67675;
    wire N__67672;
    wire N__67669;
    wire N__67666;
    wire N__67663;
    wire N__67660;
    wire N__67657;
    wire N__67654;
    wire N__67651;
    wire N__67650;
    wire N__67647;
    wire N__67644;
    wire N__67641;
    wire N__67640;
    wire N__67637;
    wire N__67634;
    wire N__67631;
    wire N__67628;
    wire N__67625;
    wire N__67622;
    wire N__67615;
    wire N__67612;
    wire N__67609;
    wire N__67606;
    wire N__67603;
    wire N__67600;
    wire N__67597;
    wire N__67594;
    wire N__67591;
    wire N__67588;
    wire N__67585;
    wire N__67582;
    wire N__67579;
    wire N__67576;
    wire N__67573;
    wire N__67570;
    wire N__67567;
    wire N__67564;
    wire N__67561;
    wire N__67558;
    wire N__67555;
    wire N__67554;
    wire N__67551;
    wire N__67548;
    wire N__67543;
    wire N__67540;
    wire N__67537;
    wire N__67534;
    wire N__67531;
    wire N__67528;
    wire N__67525;
    wire N__67524;
    wire N__67519;
    wire N__67516;
    wire N__67513;
    wire N__67510;
    wire N__67507;
    wire N__67504;
    wire N__67501;
    wire N__67498;
    wire N__67495;
    wire N__67492;
    wire N__67489;
    wire N__67486;
    wire N__67483;
    wire N__67480;
    wire N__67477;
    wire N__67474;
    wire N__67471;
    wire N__67468;
    wire N__67465;
    wire N__67462;
    wire N__67459;
    wire N__67456;
    wire N__67453;
    wire N__67450;
    wire N__67447;
    wire N__67444;
    wire N__67441;
    wire N__67438;
    wire N__67435;
    wire N__67432;
    wire N__67429;
    wire N__67426;
    wire N__67423;
    wire N__67420;
    wire N__67417;
    wire N__67414;
    wire N__67411;
    wire N__67408;
    wire N__67405;
    wire N__67402;
    wire N__67399;
    wire N__67396;
    wire N__67393;
    wire N__67390;
    wire N__67387;
    wire N__67384;
    wire N__67381;
    wire N__67378;
    wire N__67375;
    wire N__67372;
    wire N__67369;
    wire N__67366;
    wire N__67363;
    wire N__67360;
    wire N__67357;
    wire N__67354;
    wire N__67353;
    wire N__67350;
    wire N__67347;
    wire N__67344;
    wire N__67341;
    wire N__67338;
    wire N__67335;
    wire N__67330;
    wire N__67327;
    wire N__67324;
    wire N__67321;
    wire N__67318;
    wire N__67315;
    wire N__67312;
    wire N__67309;
    wire N__67306;
    wire N__67303;
    wire N__67302;
    wire N__67299;
    wire N__67296;
    wire N__67295;
    wire N__67292;
    wire N__67289;
    wire N__67286;
    wire N__67283;
    wire N__67280;
    wire N__67277;
    wire N__67270;
    wire N__67267;
    wire N__67264;
    wire N__67261;
    wire N__67258;
    wire N__67255;
    wire N__67252;
    wire N__67249;
    wire N__67246;
    wire N__67243;
    wire N__67240;
    wire N__67237;
    wire N__67236;
    wire N__67235;
    wire N__67232;
    wire N__67229;
    wire N__67226;
    wire N__67219;
    wire N__67216;
    wire N__67213;
    wire N__67210;
    wire N__67207;
    wire N__67204;
    wire N__67201;
    wire N__67198;
    wire N__67195;
    wire N__67192;
    wire N__67189;
    wire N__67186;
    wire N__67183;
    wire N__67180;
    wire N__67177;
    wire N__67174;
    wire N__67171;
    wire N__67170;
    wire N__67169;
    wire N__67166;
    wire N__67163;
    wire N__67160;
    wire N__67157;
    wire N__67154;
    wire N__67151;
    wire N__67144;
    wire N__67143;
    wire N__67140;
    wire N__67137;
    wire N__67136;
    wire N__67133;
    wire N__67130;
    wire N__67127;
    wire N__67124;
    wire N__67117;
    wire N__67114;
    wire N__67111;
    wire N__67110;
    wire N__67107;
    wire N__67106;
    wire N__67105;
    wire N__67104;
    wire N__67101;
    wire N__67100;
    wire N__67099;
    wire N__67096;
    wire N__67093;
    wire N__67088;
    wire N__67085;
    wire N__67080;
    wire N__67077;
    wire N__67072;
    wire N__67063;
    wire N__67062;
    wire N__67061;
    wire N__67058;
    wire N__67057;
    wire N__67054;
    wire N__67051;
    wire N__67048;
    wire N__67047;
    wire N__67044;
    wire N__67041;
    wire N__67038;
    wire N__67035;
    wire N__67032;
    wire N__67025;
    wire N__67018;
    wire N__67015;
    wire N__67012;
    wire N__67011;
    wire N__67008;
    wire N__67007;
    wire N__67004;
    wire N__67001;
    wire N__66998;
    wire N__66991;
    wire N__66988;
    wire N__66987;
    wire N__66986;
    wire N__66985;
    wire N__66982;
    wire N__66977;
    wire N__66974;
    wire N__66973;
    wire N__66970;
    wire N__66967;
    wire N__66964;
    wire N__66961;
    wire N__66958;
    wire N__66955;
    wire N__66946;
    wire N__66945;
    wire N__66942;
    wire N__66939;
    wire N__66938;
    wire N__66935;
    wire N__66932;
    wire N__66929;
    wire N__66926;
    wire N__66923;
    wire N__66916;
    wire N__66915;
    wire N__66914;
    wire N__66911;
    wire N__66908;
    wire N__66905;
    wire N__66904;
    wire N__66901;
    wire N__66898;
    wire N__66895;
    wire N__66894;
    wire N__66891;
    wire N__66886;
    wire N__66883;
    wire N__66880;
    wire N__66877;
    wire N__66874;
    wire N__66865;
    wire N__66862;
    wire N__66859;
    wire N__66856;
    wire N__66853;
    wire N__66850;
    wire N__66847;
    wire N__66844;
    wire N__66841;
    wire N__66838;
    wire N__66835;
    wire N__66832;
    wire N__66829;
    wire N__66826;
    wire N__66823;
    wire N__66820;
    wire N__66817;
    wire N__66814;
    wire N__66811;
    wire N__66808;
    wire N__66807;
    wire N__66806;
    wire N__66805;
    wire N__66804;
    wire N__66801;
    wire N__66800;
    wire N__66797;
    wire N__66794;
    wire N__66791;
    wire N__66784;
    wire N__66779;
    wire N__66776;
    wire N__66773;
    wire N__66770;
    wire N__66767;
    wire N__66764;
    wire N__66761;
    wire N__66756;
    wire N__66751;
    wire N__66748;
    wire N__66745;
    wire N__66742;
    wire N__66739;
    wire N__66736;
    wire N__66733;
    wire N__66730;
    wire N__66727;
    wire N__66724;
    wire N__66721;
    wire N__66718;
    wire N__66715;
    wire N__66712;
    wire N__66709;
    wire N__66706;
    wire N__66703;
    wire N__66700;
    wire N__66697;
    wire N__66694;
    wire N__66691;
    wire N__66688;
    wire N__66685;
    wire N__66682;
    wire N__66679;
    wire N__66676;
    wire N__66673;
    wire N__66670;
    wire N__66667;
    wire N__66664;
    wire N__66661;
    wire N__66658;
    wire N__66655;
    wire N__66652;
    wire N__66649;
    wire N__66646;
    wire N__66643;
    wire N__66640;
    wire N__66637;
    wire N__66634;
    wire N__66631;
    wire N__66628;
    wire N__66625;
    wire N__66622;
    wire N__66621;
    wire N__66618;
    wire N__66615;
    wire N__66612;
    wire N__66611;
    wire N__66608;
    wire N__66607;
    wire N__66604;
    wire N__66603;
    wire N__66602;
    wire N__66601;
    wire N__66600;
    wire N__66597;
    wire N__66594;
    wire N__66591;
    wire N__66588;
    wire N__66579;
    wire N__66576;
    wire N__66571;
    wire N__66562;
    wire N__66559;
    wire N__66556;
    wire N__66553;
    wire N__66550;
    wire N__66547;
    wire N__66544;
    wire N__66541;
    wire N__66540;
    wire N__66537;
    wire N__66536;
    wire N__66533;
    wire N__66530;
    wire N__66527;
    wire N__66524;
    wire N__66521;
    wire N__66516;
    wire N__66511;
    wire N__66508;
    wire N__66505;
    wire N__66502;
    wire N__66499;
    wire N__66496;
    wire N__66495;
    wire N__66492;
    wire N__66489;
    wire N__66486;
    wire N__66483;
    wire N__66480;
    wire N__66477;
    wire N__66474;
    wire N__66471;
    wire N__66466;
    wire N__66463;
    wire N__66462;
    wire N__66461;
    wire N__66460;
    wire N__66457;
    wire N__66456;
    wire N__66455;
    wire N__66454;
    wire N__66451;
    wire N__66448;
    wire N__66447;
    wire N__66444;
    wire N__66443;
    wire N__66442;
    wire N__66441;
    wire N__66438;
    wire N__66433;
    wire N__66430;
    wire N__66427;
    wire N__66424;
    wire N__66419;
    wire N__66416;
    wire N__66415;
    wire N__66412;
    wire N__66409;
    wire N__66406;
    wire N__66403;
    wire N__66398;
    wire N__66393;
    wire N__66392;
    wire N__66391;
    wire N__66388;
    wire N__66387;
    wire N__66386;
    wire N__66383;
    wire N__66380;
    wire N__66377;
    wire N__66372;
    wire N__66369;
    wire N__66366;
    wire N__66361;
    wire N__66358;
    wire N__66353;
    wire N__66334;
    wire N__66331;
    wire N__66328;
    wire N__66325;
    wire N__66322;
    wire N__66319;
    wire N__66316;
    wire N__66313;
    wire N__66310;
    wire N__66309;
    wire N__66306;
    wire N__66303;
    wire N__66302;
    wire N__66301;
    wire N__66300;
    wire N__66299;
    wire N__66296;
    wire N__66293;
    wire N__66286;
    wire N__66283;
    wire N__66278;
    wire N__66273;
    wire N__66270;
    wire N__66267;
    wire N__66262;
    wire N__66259;
    wire N__66258;
    wire N__66257;
    wire N__66254;
    wire N__66251;
    wire N__66248;
    wire N__66245;
    wire N__66244;
    wire N__66243;
    wire N__66242;
    wire N__66241;
    wire N__66238;
    wire N__66237;
    wire N__66234;
    wire N__66231;
    wire N__66226;
    wire N__66223;
    wire N__66220;
    wire N__66217;
    wire N__66214;
    wire N__66211;
    wire N__66202;
    wire N__66199;
    wire N__66196;
    wire N__66191;
    wire N__66184;
    wire N__66181;
    wire N__66178;
    wire N__66175;
    wire N__66172;
    wire N__66169;
    wire N__66166;
    wire N__66163;
    wire N__66160;
    wire N__66157;
    wire N__66154;
    wire N__66151;
    wire N__66148;
    wire N__66145;
    wire N__66142;
    wire N__66139;
    wire N__66136;
    wire N__66133;
    wire N__66130;
    wire N__66127;
    wire N__66124;
    wire N__66121;
    wire N__66118;
    wire N__66115;
    wire N__66112;
    wire N__66109;
    wire N__66106;
    wire N__66103;
    wire N__66100;
    wire N__66097;
    wire N__66094;
    wire N__66091;
    wire N__66088;
    wire N__66085;
    wire N__66082;
    wire N__66079;
    wire N__66076;
    wire N__66073;
    wire N__66070;
    wire N__66067;
    wire N__66064;
    wire N__66063;
    wire N__66062;
    wire N__66061;
    wire N__66058;
    wire N__66053;
    wire N__66050;
    wire N__66047;
    wire N__66044;
    wire N__66037;
    wire N__66036;
    wire N__66033;
    wire N__66030;
    wire N__66029;
    wire N__66028;
    wire N__66025;
    wire N__66022;
    wire N__66019;
    wire N__66016;
    wire N__66015;
    wire N__66014;
    wire N__66011;
    wire N__66008;
    wire N__66005;
    wire N__66000;
    wire N__65997;
    wire N__65992;
    wire N__65987;
    wire N__65980;
    wire N__65977;
    wire N__65974;
    wire N__65973;
    wire N__65972;
    wire N__65971;
    wire N__65970;
    wire N__65967;
    wire N__65962;
    wire N__65957;
    wire N__65954;
    wire N__65949;
    wire N__65948;
    wire N__65947;
    wire N__65944;
    wire N__65941;
    wire N__65936;
    wire N__65929;
    wire N__65926;
    wire N__65923;
    wire N__65920;
    wire N__65917;
    wire N__65914;
    wire N__65911;
    wire N__65908;
    wire N__65905;
    wire N__65904;
    wire N__65903;
    wire N__65902;
    wire N__65899;
    wire N__65896;
    wire N__65891;
    wire N__65890;
    wire N__65883;
    wire N__65882;
    wire N__65879;
    wire N__65876;
    wire N__65871;
    wire N__65866;
    wire N__65863;
    wire N__65860;
    wire N__65859;
    wire N__65856;
    wire N__65855;
    wire N__65852;
    wire N__65851;
    wire N__65848;
    wire N__65845;
    wire N__65844;
    wire N__65843;
    wire N__65838;
    wire N__65833;
    wire N__65830;
    wire N__65827;
    wire N__65822;
    wire N__65815;
    wire N__65812;
    wire N__65809;
    wire N__65806;
    wire N__65803;
    wire N__65800;
    wire N__65797;
    wire N__65794;
    wire N__65791;
    wire N__65788;
    wire N__65785;
    wire N__65782;
    wire N__65779;
    wire N__65776;
    wire N__65773;
    wire N__65770;
    wire N__65767;
    wire N__65764;
    wire N__65761;
    wire N__65758;
    wire N__65755;
    wire N__65754;
    wire N__65753;
    wire N__65752;
    wire N__65751;
    wire N__65750;
    wire N__65747;
    wire N__65746;
    wire N__65743;
    wire N__65742;
    wire N__65741;
    wire N__65740;
    wire N__65739;
    wire N__65734;
    wire N__65729;
    wire N__65728;
    wire N__65725;
    wire N__65718;
    wire N__65717;
    wire N__65716;
    wire N__65713;
    wire N__65710;
    wire N__65709;
    wire N__65706;
    wire N__65703;
    wire N__65700;
    wire N__65697;
    wire N__65692;
    wire N__65689;
    wire N__65686;
    wire N__65683;
    wire N__65680;
    wire N__65677;
    wire N__65674;
    wire N__65669;
    wire N__65662;
    wire N__65659;
    wire N__65658;
    wire N__65655;
    wire N__65652;
    wire N__65649;
    wire N__65646;
    wire N__65641;
    wire N__65638;
    wire N__65635;
    wire N__65630;
    wire N__65623;
    wire N__65614;
    wire N__65611;
    wire N__65608;
    wire N__65605;
    wire N__65604;
    wire N__65603;
    wire N__65602;
    wire N__65599;
    wire N__65596;
    wire N__65593;
    wire N__65590;
    wire N__65587;
    wire N__65584;
    wire N__65581;
    wire N__65572;
    wire N__65569;
    wire N__65568;
    wire N__65567;
    wire N__65566;
    wire N__65563;
    wire N__65560;
    wire N__65557;
    wire N__65554;
    wire N__65553;
    wire N__65552;
    wire N__65551;
    wire N__65550;
    wire N__65547;
    wire N__65544;
    wire N__65541;
    wire N__65538;
    wire N__65533;
    wire N__65530;
    wire N__65527;
    wire N__65524;
    wire N__65523;
    wire N__65518;
    wire N__65515;
    wire N__65514;
    wire N__65511;
    wire N__65508;
    wire N__65505;
    wire N__65502;
    wire N__65499;
    wire N__65496;
    wire N__65493;
    wire N__65490;
    wire N__65485;
    wire N__65482;
    wire N__65477;
    wire N__65474;
    wire N__65471;
    wire N__65458;
    wire N__65457;
    wire N__65454;
    wire N__65453;
    wire N__65450;
    wire N__65447;
    wire N__65444;
    wire N__65441;
    wire N__65440;
    wire N__65439;
    wire N__65436;
    wire N__65433;
    wire N__65430;
    wire N__65427;
    wire N__65424;
    wire N__65421;
    wire N__65418;
    wire N__65413;
    wire N__65412;
    wire N__65411;
    wire N__65410;
    wire N__65407;
    wire N__65402;
    wire N__65399;
    wire N__65392;
    wire N__65383;
    wire N__65380;
    wire N__65379;
    wire N__65376;
    wire N__65375;
    wire N__65374;
    wire N__65371;
    wire N__65370;
    wire N__65365;
    wire N__65364;
    wire N__65363;
    wire N__65362;
    wire N__65359;
    wire N__65358;
    wire N__65355;
    wire N__65352;
    wire N__65349;
    wire N__65348;
    wire N__65345;
    wire N__65342;
    wire N__65341;
    wire N__65338;
    wire N__65335;
    wire N__65332;
    wire N__65329;
    wire N__65326;
    wire N__65323;
    wire N__65320;
    wire N__65317;
    wire N__65314;
    wire N__65311;
    wire N__65310;
    wire N__65307;
    wire N__65302;
    wire N__65301;
    wire N__65294;
    wire N__65291;
    wire N__65286;
    wire N__65283;
    wire N__65280;
    wire N__65277;
    wire N__65274;
    wire N__65271;
    wire N__65268;
    wire N__65261;
    wire N__65254;
    wire N__65245;
    wire N__65242;
    wire N__65239;
    wire N__65236;
    wire N__65233;
    wire N__65230;
    wire N__65227;
    wire N__65224;
    wire N__65221;
    wire N__65218;
    wire N__65215;
    wire N__65212;
    wire N__65209;
    wire N__65206;
    wire N__65203;
    wire N__65200;
    wire N__65197;
    wire N__65194;
    wire N__65191;
    wire N__65190;
    wire N__65187;
    wire N__65186;
    wire N__65183;
    wire N__65180;
    wire N__65177;
    wire N__65174;
    wire N__65171;
    wire N__65168;
    wire N__65161;
    wire N__65158;
    wire N__65155;
    wire N__65152;
    wire N__65149;
    wire N__65146;
    wire N__65143;
    wire N__65140;
    wire N__65137;
    wire N__65134;
    wire N__65131;
    wire N__65128;
    wire N__65125;
    wire N__65122;
    wire N__65119;
    wire N__65116;
    wire N__65113;
    wire N__65110;
    wire N__65107;
    wire N__65104;
    wire N__65101;
    wire N__65098;
    wire N__65095;
    wire N__65092;
    wire N__65089;
    wire N__65086;
    wire N__65083;
    wire N__65080;
    wire N__65077;
    wire N__65074;
    wire N__65071;
    wire N__65068;
    wire N__65065;
    wire N__65064;
    wire N__65061;
    wire N__65060;
    wire N__65057;
    wire N__65054;
    wire N__65051;
    wire N__65048;
    wire N__65043;
    wire N__65040;
    wire N__65037;
    wire N__65032;
    wire N__65029;
    wire N__65028;
    wire N__65027;
    wire N__65024;
    wire N__65023;
    wire N__65022;
    wire N__65021;
    wire N__65020;
    wire N__65017;
    wire N__65014;
    wire N__65011;
    wire N__65002;
    wire N__64997;
    wire N__64990;
    wire N__64987;
    wire N__64986;
    wire N__64985;
    wire N__64984;
    wire N__64983;
    wire N__64980;
    wire N__64979;
    wire N__64978;
    wire N__64977;
    wire N__64976;
    wire N__64975;
    wire N__64968;
    wire N__64965;
    wire N__64962;
    wire N__64955;
    wire N__64952;
    wire N__64951;
    wire N__64950;
    wire N__64949;
    wire N__64948;
    wire N__64947;
    wire N__64946;
    wire N__64945;
    wire N__64944;
    wire N__64943;
    wire N__64940;
    wire N__64937;
    wire N__64934;
    wire N__64927;
    wire N__64924;
    wire N__64921;
    wire N__64918;
    wire N__64909;
    wire N__64904;
    wire N__64899;
    wire N__64894;
    wire N__64879;
    wire N__64878;
    wire N__64877;
    wire N__64876;
    wire N__64873;
    wire N__64870;
    wire N__64867;
    wire N__64864;
    wire N__64855;
    wire N__64852;
    wire N__64849;
    wire N__64846;
    wire N__64843;
    wire N__64840;
    wire N__64837;
    wire N__64834;
    wire N__64831;
    wire N__64828;
    wire N__64827;
    wire N__64824;
    wire N__64821;
    wire N__64820;
    wire N__64815;
    wire N__64812;
    wire N__64811;
    wire N__64808;
    wire N__64805;
    wire N__64802;
    wire N__64801;
    wire N__64796;
    wire N__64793;
    wire N__64790;
    wire N__64787;
    wire N__64784;
    wire N__64781;
    wire N__64774;
    wire N__64771;
    wire N__64768;
    wire N__64765;
    wire N__64762;
    wire N__64759;
    wire N__64756;
    wire N__64753;
    wire N__64750;
    wire N__64747;
    wire N__64744;
    wire N__64741;
    wire N__64738;
    wire N__64735;
    wire N__64732;
    wire N__64729;
    wire N__64726;
    wire N__64723;
    wire N__64720;
    wire N__64717;
    wire N__64714;
    wire N__64711;
    wire N__64708;
    wire N__64705;
    wire N__64702;
    wire N__64699;
    wire N__64696;
    wire N__64693;
    wire N__64690;
    wire N__64687;
    wire N__64684;
    wire N__64681;
    wire N__64678;
    wire N__64677;
    wire N__64674;
    wire N__64671;
    wire N__64666;
    wire N__64663;
    wire N__64660;
    wire N__64657;
    wire N__64654;
    wire N__64651;
    wire N__64648;
    wire N__64645;
    wire N__64642;
    wire N__64639;
    wire N__64636;
    wire N__64633;
    wire N__64630;
    wire N__64627;
    wire N__64624;
    wire N__64621;
    wire N__64618;
    wire N__64615;
    wire N__64612;
    wire N__64609;
    wire N__64606;
    wire N__64603;
    wire N__64600;
    wire N__64597;
    wire N__64594;
    wire N__64591;
    wire N__64588;
    wire N__64585;
    wire N__64582;
    wire N__64579;
    wire N__64576;
    wire N__64573;
    wire N__64570;
    wire N__64567;
    wire N__64564;
    wire N__64561;
    wire N__64558;
    wire N__64555;
    wire N__64552;
    wire N__64549;
    wire N__64546;
    wire N__64543;
    wire N__64540;
    wire N__64537;
    wire N__64534;
    wire N__64531;
    wire N__64528;
    wire N__64525;
    wire N__64522;
    wire N__64519;
    wire N__64516;
    wire N__64513;
    wire N__64510;
    wire N__64507;
    wire N__64504;
    wire N__64501;
    wire N__64498;
    wire N__64495;
    wire N__64492;
    wire N__64489;
    wire N__64486;
    wire N__64483;
    wire N__64480;
    wire N__64477;
    wire N__64474;
    wire N__64471;
    wire N__64468;
    wire N__64465;
    wire N__64462;
    wire N__64459;
    wire N__64456;
    wire N__64453;
    wire N__64450;
    wire N__64447;
    wire N__64444;
    wire N__64441;
    wire N__64438;
    wire N__64435;
    wire N__64432;
    wire N__64429;
    wire N__64426;
    wire N__64423;
    wire N__64420;
    wire N__64417;
    wire N__64414;
    wire N__64411;
    wire N__64410;
    wire N__64407;
    wire N__64404;
    wire N__64401;
    wire N__64398;
    wire N__64393;
    wire N__64390;
    wire N__64387;
    wire N__64384;
    wire N__64381;
    wire N__64378;
    wire N__64375;
    wire N__64372;
    wire N__64369;
    wire N__64366;
    wire N__64363;
    wire N__64360;
    wire N__64357;
    wire N__64354;
    wire N__64351;
    wire N__64348;
    wire N__64345;
    wire N__64342;
    wire N__64339;
    wire N__64336;
    wire N__64333;
    wire N__64330;
    wire N__64327;
    wire N__64326;
    wire N__64323;
    wire N__64320;
    wire N__64317;
    wire N__64314;
    wire N__64311;
    wire N__64308;
    wire N__64303;
    wire N__64300;
    wire N__64297;
    wire N__64294;
    wire N__64291;
    wire N__64288;
    wire N__64285;
    wire N__64282;
    wire N__64279;
    wire N__64276;
    wire N__64273;
    wire N__64270;
    wire N__64267;
    wire N__64264;
    wire N__64261;
    wire N__64258;
    wire N__64255;
    wire N__64252;
    wire N__64249;
    wire N__64246;
    wire N__64243;
    wire N__64240;
    wire N__64239;
    wire N__64236;
    wire N__64233;
    wire N__64230;
    wire N__64227;
    wire N__64222;
    wire N__64219;
    wire N__64216;
    wire N__64213;
    wire N__64210;
    wire N__64207;
    wire N__64204;
    wire N__64201;
    wire N__64198;
    wire N__64195;
    wire N__64192;
    wire N__64189;
    wire N__64186;
    wire N__64183;
    wire N__64180;
    wire N__64177;
    wire N__64174;
    wire N__64171;
    wire N__64168;
    wire N__64165;
    wire N__64162;
    wire N__64159;
    wire N__64156;
    wire N__64153;
    wire N__64150;
    wire N__64147;
    wire N__64144;
    wire N__64141;
    wire N__64138;
    wire N__64135;
    wire N__64132;
    wire N__64129;
    wire N__64126;
    wire N__64123;
    wire N__64120;
    wire N__64117;
    wire N__64114;
    wire N__64111;
    wire N__64108;
    wire N__64105;
    wire N__64102;
    wire N__64099;
    wire N__64096;
    wire N__64093;
    wire N__64090;
    wire N__64087;
    wire N__64084;
    wire N__64081;
    wire N__64080;
    wire N__64077;
    wire N__64074;
    wire N__64073;
    wire N__64070;
    wire N__64067;
    wire N__64064;
    wire N__64061;
    wire N__64058;
    wire N__64055;
    wire N__64048;
    wire N__64045;
    wire N__64042;
    wire N__64039;
    wire N__64036;
    wire N__64033;
    wire N__64030;
    wire N__64027;
    wire N__64024;
    wire N__64021;
    wire N__64018;
    wire N__64015;
    wire N__64012;
    wire N__64009;
    wire N__64006;
    wire N__64003;
    wire N__64000;
    wire N__63997;
    wire N__63994;
    wire N__63991;
    wire N__63988;
    wire N__63985;
    wire N__63982;
    wire N__63979;
    wire N__63976;
    wire N__63973;
    wire N__63970;
    wire N__63967;
    wire N__63964;
    wire N__63961;
    wire N__63958;
    wire N__63955;
    wire N__63952;
    wire N__63949;
    wire N__63946;
    wire N__63943;
    wire N__63940;
    wire N__63937;
    wire N__63934;
    wire N__63931;
    wire N__63928;
    wire N__63925;
    wire N__63922;
    wire N__63919;
    wire N__63916;
    wire N__63913;
    wire N__63910;
    wire N__63907;
    wire N__63904;
    wire N__63901;
    wire N__63898;
    wire N__63895;
    wire N__63892;
    wire N__63889;
    wire N__63886;
    wire N__63883;
    wire N__63880;
    wire N__63877;
    wire N__63874;
    wire N__63873;
    wire N__63870;
    wire N__63867;
    wire N__63864;
    wire N__63861;
    wire N__63856;
    wire N__63853;
    wire N__63850;
    wire N__63847;
    wire N__63844;
    wire N__63841;
    wire N__63838;
    wire N__63835;
    wire N__63834;
    wire N__63833;
    wire N__63832;
    wire N__63827;
    wire N__63822;
    wire N__63819;
    wire N__63818;
    wire N__63815;
    wire N__63814;
    wire N__63813;
    wire N__63812;
    wire N__63811;
    wire N__63810;
    wire N__63809;
    wire N__63806;
    wire N__63803;
    wire N__63800;
    wire N__63797;
    wire N__63794;
    wire N__63791;
    wire N__63784;
    wire N__63775;
    wire N__63766;
    wire N__63765;
    wire N__63764;
    wire N__63763;
    wire N__63762;
    wire N__63761;
    wire N__63758;
    wire N__63755;
    wire N__63754;
    wire N__63749;
    wire N__63748;
    wire N__63745;
    wire N__63738;
    wire N__63735;
    wire N__63732;
    wire N__63729;
    wire N__63722;
    wire N__63719;
    wire N__63716;
    wire N__63711;
    wire N__63706;
    wire N__63703;
    wire N__63700;
    wire N__63697;
    wire N__63694;
    wire N__63691;
    wire N__63688;
    wire N__63685;
    wire N__63682;
    wire N__63679;
    wire N__63676;
    wire N__63673;
    wire N__63670;
    wire N__63667;
    wire N__63664;
    wire N__63661;
    wire N__63658;
    wire N__63655;
    wire N__63654;
    wire N__63651;
    wire N__63648;
    wire N__63645;
    wire N__63642;
    wire N__63639;
    wire N__63634;
    wire N__63631;
    wire N__63628;
    wire N__63625;
    wire N__63622;
    wire N__63621;
    wire N__63618;
    wire N__63615;
    wire N__63612;
    wire N__63609;
    wire N__63606;
    wire N__63603;
    wire N__63598;
    wire N__63595;
    wire N__63592;
    wire N__63591;
    wire N__63590;
    wire N__63587;
    wire N__63584;
    wire N__63583;
    wire N__63580;
    wire N__63575;
    wire N__63572;
    wire N__63567;
    wire N__63562;
    wire N__63559;
    wire N__63556;
    wire N__63553;
    wire N__63550;
    wire N__63547;
    wire N__63544;
    wire N__63541;
    wire N__63538;
    wire N__63535;
    wire N__63532;
    wire N__63529;
    wire N__63526;
    wire N__63523;
    wire N__63520;
    wire N__63517;
    wire N__63514;
    wire N__63513;
    wire N__63510;
    wire N__63507;
    wire N__63504;
    wire N__63501;
    wire N__63496;
    wire N__63493;
    wire N__63490;
    wire N__63487;
    wire N__63484;
    wire N__63481;
    wire N__63478;
    wire N__63475;
    wire N__63472;
    wire N__63469;
    wire N__63466;
    wire N__63463;
    wire N__63460;
    wire N__63457;
    wire N__63454;
    wire N__63451;
    wire N__63448;
    wire N__63445;
    wire N__63442;
    wire N__63439;
    wire N__63436;
    wire N__63433;
    wire N__63430;
    wire N__63427;
    wire N__63424;
    wire N__63423;
    wire N__63420;
    wire N__63417;
    wire N__63412;
    wire N__63409;
    wire N__63408;
    wire N__63407;
    wire N__63406;
    wire N__63405;
    wire N__63402;
    wire N__63397;
    wire N__63394;
    wire N__63391;
    wire N__63386;
    wire N__63383;
    wire N__63376;
    wire N__63373;
    wire N__63370;
    wire N__63367;
    wire N__63364;
    wire N__63361;
    wire N__63358;
    wire N__63357;
    wire N__63354;
    wire N__63351;
    wire N__63348;
    wire N__63345;
    wire N__63342;
    wire N__63339;
    wire N__63336;
    wire N__63331;
    wire N__63328;
    wire N__63325;
    wire N__63322;
    wire N__63319;
    wire N__63316;
    wire N__63313;
    wire N__63310;
    wire N__63307;
    wire N__63304;
    wire N__63301;
    wire N__63298;
    wire N__63295;
    wire N__63292;
    wire N__63289;
    wire N__63286;
    wire N__63283;
    wire N__63280;
    wire N__63277;
    wire N__63274;
    wire N__63271;
    wire N__63268;
    wire N__63265;
    wire N__63262;
    wire N__63259;
    wire N__63256;
    wire N__63253;
    wire N__63252;
    wire N__63249;
    wire N__63248;
    wire N__63245;
    wire N__63242;
    wire N__63241;
    wire N__63238;
    wire N__63235;
    wire N__63232;
    wire N__63229;
    wire N__63226;
    wire N__63223;
    wire N__63214;
    wire N__63211;
    wire N__63210;
    wire N__63207;
    wire N__63204;
    wire N__63199;
    wire N__63196;
    wire N__63193;
    wire N__63192;
    wire N__63189;
    wire N__63186;
    wire N__63181;
    wire N__63178;
    wire N__63175;
    wire N__63172;
    wire N__63169;
    wire N__63166;
    wire N__63163;
    wire N__63160;
    wire N__63157;
    wire N__63154;
    wire N__63151;
    wire N__63150;
    wire N__63149;
    wire N__63146;
    wire N__63143;
    wire N__63140;
    wire N__63135;
    wire N__63132;
    wire N__63129;
    wire N__63124;
    wire N__63121;
    wire N__63118;
    wire N__63115;
    wire N__63112;
    wire N__63109;
    wire N__63106;
    wire N__63103;
    wire N__63100;
    wire N__63097;
    wire N__63094;
    wire N__63091;
    wire N__63088;
    wire N__63085;
    wire N__63082;
    wire N__63079;
    wire N__63076;
    wire N__63073;
    wire N__63070;
    wire N__63067;
    wire N__63064;
    wire N__63061;
    wire N__63058;
    wire N__63055;
    wire N__63052;
    wire N__63049;
    wire N__63046;
    wire N__63043;
    wire N__63040;
    wire N__63037;
    wire N__63034;
    wire N__63031;
    wire N__63028;
    wire N__63025;
    wire N__63022;
    wire N__63019;
    wire N__63016;
    wire N__63013;
    wire N__63010;
    wire N__63007;
    wire N__63004;
    wire N__63001;
    wire N__62998;
    wire N__62995;
    wire N__62992;
    wire N__62989;
    wire N__62986;
    wire N__62983;
    wire N__62980;
    wire N__62977;
    wire N__62974;
    wire N__62971;
    wire N__62968;
    wire N__62965;
    wire N__62962;
    wire N__62959;
    wire N__62956;
    wire N__62953;
    wire N__62950;
    wire N__62947;
    wire N__62944;
    wire N__62941;
    wire N__62938;
    wire N__62935;
    wire N__62932;
    wire N__62929;
    wire N__62926;
    wire N__62923;
    wire N__62920;
    wire N__62917;
    wire N__62914;
    wire N__62911;
    wire N__62908;
    wire N__62905;
    wire N__62902;
    wire N__62899;
    wire N__62896;
    wire N__62893;
    wire N__62890;
    wire N__62889;
    wire N__62888;
    wire N__62885;
    wire N__62882;
    wire N__62881;
    wire N__62878;
    wire N__62877;
    wire N__62872;
    wire N__62865;
    wire N__62860;
    wire N__62859;
    wire N__62858;
    wire N__62855;
    wire N__62850;
    wire N__62845;
    wire N__62842;
    wire N__62839;
    wire N__62836;
    wire N__62833;
    wire N__62830;
    wire N__62827;
    wire N__62824;
    wire N__62821;
    wire N__62818;
    wire N__62815;
    wire N__62812;
    wire N__62809;
    wire N__62806;
    wire N__62803;
    wire N__62800;
    wire N__62797;
    wire N__62794;
    wire N__62791;
    wire N__62788;
    wire N__62785;
    wire N__62782;
    wire N__62779;
    wire N__62776;
    wire N__62773;
    wire N__62770;
    wire N__62767;
    wire N__62764;
    wire N__62761;
    wire N__62758;
    wire N__62755;
    wire N__62752;
    wire N__62749;
    wire N__62746;
    wire N__62743;
    wire N__62740;
    wire N__62737;
    wire N__62734;
    wire N__62731;
    wire N__62728;
    wire N__62725;
    wire N__62722;
    wire N__62721;
    wire N__62720;
    wire N__62717;
    wire N__62714;
    wire N__62711;
    wire N__62704;
    wire N__62703;
    wire N__62702;
    wire N__62699;
    wire N__62698;
    wire N__62697;
    wire N__62696;
    wire N__62693;
    wire N__62690;
    wire N__62687;
    wire N__62680;
    wire N__62671;
    wire N__62668;
    wire N__62665;
    wire N__62662;
    wire N__62659;
    wire N__62656;
    wire N__62653;
    wire N__62650;
    wire N__62647;
    wire N__62644;
    wire N__62641;
    wire N__62638;
    wire N__62635;
    wire N__62632;
    wire N__62629;
    wire N__62626;
    wire N__62623;
    wire N__62620;
    wire N__62617;
    wire N__62614;
    wire N__62611;
    wire N__62610;
    wire N__62607;
    wire N__62604;
    wire N__62601;
    wire N__62598;
    wire N__62593;
    wire N__62590;
    wire N__62589;
    wire N__62588;
    wire N__62587;
    wire N__62586;
    wire N__62585;
    wire N__62582;
    wire N__62577;
    wire N__62574;
    wire N__62569;
    wire N__62566;
    wire N__62561;
    wire N__62558;
    wire N__62555;
    wire N__62552;
    wire N__62549;
    wire N__62542;
    wire N__62539;
    wire N__62536;
    wire N__62533;
    wire N__62530;
    wire N__62527;
    wire N__62524;
    wire N__62521;
    wire N__62518;
    wire N__62515;
    wire N__62512;
    wire N__62509;
    wire N__62506;
    wire N__62505;
    wire N__62500;
    wire N__62497;
    wire N__62494;
    wire N__62491;
    wire N__62488;
    wire N__62485;
    wire N__62482;
    wire N__62479;
    wire N__62476;
    wire N__62473;
    wire N__62470;
    wire N__62467;
    wire N__62464;
    wire N__62461;
    wire N__62458;
    wire N__62455;
    wire N__62452;
    wire N__62449;
    wire N__62448;
    wire N__62447;
    wire N__62444;
    wire N__62441;
    wire N__62438;
    wire N__62431;
    wire N__62428;
    wire N__62425;
    wire N__62424;
    wire N__62423;
    wire N__62420;
    wire N__62415;
    wire N__62410;
    wire N__62407;
    wire N__62404;
    wire N__62403;
    wire N__62402;
    wire N__62401;
    wire N__62400;
    wire N__62397;
    wire N__62392;
    wire N__62389;
    wire N__62386;
    wire N__62381;
    wire N__62374;
    wire N__62373;
    wire N__62372;
    wire N__62371;
    wire N__62370;
    wire N__62367;
    wire N__62362;
    wire N__62359;
    wire N__62358;
    wire N__62355;
    wire N__62352;
    wire N__62349;
    wire N__62346;
    wire N__62345;
    wire N__62344;
    wire N__62341;
    wire N__62336;
    wire N__62333;
    wire N__62330;
    wire N__62325;
    wire N__62322;
    wire N__62319;
    wire N__62308;
    wire N__62305;
    wire N__62304;
    wire N__62303;
    wire N__62302;
    wire N__62299;
    wire N__62296;
    wire N__62295;
    wire N__62294;
    wire N__62289;
    wire N__62284;
    wire N__62279;
    wire N__62276;
    wire N__62269;
    wire N__62268;
    wire N__62263;
    wire N__62260;
    wire N__62257;
    wire N__62254;
    wire N__62251;
    wire N__62250;
    wire N__62245;
    wire N__62242;
    wire N__62239;
    wire N__62236;
    wire N__62235;
    wire N__62232;
    wire N__62229;
    wire N__62226;
    wire N__62221;
    wire N__62218;
    wire N__62215;
    wire N__62212;
    wire N__62209;
    wire N__62206;
    wire N__62203;
    wire N__62200;
    wire N__62197;
    wire N__62194;
    wire N__62191;
    wire N__62188;
    wire N__62185;
    wire N__62182;
    wire N__62181;
    wire N__62180;
    wire N__62177;
    wire N__62174;
    wire N__62171;
    wire N__62168;
    wire N__62165;
    wire N__62162;
    wire N__62157;
    wire N__62152;
    wire N__62151;
    wire N__62148;
    wire N__62145;
    wire N__62140;
    wire N__62137;
    wire N__62134;
    wire N__62131;
    wire N__62130;
    wire N__62129;
    wire N__62126;
    wire N__62125;
    wire N__62122;
    wire N__62119;
    wire N__62116;
    wire N__62113;
    wire N__62110;
    wire N__62107;
    wire N__62102;
    wire N__62097;
    wire N__62094;
    wire N__62091;
    wire N__62086;
    wire N__62083;
    wire N__62080;
    wire N__62077;
    wire N__62074;
    wire N__62071;
    wire N__62068;
    wire N__62065;
    wire N__62062;
    wire N__62059;
    wire N__62056;
    wire N__62053;
    wire N__62050;
    wire N__62047;
    wire N__62044;
    wire N__62041;
    wire N__62038;
    wire N__62037;
    wire N__62036;
    wire N__62033;
    wire N__62030;
    wire N__62027;
    wire N__62022;
    wire N__62019;
    wire N__62016;
    wire N__62011;
    wire N__62008;
    wire N__62005;
    wire N__62004;
    wire N__62001;
    wire N__62000;
    wire N__61999;
    wire N__61998;
    wire N__61995;
    wire N__61992;
    wire N__61991;
    wire N__61986;
    wire N__61983;
    wire N__61980;
    wire N__61977;
    wire N__61976;
    wire N__61975;
    wire N__61974;
    wire N__61973;
    wire N__61972;
    wire N__61971;
    wire N__61968;
    wire N__61965;
    wire N__61960;
    wire N__61957;
    wire N__61952;
    wire N__61943;
    wire N__61940;
    wire N__61935;
    wire N__61932;
    wire N__61929;
    wire N__61924;
    wire N__61921;
    wire N__61912;
    wire N__61909;
    wire N__61906;
    wire N__61903;
    wire N__61900;
    wire N__61897;
    wire N__61894;
    wire N__61891;
    wire N__61888;
    wire N__61885;
    wire N__61882;
    wire N__61879;
    wire N__61876;
    wire N__61873;
    wire N__61870;
    wire N__61867;
    wire N__61864;
    wire N__61861;
    wire N__61858;
    wire N__61855;
    wire N__61852;
    wire N__61849;
    wire N__61846;
    wire N__61843;
    wire N__61840;
    wire N__61837;
    wire N__61834;
    wire N__61831;
    wire N__61828;
    wire N__61825;
    wire N__61822;
    wire N__61821;
    wire N__61820;
    wire N__61819;
    wire N__61816;
    wire N__61811;
    wire N__61808;
    wire N__61805;
    wire N__61802;
    wire N__61795;
    wire N__61792;
    wire N__61789;
    wire N__61788;
    wire N__61787;
    wire N__61782;
    wire N__61781;
    wire N__61778;
    wire N__61777;
    wire N__61776;
    wire N__61773;
    wire N__61770;
    wire N__61765;
    wire N__61762;
    wire N__61759;
    wire N__61756;
    wire N__61751;
    wire N__61748;
    wire N__61741;
    wire N__61738;
    wire N__61735;
    wire N__61732;
    wire N__61731;
    wire N__61730;
    wire N__61727;
    wire N__61722;
    wire N__61717;
    wire N__61714;
    wire N__61711;
    wire N__61708;
    wire N__61705;
    wire N__61702;
    wire N__61699;
    wire N__61696;
    wire N__61693;
    wire N__61690;
    wire N__61687;
    wire N__61684;
    wire N__61681;
    wire N__61678;
    wire N__61675;
    wire N__61672;
    wire N__61669;
    wire N__61666;
    wire N__61663;
    wire N__61660;
    wire N__61657;
    wire N__61654;
    wire N__61651;
    wire N__61648;
    wire N__61645;
    wire N__61642;
    wire N__61641;
    wire N__61638;
    wire N__61635;
    wire N__61632;
    wire N__61627;
    wire N__61624;
    wire N__61621;
    wire N__61618;
    wire N__61615;
    wire N__61612;
    wire N__61609;
    wire N__61606;
    wire N__61603;
    wire N__61600;
    wire N__61597;
    wire N__61594;
    wire N__61591;
    wire N__61588;
    wire N__61585;
    wire N__61582;
    wire N__61579;
    wire N__61576;
    wire N__61573;
    wire N__61570;
    wire N__61567;
    wire N__61564;
    wire N__61561;
    wire N__61558;
    wire N__61555;
    wire N__61552;
    wire N__61549;
    wire N__61546;
    wire N__61543;
    wire N__61540;
    wire N__61537;
    wire N__61534;
    wire N__61531;
    wire N__61528;
    wire N__61525;
    wire N__61522;
    wire N__61519;
    wire N__61516;
    wire N__61513;
    wire N__61510;
    wire N__61507;
    wire N__61504;
    wire N__61501;
    wire N__61498;
    wire N__61495;
    wire N__61492;
    wire N__61489;
    wire N__61486;
    wire N__61483;
    wire N__61480;
    wire N__61477;
    wire N__61474;
    wire N__61471;
    wire N__61468;
    wire N__61465;
    wire N__61462;
    wire N__61459;
    wire N__61456;
    wire N__61455;
    wire N__61452;
    wire N__61449;
    wire N__61446;
    wire N__61443;
    wire N__61438;
    wire N__61435;
    wire N__61432;
    wire N__61429;
    wire N__61428;
    wire N__61425;
    wire N__61424;
    wire N__61421;
    wire N__61418;
    wire N__61415;
    wire N__61412;
    wire N__61407;
    wire N__61402;
    wire N__61399;
    wire N__61396;
    wire N__61393;
    wire N__61390;
    wire N__61387;
    wire N__61384;
    wire N__61381;
    wire N__61378;
    wire N__61375;
    wire N__61372;
    wire N__61369;
    wire N__61366;
    wire N__61363;
    wire N__61360;
    wire N__61357;
    wire N__61354;
    wire N__61351;
    wire N__61348;
    wire N__61345;
    wire N__61342;
    wire N__61339;
    wire N__61336;
    wire N__61333;
    wire N__61330;
    wire N__61327;
    wire N__61324;
    wire N__61321;
    wire N__61318;
    wire N__61315;
    wire N__61312;
    wire N__61309;
    wire N__61306;
    wire N__61303;
    wire N__61300;
    wire N__61297;
    wire N__61294;
    wire N__61291;
    wire N__61288;
    wire N__61285;
    wire N__61282;
    wire N__61279;
    wire N__61276;
    wire N__61273;
    wire N__61270;
    wire N__61267;
    wire N__61264;
    wire N__61261;
    wire N__61258;
    wire N__61255;
    wire N__61252;
    wire N__61249;
    wire N__61246;
    wire N__61243;
    wire N__61240;
    wire N__61237;
    wire N__61234;
    wire N__61231;
    wire N__61228;
    wire N__61227;
    wire N__61226;
    wire N__61223;
    wire N__61220;
    wire N__61217;
    wire N__61210;
    wire N__61207;
    wire N__61204;
    wire N__61201;
    wire N__61198;
    wire N__61195;
    wire N__61192;
    wire N__61189;
    wire N__61186;
    wire N__61183;
    wire N__61180;
    wire N__61177;
    wire N__61174;
    wire N__61171;
    wire N__61168;
    wire N__61165;
    wire N__61162;
    wire N__61159;
    wire N__61156;
    wire N__61153;
    wire N__61150;
    wire N__61147;
    wire N__61146;
    wire N__61143;
    wire N__61140;
    wire N__61137;
    wire N__61134;
    wire N__61129;
    wire N__61126;
    wire N__61123;
    wire N__61120;
    wire N__61117;
    wire N__61114;
    wire N__61111;
    wire N__61108;
    wire N__61105;
    wire N__61102;
    wire N__61099;
    wire N__61096;
    wire N__61095;
    wire N__61094;
    wire N__61093;
    wire N__61090;
    wire N__61089;
    wire N__61084;
    wire N__61081;
    wire N__61076;
    wire N__61069;
    wire N__61066;
    wire N__61063;
    wire N__61060;
    wire N__61057;
    wire N__61054;
    wire N__61051;
    wire N__61048;
    wire N__61047;
    wire N__61046;
    wire N__61043;
    wire N__61040;
    wire N__61037;
    wire N__61034;
    wire N__61029;
    wire N__61024;
    wire N__61021;
    wire N__61018;
    wire N__61015;
    wire N__61012;
    wire N__61009;
    wire N__61006;
    wire N__61003;
    wire N__61000;
    wire N__60999;
    wire N__60998;
    wire N__60995;
    wire N__60990;
    wire N__60985;
    wire N__60984;
    wire N__60983;
    wire N__60978;
    wire N__60975;
    wire N__60974;
    wire N__60973;
    wire N__60970;
    wire N__60967;
    wire N__60962;
    wire N__60961;
    wire N__60960;
    wire N__60959;
    wire N__60952;
    wire N__60945;
    wire N__60940;
    wire N__60937;
    wire N__60934;
    wire N__60931;
    wire N__60928;
    wire N__60925;
    wire N__60922;
    wire N__60919;
    wire N__60916;
    wire N__60913;
    wire N__60910;
    wire N__60907;
    wire N__60904;
    wire N__60901;
    wire N__60898;
    wire N__60895;
    wire N__60892;
    wire N__60891;
    wire N__60890;
    wire N__60887;
    wire N__60884;
    wire N__60881;
    wire N__60874;
    wire N__60871;
    wire N__60868;
    wire N__60865;
    wire N__60862;
    wire N__60859;
    wire N__60856;
    wire N__60853;
    wire N__60850;
    wire N__60847;
    wire N__60844;
    wire N__60841;
    wire N__60838;
    wire N__60835;
    wire N__60832;
    wire N__60829;
    wire N__60826;
    wire N__60823;
    wire N__60820;
    wire N__60817;
    wire N__60814;
    wire N__60811;
    wire N__60810;
    wire N__60807;
    wire N__60804;
    wire N__60801;
    wire N__60800;
    wire N__60797;
    wire N__60794;
    wire N__60791;
    wire N__60788;
    wire N__60783;
    wire N__60778;
    wire N__60777;
    wire N__60776;
    wire N__60775;
    wire N__60772;
    wire N__60769;
    wire N__60766;
    wire N__60765;
    wire N__60762;
    wire N__60759;
    wire N__60756;
    wire N__60755;
    wire N__60754;
    wire N__60753;
    wire N__60748;
    wire N__60745;
    wire N__60742;
    wire N__60739;
    wire N__60736;
    wire N__60733;
    wire N__60732;
    wire N__60731;
    wire N__60730;
    wire N__60727;
    wire N__60724;
    wire N__60719;
    wire N__60716;
    wire N__60709;
    wire N__60706;
    wire N__60705;
    wire N__60702;
    wire N__60699;
    wire N__60696;
    wire N__60693;
    wire N__60688;
    wire N__60683;
    wire N__60670;
    wire N__60667;
    wire N__60664;
    wire N__60661;
    wire N__60658;
    wire N__60655;
    wire N__60652;
    wire N__60651;
    wire N__60650;
    wire N__60649;
    wire N__60644;
    wire N__60641;
    wire N__60638;
    wire N__60635;
    wire N__60632;
    wire N__60627;
    wire N__60624;
    wire N__60621;
    wire N__60616;
    wire N__60613;
    wire N__60610;
    wire N__60607;
    wire N__60604;
    wire N__60601;
    wire N__60598;
    wire N__60595;
    wire N__60592;
    wire N__60589;
    wire N__60586;
    wire N__60583;
    wire N__60580;
    wire N__60577;
    wire N__60574;
    wire N__60571;
    wire N__60568;
    wire N__60565;
    wire N__60562;
    wire N__60559;
    wire N__60556;
    wire N__60553;
    wire N__60550;
    wire N__60547;
    wire N__60544;
    wire N__60541;
    wire N__60538;
    wire N__60535;
    wire N__60534;
    wire N__60531;
    wire N__60530;
    wire N__60529;
    wire N__60528;
    wire N__60525;
    wire N__60522;
    wire N__60519;
    wire N__60516;
    wire N__60515;
    wire N__60512;
    wire N__60509;
    wire N__60506;
    wire N__60505;
    wire N__60504;
    wire N__60501;
    wire N__60498;
    wire N__60497;
    wire N__60496;
    wire N__60493;
    wire N__60488;
    wire N__60485;
    wire N__60480;
    wire N__60477;
    wire N__60474;
    wire N__60467;
    wire N__60460;
    wire N__60451;
    wire N__60450;
    wire N__60449;
    wire N__60448;
    wire N__60445;
    wire N__60442;
    wire N__60439;
    wire N__60436;
    wire N__60433;
    wire N__60430;
    wire N__60427;
    wire N__60424;
    wire N__60419;
    wire N__60418;
    wire N__60417;
    wire N__60416;
    wire N__60415;
    wire N__60414;
    wire N__60409;
    wire N__60406;
    wire N__60397;
    wire N__60394;
    wire N__60385;
    wire N__60382;
    wire N__60379;
    wire N__60376;
    wire N__60375;
    wire N__60372;
    wire N__60369;
    wire N__60364;
    wire N__60361;
    wire N__60358;
    wire N__60355;
    wire N__60354;
    wire N__60351;
    wire N__60348;
    wire N__60345;
    wire N__60342;
    wire N__60337;
    wire N__60334;
    wire N__60333;
    wire N__60332;
    wire N__60329;
    wire N__60328;
    wire N__60327;
    wire N__60324;
    wire N__60323;
    wire N__60322;
    wire N__60321;
    wire N__60320;
    wire N__60319;
    wire N__60316;
    wire N__60315;
    wire N__60314;
    wire N__60311;
    wire N__60308;
    wire N__60303;
    wire N__60302;
    wire N__60299;
    wire N__60298;
    wire N__60295;
    wire N__60288;
    wire N__60285;
    wire N__60282;
    wire N__60279;
    wire N__60272;
    wire N__60269;
    wire N__60264;
    wire N__60261;
    wire N__60258;
    wire N__60255;
    wire N__60248;
    wire N__60235;
    wire N__60232;
    wire N__60229;
    wire N__60226;
    wire N__60223;
    wire N__60220;
    wire N__60217;
    wire N__60214;
    wire N__60211;
    wire N__60208;
    wire N__60205;
    wire N__60202;
    wire N__60199;
    wire N__60196;
    wire N__60193;
    wire N__60190;
    wire N__60187;
    wire N__60184;
    wire N__60181;
    wire N__60178;
    wire N__60175;
    wire N__60172;
    wire N__60169;
    wire N__60166;
    wire N__60165;
    wire N__60164;
    wire N__60161;
    wire N__60158;
    wire N__60155;
    wire N__60150;
    wire N__60147;
    wire N__60144;
    wire N__60139;
    wire N__60136;
    wire N__60133;
    wire N__60132;
    wire N__60131;
    wire N__60128;
    wire N__60125;
    wire N__60122;
    wire N__60121;
    wire N__60118;
    wire N__60113;
    wire N__60110;
    wire N__60103;
    wire N__60100;
    wire N__60097;
    wire N__60094;
    wire N__60091;
    wire N__60088;
    wire N__60085;
    wire N__60082;
    wire N__60079;
    wire N__60076;
    wire N__60073;
    wire N__60070;
    wire N__60067;
    wire N__60064;
    wire N__60061;
    wire N__60058;
    wire N__60055;
    wire N__60052;
    wire N__60051;
    wire N__60048;
    wire N__60045;
    wire N__60040;
    wire N__60037;
    wire N__60034;
    wire N__60031;
    wire N__60028;
    wire N__60025;
    wire N__60022;
    wire N__60019;
    wire N__60016;
    wire N__60013;
    wire N__60010;
    wire N__60007;
    wire N__60004;
    wire N__60001;
    wire N__59998;
    wire N__59995;
    wire N__59992;
    wire N__59989;
    wire N__59988;
    wire N__59985;
    wire N__59982;
    wire N__59977;
    wire N__59974;
    wire N__59971;
    wire N__59970;
    wire N__59967;
    wire N__59964;
    wire N__59959;
    wire N__59956;
    wire N__59953;
    wire N__59950;
    wire N__59947;
    wire N__59944;
    wire N__59941;
    wire N__59938;
    wire N__59935;
    wire N__59932;
    wire N__59929;
    wire N__59926;
    wire N__59923;
    wire N__59920;
    wire N__59917;
    wire N__59914;
    wire N__59911;
    wire N__59908;
    wire N__59905;
    wire N__59902;
    wire N__59899;
    wire N__59896;
    wire N__59893;
    wire N__59890;
    wire N__59887;
    wire N__59884;
    wire N__59881;
    wire N__59878;
    wire N__59875;
    wire N__59872;
    wire N__59869;
    wire N__59866;
    wire N__59863;
    wire N__59862;
    wire N__59859;
    wire N__59856;
    wire N__59853;
    wire N__59850;
    wire N__59847;
    wire N__59844;
    wire N__59839;
    wire N__59836;
    wire N__59833;
    wire N__59830;
    wire N__59827;
    wire N__59824;
    wire N__59821;
    wire N__59818;
    wire N__59815;
    wire N__59812;
    wire N__59809;
    wire N__59806;
    wire N__59803;
    wire N__59800;
    wire N__59797;
    wire N__59794;
    wire N__59791;
    wire N__59788;
    wire N__59785;
    wire N__59782;
    wire N__59779;
    wire N__59776;
    wire N__59773;
    wire N__59770;
    wire N__59767;
    wire N__59764;
    wire N__59761;
    wire N__59758;
    wire N__59755;
    wire N__59752;
    wire N__59749;
    wire N__59746;
    wire N__59743;
    wire N__59740;
    wire N__59737;
    wire N__59734;
    wire N__59731;
    wire N__59728;
    wire N__59725;
    wire N__59722;
    wire N__59719;
    wire N__59716;
    wire N__59713;
    wire N__59710;
    wire N__59707;
    wire N__59704;
    wire N__59701;
    wire N__59698;
    wire N__59695;
    wire N__59692;
    wire N__59689;
    wire N__59686;
    wire N__59683;
    wire N__59680;
    wire N__59677;
    wire N__59674;
    wire N__59671;
    wire N__59668;
    wire N__59665;
    wire N__59662;
    wire N__59659;
    wire N__59656;
    wire N__59653;
    wire N__59650;
    wire N__59647;
    wire N__59644;
    wire N__59641;
    wire N__59638;
    wire N__59635;
    wire N__59632;
    wire N__59629;
    wire N__59626;
    wire N__59623;
    wire N__59620;
    wire N__59617;
    wire N__59614;
    wire N__59611;
    wire N__59608;
    wire N__59605;
    wire N__59602;
    wire N__59599;
    wire N__59596;
    wire N__59593;
    wire N__59590;
    wire N__59587;
    wire N__59584;
    wire N__59581;
    wire N__59578;
    wire N__59575;
    wire N__59574;
    wire N__59573;
    wire N__59572;
    wire N__59569;
    wire N__59566;
    wire N__59563;
    wire N__59560;
    wire N__59555;
    wire N__59552;
    wire N__59549;
    wire N__59542;
    wire N__59539;
    wire N__59536;
    wire N__59533;
    wire N__59530;
    wire N__59527;
    wire N__59524;
    wire N__59521;
    wire N__59518;
    wire N__59515;
    wire N__59512;
    wire N__59509;
    wire N__59506;
    wire N__59503;
    wire N__59500;
    wire N__59497;
    wire N__59494;
    wire N__59491;
    wire N__59488;
    wire N__59485;
    wire N__59482;
    wire N__59479;
    wire N__59476;
    wire N__59473;
    wire N__59470;
    wire N__59467;
    wire N__59464;
    wire N__59461;
    wire N__59458;
    wire N__59455;
    wire N__59452;
    wire N__59449;
    wire N__59446;
    wire N__59443;
    wire N__59440;
    wire N__59437;
    wire N__59434;
    wire N__59431;
    wire N__59428;
    wire N__59425;
    wire N__59422;
    wire N__59419;
    wire N__59416;
    wire N__59413;
    wire N__59410;
    wire N__59407;
    wire N__59404;
    wire N__59401;
    wire N__59398;
    wire N__59395;
    wire N__59392;
    wire N__59389;
    wire N__59386;
    wire N__59383;
    wire N__59380;
    wire N__59377;
    wire N__59374;
    wire N__59371;
    wire N__59368;
    wire N__59365;
    wire N__59362;
    wire N__59359;
    wire N__59356;
    wire N__59353;
    wire N__59350;
    wire N__59347;
    wire N__59344;
    wire N__59341;
    wire N__59338;
    wire N__59335;
    wire N__59332;
    wire N__59329;
    wire N__59326;
    wire N__59323;
    wire N__59320;
    wire N__59317;
    wire N__59314;
    wire N__59311;
    wire N__59308;
    wire N__59307;
    wire N__59304;
    wire N__59301;
    wire N__59296;
    wire N__59293;
    wire N__59290;
    wire N__59289;
    wire N__59288;
    wire N__59285;
    wire N__59284;
    wire N__59283;
    wire N__59282;
    wire N__59281;
    wire N__59280;
    wire N__59275;
    wire N__59272;
    wire N__59263;
    wire N__59260;
    wire N__59251;
    wire N__59250;
    wire N__59247;
    wire N__59246;
    wire N__59243;
    wire N__59242;
    wire N__59239;
    wire N__59236;
    wire N__59235;
    wire N__59234;
    wire N__59231;
    wire N__59228;
    wire N__59225;
    wire N__59218;
    wire N__59215;
    wire N__59206;
    wire N__59205;
    wire N__59204;
    wire N__59201;
    wire N__59198;
    wire N__59195;
    wire N__59194;
    wire N__59189;
    wire N__59186;
    wire N__59183;
    wire N__59180;
    wire N__59175;
    wire N__59170;
    wire N__59167;
    wire N__59164;
    wire N__59161;
    wire N__59158;
    wire N__59155;
    wire N__59152;
    wire N__59151;
    wire N__59148;
    wire N__59145;
    wire N__59140;
    wire N__59137;
    wire N__59134;
    wire N__59131;
    wire N__59128;
    wire N__59125;
    wire N__59122;
    wire N__59119;
    wire N__59116;
    wire N__59113;
    wire N__59110;
    wire N__59107;
    wire N__59104;
    wire N__59101;
    wire N__59098;
    wire N__59095;
    wire N__59092;
    wire N__59089;
    wire N__59086;
    wire N__59083;
    wire N__59080;
    wire N__59077;
    wire N__59074;
    wire N__59071;
    wire N__59068;
    wire N__59065;
    wire N__59062;
    wire N__59059;
    wire N__59056;
    wire N__59053;
    wire N__59050;
    wire N__59047;
    wire N__59044;
    wire N__59041;
    wire N__59038;
    wire N__59035;
    wire N__59032;
    wire N__59029;
    wire N__59026;
    wire N__59023;
    wire N__59020;
    wire N__59017;
    wire N__59014;
    wire N__59011;
    wire N__59008;
    wire N__59005;
    wire N__59002;
    wire N__58999;
    wire N__58996;
    wire N__58993;
    wire N__58990;
    wire N__58987;
    wire N__58984;
    wire N__58981;
    wire N__58978;
    wire N__58975;
    wire N__58972;
    wire N__58969;
    wire N__58966;
    wire N__58963;
    wire N__58960;
    wire N__58957;
    wire N__58954;
    wire N__58951;
    wire N__58948;
    wire N__58945;
    wire N__58942;
    wire N__58939;
    wire N__58936;
    wire N__58933;
    wire N__58930;
    wire N__58927;
    wire N__58924;
    wire N__58921;
    wire N__58920;
    wire N__58919;
    wire N__58918;
    wire N__58917;
    wire N__58916;
    wire N__58913;
    wire N__58904;
    wire N__58903;
    wire N__58900;
    wire N__58895;
    wire N__58892;
    wire N__58885;
    wire N__58882;
    wire N__58879;
    wire N__58876;
    wire N__58873;
    wire N__58870;
    wire N__58867;
    wire N__58864;
    wire N__58861;
    wire N__58858;
    wire N__58855;
    wire N__58852;
    wire N__58849;
    wire N__58846;
    wire N__58843;
    wire N__58840;
    wire N__58837;
    wire N__58834;
    wire N__58831;
    wire N__58828;
    wire N__58825;
    wire N__58822;
    wire N__58819;
    wire N__58816;
    wire N__58813;
    wire N__58810;
    wire N__58809;
    wire N__58804;
    wire N__58803;
    wire N__58802;
    wire N__58801;
    wire N__58800;
    wire N__58797;
    wire N__58794;
    wire N__58791;
    wire N__58788;
    wire N__58787;
    wire N__58786;
    wire N__58785;
    wire N__58782;
    wire N__58779;
    wire N__58776;
    wire N__58773;
    wire N__58770;
    wire N__58767;
    wire N__58762;
    wire N__58755;
    wire N__58744;
    wire N__58741;
    wire N__58738;
    wire N__58735;
    wire N__58732;
    wire N__58729;
    wire N__58726;
    wire N__58723;
    wire N__58722;
    wire N__58719;
    wire N__58718;
    wire N__58715;
    wire N__58712;
    wire N__58709;
    wire N__58706;
    wire N__58703;
    wire N__58700;
    wire N__58697;
    wire N__58690;
    wire N__58687;
    wire N__58684;
    wire N__58681;
    wire N__58678;
    wire N__58675;
    wire N__58672;
    wire N__58669;
    wire N__58666;
    wire N__58663;
    wire N__58660;
    wire N__58657;
    wire N__58654;
    wire N__58651;
    wire N__58648;
    wire N__58645;
    wire N__58642;
    wire N__58639;
    wire N__58636;
    wire N__58633;
    wire N__58630;
    wire N__58627;
    wire N__58624;
    wire N__58621;
    wire N__58618;
    wire N__58615;
    wire N__58612;
    wire N__58609;
    wire N__58606;
    wire N__58603;
    wire N__58600;
    wire N__58597;
    wire N__58594;
    wire N__58591;
    wire N__58588;
    wire N__58585;
    wire N__58582;
    wire N__58579;
    wire N__58576;
    wire N__58573;
    wire N__58570;
    wire N__58567;
    wire N__58564;
    wire N__58561;
    wire N__58558;
    wire N__58555;
    wire N__58552;
    wire N__58551;
    wire N__58548;
    wire N__58545;
    wire N__58540;
    wire N__58537;
    wire N__58534;
    wire N__58531;
    wire N__58528;
    wire N__58525;
    wire N__58522;
    wire N__58519;
    wire N__58516;
    wire N__58513;
    wire N__58510;
    wire N__58507;
    wire N__58504;
    wire N__58501;
    wire N__58498;
    wire N__58495;
    wire N__58492;
    wire N__58489;
    wire N__58486;
    wire N__58483;
    wire N__58480;
    wire N__58477;
    wire N__58474;
    wire N__58471;
    wire N__58468;
    wire N__58465;
    wire N__58462;
    wire N__58459;
    wire N__58456;
    wire N__58453;
    wire N__58450;
    wire N__58447;
    wire N__58444;
    wire N__58441;
    wire N__58438;
    wire N__58435;
    wire N__58432;
    wire N__58429;
    wire N__58426;
    wire N__58423;
    wire N__58420;
    wire N__58417;
    wire N__58414;
    wire N__58413;
    wire N__58410;
    wire N__58407;
    wire N__58402;
    wire N__58399;
    wire N__58396;
    wire N__58393;
    wire N__58390;
    wire N__58387;
    wire N__58384;
    wire N__58381;
    wire N__58378;
    wire N__58375;
    wire N__58372;
    wire N__58369;
    wire N__58366;
    wire N__58363;
    wire N__58360;
    wire N__58359;
    wire N__58356;
    wire N__58353;
    wire N__58348;
    wire N__58345;
    wire N__58342;
    wire N__58339;
    wire N__58336;
    wire N__58333;
    wire N__58330;
    wire N__58327;
    wire N__58324;
    wire N__58321;
    wire N__58318;
    wire N__58315;
    wire N__58312;
    wire N__58309;
    wire N__58306;
    wire N__58303;
    wire N__58300;
    wire N__58297;
    wire N__58294;
    wire N__58291;
    wire N__58288;
    wire N__58285;
    wire N__58282;
    wire N__58279;
    wire N__58276;
    wire N__58273;
    wire N__58270;
    wire N__58267;
    wire N__58264;
    wire N__58261;
    wire N__58258;
    wire N__58255;
    wire N__58252;
    wire N__58249;
    wire N__58246;
    wire N__58243;
    wire N__58240;
    wire N__58237;
    wire N__58236;
    wire N__58235;
    wire N__58232;
    wire N__58229;
    wire N__58226;
    wire N__58223;
    wire N__58220;
    wire N__58217;
    wire N__58210;
    wire N__58207;
    wire N__58204;
    wire N__58201;
    wire N__58198;
    wire N__58195;
    wire N__58192;
    wire N__58189;
    wire N__58186;
    wire N__58183;
    wire N__58180;
    wire N__58177;
    wire N__58174;
    wire N__58171;
    wire N__58168;
    wire N__58165;
    wire N__58162;
    wire N__58159;
    wire N__58156;
    wire N__58153;
    wire N__58150;
    wire N__58147;
    wire N__58144;
    wire N__58141;
    wire N__58138;
    wire N__58135;
    wire N__58132;
    wire N__58129;
    wire N__58126;
    wire N__58123;
    wire N__58120;
    wire N__58117;
    wire N__58114;
    wire N__58111;
    wire N__58108;
    wire N__58105;
    wire N__58102;
    wire N__58099;
    wire N__58096;
    wire N__58093;
    wire N__58090;
    wire N__58087;
    wire N__58084;
    wire N__58081;
    wire N__58078;
    wire N__58075;
    wire N__58072;
    wire N__58069;
    wire N__58066;
    wire N__58063;
    wire N__58060;
    wire N__58059;
    wire N__58056;
    wire N__58055;
    wire N__58052;
    wire N__58049;
    wire N__58046;
    wire N__58043;
    wire N__58040;
    wire N__58037;
    wire N__58034;
    wire N__58027;
    wire N__58024;
    wire N__58021;
    wire N__58018;
    wire N__58015;
    wire N__58012;
    wire N__58009;
    wire N__58006;
    wire N__58003;
    wire N__58000;
    wire N__57999;
    wire N__57996;
    wire N__57993;
    wire N__57990;
    wire N__57987;
    wire N__57982;
    wire N__57979;
    wire N__57976;
    wire N__57973;
    wire N__57970;
    wire N__57967;
    wire N__57964;
    wire N__57961;
    wire N__57958;
    wire N__57955;
    wire N__57952;
    wire N__57949;
    wire N__57946;
    wire N__57943;
    wire N__57940;
    wire N__57937;
    wire N__57934;
    wire N__57931;
    wire N__57928;
    wire N__57925;
    wire N__57922;
    wire N__57919;
    wire N__57916;
    wire N__57913;
    wire N__57910;
    wire N__57907;
    wire N__57904;
    wire N__57901;
    wire N__57898;
    wire N__57895;
    wire N__57892;
    wire N__57889;
    wire N__57886;
    wire N__57883;
    wire N__57880;
    wire N__57877;
    wire N__57874;
    wire N__57871;
    wire N__57868;
    wire N__57865;
    wire N__57862;
    wire N__57859;
    wire N__57856;
    wire N__57853;
    wire N__57850;
    wire N__57847;
    wire N__57844;
    wire N__57841;
    wire N__57838;
    wire N__57835;
    wire N__57832;
    wire N__57829;
    wire N__57826;
    wire N__57823;
    wire N__57820;
    wire N__57817;
    wire N__57814;
    wire N__57811;
    wire N__57808;
    wire N__57805;
    wire N__57802;
    wire N__57799;
    wire N__57796;
    wire N__57793;
    wire N__57790;
    wire N__57787;
    wire N__57784;
    wire N__57781;
    wire N__57778;
    wire N__57775;
    wire N__57772;
    wire N__57769;
    wire N__57766;
    wire N__57763;
    wire N__57760;
    wire N__57759;
    wire N__57756;
    wire N__57753;
    wire N__57752;
    wire N__57749;
    wire N__57746;
    wire N__57743;
    wire N__57738;
    wire N__57735;
    wire N__57732;
    wire N__57729;
    wire N__57724;
    wire N__57721;
    wire N__57718;
    wire N__57715;
    wire N__57712;
    wire N__57709;
    wire N__57706;
    wire N__57703;
    wire N__57700;
    wire N__57697;
    wire N__57694;
    wire N__57691;
    wire N__57688;
    wire N__57685;
    wire N__57682;
    wire N__57679;
    wire N__57676;
    wire N__57673;
    wire N__57670;
    wire N__57667;
    wire N__57664;
    wire N__57661;
    wire N__57658;
    wire N__57655;
    wire N__57652;
    wire N__57649;
    wire N__57646;
    wire N__57643;
    wire N__57640;
    wire N__57637;
    wire N__57634;
    wire N__57631;
    wire N__57628;
    wire N__57625;
    wire N__57624;
    wire N__57621;
    wire N__57618;
    wire N__57617;
    wire N__57616;
    wire N__57613;
    wire N__57612;
    wire N__57609;
    wire N__57606;
    wire N__57605;
    wire N__57602;
    wire N__57601;
    wire N__57600;
    wire N__57597;
    wire N__57594;
    wire N__57589;
    wire N__57586;
    wire N__57583;
    wire N__57578;
    wire N__57577;
    wire N__57576;
    wire N__57573;
    wire N__57570;
    wire N__57561;
    wire N__57556;
    wire N__57547;
    wire N__57546;
    wire N__57543;
    wire N__57540;
    wire N__57535;
    wire N__57532;
    wire N__57529;
    wire N__57526;
    wire N__57523;
    wire N__57520;
    wire N__57517;
    wire N__57514;
    wire N__57511;
    wire N__57508;
    wire N__57505;
    wire N__57502;
    wire N__57499;
    wire N__57496;
    wire N__57493;
    wire N__57490;
    wire N__57487;
    wire N__57484;
    wire N__57481;
    wire N__57478;
    wire N__57475;
    wire N__57472;
    wire N__57469;
    wire N__57466;
    wire N__57463;
    wire N__57460;
    wire N__57457;
    wire N__57454;
    wire N__57451;
    wire N__57448;
    wire N__57445;
    wire N__57442;
    wire N__57439;
    wire N__57436;
    wire N__57433;
    wire N__57430;
    wire N__57427;
    wire N__57424;
    wire N__57421;
    wire N__57420;
    wire N__57417;
    wire N__57414;
    wire N__57411;
    wire N__57408;
    wire N__57403;
    wire N__57400;
    wire N__57397;
    wire N__57394;
    wire N__57391;
    wire N__57388;
    wire N__57385;
    wire N__57382;
    wire N__57379;
    wire N__57376;
    wire N__57373;
    wire N__57370;
    wire N__57367;
    wire N__57364;
    wire N__57361;
    wire N__57358;
    wire N__57355;
    wire N__57352;
    wire N__57349;
    wire N__57348;
    wire N__57345;
    wire N__57342;
    wire N__57341;
    wire N__57340;
    wire N__57335;
    wire N__57332;
    wire N__57329;
    wire N__57326;
    wire N__57321;
    wire N__57316;
    wire N__57313;
    wire N__57310;
    wire N__57307;
    wire N__57304;
    wire N__57301;
    wire N__57298;
    wire N__57295;
    wire N__57292;
    wire N__57289;
    wire N__57286;
    wire N__57283;
    wire N__57280;
    wire N__57277;
    wire N__57274;
    wire N__57271;
    wire N__57270;
    wire N__57267;
    wire N__57264;
    wire N__57261;
    wire N__57258;
    wire N__57253;
    wire N__57250;
    wire N__57247;
    wire N__57246;
    wire N__57245;
    wire N__57242;
    wire N__57239;
    wire N__57236;
    wire N__57235;
    wire N__57234;
    wire N__57227;
    wire N__57224;
    wire N__57221;
    wire N__57220;
    wire N__57219;
    wire N__57218;
    wire N__57213;
    wire N__57210;
    wire N__57207;
    wire N__57202;
    wire N__57199;
    wire N__57194;
    wire N__57191;
    wire N__57188;
    wire N__57185;
    wire N__57182;
    wire N__57179;
    wire N__57176;
    wire N__57169;
    wire N__57166;
    wire N__57165;
    wire N__57162;
    wire N__57159;
    wire N__57154;
    wire N__57153;
    wire N__57152;
    wire N__57151;
    wire N__57148;
    wire N__57145;
    wire N__57140;
    wire N__57133;
    wire N__57130;
    wire N__57127;
    wire N__57124;
    wire N__57121;
    wire N__57118;
    wire N__57115;
    wire N__57112;
    wire N__57109;
    wire N__57106;
    wire N__57103;
    wire N__57100;
    wire N__57097;
    wire N__57094;
    wire N__57091;
    wire N__57088;
    wire N__57085;
    wire N__57082;
    wire N__57079;
    wire N__57076;
    wire N__57073;
    wire N__57070;
    wire N__57067;
    wire N__57064;
    wire N__57061;
    wire N__57058;
    wire N__57055;
    wire N__57052;
    wire N__57049;
    wire N__57046;
    wire N__57043;
    wire N__57040;
    wire N__57037;
    wire N__57034;
    wire N__57031;
    wire N__57028;
    wire N__57027;
    wire N__57026;
    wire N__57025;
    wire N__57024;
    wire N__57023;
    wire N__57020;
    wire N__57019;
    wire N__57010;
    wire N__57007;
    wire N__57004;
    wire N__57001;
    wire N__56998;
    wire N__56989;
    wire N__56986;
    wire N__56983;
    wire N__56982;
    wire N__56981;
    wire N__56980;
    wire N__56977;
    wire N__56974;
    wire N__56969;
    wire N__56968;
    wire N__56961;
    wire N__56958;
    wire N__56955;
    wire N__56950;
    wire N__56947;
    wire N__56944;
    wire N__56941;
    wire N__56938;
    wire N__56935;
    wire N__56932;
    wire N__56929;
    wire N__56926;
    wire N__56925;
    wire N__56922;
    wire N__56921;
    wire N__56918;
    wire N__56915;
    wire N__56912;
    wire N__56909;
    wire N__56906;
    wire N__56903;
    wire N__56898;
    wire N__56895;
    wire N__56890;
    wire N__56887;
    wire N__56884;
    wire N__56881;
    wire N__56878;
    wire N__56875;
    wire N__56872;
    wire N__56869;
    wire N__56866;
    wire N__56863;
    wire N__56860;
    wire N__56857;
    wire N__56854;
    wire N__56851;
    wire N__56848;
    wire N__56845;
    wire N__56842;
    wire N__56839;
    wire N__56836;
    wire N__56833;
    wire N__56830;
    wire N__56827;
    wire N__56824;
    wire N__56821;
    wire N__56818;
    wire N__56815;
    wire N__56812;
    wire N__56809;
    wire N__56806;
    wire N__56803;
    wire N__56800;
    wire N__56797;
    wire N__56794;
    wire N__56791;
    wire N__56788;
    wire N__56785;
    wire N__56782;
    wire N__56779;
    wire N__56776;
    wire N__56773;
    wire N__56770;
    wire N__56767;
    wire N__56764;
    wire N__56761;
    wire N__56758;
    wire N__56755;
    wire N__56752;
    wire N__56749;
    wire N__56746;
    wire N__56743;
    wire N__56740;
    wire N__56737;
    wire N__56734;
    wire N__56731;
    wire N__56728;
    wire N__56725;
    wire N__56724;
    wire N__56721;
    wire N__56718;
    wire N__56713;
    wire N__56710;
    wire N__56707;
    wire N__56704;
    wire N__56701;
    wire N__56698;
    wire N__56695;
    wire N__56692;
    wire N__56691;
    wire N__56688;
    wire N__56687;
    wire N__56684;
    wire N__56683;
    wire N__56680;
    wire N__56677;
    wire N__56674;
    wire N__56671;
    wire N__56668;
    wire N__56665;
    wire N__56660;
    wire N__56657;
    wire N__56652;
    wire N__56647;
    wire N__56644;
    wire N__56641;
    wire N__56638;
    wire N__56635;
    wire N__56634;
    wire N__56633;
    wire N__56630;
    wire N__56625;
    wire N__56622;
    wire N__56619;
    wire N__56616;
    wire N__56613;
    wire N__56608;
    wire N__56605;
    wire N__56602;
    wire N__56599;
    wire N__56596;
    wire N__56593;
    wire N__56590;
    wire N__56587;
    wire N__56584;
    wire N__56581;
    wire N__56578;
    wire N__56575;
    wire N__56572;
    wire N__56569;
    wire N__56566;
    wire N__56563;
    wire N__56560;
    wire N__56557;
    wire N__56554;
    wire N__56551;
    wire N__56548;
    wire N__56545;
    wire N__56542;
    wire N__56539;
    wire N__56536;
    wire N__56533;
    wire N__56530;
    wire N__56527;
    wire N__56524;
    wire N__56521;
    wire N__56518;
    wire N__56515;
    wire N__56512;
    wire N__56509;
    wire N__56506;
    wire N__56503;
    wire N__56500;
    wire N__56497;
    wire N__56494;
    wire N__56491;
    wire N__56488;
    wire N__56485;
    wire N__56482;
    wire N__56479;
    wire N__56476;
    wire N__56473;
    wire N__56470;
    wire N__56467;
    wire N__56464;
    wire N__56461;
    wire N__56458;
    wire N__56455;
    wire N__56452;
    wire N__56449;
    wire N__56446;
    wire N__56443;
    wire N__56440;
    wire N__56437;
    wire N__56434;
    wire N__56431;
    wire N__56428;
    wire N__56425;
    wire N__56422;
    wire N__56419;
    wire N__56416;
    wire N__56413;
    wire N__56410;
    wire N__56407;
    wire N__56404;
    wire N__56401;
    wire N__56398;
    wire N__56395;
    wire N__56392;
    wire N__56389;
    wire N__56386;
    wire N__56383;
    wire N__56380;
    wire N__56377;
    wire N__56374;
    wire N__56373;
    wire N__56370;
    wire N__56367;
    wire N__56364;
    wire N__56361;
    wire N__56358;
    wire N__56355;
    wire N__56352;
    wire N__56349;
    wire N__56344;
    wire N__56341;
    wire N__56338;
    wire N__56335;
    wire N__56332;
    wire N__56329;
    wire N__56326;
    wire N__56323;
    wire N__56320;
    wire N__56317;
    wire N__56314;
    wire N__56311;
    wire N__56308;
    wire N__56305;
    wire N__56302;
    wire N__56299;
    wire N__56296;
    wire N__56293;
    wire N__56290;
    wire N__56287;
    wire N__56284;
    wire N__56281;
    wire N__56280;
    wire N__56279;
    wire N__56276;
    wire N__56273;
    wire N__56270;
    wire N__56267;
    wire N__56264;
    wire N__56261;
    wire N__56258;
    wire N__56253;
    wire N__56248;
    wire N__56245;
    wire N__56242;
    wire N__56239;
    wire N__56238;
    wire N__56233;
    wire N__56230;
    wire N__56227;
    wire N__56224;
    wire N__56221;
    wire N__56218;
    wire N__56215;
    wire N__56212;
    wire N__56209;
    wire N__56206;
    wire N__56205;
    wire N__56202;
    wire N__56199;
    wire N__56198;
    wire N__56195;
    wire N__56192;
    wire N__56189;
    wire N__56186;
    wire N__56183;
    wire N__56180;
    wire N__56175;
    wire N__56172;
    wire N__56167;
    wire N__56164;
    wire N__56161;
    wire N__56158;
    wire N__56157;
    wire N__56154;
    wire N__56153;
    wire N__56150;
    wire N__56147;
    wire N__56144;
    wire N__56141;
    wire N__56140;
    wire N__56135;
    wire N__56132;
    wire N__56129;
    wire N__56122;
    wire N__56119;
    wire N__56116;
    wire N__56115;
    wire N__56112;
    wire N__56111;
    wire N__56108;
    wire N__56105;
    wire N__56102;
    wire N__56095;
    wire N__56092;
    wire N__56089;
    wire N__56088;
    wire N__56085;
    wire N__56082;
    wire N__56079;
    wire N__56074;
    wire N__56071;
    wire N__56068;
    wire N__56065;
    wire N__56062;
    wire N__56059;
    wire N__56056;
    wire N__56053;
    wire N__56050;
    wire N__56047;
    wire N__56044;
    wire N__56041;
    wire N__56038;
    wire N__56035;
    wire N__56032;
    wire N__56029;
    wire N__56026;
    wire N__56023;
    wire N__56020;
    wire N__56017;
    wire N__56014;
    wire N__56011;
    wire N__56008;
    wire N__56005;
    wire N__56002;
    wire N__55999;
    wire N__55996;
    wire N__55993;
    wire N__55990;
    wire N__55987;
    wire N__55984;
    wire N__55981;
    wire N__55978;
    wire N__55977;
    wire N__55974;
    wire N__55971;
    wire N__55966;
    wire N__55963;
    wire N__55960;
    wire N__55957;
    wire N__55954;
    wire N__55951;
    wire N__55948;
    wire N__55945;
    wire N__55942;
    wire N__55939;
    wire N__55936;
    wire N__55933;
    wire N__55930;
    wire N__55927;
    wire N__55924;
    wire N__55921;
    wire N__55918;
    wire N__55915;
    wire N__55912;
    wire N__55909;
    wire N__55906;
    wire N__55903;
    wire N__55900;
    wire N__55897;
    wire N__55894;
    wire N__55891;
    wire N__55888;
    wire N__55885;
    wire N__55882;
    wire N__55879;
    wire N__55876;
    wire N__55873;
    wire N__55870;
    wire N__55867;
    wire N__55864;
    wire N__55861;
    wire N__55858;
    wire N__55855;
    wire N__55852;
    wire N__55849;
    wire N__55846;
    wire N__55843;
    wire N__55840;
    wire N__55837;
    wire N__55836;
    wire N__55833;
    wire N__55832;
    wire N__55829;
    wire N__55826;
    wire N__55823;
    wire N__55816;
    wire N__55813;
    wire N__55810;
    wire N__55807;
    wire N__55804;
    wire N__55801;
    wire N__55798;
    wire N__55795;
    wire N__55792;
    wire N__55789;
    wire N__55786;
    wire N__55783;
    wire N__55780;
    wire N__55777;
    wire N__55774;
    wire N__55771;
    wire N__55768;
    wire N__55765;
    wire N__55762;
    wire N__55759;
    wire N__55756;
    wire N__55753;
    wire N__55750;
    wire N__55747;
    wire N__55744;
    wire N__55741;
    wire N__55738;
    wire N__55735;
    wire N__55732;
    wire N__55731;
    wire N__55730;
    wire N__55725;
    wire N__55724;
    wire N__55721;
    wire N__55720;
    wire N__55719;
    wire N__55716;
    wire N__55711;
    wire N__55710;
    wire N__55709;
    wire N__55704;
    wire N__55701;
    wire N__55698;
    wire N__55695;
    wire N__55692;
    wire N__55689;
    wire N__55686;
    wire N__55683;
    wire N__55680;
    wire N__55669;
    wire N__55666;
    wire N__55663;
    wire N__55660;
    wire N__55657;
    wire N__55654;
    wire N__55651;
    wire N__55648;
    wire N__55645;
    wire N__55642;
    wire N__55641;
    wire N__55640;
    wire N__55637;
    wire N__55634;
    wire N__55631;
    wire N__55626;
    wire N__55623;
    wire N__55618;
    wire N__55615;
    wire N__55614;
    wire N__55611;
    wire N__55608;
    wire N__55603;
    wire N__55600;
    wire N__55597;
    wire N__55594;
    wire N__55591;
    wire N__55588;
    wire N__55585;
    wire N__55582;
    wire N__55579;
    wire N__55576;
    wire N__55573;
    wire N__55570;
    wire N__55567;
    wire N__55564;
    wire N__55561;
    wire N__55558;
    wire N__55555;
    wire N__55552;
    wire N__55549;
    wire N__55546;
    wire N__55543;
    wire N__55540;
    wire N__55537;
    wire N__55534;
    wire N__55531;
    wire N__55528;
    wire N__55525;
    wire N__55522;
    wire N__55519;
    wire N__55516;
    wire N__55513;
    wire N__55510;
    wire N__55507;
    wire N__55504;
    wire N__55501;
    wire N__55498;
    wire N__55495;
    wire N__55492;
    wire N__55489;
    wire N__55486;
    wire N__55483;
    wire N__55480;
    wire N__55477;
    wire N__55474;
    wire N__55471;
    wire N__55468;
    wire N__55465;
    wire N__55462;
    wire N__55459;
    wire N__55456;
    wire N__55453;
    wire N__55450;
    wire N__55447;
    wire N__55444;
    wire N__55441;
    wire N__55438;
    wire N__55435;
    wire N__55432;
    wire N__55429;
    wire N__55426;
    wire N__55423;
    wire N__55420;
    wire N__55417;
    wire N__55414;
    wire N__55411;
    wire N__55408;
    wire N__55405;
    wire N__55402;
    wire N__55399;
    wire N__55396;
    wire N__55393;
    wire N__55390;
    wire N__55387;
    wire N__55384;
    wire N__55381;
    wire N__55378;
    wire N__55377;
    wire N__55376;
    wire N__55375;
    wire N__55366;
    wire N__55363;
    wire N__55360;
    wire N__55357;
    wire N__55354;
    wire N__55351;
    wire N__55348;
    wire N__55345;
    wire N__55342;
    wire N__55339;
    wire N__55336;
    wire N__55333;
    wire N__55330;
    wire N__55327;
    wire N__55324;
    wire N__55321;
    wire N__55318;
    wire N__55315;
    wire N__55312;
    wire N__55309;
    wire N__55306;
    wire N__55303;
    wire N__55300;
    wire N__55297;
    wire N__55294;
    wire N__55291;
    wire N__55288;
    wire N__55285;
    wire N__55282;
    wire N__55279;
    wire N__55276;
    wire N__55273;
    wire N__55270;
    wire N__55267;
    wire N__55264;
    wire N__55261;
    wire N__55258;
    wire N__55255;
    wire N__55252;
    wire N__55249;
    wire N__55246;
    wire N__55243;
    wire N__55240;
    wire N__55237;
    wire N__55234;
    wire N__55231;
    wire N__55228;
    wire N__55225;
    wire N__55222;
    wire N__55219;
    wire N__55216;
    wire N__55213;
    wire N__55210;
    wire N__55207;
    wire N__55204;
    wire N__55201;
    wire N__55198;
    wire N__55195;
    wire N__55192;
    wire N__55189;
    wire N__55186;
    wire N__55183;
    wire N__55180;
    wire N__55177;
    wire N__55174;
    wire N__55171;
    wire N__55168;
    wire N__55165;
    wire N__55162;
    wire N__55159;
    wire N__55156;
    wire N__55153;
    wire N__55150;
    wire N__55147;
    wire N__55144;
    wire N__55141;
    wire N__55138;
    wire N__55135;
    wire N__55132;
    wire N__55129;
    wire N__55126;
    wire N__55123;
    wire N__55120;
    wire N__55117;
    wire N__55114;
    wire N__55111;
    wire N__55108;
    wire N__55105;
    wire N__55102;
    wire N__55099;
    wire N__55096;
    wire N__55093;
    wire N__55090;
    wire N__55087;
    wire N__55084;
    wire N__55081;
    wire N__55078;
    wire N__55075;
    wire N__55072;
    wire N__55069;
    wire N__55066;
    wire N__55063;
    wire N__55060;
    wire N__55057;
    wire N__55054;
    wire N__55051;
    wire N__55048;
    wire N__55045;
    wire N__55042;
    wire N__55039;
    wire N__55036;
    wire N__55033;
    wire N__55030;
    wire N__55027;
    wire N__55024;
    wire N__55021;
    wire N__55018;
    wire N__55015;
    wire N__55012;
    wire N__55009;
    wire N__55006;
    wire N__55005;
    wire N__55002;
    wire N__54999;
    wire N__54994;
    wire N__54991;
    wire N__54988;
    wire N__54985;
    wire N__54982;
    wire N__54979;
    wire N__54976;
    wire N__54973;
    wire N__54970;
    wire N__54967;
    wire N__54964;
    wire N__54961;
    wire N__54958;
    wire N__54955;
    wire N__54952;
    wire N__54949;
    wire N__54946;
    wire N__54943;
    wire N__54940;
    wire N__54937;
    wire N__54934;
    wire N__54931;
    wire N__54928;
    wire N__54925;
    wire N__54922;
    wire N__54919;
    wire N__54916;
    wire N__54913;
    wire N__54910;
    wire N__54907;
    wire N__54904;
    wire N__54901;
    wire N__54898;
    wire N__54895;
    wire N__54892;
    wire N__54889;
    wire N__54886;
    wire N__54883;
    wire N__54880;
    wire N__54877;
    wire N__54874;
    wire N__54871;
    wire N__54868;
    wire N__54865;
    wire N__54862;
    wire N__54859;
    wire N__54856;
    wire N__54853;
    wire N__54850;
    wire N__54847;
    wire N__54844;
    wire N__54841;
    wire N__54838;
    wire N__54835;
    wire N__54832;
    wire N__54829;
    wire N__54826;
    wire N__54823;
    wire N__54820;
    wire N__54817;
    wire N__54814;
    wire N__54811;
    wire N__54808;
    wire N__54805;
    wire N__54802;
    wire N__54799;
    wire N__54796;
    wire N__54793;
    wire N__54790;
    wire N__54787;
    wire N__54784;
    wire N__54781;
    wire N__54778;
    wire N__54775;
    wire N__54772;
    wire N__54769;
    wire N__54766;
    wire N__54763;
    wire N__54760;
    wire N__54757;
    wire N__54754;
    wire N__54751;
    wire N__54748;
    wire N__54745;
    wire N__54742;
    wire N__54739;
    wire N__54736;
    wire N__54733;
    wire N__54730;
    wire N__54727;
    wire N__54724;
    wire N__54721;
    wire N__54718;
    wire N__54715;
    wire N__54712;
    wire N__54709;
    wire N__54706;
    wire N__54703;
    wire N__54700;
    wire N__54697;
    wire N__54694;
    wire N__54691;
    wire N__54688;
    wire N__54685;
    wire N__54682;
    wire N__54679;
    wire N__54676;
    wire N__54673;
    wire N__54670;
    wire N__54669;
    wire N__54666;
    wire N__54663;
    wire N__54658;
    wire N__54657;
    wire N__54654;
    wire N__54651;
    wire N__54650;
    wire N__54647;
    wire N__54644;
    wire N__54641;
    wire N__54638;
    wire N__54635;
    wire N__54632;
    wire N__54625;
    wire N__54622;
    wire N__54619;
    wire N__54616;
    wire N__54613;
    wire N__54610;
    wire N__54607;
    wire N__54604;
    wire N__54601;
    wire N__54598;
    wire N__54595;
    wire N__54592;
    wire N__54589;
    wire N__54586;
    wire N__54583;
    wire N__54580;
    wire N__54577;
    wire N__54576;
    wire N__54573;
    wire N__54570;
    wire N__54569;
    wire N__54566;
    wire N__54563;
    wire N__54560;
    wire N__54557;
    wire N__54554;
    wire N__54551;
    wire N__54544;
    wire N__54541;
    wire N__54538;
    wire N__54535;
    wire N__54532;
    wire N__54529;
    wire N__54526;
    wire N__54523;
    wire N__54520;
    wire N__54517;
    wire N__54514;
    wire N__54511;
    wire N__54508;
    wire N__54505;
    wire N__54502;
    wire N__54499;
    wire N__54496;
    wire N__54493;
    wire N__54490;
    wire N__54487;
    wire N__54484;
    wire N__54481;
    wire N__54478;
    wire N__54475;
    wire N__54474;
    wire N__54473;
    wire N__54472;
    wire N__54469;
    wire N__54468;
    wire N__54461;
    wire N__54460;
    wire N__54457;
    wire N__54454;
    wire N__54451;
    wire N__54448;
    wire N__54445;
    wire N__54440;
    wire N__54433;
    wire N__54430;
    wire N__54427;
    wire N__54424;
    wire N__54421;
    wire N__54418;
    wire N__54415;
    wire N__54412;
    wire N__54409;
    wire N__54406;
    wire N__54403;
    wire N__54400;
    wire N__54397;
    wire N__54394;
    wire N__54391;
    wire N__54388;
    wire N__54385;
    wire N__54382;
    wire N__54379;
    wire N__54376;
    wire N__54373;
    wire N__54370;
    wire N__54369;
    wire N__54366;
    wire N__54365;
    wire N__54362;
    wire N__54361;
    wire N__54356;
    wire N__54355;
    wire N__54354;
    wire N__54351;
    wire N__54348;
    wire N__54345;
    wire N__54342;
    wire N__54341;
    wire N__54340;
    wire N__54337;
    wire N__54334;
    wire N__54327;
    wire N__54324;
    wire N__54321;
    wire N__54310;
    wire N__54309;
    wire N__54308;
    wire N__54307;
    wire N__54306;
    wire N__54301;
    wire N__54300;
    wire N__54299;
    wire N__54298;
    wire N__54297;
    wire N__54296;
    wire N__54293;
    wire N__54290;
    wire N__54287;
    wire N__54284;
    wire N__54281;
    wire N__54278;
    wire N__54275;
    wire N__54272;
    wire N__54269;
    wire N__54266;
    wire N__54263;
    wire N__54258;
    wire N__54255;
    wire N__54252;
    wire N__54235;
    wire N__54234;
    wire N__54233;
    wire N__54232;
    wire N__54231;
    wire N__54230;
    wire N__54229;
    wire N__54228;
    wire N__54225;
    wire N__54222;
    wire N__54219;
    wire N__54216;
    wire N__54213;
    wire N__54206;
    wire N__54205;
    wire N__54200;
    wire N__54195;
    wire N__54190;
    wire N__54187;
    wire N__54186;
    wire N__54181;
    wire N__54180;
    wire N__54179;
    wire N__54176;
    wire N__54173;
    wire N__54170;
    wire N__54167;
    wire N__54162;
    wire N__54151;
    wire N__54148;
    wire N__54145;
    wire N__54142;
    wire N__54139;
    wire N__54136;
    wire N__54133;
    wire N__54130;
    wire N__54127;
    wire N__54124;
    wire N__54121;
    wire N__54118;
    wire N__54115;
    wire N__54112;
    wire N__54109;
    wire N__54106;
    wire N__54103;
    wire N__54100;
    wire N__54097;
    wire N__54094;
    wire N__54091;
    wire N__54088;
    wire N__54085;
    wire N__54082;
    wire N__54081;
    wire N__54078;
    wire N__54075;
    wire N__54072;
    wire N__54071;
    wire N__54068;
    wire N__54065;
    wire N__54062;
    wire N__54059;
    wire N__54054;
    wire N__54049;
    wire N__54046;
    wire N__54043;
    wire N__54040;
    wire N__54037;
    wire N__54034;
    wire N__54031;
    wire N__54028;
    wire N__54025;
    wire N__54022;
    wire N__54019;
    wire N__54016;
    wire N__54013;
    wire N__54010;
    wire N__54007;
    wire N__54004;
    wire N__54001;
    wire N__53998;
    wire N__53995;
    wire N__53994;
    wire N__53991;
    wire N__53988;
    wire N__53987;
    wire N__53986;
    wire N__53983;
    wire N__53980;
    wire N__53977;
    wire N__53974;
    wire N__53971;
    wire N__53968;
    wire N__53965;
    wire N__53962;
    wire N__53953;
    wire N__53950;
    wire N__53947;
    wire N__53944;
    wire N__53941;
    wire N__53938;
    wire N__53935;
    wire N__53934;
    wire N__53933;
    wire N__53930;
    wire N__53925;
    wire N__53920;
    wire N__53919;
    wire N__53916;
    wire N__53913;
    wire N__53908;
    wire N__53905;
    wire N__53902;
    wire N__53899;
    wire N__53896;
    wire N__53893;
    wire N__53890;
    wire N__53887;
    wire N__53884;
    wire N__53881;
    wire N__53878;
    wire N__53875;
    wire N__53872;
    wire N__53869;
    wire N__53866;
    wire N__53863;
    wire N__53860;
    wire N__53857;
    wire N__53854;
    wire N__53851;
    wire N__53848;
    wire N__53845;
    wire N__53842;
    wire N__53839;
    wire N__53836;
    wire N__53833;
    wire N__53830;
    wire N__53827;
    wire N__53826;
    wire N__53823;
    wire N__53822;
    wire N__53819;
    wire N__53816;
    wire N__53813;
    wire N__53806;
    wire N__53805;
    wire N__53804;
    wire N__53803;
    wire N__53802;
    wire N__53797;
    wire N__53794;
    wire N__53789;
    wire N__53786;
    wire N__53781;
    wire N__53778;
    wire N__53775;
    wire N__53770;
    wire N__53767;
    wire N__53766;
    wire N__53763;
    wire N__53762;
    wire N__53761;
    wire N__53760;
    wire N__53757;
    wire N__53756;
    wire N__53753;
    wire N__53750;
    wire N__53747;
    wire N__53740;
    wire N__53737;
    wire N__53728;
    wire N__53727;
    wire N__53726;
    wire N__53725;
    wire N__53724;
    wire N__53723;
    wire N__53722;
    wire N__53717;
    wire N__53714;
    wire N__53709;
    wire N__53704;
    wire N__53703;
    wire N__53702;
    wire N__53701;
    wire N__53696;
    wire N__53693;
    wire N__53690;
    wire N__53685;
    wire N__53682;
    wire N__53677;
    wire N__53676;
    wire N__53671;
    wire N__53668;
    wire N__53665;
    wire N__53662;
    wire N__53659;
    wire N__53656;
    wire N__53647;
    wire N__53644;
    wire N__53643;
    wire N__53640;
    wire N__53639;
    wire N__53636;
    wire N__53633;
    wire N__53630;
    wire N__53627;
    wire N__53624;
    wire N__53619;
    wire N__53616;
    wire N__53613;
    wire N__53608;
    wire N__53605;
    wire N__53602;
    wire N__53599;
    wire N__53596;
    wire N__53593;
    wire N__53590;
    wire N__53587;
    wire N__53584;
    wire N__53581;
    wire N__53580;
    wire N__53579;
    wire N__53576;
    wire N__53573;
    wire N__53570;
    wire N__53563;
    wire N__53560;
    wire N__53557;
    wire N__53554;
    wire N__53551;
    wire N__53548;
    wire N__53545;
    wire N__53542;
    wire N__53539;
    wire N__53536;
    wire N__53533;
    wire N__53530;
    wire N__53527;
    wire N__53524;
    wire N__53521;
    wire N__53518;
    wire N__53515;
    wire N__53512;
    wire N__53509;
    wire N__53506;
    wire N__53503;
    wire N__53500;
    wire N__53497;
    wire N__53494;
    wire N__53491;
    wire N__53488;
    wire N__53485;
    wire N__53482;
    wire N__53479;
    wire N__53476;
    wire N__53473;
    wire N__53470;
    wire N__53467;
    wire N__53464;
    wire N__53461;
    wire N__53458;
    wire N__53455;
    wire N__53452;
    wire N__53449;
    wire N__53446;
    wire N__53443;
    wire N__53440;
    wire N__53437;
    wire N__53434;
    wire N__53433;
    wire N__53430;
    wire N__53427;
    wire N__53426;
    wire N__53423;
    wire N__53420;
    wire N__53419;
    wire N__53416;
    wire N__53413;
    wire N__53410;
    wire N__53407;
    wire N__53404;
    wire N__53395;
    wire N__53392;
    wire N__53389;
    wire N__53388;
    wire N__53383;
    wire N__53380;
    wire N__53377;
    wire N__53374;
    wire N__53371;
    wire N__53368;
    wire N__53365;
    wire N__53362;
    wire N__53359;
    wire N__53356;
    wire N__53353;
    wire N__53350;
    wire N__53347;
    wire N__53344;
    wire N__53341;
    wire N__53338;
    wire N__53337;
    wire N__53334;
    wire N__53333;
    wire N__53330;
    wire N__53327;
    wire N__53324;
    wire N__53321;
    wire N__53316;
    wire N__53311;
    wire N__53308;
    wire N__53305;
    wire N__53302;
    wire N__53299;
    wire N__53296;
    wire N__53293;
    wire N__53290;
    wire N__53287;
    wire N__53284;
    wire N__53281;
    wire N__53278;
    wire N__53275;
    wire N__53272;
    wire N__53269;
    wire N__53266;
    wire N__53263;
    wire N__53260;
    wire N__53257;
    wire N__53254;
    wire N__53251;
    wire N__53248;
    wire N__53245;
    wire N__53242;
    wire N__53239;
    wire N__53236;
    wire N__53233;
    wire N__53230;
    wire N__53227;
    wire N__53224;
    wire N__53221;
    wire N__53218;
    wire N__53215;
    wire N__53212;
    wire N__53209;
    wire N__53206;
    wire N__53203;
    wire N__53200;
    wire N__53197;
    wire N__53194;
    wire N__53191;
    wire N__53188;
    wire N__53185;
    wire N__53182;
    wire N__53179;
    wire N__53176;
    wire N__53175;
    wire N__53172;
    wire N__53169;
    wire N__53166;
    wire N__53163;
    wire N__53158;
    wire N__53155;
    wire N__53152;
    wire N__53149;
    wire N__53146;
    wire N__53143;
    wire N__53140;
    wire N__53137;
    wire N__53134;
    wire N__53131;
    wire N__53128;
    wire N__53125;
    wire N__53122;
    wire N__53119;
    wire N__53116;
    wire N__53113;
    wire N__53110;
    wire N__53107;
    wire N__53104;
    wire N__53103;
    wire N__53100;
    wire N__53099;
    wire N__53096;
    wire N__53095;
    wire N__53092;
    wire N__53089;
    wire N__53086;
    wire N__53085;
    wire N__53082;
    wire N__53079;
    wire N__53076;
    wire N__53073;
    wire N__53070;
    wire N__53059;
    wire N__53056;
    wire N__53053;
    wire N__53050;
    wire N__53047;
    wire N__53044;
    wire N__53041;
    wire N__53038;
    wire N__53035;
    wire N__53032;
    wire N__53029;
    wire N__53026;
    wire N__53023;
    wire N__53020;
    wire N__53017;
    wire N__53014;
    wire N__53011;
    wire N__53008;
    wire N__53005;
    wire N__53004;
    wire N__53003;
    wire N__53000;
    wire N__52997;
    wire N__52994;
    wire N__52987;
    wire N__52984;
    wire N__52981;
    wire N__52978;
    wire N__52975;
    wire N__52972;
    wire N__52969;
    wire N__52966;
    wire N__52963;
    wire N__52960;
    wire N__52957;
    wire N__52954;
    wire N__52953;
    wire N__52952;
    wire N__52949;
    wire N__52946;
    wire N__52943;
    wire N__52936;
    wire N__52933;
    wire N__52932;
    wire N__52931;
    wire N__52930;
    wire N__52929;
    wire N__52928;
    wire N__52927;
    wire N__52924;
    wire N__52921;
    wire N__52918;
    wire N__52917;
    wire N__52914;
    wire N__52913;
    wire N__52912;
    wire N__52911;
    wire N__52910;
    wire N__52905;
    wire N__52902;
    wire N__52899;
    wire N__52892;
    wire N__52889;
    wire N__52884;
    wire N__52879;
    wire N__52876;
    wire N__52861;
    wire N__52858;
    wire N__52855;
    wire N__52852;
    wire N__52849;
    wire N__52846;
    wire N__52843;
    wire N__52840;
    wire N__52837;
    wire N__52836;
    wire N__52833;
    wire N__52830;
    wire N__52829;
    wire N__52826;
    wire N__52823;
    wire N__52820;
    wire N__52817;
    wire N__52814;
    wire N__52811;
    wire N__52804;
    wire N__52801;
    wire N__52798;
    wire N__52795;
    wire N__52792;
    wire N__52789;
    wire N__52786;
    wire N__52783;
    wire N__52780;
    wire N__52777;
    wire N__52774;
    wire N__52771;
    wire N__52768;
    wire N__52765;
    wire N__52762;
    wire N__52759;
    wire N__52756;
    wire N__52753;
    wire N__52750;
    wire N__52747;
    wire N__52744;
    wire N__52741;
    wire N__52738;
    wire N__52735;
    wire N__52732;
    wire N__52729;
    wire N__52726;
    wire N__52723;
    wire N__52720;
    wire N__52717;
    wire N__52714;
    wire N__52711;
    wire N__52708;
    wire N__52705;
    wire N__52702;
    wire N__52699;
    wire N__52696;
    wire N__52693;
    wire N__52690;
    wire N__52687;
    wire N__52684;
    wire N__52681;
    wire N__52678;
    wire N__52677;
    wire N__52676;
    wire N__52673;
    wire N__52670;
    wire N__52667;
    wire N__52664;
    wire N__52659;
    wire N__52656;
    wire N__52653;
    wire N__52650;
    wire N__52647;
    wire N__52642;
    wire N__52641;
    wire N__52638;
    wire N__52635;
    wire N__52632;
    wire N__52629;
    wire N__52626;
    wire N__52621;
    wire N__52618;
    wire N__52615;
    wire N__52612;
    wire N__52609;
    wire N__52606;
    wire N__52603;
    wire N__52600;
    wire N__52597;
    wire N__52594;
    wire N__52591;
    wire N__52588;
    wire N__52585;
    wire N__52582;
    wire N__52579;
    wire N__52576;
    wire N__52573;
    wire N__52570;
    wire N__52567;
    wire N__52564;
    wire N__52561;
    wire N__52560;
    wire N__52559;
    wire N__52558;
    wire N__52557;
    wire N__52554;
    wire N__52551;
    wire N__52544;
    wire N__52543;
    wire N__52540;
    wire N__52535;
    wire N__52532;
    wire N__52529;
    wire N__52526;
    wire N__52519;
    wire N__52516;
    wire N__52513;
    wire N__52510;
    wire N__52507;
    wire N__52504;
    wire N__52501;
    wire N__52498;
    wire N__52495;
    wire N__52492;
    wire N__52489;
    wire N__52486;
    wire N__52483;
    wire N__52480;
    wire N__52477;
    wire N__52474;
    wire N__52471;
    wire N__52468;
    wire N__52465;
    wire N__52464;
    wire N__52461;
    wire N__52458;
    wire N__52455;
    wire N__52452;
    wire N__52449;
    wire N__52446;
    wire N__52441;
    wire N__52440;
    wire N__52439;
    wire N__52438;
    wire N__52435;
    wire N__52432;
    wire N__52431;
    wire N__52430;
    wire N__52429;
    wire N__52426;
    wire N__52423;
    wire N__52418;
    wire N__52415;
    wire N__52410;
    wire N__52407;
    wire N__52396;
    wire N__52393;
    wire N__52390;
    wire N__52387;
    wire N__52384;
    wire N__52381;
    wire N__52378;
    wire N__52375;
    wire N__52372;
    wire N__52369;
    wire N__52366;
    wire N__52363;
    wire N__52360;
    wire N__52357;
    wire N__52354;
    wire N__52351;
    wire N__52348;
    wire N__52347;
    wire N__52344;
    wire N__52341;
    wire N__52336;
    wire N__52333;
    wire N__52330;
    wire N__52327;
    wire N__52324;
    wire N__52321;
    wire N__52318;
    wire N__52315;
    wire N__52312;
    wire N__52311;
    wire N__52308;
    wire N__52305;
    wire N__52300;
    wire N__52299;
    wire N__52298;
    wire N__52295;
    wire N__52290;
    wire N__52285;
    wire N__52282;
    wire N__52279;
    wire N__52276;
    wire N__52273;
    wire N__52270;
    wire N__52267;
    wire N__52264;
    wire N__52261;
    wire N__52258;
    wire N__52255;
    wire N__52252;
    wire N__52249;
    wire N__52246;
    wire N__52243;
    wire N__52240;
    wire N__52237;
    wire N__52234;
    wire N__52231;
    wire N__52228;
    wire N__52225;
    wire N__52222;
    wire N__52219;
    wire N__52216;
    wire N__52213;
    wire N__52210;
    wire N__52207;
    wire N__52206;
    wire N__52203;
    wire N__52202;
    wire N__52201;
    wire N__52198;
    wire N__52197;
    wire N__52194;
    wire N__52191;
    wire N__52188;
    wire N__52185;
    wire N__52182;
    wire N__52177;
    wire N__52174;
    wire N__52171;
    wire N__52168;
    wire N__52165;
    wire N__52162;
    wire N__52157;
    wire N__52150;
    wire N__52147;
    wire N__52144;
    wire N__52143;
    wire N__52140;
    wire N__52137;
    wire N__52134;
    wire N__52131;
    wire N__52130;
    wire N__52127;
    wire N__52124;
    wire N__52121;
    wire N__52114;
    wire N__52111;
    wire N__52108;
    wire N__52105;
    wire N__52102;
    wire N__52099;
    wire N__52096;
    wire N__52093;
    wire N__52090;
    wire N__52087;
    wire N__52084;
    wire N__52081;
    wire N__52078;
    wire N__52075;
    wire N__52072;
    wire N__52069;
    wire N__52066;
    wire N__52063;
    wire N__52060;
    wire N__52057;
    wire N__52054;
    wire N__52051;
    wire N__52048;
    wire N__52045;
    wire N__52042;
    wire N__52039;
    wire N__52036;
    wire N__52033;
    wire N__52030;
    wire N__52027;
    wire N__52024;
    wire N__52021;
    wire N__52020;
    wire N__52017;
    wire N__52016;
    wire N__52015;
    wire N__52012;
    wire N__52009;
    wire N__52008;
    wire N__52007;
    wire N__52006;
    wire N__52003;
    wire N__52000;
    wire N__51997;
    wire N__51994;
    wire N__51987;
    wire N__51976;
    wire N__51973;
    wire N__51970;
    wire N__51967;
    wire N__51964;
    wire N__51961;
    wire N__51958;
    wire N__51955;
    wire N__51952;
    wire N__51949;
    wire N__51946;
    wire N__51943;
    wire N__51940;
    wire N__51937;
    wire N__51934;
    wire N__51931;
    wire N__51928;
    wire N__51925;
    wire N__51922;
    wire N__51919;
    wire N__51916;
    wire N__51913;
    wire N__51910;
    wire N__51907;
    wire N__51904;
    wire N__51901;
    wire N__51898;
    wire N__51895;
    wire N__51892;
    wire N__51889;
    wire N__51888;
    wire N__51885;
    wire N__51882;
    wire N__51879;
    wire N__51876;
    wire N__51873;
    wire N__51870;
    wire N__51865;
    wire N__51862;
    wire N__51859;
    wire N__51856;
    wire N__51853;
    wire N__51850;
    wire N__51847;
    wire N__51844;
    wire N__51841;
    wire N__51838;
    wire N__51835;
    wire N__51832;
    wire N__51829;
    wire N__51826;
    wire N__51823;
    wire N__51820;
    wire N__51817;
    wire N__51814;
    wire N__51811;
    wire N__51808;
    wire N__51805;
    wire N__51802;
    wire N__51799;
    wire N__51796;
    wire N__51793;
    wire N__51790;
    wire N__51787;
    wire N__51784;
    wire N__51781;
    wire N__51778;
    wire N__51775;
    wire N__51772;
    wire N__51769;
    wire N__51766;
    wire N__51763;
    wire N__51760;
    wire N__51757;
    wire N__51754;
    wire N__51751;
    wire N__51750;
    wire N__51747;
    wire N__51746;
    wire N__51745;
    wire N__51742;
    wire N__51739;
    wire N__51734;
    wire N__51727;
    wire N__51724;
    wire N__51721;
    wire N__51718;
    wire N__51715;
    wire N__51712;
    wire N__51709;
    wire N__51706;
    wire N__51703;
    wire N__51702;
    wire N__51699;
    wire N__51696;
    wire N__51691;
    wire N__51690;
    wire N__51687;
    wire N__51684;
    wire N__51681;
    wire N__51678;
    wire N__51675;
    wire N__51670;
    wire N__51667;
    wire N__51664;
    wire N__51661;
    wire N__51658;
    wire N__51655;
    wire N__51652;
    wire N__51649;
    wire N__51646;
    wire N__51643;
    wire N__51640;
    wire N__51637;
    wire N__51634;
    wire N__51631;
    wire N__51628;
    wire N__51625;
    wire N__51622;
    wire N__51619;
    wire N__51616;
    wire N__51613;
    wire N__51610;
    wire N__51607;
    wire N__51604;
    wire N__51601;
    wire N__51598;
    wire N__51595;
    wire N__51592;
    wire N__51589;
    wire N__51586;
    wire N__51583;
    wire N__51580;
    wire N__51577;
    wire N__51574;
    wire N__51571;
    wire N__51568;
    wire N__51565;
    wire N__51562;
    wire N__51559;
    wire N__51556;
    wire N__51553;
    wire N__51550;
    wire N__51549;
    wire N__51546;
    wire N__51543;
    wire N__51540;
    wire N__51537;
    wire N__51534;
    wire N__51531;
    wire N__51528;
    wire N__51525;
    wire N__51520;
    wire N__51517;
    wire N__51514;
    wire N__51511;
    wire N__51508;
    wire N__51505;
    wire N__51502;
    wire N__51499;
    wire N__51496;
    wire N__51493;
    wire N__51490;
    wire N__51487;
    wire N__51484;
    wire N__51481;
    wire N__51478;
    wire N__51475;
    wire N__51472;
    wire N__51469;
    wire N__51466;
    wire N__51463;
    wire N__51460;
    wire N__51457;
    wire N__51456;
    wire N__51453;
    wire N__51450;
    wire N__51449;
    wire N__51444;
    wire N__51441;
    wire N__51438;
    wire N__51435;
    wire N__51430;
    wire N__51427;
    wire N__51424;
    wire N__51421;
    wire N__51418;
    wire N__51415;
    wire N__51412;
    wire N__51409;
    wire N__51406;
    wire N__51403;
    wire N__51400;
    wire N__51397;
    wire N__51394;
    wire N__51391;
    wire N__51388;
    wire N__51385;
    wire N__51382;
    wire N__51379;
    wire N__51376;
    wire N__51373;
    wire N__51372;
    wire N__51371;
    wire N__51370;
    wire N__51367;
    wire N__51364;
    wire N__51359;
    wire N__51358;
    wire N__51355;
    wire N__51352;
    wire N__51349;
    wire N__51348;
    wire N__51345;
    wire N__51340;
    wire N__51337;
    wire N__51334;
    wire N__51325;
    wire N__51324;
    wire N__51321;
    wire N__51318;
    wire N__51315;
    wire N__51310;
    wire N__51307;
    wire N__51304;
    wire N__51301;
    wire N__51298;
    wire N__51295;
    wire N__51292;
    wire N__51289;
    wire N__51286;
    wire N__51285;
    wire N__51282;
    wire N__51279;
    wire N__51274;
    wire N__51271;
    wire N__51268;
    wire N__51265;
    wire N__51264;
    wire N__51263;
    wire N__51262;
    wire N__51259;
    wire N__51252;
    wire N__51247;
    wire N__51244;
    wire N__51241;
    wire N__51238;
    wire N__51235;
    wire N__51232;
    wire N__51229;
    wire N__51226;
    wire N__51223;
    wire N__51220;
    wire N__51217;
    wire N__51216;
    wire N__51213;
    wire N__51212;
    wire N__51209;
    wire N__51204;
    wire N__51199;
    wire N__51196;
    wire N__51193;
    wire N__51190;
    wire N__51187;
    wire N__51184;
    wire N__51181;
    wire N__51178;
    wire N__51175;
    wire N__51172;
    wire N__51169;
    wire N__51166;
    wire N__51163;
    wire N__51160;
    wire N__51157;
    wire N__51154;
    wire N__51151;
    wire N__51148;
    wire N__51145;
    wire N__51142;
    wire N__51139;
    wire N__51136;
    wire N__51133;
    wire N__51130;
    wire N__51127;
    wire N__51124;
    wire N__51121;
    wire N__51118;
    wire N__51115;
    wire N__51112;
    wire N__51109;
    wire N__51106;
    wire N__51103;
    wire N__51100;
    wire N__51097;
    wire N__51094;
    wire N__51091;
    wire N__51088;
    wire N__51085;
    wire N__51082;
    wire N__51079;
    wire N__51076;
    wire N__51073;
    wire N__51070;
    wire N__51067;
    wire N__51064;
    wire N__51061;
    wire N__51058;
    wire N__51055;
    wire N__51052;
    wire N__51049;
    wire N__51046;
    wire N__51043;
    wire N__51040;
    wire N__51037;
    wire N__51034;
    wire N__51031;
    wire N__51028;
    wire N__51025;
    wire N__51022;
    wire N__51019;
    wire N__51016;
    wire N__51013;
    wire N__51010;
    wire N__51007;
    wire N__51004;
    wire N__51001;
    wire N__50998;
    wire N__50995;
    wire N__50992;
    wire N__50989;
    wire N__50986;
    wire N__50983;
    wire N__50980;
    wire N__50977;
    wire N__50974;
    wire N__50971;
    wire N__50968;
    wire N__50965;
    wire N__50962;
    wire N__50959;
    wire N__50956;
    wire N__50953;
    wire N__50950;
    wire N__50947;
    wire N__50944;
    wire N__50941;
    wire N__50938;
    wire N__50935;
    wire N__50932;
    wire N__50929;
    wire N__50926;
    wire N__50923;
    wire N__50920;
    wire N__50919;
    wire N__50916;
    wire N__50913;
    wire N__50910;
    wire N__50907;
    wire N__50902;
    wire N__50899;
    wire N__50896;
    wire N__50893;
    wire N__50890;
    wire N__50887;
    wire N__50884;
    wire N__50881;
    wire N__50878;
    wire N__50875;
    wire N__50872;
    wire N__50869;
    wire N__50866;
    wire N__50863;
    wire N__50860;
    wire N__50857;
    wire N__50854;
    wire N__50853;
    wire N__50852;
    wire N__50849;
    wire N__50846;
    wire N__50843;
    wire N__50840;
    wire N__50835;
    wire N__50832;
    wire N__50829;
    wire N__50826;
    wire N__50823;
    wire N__50818;
    wire N__50817;
    wire N__50816;
    wire N__50815;
    wire N__50814;
    wire N__50811;
    wire N__50806;
    wire N__50805;
    wire N__50804;
    wire N__50801;
    wire N__50798;
    wire N__50793;
    wire N__50788;
    wire N__50779;
    wire N__50778;
    wire N__50777;
    wire N__50776;
    wire N__50775;
    wire N__50772;
    wire N__50771;
    wire N__50768;
    wire N__50767;
    wire N__50764;
    wire N__50761;
    wire N__50758;
    wire N__50753;
    wire N__50750;
    wire N__50747;
    wire N__50738;
    wire N__50731;
    wire N__50728;
    wire N__50725;
    wire N__50722;
    wire N__50719;
    wire N__50718;
    wire N__50717;
    wire N__50714;
    wire N__50711;
    wire N__50710;
    wire N__50707;
    wire N__50704;
    wire N__50703;
    wire N__50702;
    wire N__50699;
    wire N__50696;
    wire N__50695;
    wire N__50692;
    wire N__50689;
    wire N__50684;
    wire N__50681;
    wire N__50676;
    wire N__50669;
    wire N__50666;
    wire N__50663;
    wire N__50660;
    wire N__50657;
    wire N__50650;
    wire N__50647;
    wire N__50644;
    wire N__50643;
    wire N__50640;
    wire N__50637;
    wire N__50634;
    wire N__50629;
    wire N__50626;
    wire N__50623;
    wire N__50620;
    wire N__50617;
    wire N__50614;
    wire N__50611;
    wire N__50608;
    wire N__50605;
    wire N__50602;
    wire N__50599;
    wire N__50596;
    wire N__50593;
    wire N__50592;
    wire N__50589;
    wire N__50586;
    wire N__50581;
    wire N__50578;
    wire N__50575;
    wire N__50572;
    wire N__50569;
    wire N__50566;
    wire N__50563;
    wire N__50560;
    wire N__50557;
    wire N__50556;
    wire N__50551;
    wire N__50550;
    wire N__50549;
    wire N__50548;
    wire N__50547;
    wire N__50546;
    wire N__50543;
    wire N__50538;
    wire N__50535;
    wire N__50532;
    wire N__50529;
    wire N__50522;
    wire N__50519;
    wire N__50512;
    wire N__50509;
    wire N__50508;
    wire N__50507;
    wire N__50504;
    wire N__50503;
    wire N__50502;
    wire N__50501;
    wire N__50496;
    wire N__50493;
    wire N__50490;
    wire N__50487;
    wire N__50486;
    wire N__50483;
    wire N__50480;
    wire N__50473;
    wire N__50470;
    wire N__50461;
    wire N__50458;
    wire N__50455;
    wire N__50452;
    wire N__50451;
    wire N__50448;
    wire N__50445;
    wire N__50442;
    wire N__50439;
    wire N__50434;
    wire N__50431;
    wire N__50430;
    wire N__50429;
    wire N__50428;
    wire N__50423;
    wire N__50422;
    wire N__50421;
    wire N__50420;
    wire N__50417;
    wire N__50414;
    wire N__50411;
    wire N__50404;
    wire N__50395;
    wire N__50392;
    wire N__50389;
    wire N__50386;
    wire N__50383;
    wire N__50380;
    wire N__50377;
    wire N__50374;
    wire N__50373;
    wire N__50370;
    wire N__50367;
    wire N__50366;
    wire N__50365;
    wire N__50362;
    wire N__50359;
    wire N__50356;
    wire N__50353;
    wire N__50344;
    wire N__50341;
    wire N__50338;
    wire N__50335;
    wire N__50332;
    wire N__50329;
    wire N__50326;
    wire N__50323;
    wire N__50320;
    wire N__50317;
    wire N__50314;
    wire N__50311;
    wire N__50310;
    wire N__50307;
    wire N__50304;
    wire N__50299;
    wire N__50296;
    wire N__50293;
    wire N__50290;
    wire N__50287;
    wire N__50284;
    wire N__50281;
    wire N__50278;
    wire N__50275;
    wire N__50272;
    wire N__50269;
    wire N__50266;
    wire N__50263;
    wire N__50260;
    wire N__50257;
    wire N__50254;
    wire N__50251;
    wire N__50248;
    wire N__50245;
    wire N__50242;
    wire N__50239;
    wire N__50236;
    wire N__50233;
    wire N__50230;
    wire N__50227;
    wire N__50224;
    wire N__50221;
    wire N__50218;
    wire N__50215;
    wire N__50212;
    wire N__50209;
    wire N__50206;
    wire N__50203;
    wire N__50202;
    wire N__50199;
    wire N__50196;
    wire N__50193;
    wire N__50190;
    wire N__50187;
    wire N__50184;
    wire N__50179;
    wire N__50176;
    wire N__50173;
    wire N__50170;
    wire N__50167;
    wire N__50164;
    wire N__50161;
    wire N__50158;
    wire N__50155;
    wire N__50152;
    wire N__50149;
    wire N__50146;
    wire N__50143;
    wire N__50140;
    wire N__50137;
    wire N__50134;
    wire N__50131;
    wire N__50128;
    wire N__50125;
    wire N__50122;
    wire N__50119;
    wire N__50118;
    wire N__50115;
    wire N__50112;
    wire N__50109;
    wire N__50106;
    wire N__50103;
    wire N__50100;
    wire N__50095;
    wire N__50092;
    wire N__50089;
    wire N__50086;
    wire N__50083;
    wire N__50080;
    wire N__50077;
    wire N__50074;
    wire N__50071;
    wire N__50068;
    wire N__50065;
    wire N__50062;
    wire N__50059;
    wire N__50056;
    wire N__50053;
    wire N__50050;
    wire N__50047;
    wire N__50044;
    wire N__50041;
    wire N__50038;
    wire N__50037;
    wire N__50034;
    wire N__50031;
    wire N__50028;
    wire N__50025;
    wire N__50020;
    wire N__50017;
    wire N__50014;
    wire N__50011;
    wire N__50008;
    wire N__50005;
    wire N__50002;
    wire N__49999;
    wire N__49996;
    wire N__49993;
    wire N__49990;
    wire N__49987;
    wire N__49986;
    wire N__49983;
    wire N__49980;
    wire N__49977;
    wire N__49974;
    wire N__49969;
    wire N__49966;
    wire N__49963;
    wire N__49960;
    wire N__49957;
    wire N__49954;
    wire N__49953;
    wire N__49952;
    wire N__49949;
    wire N__49946;
    wire N__49943;
    wire N__49940;
    wire N__49937;
    wire N__49934;
    wire N__49931;
    wire N__49928;
    wire N__49925;
    wire N__49918;
    wire N__49915;
    wire N__49912;
    wire N__49909;
    wire N__49906;
    wire N__49903;
    wire N__49900;
    wire N__49897;
    wire N__49894;
    wire N__49891;
    wire N__49888;
    wire N__49885;
    wire N__49882;
    wire N__49881;
    wire N__49878;
    wire N__49877;
    wire N__49874;
    wire N__49871;
    wire N__49868;
    wire N__49865;
    wire N__49860;
    wire N__49855;
    wire N__49852;
    wire N__49849;
    wire N__49846;
    wire N__49843;
    wire N__49840;
    wire N__49837;
    wire N__49834;
    wire N__49831;
    wire N__49828;
    wire N__49825;
    wire N__49822;
    wire N__49819;
    wire N__49816;
    wire N__49813;
    wire N__49810;
    wire N__49807;
    wire N__49804;
    wire N__49801;
    wire N__49798;
    wire N__49795;
    wire N__49792;
    wire N__49789;
    wire N__49786;
    wire N__49783;
    wire N__49780;
    wire N__49777;
    wire N__49774;
    wire N__49771;
    wire N__49768;
    wire N__49765;
    wire N__49762;
    wire N__49759;
    wire N__49756;
    wire N__49753;
    wire N__49750;
    wire N__49747;
    wire N__49744;
    wire N__49741;
    wire N__49738;
    wire N__49735;
    wire N__49732;
    wire N__49729;
    wire N__49726;
    wire N__49723;
    wire N__49720;
    wire N__49717;
    wire N__49714;
    wire N__49711;
    wire N__49708;
    wire N__49705;
    wire N__49702;
    wire N__49699;
    wire N__49696;
    wire N__49693;
    wire N__49690;
    wire N__49687;
    wire N__49684;
    wire N__49681;
    wire N__49678;
    wire N__49677;
    wire N__49676;
    wire N__49675;
    wire N__49672;
    wire N__49669;
    wire N__49666;
    wire N__49663;
    wire N__49654;
    wire N__49651;
    wire N__49648;
    wire N__49645;
    wire N__49642;
    wire N__49639;
    wire N__49636;
    wire N__49633;
    wire N__49630;
    wire N__49627;
    wire N__49624;
    wire N__49621;
    wire N__49618;
    wire N__49615;
    wire N__49612;
    wire N__49609;
    wire N__49606;
    wire N__49603;
    wire N__49600;
    wire N__49597;
    wire N__49596;
    wire N__49593;
    wire N__49590;
    wire N__49585;
    wire N__49582;
    wire N__49579;
    wire N__49576;
    wire N__49573;
    wire N__49570;
    wire N__49569;
    wire N__49568;
    wire N__49565;
    wire N__49562;
    wire N__49559;
    wire N__49556;
    wire N__49553;
    wire N__49550;
    wire N__49547;
    wire N__49544;
    wire N__49541;
    wire N__49534;
    wire N__49531;
    wire N__49528;
    wire N__49525;
    wire N__49522;
    wire N__49521;
    wire N__49518;
    wire N__49515;
    wire N__49512;
    wire N__49509;
    wire N__49504;
    wire N__49501;
    wire N__49498;
    wire N__49495;
    wire N__49492;
    wire N__49489;
    wire N__49488;
    wire N__49485;
    wire N__49482;
    wire N__49477;
    wire N__49476;
    wire N__49475;
    wire N__49474;
    wire N__49473;
    wire N__49470;
    wire N__49465;
    wire N__49464;
    wire N__49459;
    wire N__49458;
    wire N__49457;
    wire N__49452;
    wire N__49449;
    wire N__49446;
    wire N__49441;
    wire N__49438;
    wire N__49435;
    wire N__49426;
    wire N__49423;
    wire N__49420;
    wire N__49417;
    wire N__49414;
    wire N__49411;
    wire N__49408;
    wire N__49405;
    wire N__49402;
    wire N__49399;
    wire N__49396;
    wire N__49395;
    wire N__49394;
    wire N__49391;
    wire N__49388;
    wire N__49385;
    wire N__49382;
    wire N__49379;
    wire N__49376;
    wire N__49369;
    wire N__49368;
    wire N__49367;
    wire N__49364;
    wire N__49361;
    wire N__49358;
    wire N__49355;
    wire N__49352;
    wire N__49345;
    wire N__49342;
    wire N__49341;
    wire N__49340;
    wire N__49337;
    wire N__49336;
    wire N__49331;
    wire N__49328;
    wire N__49325;
    wire N__49318;
    wire N__49317;
    wire N__49314;
    wire N__49311;
    wire N__49310;
    wire N__49305;
    wire N__49304;
    wire N__49303;
    wire N__49300;
    wire N__49297;
    wire N__49294;
    wire N__49291;
    wire N__49282;
    wire N__49279;
    wire N__49276;
    wire N__49273;
    wire N__49272;
    wire N__49269;
    wire N__49266;
    wire N__49263;
    wire N__49260;
    wire N__49255;
    wire N__49252;
    wire N__49249;
    wire N__49246;
    wire N__49243;
    wire N__49240;
    wire N__49237;
    wire N__49234;
    wire N__49231;
    wire N__49228;
    wire N__49225;
    wire N__49222;
    wire N__49219;
    wire N__49216;
    wire N__49213;
    wire N__49210;
    wire N__49207;
    wire N__49204;
    wire N__49201;
    wire N__49198;
    wire N__49195;
    wire N__49192;
    wire N__49189;
    wire N__49186;
    wire N__49183;
    wire N__49180;
    wire N__49177;
    wire N__49174;
    wire N__49171;
    wire N__49168;
    wire N__49165;
    wire N__49162;
    wire N__49159;
    wire N__49156;
    wire N__49153;
    wire N__49150;
    wire N__49147;
    wire N__49144;
    wire N__49141;
    wire N__49138;
    wire N__49135;
    wire N__49132;
    wire N__49129;
    wire N__49126;
    wire N__49123;
    wire N__49120;
    wire N__49117;
    wire N__49114;
    wire N__49111;
    wire N__49108;
    wire N__49105;
    wire N__49102;
    wire N__49099;
    wire N__49096;
    wire N__49093;
    wire N__49090;
    wire N__49087;
    wire N__49084;
    wire N__49081;
    wire N__49078;
    wire N__49075;
    wire N__49072;
    wire N__49069;
    wire N__49066;
    wire N__49063;
    wire N__49060;
    wire N__49057;
    wire N__49054;
    wire N__49051;
    wire N__49048;
    wire N__49045;
    wire N__49042;
    wire N__49039;
    wire N__49036;
    wire N__49033;
    wire N__49030;
    wire N__49027;
    wire N__49024;
    wire N__49021;
    wire N__49018;
    wire N__49015;
    wire N__49012;
    wire N__49009;
    wire N__49006;
    wire N__49003;
    wire N__49000;
    wire N__48997;
    wire N__48994;
    wire N__48991;
    wire N__48988;
    wire N__48985;
    wire N__48982;
    wire N__48979;
    wire N__48976;
    wire N__48973;
    wire N__48970;
    wire N__48967;
    wire N__48964;
    wire N__48961;
    wire N__48958;
    wire N__48955;
    wire N__48952;
    wire N__48949;
    wire N__48946;
    wire N__48943;
    wire N__48940;
    wire N__48937;
    wire N__48934;
    wire N__48931;
    wire N__48928;
    wire N__48925;
    wire N__48922;
    wire N__48919;
    wire N__48916;
    wire N__48913;
    wire N__48910;
    wire N__48907;
    wire N__48904;
    wire N__48901;
    wire N__48898;
    wire N__48895;
    wire N__48892;
    wire N__48889;
    wire N__48886;
    wire N__48883;
    wire N__48880;
    wire N__48877;
    wire N__48874;
    wire N__48871;
    wire N__48868;
    wire N__48865;
    wire N__48862;
    wire N__48859;
    wire N__48856;
    wire N__48853;
    wire N__48850;
    wire N__48847;
    wire N__48844;
    wire N__48841;
    wire N__48838;
    wire N__48835;
    wire N__48832;
    wire N__48829;
    wire N__48826;
    wire N__48823;
    wire N__48820;
    wire N__48817;
    wire N__48816;
    wire N__48813;
    wire N__48812;
    wire N__48809;
    wire N__48806;
    wire N__48803;
    wire N__48798;
    wire N__48795;
    wire N__48790;
    wire N__48787;
    wire N__48784;
    wire N__48781;
    wire N__48778;
    wire N__48775;
    wire N__48772;
    wire N__48769;
    wire N__48766;
    wire N__48763;
    wire N__48760;
    wire N__48757;
    wire N__48754;
    wire N__48751;
    wire N__48748;
    wire N__48745;
    wire N__48742;
    wire N__48739;
    wire N__48736;
    wire N__48733;
    wire N__48730;
    wire N__48727;
    wire N__48726;
    wire N__48723;
    wire N__48720;
    wire N__48715;
    wire N__48712;
    wire N__48709;
    wire N__48706;
    wire N__48703;
    wire N__48700;
    wire N__48697;
    wire N__48694;
    wire N__48691;
    wire N__48688;
    wire N__48685;
    wire N__48682;
    wire N__48679;
    wire N__48676;
    wire N__48673;
    wire N__48670;
    wire N__48667;
    wire N__48664;
    wire N__48661;
    wire N__48658;
    wire N__48655;
    wire N__48652;
    wire N__48649;
    wire N__48646;
    wire N__48643;
    wire N__48640;
    wire N__48637;
    wire N__48634;
    wire N__48631;
    wire N__48628;
    wire N__48625;
    wire N__48622;
    wire N__48619;
    wire N__48616;
    wire N__48613;
    wire N__48610;
    wire N__48607;
    wire N__48604;
    wire N__48601;
    wire N__48598;
    wire N__48595;
    wire N__48592;
    wire N__48589;
    wire N__48586;
    wire N__48583;
    wire N__48580;
    wire N__48577;
    wire N__48574;
    wire N__48571;
    wire N__48568;
    wire N__48565;
    wire N__48562;
    wire N__48559;
    wire N__48556;
    wire N__48553;
    wire N__48550;
    wire N__48547;
    wire N__48544;
    wire N__48541;
    wire N__48538;
    wire N__48535;
    wire N__48532;
    wire N__48529;
    wire N__48526;
    wire N__48523;
    wire N__48520;
    wire N__48517;
    wire N__48514;
    wire N__48511;
    wire N__48508;
    wire N__48505;
    wire N__48502;
    wire N__48499;
    wire N__48496;
    wire N__48493;
    wire N__48490;
    wire N__48487;
    wire N__48484;
    wire N__48481;
    wire N__48478;
    wire N__48475;
    wire N__48472;
    wire N__48471;
    wire N__48470;
    wire N__48467;
    wire N__48464;
    wire N__48461;
    wire N__48454;
    wire N__48451;
    wire N__48448;
    wire N__48445;
    wire N__48442;
    wire N__48439;
    wire N__48436;
    wire N__48433;
    wire N__48430;
    wire N__48427;
    wire N__48424;
    wire N__48421;
    wire N__48418;
    wire N__48415;
    wire N__48412;
    wire N__48409;
    wire N__48406;
    wire N__48403;
    wire N__48400;
    wire N__48397;
    wire N__48394;
    wire N__48391;
    wire N__48388;
    wire N__48385;
    wire N__48382;
    wire N__48379;
    wire N__48376;
    wire N__48373;
    wire N__48370;
    wire N__48367;
    wire N__48364;
    wire N__48361;
    wire N__48358;
    wire N__48355;
    wire N__48352;
    wire N__48349;
    wire N__48346;
    wire N__48343;
    wire N__48340;
    wire N__48337;
    wire N__48334;
    wire N__48331;
    wire N__48328;
    wire N__48325;
    wire N__48322;
    wire N__48319;
    wire N__48316;
    wire N__48313;
    wire N__48310;
    wire N__48307;
    wire N__48304;
    wire N__48301;
    wire N__48298;
    wire N__48295;
    wire N__48292;
    wire N__48289;
    wire N__48286;
    wire N__48283;
    wire N__48280;
    wire N__48277;
    wire N__48274;
    wire N__48271;
    wire N__48268;
    wire N__48265;
    wire N__48262;
    wire N__48259;
    wire N__48256;
    wire N__48253;
    wire N__48250;
    wire N__48247;
    wire N__48244;
    wire N__48241;
    wire N__48238;
    wire N__48235;
    wire N__48234;
    wire N__48233;
    wire N__48230;
    wire N__48227;
    wire N__48224;
    wire N__48221;
    wire N__48218;
    wire N__48215;
    wire N__48208;
    wire N__48205;
    wire N__48202;
    wire N__48199;
    wire N__48196;
    wire N__48193;
    wire N__48190;
    wire N__48187;
    wire N__48184;
    wire N__48181;
    wire N__48178;
    wire N__48175;
    wire N__48172;
    wire N__48169;
    wire N__48166;
    wire N__48163;
    wire N__48160;
    wire N__48157;
    wire N__48154;
    wire N__48151;
    wire N__48148;
    wire N__48145;
    wire VCCG0;
    wire GNDG0;
    wire N_4015_i;
    wire shift_srl_3Z0Z_10;
    wire shift_srl_3Z0Z_11;
    wire shift_srl_3Z0Z_12;
    wire shift_srl_3Z0Z_8;
    wire shift_srl_3Z0Z_9;
    wire shift_srl_3Z0Z_5;
    wire shift_srl_3Z0Z_6;
    wire shift_srl_3Z0Z_7;
    wire shift_srl_3Z0Z_13;
    wire shift_srl_3Z0Z_14;
    wire shift_srl_3Z0Z_3;
    wire shift_srl_3Z0Z_4;
    wire rco_c_3;
    wire rco_c_3_cascade_;
    wire shift_srl_3Z0Z_0;
    wire shift_srl_3Z0Z_1;
    wire shift_srl_3Z0Z_2;
    wire clk_en_3;
    wire shift_srl_4Z0Z_0;
    wire shift_srl_4Z0Z_1;
    wire shift_srl_4Z0Z_2;
    wire shift_srl_4Z0Z_3;
    wire shift_srl_4Z0Z_4;
    wire shift_srl_4Z0Z_5;
    wire shift_srl_4Z0Z_6;
    wire shift_srl_6Z0Z_14;
    wire shift_srl_6Z0Z_13;
    wire shift_srl_6Z0Z_12;
    wire shift_srl_6Z0Z_11;
    wire shift_srl_6Z0Z_10;
    wire shift_srl_6Z0Z_9;
    wire shift_srl_5Z0Z_10;
    wire shift_srl_5Z0Z_11;
    wire shift_srl_5Z0Z_12;
    wire shift_srl_5Z0Z_13;
    wire shift_srl_5Z0Z_14;
    wire shift_srl_5Z0Z_9;
    wire shift_srl_5Z0Z_8;
    wire rco_c_5;
    wire rco_c_5_cascade_;
    wire rco_c_4;
    wire rco_c_4_cascade_;
    wire shift_srl_5Z0Z_4;
    wire shift_srl_5Z0Z_5;
    wire shift_srl_5Z0Z_6;
    wire shift_srl_5Z0Z_7;
    wire shift_srl_5Z0Z_3;
    wire shift_srl_5Z0Z_0;
    wire shift_srl_5Z0Z_1;
    wire shift_srl_5Z0Z_2;
    wire clk_en_5;
    wire shift_srl_130Z0Z_8;
    wire shift_srl_130Z0Z_6;
    wire shift_srl_130Z0Z_7;
    wire shift_srl_137Z0Z_0;
    wire shift_srl_137Z0Z_1;
    wire shift_srl_137Z0Z_2;
    wire shift_srl_137Z0Z_3;
    wire shift_srl_137Z0Z_4;
    wire shift_srl_137Z0Z_5;
    wire shift_srl_137Z0Z_6;
    wire shift_srl_22Z0Z_3;
    wire shift_srl_22Z0Z_4;
    wire shift_srl_22Z0Z_5;
    wire shift_srl_22Z0Z_6;
    wire shift_srl_22Z0Z_0;
    wire shift_srl_13Z0Z_2;
    wire shift_srl_13Z0Z_3;
    wire shift_srl_13Z0Z_0;
    wire shift_srl_13Z0Z_1;
    wire shift_srl_13Z0Z_4;
    wire shift_srl_13Z0Z_5;
    wire shift_srl_13Z0Z_6;
    wire shift_srl_12Z0Z_7;
    wire shift_srl_12Z0Z_6;
    wire shift_srl_12Z0Z_0;
    wire shift_srl_12Z0Z_1;
    wire shift_srl_12Z0Z_2;
    wire shift_srl_12Z0Z_3;
    wire shift_srl_12Z0Z_4;
    wire shift_srl_12Z0Z_5;
    wire shift_srl_4Z0Z_10;
    wire shift_srl_4Z0Z_11;
    wire shift_srl_4Z0Z_12;
    wire shift_srl_4Z0Z_13;
    wire shift_srl_4Z0Z_14;
    wire shift_srl_4Z0Z_9;
    wire shift_srl_4Z0Z_7;
    wire shift_srl_4Z0Z_8;
    wire clk_en_4;
    wire shift_srl_6Z0Z_8;
    wire shift_srl_6Z0Z_7;
    wire shift_srl_6Z0Z_0;
    wire shift_srl_6Z0Z_1;
    wire shift_srl_6Z0Z_2;
    wire shift_srl_6Z0Z_3;
    wire shift_srl_6Z0Z_4;
    wire shift_srl_6Z0Z_5;
    wire shift_srl_6Z0Z_6;
    wire clk_en_6;
    wire rco_c_6;
    wire rco_c_6_cascade_;
    wire shift_srl_7Z0Z_0;
    wire shift_srl_7Z0Z_1;
    wire shift_srl_7Z0Z_2;
    wire shift_srl_7Z0Z_3;
    wire shift_srl_7Z0Z_4;
    wire shift_srl_7Z0Z_5;
    wire shift_srl_129Z0Z_8;
    wire shift_srl_130Z0Z_0;
    wire shift_srl_130Z0Z_1;
    wire shift_srl_130Z0Z_2;
    wire shift_srl_130Z0Z_3;
    wire shift_srl_130Z0Z_4;
    wire shift_srl_130Z0Z_5;
    wire shift_srl_129_RNIDM4DZ0Z_15_cascade_;
    wire g0_11_cascade_;
    wire g0_16_0;
    wire g0_17_cascade_;
    wire shift_srl_136Z0Z_10;
    wire shift_srl_136Z0Z_11;
    wire shift_srl_136Z0Z_12;
    wire shift_srl_136Z0Z_13;
    wire shift_srl_136Z0Z_14;
    wire shift_srl_136Z0Z_9;
    wire shift_srl_136Z0Z_8;
    wire shift_srl_136Z0Z_0;
    wire shift_srl_136Z0Z_1;
    wire shift_srl_136Z0Z_2;
    wire shift_srl_136Z0Z_3;
    wire shift_srl_136Z0Z_4;
    wire shift_srl_136Z0Z_5;
    wire shift_srl_136Z0Z_6;
    wire shift_srl_136Z0Z_7;
    wire shift_srl_138Z0Z_1;
    wire shift_srl_138Z0Z_2;
    wire shift_srl_138Z0Z_3;
    wire shift_srl_138Z0Z_4;
    wire shift_srl_138Z0Z_0;
    wire shift_srl_138Z0Z_10;
    wire shift_srl_22Z0Z_1;
    wire shift_srl_22Z0Z_2;
    wire shift_srl_15Z0Z_0;
    wire shift_srl_15Z0Z_1;
    wire shift_srl_15Z0Z_2;
    wire shift_srl_15Z0Z_3;
    wire shift_srl_15Z0Z_4;
    wire shift_srl_15Z0Z_5;
    wire shift_srl_15Z0Z_6;
    wire shift_srl_14Z0Z_10;
    wire shift_srl_14Z0Z_11;
    wire shift_srl_14Z0Z_5;
    wire shift_srl_14Z0Z_6;
    wire shift_srl_14Z0Z_9;
    wire shift_srl_14Z0Z_7;
    wire shift_srl_14Z0Z_8;
    wire shift_srl_13Z0Z_10;
    wire shift_srl_13Z0Z_11;
    wire shift_srl_13Z0Z_12;
    wire shift_srl_13Z0Z_13;
    wire shift_srl_13Z0Z_14;
    wire shift_srl_13Z0Z_9;
    wire shift_srl_13Z0Z_7;
    wire shift_srl_13Z0Z_8;
    wire shift_srl_12Z0Z_14;
    wire shift_srl_12Z0Z_13;
    wire shift_srl_12Z0Z_12;
    wire shift_srl_12Z0Z_11;
    wire shift_srl_12Z0Z_10;
    wire shift_srl_12Z0Z_8;
    wire shift_srl_12Z0Z_9;
    wire clk_en_12;
    wire shift_srl_6Z0Z_15;
    wire shift_srl_5Z0Z_15;
    wire shift_srl_4Z0Z_15;
    wire shift_srl_6_RNI00BHZ0Z_15_cascade_;
    wire shift_srl_7_RNI00TC1Z0Z_15_cascade_;
    wire rco_c_13;
    wire rco_c_13_cascade_;
    wire rco_c_16_cascade_;
    wire rco_c_16;
    wire rco_c_19;
    wire rco_c_12_cascade_;
    wire clk_en_13;
    wire rco_int_0_a2_sx_12;
    wire rco_c_12;
    wire rco_int_0_a2_sx_11;
    wire shift_srl_6_RNI00BHZ0Z_15;
    wire shift_srl_3Z0Z_15;
    wire rco_c_7_cascade_;
    wire shift_srl_21Z0Z_10;
    wire shift_srl_21Z0Z_11;
    wire shift_srl_21Z0Z_12;
    wire shift_srl_21Z0Z_13;
    wire shift_srl_21Z0Z_14;
    wire shift_srl_21Z0Z_9;
    wire shift_srl_21Z0Z_8;
    wire shift_srl_7Z0Z_10;
    wire shift_srl_7Z0Z_11;
    wire shift_srl_7Z0Z_12;
    wire shift_srl_7Z0Z_13;
    wire shift_srl_7Z0Z_14;
    wire shift_srl_7Z0Z_9;
    wire shift_srl_7Z0Z_8;
    wire shift_srl_7Z0Z_6;
    wire shift_srl_7Z0Z_7;
    wire clk_en_7;
    wire shift_srl_18Z0Z_10;
    wire shift_srl_18Z0Z_11;
    wire shift_srl_18Z0Z_12;
    wire shift_srl_18Z0Z_13;
    wire shift_srl_18Z0Z_14;
    wire shift_srl_18Z0Z_9;
    wire shift_srl_18Z0Z_8;
    wire shift_srl_129Z0Z_0;
    wire shift_srl_129Z0Z_1;
    wire shift_srl_129Z0Z_2;
    wire shift_srl_129Z0Z_3;
    wire shift_srl_129Z0Z_4;
    wire shift_srl_129Z0Z_5;
    wire shift_srl_129Z0Z_6;
    wire shift_srl_129Z0Z_7;
    wire g0_8_1;
    wire shift_srl_130Z0Z_14;
    wire shift_srl_130Z0Z_13;
    wire shift_srl_130Z0Z_12;
    wire shift_srl_130Z0Z_11;
    wire shift_srl_130Z0Z_9;
    wire shift_srl_130Z0Z_10;
    wire clk_en_130;
    wire shift_srl_137Z0Z_10;
    wire shift_srl_137Z0Z_11;
    wire shift_srl_137Z0Z_12;
    wire shift_srl_137Z0Z_13;
    wire shift_srl_137Z0Z_14;
    wire shift_srl_137Z0Z_9;
    wire shift_srl_137Z0Z_7;
    wire shift_srl_137Z0Z_8;
    wire clk_en_137;
    wire g0_4_0_cascade_;
    wire g0_13_cascade_;
    wire g0_15_0;
    wire g0_16_1_cascade_;
    wire clk_en_136;
    wire g0_8_0_cascade_;
    wire shift_srl_138Z0Z_9;
    wire shift_srl_138Z0Z_11;
    wire shift_srl_138Z0Z_12;
    wire shift_srl_138Z0Z_13;
    wire shift_srl_138Z0Z_14;
    wire shift_srl_138Z0Z_5;
    wire shift_srl_138Z0Z_6;
    wire shift_srl_138Z0Z_7;
    wire shift_srl_138Z0Z_8;
    wire clk_en_138;
    wire rco_c_124;
    wire shift_srl_15Z0Z_10;
    wire shift_srl_15Z0Z_11;
    wire shift_srl_15Z0Z_12;
    wire shift_srl_15Z0Z_13;
    wire shift_srl_15Z0Z_14;
    wire shift_srl_15Z0Z_9;
    wire shift_srl_15Z0Z_7;
    wire shift_srl_15Z0Z_8;
    wire clk_en_15;
    wire shift_srl_14Z0Z_0;
    wire shift_srl_14Z0Z_1;
    wire shift_srl_14Z0Z_2;
    wire shift_srl_14Z0Z_3;
    wire shift_srl_14Z0Z_4;
    wire shift_srl_14Z0Z_12;
    wire shift_srl_14Z0Z_13;
    wire shift_srl_14Z0Z_14;
    wire clk_en_14;
    wire shift_srl_11Z0Z_14;
    wire shift_srl_11Z0Z_13;
    wire shift_srl_11Z0Z_12;
    wire shift_srl_11Z0Z_11;
    wire shift_srl_11Z0Z_10;
    wire shift_srl_11Z0Z_9;
    wire shift_srl_16Z0Z_10;
    wire shift_srl_16Z0Z_11;
    wire shift_srl_16Z0Z_12;
    wire shift_srl_16Z0Z_13;
    wire shift_srl_16Z0Z_14;
    wire rco_c_11;
    wire rco_c_14_cascade_;
    wire rco_c_17_cascade_;
    wire rco_c_20;
    wire rco_c_17;
    wire rco_c_14;
    wire rco_int_0_a2_21_m6_0_a2_s_6_cascade_;
    wire rco_c_18;
    wire rco_c_18_cascade_;
    wire shift_srl_15Z0Z_15;
    wire rco_int_0_a2_sx_15_cascade_;
    wire shift_srl_14Z0Z_15;
    wire rco_c_15;
    wire rco_c_15_cascade_;
    wire shift_srl_16Z0Z_15;
    wire shift_srl_12Z0Z_15;
    wire shift_srl_13Z0Z_15;
    wire rco_int_0_a2_sx_13;
    wire shift_srl_18Z0Z_15;
    wire shift_srl_18Z0Z_0;
    wire shift_srl_21Z0Z_15;
    wire shift_srl_21Z0Z_0;
    wire shift_srl_21Z0Z_1;
    wire shift_srl_21Z0Z_2;
    wire shift_srl_21Z0Z_3;
    wire shift_srl_21Z0Z_4;
    wire shift_srl_21Z0Z_5;
    wire shift_srl_21Z0Z_6;
    wire shift_srl_21Z0Z_7;
    wire clk_en_21;
    wire shift_srl_18Z0Z_1;
    wire shift_srl_18Z0Z_2;
    wire shift_srl_18Z0Z_3;
    wire shift_srl_18Z0Z_4;
    wire shift_srl_18Z0Z_5;
    wire shift_srl_18Z0Z_6;
    wire shift_srl_18Z0Z_7;
    wire clk_en_18;
    wire shift_srl_133Z0Z_13;
    wire shift_srl_133Z0Z_12;
    wire shift_srl_133Z0Z_11;
    wire shift_srl_131Z0Z_2;
    wire shift_srl_131Z0Z_3;
    wire shift_srl_131Z0Z_4;
    wire shift_srl_131Z0Z_5;
    wire shift_srl_131Z0Z_6;
    wire shift_srl_131Z0Z_7;
    wire rco_obuf_RNO_0Z0Z_131_cascade_;
    wire rco_c_131;
    wire rco_c_130;
    wire g0_2_0;
    wire rco_c_123_cascade_;
    wire clk_en_133;
    wire g0_2_1;
    wire g0_11_0;
    wire g0_6;
    wire shift_srl_129Z0Z_13;
    wire shift_srl_129Z0Z_12;
    wire shift_srl_129Z0Z_11;
    wire shift_srl_129Z0Z_9;
    wire shift_srl_129Z0Z_10;
    wire shift_srl_134Z0Z_10;
    wire shift_srl_134Z0Z_11;
    wire shift_srl_134Z0Z_12;
    wire shift_srl_134Z0Z_13;
    wire shift_srl_134Z0Z_14;
    wire shift_srl_134Z0Z_9;
    wire shift_srl_134Z0Z_8;
    wire rco_c_137;
    wire shift_srl_138Z0Z_15;
    wire shift_srl_133_fast_RNIML0IZ0Z_15_cascade_;
    wire rco_c_136;
    wire shift_srl_133Z0Z_14;
    wire shift_srl_133_fastZ0Z_15;
    wire shift_srl_137Z0Z_15;
    wire g0_7;
    wire rco_c_134;
    wire shift_srl_133_fast_RNIML0IZ0Z_15;
    wire rco_c_135;
    wire rco_c_125;
    wire shift_srl_22Z0Z_10;
    wire shift_srl_22Z0Z_11;
    wire shift_srl_22Z0Z_12;
    wire shift_srl_22Z0Z_13;
    wire shift_srl_22Z0Z_7;
    wire shift_srl_22Z0Z_14;
    wire shift_srl_22Z0Z_8;
    wire shift_srl_22Z0Z_9;
    wire shift_srl_11Z0Z_15;
    wire shift_srl_11Z0Z_0;
    wire shift_srl_11Z0Z_1;
    wire shift_srl_11Z0Z_2;
    wire shift_srl_11Z0Z_3;
    wire shift_srl_11Z0Z_4;
    wire shift_srl_11Z0Z_7;
    wire shift_srl_11Z0Z_8;
    wire shift_srl_11Z0Z_5;
    wire shift_srl_11Z0Z_6;
    wire clk_en_11;
    wire shift_srl_16Z0Z_0;
    wire shift_srl_16Z0Z_1;
    wire shift_srl_16Z0Z_7;
    wire shift_srl_16Z0Z_2;
    wire shift_srl_16Z0Z_3;
    wire shift_srl_16Z0Z_4;
    wire shift_srl_16Z0Z_5;
    wire shift_srl_16Z0Z_6;
    wire shift_srl_16Z0Z_8;
    wire shift_srl_16Z0Z_9;
    wire clk_en_16;
    wire shift_srl_20Z0Z_1;
    wire shift_srl_20Z0Z_2;
    wire shift_srl_20Z0Z_0;
    wire shift_srl_20Z0Z_3;
    wire shift_srl_20Z0Z_4;
    wire shift_srl_20Z0Z_5;
    wire shift_srl_20Z0Z_6;
    wire shift_srl_20Z0Z_10;
    wire shift_srl_20Z0Z_9;
    wire shift_srl_20Z0Z_13;
    wire shift_srl_20Z0Z_14;
    wire shift_srl_20Z0Z_15;
    wire shift_srl_20Z0Z_11;
    wire shift_srl_20Z0Z_12;
    wire shift_srl_20Z0Z_7;
    wire shift_srl_20Z0Z_8;
    wire clk_en_20;
    wire rco_c_7;
    wire shift_srl_8Z0Z_0;
    wire shift_srl_8Z0Z_1;
    wire shift_srl_8Z0Z_2;
    wire shift_srl_8Z0Z_3;
    wire shift_srl_8Z0Z_6;
    wire shift_srl_8Z0Z_4;
    wire shift_srl_8Z0Z_5;
    wire shift_srl_8Z0Z_7;
    wire shift_srl_133Z0Z_4;
    wire shift_srl_133Z0Z_5;
    wire shift_srl_133Z0Z_6;
    wire shift_srl_133Z0Z_7;
    wire shift_srl_133Z0Z_10;
    wire shift_srl_133Z0Z_8;
    wire shift_srl_133Z0Z_9;
    wire shift_srl_132Z0Z_10;
    wire shift_srl_132Z0Z_11;
    wire shift_srl_132Z0Z_12;
    wire shift_srl_132Z0Z_13;
    wire shift_srl_132Z0Z_9;
    wire shift_srl_132Z0Z_8;
    wire shift_srl_131Z0Z_10;
    wire shift_srl_131Z0Z_11;
    wire shift_srl_131Z0Z_12;
    wire shift_srl_131Z0Z_13;
    wire shift_srl_131Z0Z_14;
    wire shift_srl_131Z0Z_8;
    wire shift_srl_131Z0Z_9;
    wire shift_srl_131Z0Z_0;
    wire shift_srl_131Z0Z_1;
    wire clk_en_131;
    wire shift_srl_134Z0Z_15;
    wire g0_2_cascade_;
    wire g0_13_0_cascade_;
    wire g0_10_1_cascade_;
    wire g0_14_0;
    wire g0_12_1;
    wire shift_srl_135Z0Z_11;
    wire shift_srl_135Z0Z_12;
    wire shift_srl_135Z0Z_13;
    wire shift_srl_135Z0Z_14;
    wire shift_srl_135Z0Z_9;
    wire shift_srl_135Z0Z_10;
    wire shift_srl_2Z0Z_10;
    wire shift_srl_2Z0Z_11;
    wire shift_srl_2Z0Z_12;
    wire shift_srl_2Z0Z_8;
    wire shift_srl_2Z0Z_9;
    wire shift_srl_2Z0Z_2;
    wire shift_srl_2Z0Z_0;
    wire shift_srl_2Z0Z_1;
    wire shift_srl_2Z0Z_13;
    wire shift_srl_2Z0Z_3;
    wire shift_srl_2Z0Z_4;
    wire shift_srl_2Z0Z_5;
    wire shift_srl_2Z0Z_6;
    wire shift_srl_2Z0Z_7;
    wire N_701;
    wire shift_srl_10_RNIQHCJ1Z0Z_15_cascade_;
    wire rco_c_21;
    wire rco_c_21_cascade_;
    wire shift_srl_2Z0Z_14;
    wire shift_srl_7_RNI00TC1Z0Z_15;
    wire N_453_cascade_;
    wire rco_c_10;
    wire shift_srl_2Z0Z_15;
    wire N_453_i;
    wire shift_srl_23Z0Z_10;
    wire shift_srl_23Z0Z_11;
    wire shift_srl_23Z0Z_12;
    wire shift_srl_23Z0Z_13;
    wire shift_srl_23Z0Z_9;
    wire shift_srl_23Z0Z_8;
    wire shift_srl_23Z0Z_7;
    wire shift_srl_19Z0Z_10;
    wire shift_srl_19Z0Z_6;
    wire shift_srl_19Z0Z_14;
    wire shift_srl_19Z0Z_9;
    wire shift_srl_19Z0Z_7;
    wire shift_srl_19Z0Z_8;
    wire shift_srl_19Z0Z_15;
    wire shift_srl_19Z0Z_0;
    wire shift_srl_19Z0Z_1;
    wire shift_srl_19Z0Z_2;
    wire shift_srl_19Z0Z_3;
    wire shift_srl_19Z0Z_4;
    wire shift_srl_19Z0Z_5;
    wire shift_srl_19Z0Z_11;
    wire shift_srl_19Z0Z_12;
    wire shift_srl_19Z0Z_13;
    wire clk_en_19;
    wire shift_srl_17Z0Z_15;
    wire shift_srl_17Z0Z_0;
    wire shift_srl_17Z0Z_1;
    wire shift_srl_17Z0Z_2;
    wire shift_srl_17Z0Z_3;
    wire shift_srl_17Z0Z_4;
    wire shift_srl_17Z0Z_5;
    wire shift_srl_17Z0Z_6;
    wire shift_srl_17Z0Z_10;
    wire shift_srl_17Z0Z_11;
    wire shift_srl_17Z0Z_12;
    wire shift_srl_17Z0Z_13;
    wire shift_srl_17Z0Z_14;
    wire shift_srl_17Z0Z_9;
    wire shift_srl_17Z0Z_7;
    wire shift_srl_17Z0Z_8;
    wire clk_en_17;
    wire rco_c_8;
    wire shift_srl_9Z0Z_0;
    wire shift_srl_9Z0Z_1;
    wire shift_srl_9Z0Z_2;
    wire shift_srl_9Z0Z_3;
    wire shift_srl_9Z0Z_4;
    wire shift_srl_9Z0Z_5;
    wire shift_srl_8Z0Z_10;
    wire shift_srl_8Z0Z_11;
    wire shift_srl_8Z0Z_12;
    wire shift_srl_8Z0Z_13;
    wire shift_srl_8Z0Z_14;
    wire shift_srl_8Z0Z_8;
    wire shift_srl_8Z0Z_9;
    wire clk_en_8;
    wire shift_srl_128Z0Z_7;
    wire shift_srl_132Z0Z_0;
    wire shift_srl_132Z0Z_1;
    wire shift_srl_132Z0Z_2;
    wire shift_srl_132Z0Z_3;
    wire shift_srl_132Z0Z_4;
    wire shift_srl_132Z0Z_5;
    wire shift_srl_132Z0Z_6;
    wire shift_srl_132Z0Z_7;
    wire shift_srl_132Z0Z_14;
    wire g0_43_1_cascade_;
    wire clk_en_132;
    wire shift_srl_130Z0Z_15;
    wire shift_srl_132_RNI731TZ0Z_15_cascade_;
    wire rco_int_0_a3_0_a2_0_132_cascade_;
    wire shift_srl_134Z0Z_0;
    wire shift_srl_134Z0Z_1;
    wire shift_srl_134Z0Z_2;
    wire shift_srl_134Z0Z_3;
    wire shift_srl_134Z0Z_4;
    wire shift_srl_134Z0Z_5;
    wire shift_srl_134Z0Z_6;
    wire shift_srl_134Z0Z_7;
    wire clk_en_134;
    wire g0_10_0;
    wire g0_9_2_cascade_;
    wire g0_11_1;
    wire g0_12_0_cascade_;
    wire g0_16_2;
    wire shift_srl_135Z0Z_8;
    wire shift_srl_135Z0Z_15;
    wire shift_srl_135Z0Z_2;
    wire shift_srl_135Z0Z_3;
    wire shift_srl_135Z0Z_4;
    wire shift_srl_135Z0Z_0;
    wire shift_srl_135Z0Z_1;
    wire shift_srl_135Z0Z_5;
    wire shift_srl_135Z0Z_6;
    wire shift_srl_135Z0Z_7;
    wire clk_en_135;
    wire shift_srl_116Z0Z_0;
    wire shift_srl_116Z0Z_1;
    wire shift_srl_116Z0Z_2;
    wire shift_srl_116Z0Z_3;
    wire shift_srl_116Z0Z_4;
    wire shift_srl_116Z0Z_5;
    wire shift_srl_116Z0Z_6;
    wire shift_srl_116Z0Z_7;
    wire rco_c_113;
    wire shift_srl_107Z0Z_0;
    wire rco_c_164;
    wire shift_srl_1Z0Z_7;
    wire shift_srl_1Z0Z_6;
    wire shift_srl_1Z0Z_5;
    wire shift_srl_1Z0Z_4;
    wire N_12_i;
    wire shift_srl_1Z0Z_13;
    wire shift_srl_1Z0Z_12;
    wire shift_srl_1Z0Z_11;
    wire shift_srl_1Z0Z_10;
    wire shift_srl_1Z0Z_8;
    wire shift_srl_1Z0Z_9;
    wire shift_srl_1Z0Z_14;
    wire shift_srl_22Z0Z_15;
    wire shift_srl_23Z0Z_14;
    wire shift_srl_23Z0Z_15;
    wire shift_srl_23Z0Z_0;
    wire shift_srl_23Z0Z_1;
    wire shift_srl_23Z0Z_2;
    wire shift_srl_23Z0Z_3;
    wire shift_srl_23Z0Z_4;
    wire shift_srl_23Z0Z_5;
    wire shift_srl_23Z0Z_6;
    wire N_702;
    wire rco_c_155;
    wire rco_c_154;
    wire rco_c_156;
    wire rco_c_159;
    wire rco_c_160;
    wire rco_c_161;
    wire shift_srl_154Z0Z_0;
    wire shift_srl_154Z0Z_1;
    wire shift_srl_154Z0Z_2;
    wire rco_c_26;
    wire shift_srl_8Z0Z_15;
    wire rco_int_0_a2_0_9;
    wire shift_srl_7Z0Z_15;
    wire N_453;
    wire rco_int_0_a2_0_9_cascade_;
    wire rco_int_0_a2_out_1;
    wire rco_c_9_cascade_;
    wire N_4016_i_cascade_;
    wire rco_c_25;
    wire shift_srl_9Z0Z_15;
    wire shift_srl_9Z0Z_10;
    wire shift_srl_9Z0Z_11;
    wire shift_srl_9Z0Z_12;
    wire shift_srl_9Z0Z_13;
    wire shift_srl_9Z0Z_14;
    wire shift_srl_9Z0Z_9;
    wire shift_srl_9Z0Z_8;
    wire shift_srl_9Z0Z_6;
    wire shift_srl_9Z0Z_7;
    wire clk_en_9;
    wire shift_srl_128Z0Z_0;
    wire shift_srl_128Z0Z_1;
    wire shift_srl_128Z0Z_2;
    wire shift_srl_128Z0Z_3;
    wire shift_srl_128Z0Z_4;
    wire shift_srl_128Z0Z_5;
    wire shift_srl_128Z0Z_6;
    wire shift_srl_129Z0Z_14;
    wire clk_en_129;
    wire shift_srl_132Z0Z_15;
    wire shift_srl_131Z0Z_15;
    wire shift_srl_129Z0Z_15;
    wire g0_3;
    wire shift_srl_128Z0Z_14;
    wire shift_srl_128Z0Z_13;
    wire shift_srl_128Z0Z_12;
    wire shift_srl_128Z0Z_11;
    wire shift_srl_128Z0Z_10;
    wire shift_srl_128Z0Z_8;
    wire shift_srl_128Z0Z_9;
    wire g0_9_3;
    wire rco_int_0_a2_0_a2_1_1_sx_145;
    wire shift_srl_136Z0Z_15;
    wire g0_10;
    wire shift_srl_116Z0Z_14;
    wire shift_srl_116Z0Z_13;
    wire shift_srl_116Z0Z_12;
    wire shift_srl_116Z0Z_11;
    wire shift_srl_116Z0Z_10;
    wire shift_srl_116Z0Z_8;
    wire shift_srl_116Z0Z_9;
    wire clk_en_116;
    wire shift_srl_112Z0Z_0;
    wire shift_srl_112Z0Z_1;
    wire shift_srl_112Z0Z_2;
    wire shift_srl_112Z0Z_3;
    wire shift_srl_112Z0Z_4;
    wire shift_srl_112Z0Z_5;
    wire shift_srl_112Z0Z_6;
    wire shift_srl_123Z0Z_4;
    wire shift_srl_123Z0Z_5;
    wire shift_srl_123Z0Z_3;
    wire shift_srl_107Z0Z_3;
    wire shift_srl_107Z0Z_4;
    wire shift_srl_107Z0Z_5;
    wire shift_srl_107Z0Z_6;
    wire shift_srl_107Z0Z_1;
    wire shift_srl_107Z0Z_2;
    wire rco_c_151;
    wire shift_srl_1Z0Z_0;
    wire shift_srl_1Z0Z_1;
    wire shift_srl_1Z0Z_2;
    wire shift_srl_1Z0Z_3;
    wire N_10_i;
    wire shift_srl_10Z0Z_10;
    wire shift_srl_10Z0Z_11;
    wire shift_srl_10Z0Z_12;
    wire shift_srl_10Z0Z_13;
    wire shift_srl_10Z0Z_14;
    wire shift_srl_10Z0Z_9;
    wire shift_srl_10Z0Z_8;
    wire shift_srl_150Z0Z_0;
    wire shift_srl_150Z0Z_1;
    wire shift_srl_150Z0Z_2;
    wire shift_srl_150Z0Z_3;
    wire shift_srl_150Z0Z_4;
    wire shift_srl_150Z0Z_5;
    wire shift_srl_150Z0Z_6;
    wire shift_srl_150Z0Z_10;
    wire shift_srl_150Z0Z_11;
    wire shift_srl_150Z0Z_12;
    wire shift_srl_150Z0Z_13;
    wire shift_srl_150Z0Z_14;
    wire shift_srl_150Z0Z_9;
    wire shift_srl_150Z0Z_7;
    wire shift_srl_150Z0Z_8;
    wire shift_srl_147Z0Z_5;
    wire shift_srl_147Z0Z_6;
    wire shift_srl_146Z0Z_5;
    wire shift_srl_146Z0Z_3;
    wire shift_srl_146Z0Z_4;
    wire shift_srl_146Z0Z_10;
    wire shift_srl_146Z0Z_11;
    wire shift_srl_146Z0Z_12;
    wire shift_srl_146Z0Z_13;
    wire shift_srl_146Z0Z_9;
    wire shift_srl_146Z0Z_8;
    wire shift_srl_146Z0Z_6;
    wire shift_srl_146Z0Z_7;
    wire shift_srl_27Z0Z_0;
    wire shift_srl_27Z0Z_1;
    wire shift_srl_27Z0Z_2;
    wire shift_srl_27Z0Z_3;
    wire shift_srl_27Z0Z_4;
    wire shift_srl_27Z0Z_5;
    wire shift_srl_27Z0Z_6;
    wire shift_srl_27Z0Z_10;
    wire shift_srl_27Z0Z_11;
    wire shift_srl_27Z0Z_12;
    wire shift_srl_27Z0Z_7;
    wire shift_srl_27Z0Z_13;
    wire shift_srl_27Z0Z_14;
    wire shift_srl_27Z0Z_8;
    wire shift_srl_27Z0Z_9;
    wire clk_en_27;
    wire shift_srl_149Z0Z_10;
    wire shift_srl_149Z0Z_11;
    wire shift_srl_149Z0Z_12;
    wire shift_srl_149Z0Z_13;
    wire shift_srl_149Z0Z_14;
    wire shift_srl_149Z0Z_9;
    wire shift_srl_149Z0Z_8;
    wire shift_srl_149Z0Z_0;
    wire shift_srl_149Z0Z_1;
    wire shift_srl_149Z0Z_2;
    wire shift_srl_149Z0Z_3;
    wire shift_srl_149Z0Z_4;
    wire shift_srl_149Z0Z_5;
    wire shift_srl_149Z0Z_6;
    wire shift_srl_149Z0Z_7;
    wire shift_srl_123Z0Z_10;
    wire shift_srl_123Z0Z_11;
    wire shift_srl_123Z0Z_12;
    wire shift_srl_123Z0Z_13;
    wire shift_srl_123Z0Z_9;
    wire shift_srl_123Z0Z_8;
    wire shift_srl_123Z0Z_6;
    wire shift_srl_123Z0Z_7;
    wire clk_en_0_a3_0_a2_sx_123_cascade_;
    wire clk_en_0_a3_0_a2_sx_125_cascade_;
    wire shift_srl_118Z0Z_14;
    wire shift_srl_118Z0Z_13;
    wire shift_srl_118Z0Z_12;
    wire shift_srl_125Z0Z_0;
    wire shift_srl_125Z0Z_1;
    wire shift_srl_125Z0Z_2;
    wire shift_srl_125Z0Z_3;
    wire shift_srl_125Z0Z_4;
    wire shift_srl_125Z0Z_5;
    wire shift_srl_125Z0Z_6;
    wire shift_srl_113Z0Z_7;
    wire shift_srl_113Z0Z_6;
    wire shift_srl_113Z0Z_0;
    wire shift_srl_113Z0Z_1;
    wire shift_srl_113Z0Z_2;
    wire shift_srl_113Z0Z_3;
    wire shift_srl_113Z0Z_4;
    wire shift_srl_113Z0Z_5;
    wire shift_srl_110Z0Z_10;
    wire shift_srl_110Z0Z_11;
    wire shift_srl_110Z0Z_12;
    wire shift_srl_110Z0Z_13;
    wire shift_srl_110Z0Z_9;
    wire rco_c_122;
    wire shift_srl_133Z0Z_0;
    wire shift_srl_133Z0Z_1;
    wire shift_srl_133Z0Z_2;
    wire shift_srl_133Z0Z_3;
    wire clk_en_g_133;
    wire shift_srl_105Z0Z_6;
    wire shift_srl_105Z0Z_5;
    wire shift_srl_106Z0Z_2;
    wire shift_srl_106Z0Z_3;
    wire shift_srl_106Z0Z_4;
    wire shift_srl_106Z0Z_5;
    wire shift_srl_106Z0Z_6;
    wire shift_srl_106Z0Z_7;
    wire shift_srl_118Z0Z_10;
    wire shift_srl_118Z0Z_11;
    wire shift_srl_118Z0Z_9;
    wire shift_srl_118Z0Z_8;
    wire rco_c_108;
    wire rco_c_108_cascade_;
    wire rco_c_109;
    wire rco_c_107;
    wire shift_srl_0Z0Z_0;
    wire shift_srl_0Z0Z_1;
    wire shift_srl_0Z0Z_2;
    wire shift_srl_0Z0Z_3;
    wire shift_srl_0Z0Z_4;
    wire shift_srl_0Z0Z_7;
    wire shift_srl_0Z0Z_5;
    wire shift_srl_0Z0Z_6;
    wire shift_srl_0Z0Z_8;
    wire shift_srl_0Z0Z_9;
    wire rco_c_152;
    wire shift_srl_10Z0Z_4;
    wire shift_srl_10Z0Z_7;
    wire shift_srl_10Z0Z_5;
    wire shift_srl_10Z0Z_6;
    wire shift_srl_10Z0Z_15;
    wire shift_srl_10Z0Z_0;
    wire shift_srl_10Z0Z_1;
    wire shift_srl_10Z0Z_2;
    wire shift_srl_10Z0Z_3;
    wire clk_en_10;
    wire shift_srl_149_RNIU42SZ0Z_15_cascade_;
    wire clk_en_150;
    wire shift_srl_147Z0Z_14;
    wire shift_srl_147Z0Z_13;
    wire shift_srl_147Z0Z_12;
    wire shift_srl_147Z0Z_11;
    wire shift_srl_147Z0Z_10;
    wire shift_srl_147Z0Z_0;
    wire shift_srl_147Z0Z_1;
    wire shift_srl_147Z0Z_2;
    wire shift_srl_147Z0Z_3;
    wire shift_srl_147Z0Z_4;
    wire shift_srl_147Z0Z_9;
    wire shift_srl_147Z0Z_7;
    wire shift_srl_147Z0Z_8;
    wire clk_en_147;
    wire shift_srl_146Z0Z_0;
    wire shift_srl_146Z0Z_1;
    wire shift_srl_146Z0Z_2;
    wire shift_srl_160Z0Z_10;
    wire shift_srl_160Z0Z_3;
    wire shift_srl_160Z0Z_1;
    wire shift_srl_160Z0Z_2;
    wire shift_srl_160Z0Z_9;
    wire shift_srl_160Z0Z_8;
    wire shift_srl_160Z0Z_14;
    wire shift_srl_160Z0Z_7;
    wire shift_srl_160Z0Z_0;
    wire shift_srl_160Z0Z_11;
    wire shift_srl_160Z0Z_4;
    wire shift_srl_160Z0Z_5;
    wire shift_srl_160Z0Z_6;
    wire shift_srl_160Z0Z_12;
    wire shift_srl_160Z0Z_13;
    wire shift_srl_161Z0Z_10;
    wire shift_srl_161Z0Z_11;
    wire shift_srl_161Z0Z_12;
    wire shift_srl_161Z0Z_13;
    wire shift_srl_161Z0Z_14;
    wire shift_srl_161Z0Z_9;
    wire shift_srl_161Z0Z_8;
    wire rco_c_148;
    wire rco_c_147;
    wire clk_en_0_a3_0_a2_sx_149_cascade_;
    wire clk_en_149;
    wire shift_srl_146Z0Z_14;
    wire clk_en_146;
    wire shift_srl_149Z0Z_15;
    wire shift_srl_150Z0Z_15;
    wire shift_srl_150_RNIPH7TZ0Z_15_cascade_;
    wire shift_srl_146_RNIVSUTZ0Z_15_cascade_;
    wire shift_srl_126Z0Z_10;
    wire shift_srl_126Z0Z_11;
    wire shift_srl_126Z0Z_9;
    wire shift_srl_126Z0Z_7;
    wire shift_srl_126Z0Z_8;
    wire clk_en_0_a2_0_a2_sx_128_cascade_;
    wire clk_en_128;
    wire shift_srl_123Z0Z_14;
    wire shift_srl_123Z0Z_15;
    wire shift_srl_123Z0Z_0;
    wire shift_srl_123Z0Z_1;
    wire shift_srl_123Z0Z_2;
    wire clk_en_123;
    wire shift_srl_121Z0Z_10;
    wire shift_srl_121Z0Z_11;
    wire shift_srl_121Z0Z_12;
    wire shift_srl_121Z0Z_13;
    wire shift_srl_121Z0Z_14;
    wire shift_srl_121Z0Z_9;
    wire shift_srl_121Z0Z_8;
    wire shift_srl_125Z0Z_10;
    wire shift_srl_125Z0Z_11;
    wire shift_srl_125Z0Z_12;
    wire shift_srl_125Z0Z_13;
    wire shift_srl_125Z0Z_14;
    wire shift_srl_125Z0Z_9;
    wire shift_srl_125Z0Z_7;
    wire shift_srl_125Z0Z_8;
    wire clk_en_125;
    wire g0_9_1_cascade_;
    wire g0_14;
    wire g0_9_0;
    wire g0_8_2;
    wire clk_en_0_a3_0_a2_sx_110_cascade_;
    wire clk_en_0_a3_0_a2_1_110;
    wire shift_srl_108Z0Z_14;
    wire shift_srl_108Z0Z_13;
    wire shift_srl_108Z0Z_12;
    wire shift_srl_110Z0Z_0;
    wire shift_srl_110Z0Z_1;
    wire shift_srl_110Z0Z_2;
    wire shift_srl_110Z0Z_3;
    wire shift_srl_110Z0Z_4;
    wire shift_srl_110Z0Z_5;
    wire shift_srl_110Z0Z_8;
    wire shift_srl_110Z0Z_6;
    wire shift_srl_110Z0Z_7;
    wire shift_srl_107Z0Z_10;
    wire shift_srl_107Z0Z_11;
    wire shift_srl_107Z0Z_12;
    wire shift_srl_107Z0Z_13;
    wire shift_srl_107Z0Z_14;
    wire shift_srl_107Z0Z_9;
    wire shift_srl_107Z0Z_7;
    wire shift_srl_107Z0Z_8;
    wire clk_en_107;
    wire rco_c_106;
    wire shift_srl_106_RNIPC6S1Z0Z_15;
    wire shift_srl_106_RNIPC6S1Z0Z_15_cascade_;
    wire rco_int_0_a3_0_a2_out_0_cascade_;
    wire clk_en_0_a3_0_a2_sx_109;
    wire shift_srl_106Z0Z_10;
    wire shift_srl_106Z0Z_11;
    wire shift_srl_106Z0Z_12;
    wire shift_srl_106Z0Z_13;
    wire shift_srl_106Z0Z_14;
    wire shift_srl_106Z0Z_8;
    wire shift_srl_106Z0Z_9;
    wire shift_srl_106Z0Z_0;
    wire shift_srl_106Z0Z_1;
    wire clk_en_106;
    wire shift_srl_108Z0Z_0;
    wire shift_srl_108Z0Z_1;
    wire shift_srl_108Z0Z_2;
    wire shift_srl_108Z0Z_3;
    wire shift_srl_108Z0Z_4;
    wire shift_srl_108Z0Z_5;
    wire shift_srl_108Z0Z_6;
    wire shift_srl_108Z0Z_10;
    wire shift_srl_108Z0Z_11;
    wire shift_srl_108Z0Z_9;
    wire shift_srl_108Z0Z_7;
    wire shift_srl_108Z0Z_8;
    wire clk_en_108;
    wire shift_srl_0Z0Z_10;
    wire shift_srl_0Z0Z_11;
    wire shift_srl_0Z0Z_12;
    wire shift_srl_0Z0Z_13;
    wire shift_srl_0Z0Z_14;
    wire shift_srl_148Z0Z_10;
    wire shift_srl_148Z0Z_11;
    wire shift_srl_148Z0Z_12;
    wire shift_srl_148Z0Z_13;
    wire shift_srl_148Z0Z_14;
    wire shift_srl_148Z0Z_9;
    wire shift_srl_148Z0Z_8;
    wire shift_srl_147Z0Z_15;
    wire shift_srl_148Z0Z_15;
    wire shift_srl_148Z0Z_0;
    wire shift_srl_148Z0Z_1;
    wire en_in_c;
    wire shift_srl_1Z0Z_15;
    wire N_452_i;
    wire shift_srl_154Z0Z_10;
    wire shift_srl_154Z0Z_9;
    wire shift_srl_154Z0Z_8;
    wire shift_srl_154Z0Z_7;
    wire shift_srl_154Z0Z_6;
    wire shift_srl_154Z0Z_5;
    wire shift_srl_154Z0Z_3;
    wire shift_srl_154Z0Z_4;
    wire shift_srl_157Z0Z_10;
    wire shift_srl_157Z0Z_11;
    wire shift_srl_157Z0Z_5;
    wire shift_srl_157Z0Z_9;
    wire shift_srl_157Z0Z_8;
    wire clk_en_160;
    wire shift_srl_154Z0Z_14;
    wire shift_srl_154Z0Z_13;
    wire shift_srl_154Z0Z_11;
    wire shift_srl_154Z0Z_12;
    wire clk_en_154;
    wire shift_srl_161Z0Z_0;
    wire shift_srl_161Z0Z_1;
    wire shift_srl_161Z0Z_2;
    wire shift_srl_161Z0Z_3;
    wire shift_srl_161Z0Z_4;
    wire shift_srl_161Z0Z_5;
    wire shift_srl_161Z0Z_6;
    wire shift_srl_161Z0Z_7;
    wire clk_en_161;
    wire shift_srl_124Z0Z_10;
    wire shift_srl_124Z0Z_11;
    wire shift_srl_124Z0Z_12;
    wire shift_srl_124Z0Z_13;
    wire shift_srl_124Z0Z_9;
    wire shift_srl_124Z0Z_8;
    wire shift_srl_126Z0Z_12;
    wire shift_srl_126Z0Z_0;
    wire shift_srl_126Z0Z_1;
    wire shift_srl_126Z0Z_2;
    wire shift_srl_126Z0Z_3;
    wire shift_srl_126Z0Z_4;
    wire shift_srl_126Z0Z_5;
    wire shift_srl_126Z0Z_6;
    wire shift_srl_126Z0Z_13;
    wire shift_srl_126Z0Z_14;
    wire rco_c_126;
    wire rco_c_123;
    wire clk_en_126;
    wire shift_srl_124Z0Z_14;
    wire rco_int_0_a2_1_a2_0_127_cascade_;
    wire rco_int_0_a2_0_a2_1_sx_sx_145;
    wire rco_int_0_a2_0_a2_1_sx_145_cascade_;
    wire shift_srl_122Z0Z_10;
    wire shift_srl_122Z0Z_11;
    wire shift_srl_122Z0Z_12;
    wire shift_srl_122Z0Z_13;
    wire shift_srl_122Z0Z_14;
    wire shift_srl_122Z0Z_9;
    wire shift_srl_122Z0Z_8;
    wire shift_srl_113Z0Z_14;
    wire shift_srl_113Z0Z_13;
    wire shift_srl_113Z0Z_12;
    wire shift_srl_113Z0Z_11;
    wire shift_srl_113Z0Z_10;
    wire shift_srl_113Z0Z_8;
    wire shift_srl_113Z0Z_9;
    wire clk_en_113;
    wire shift_srl_112Z0Z_10;
    wire shift_srl_112Z0Z_11;
    wire shift_srl_112Z0Z_12;
    wire shift_srl_112Z0Z_13;
    wire shift_srl_112Z0Z_14;
    wire shift_srl_112Z0Z_9;
    wire shift_srl_112Z0Z_7;
    wire shift_srl_112Z0Z_8;
    wire shift_srl_109Z0Z_10;
    wire shift_srl_109Z0Z_11;
    wire shift_srl_109Z0Z_12;
    wire shift_srl_109Z0Z_13;
    wire shift_srl_109Z0Z_14;
    wire shift_srl_109Z0Z_9;
    wire shift_srl_109Z0Z_8;
    wire shift_srl_109Z0Z_0;
    wire shift_srl_109Z0Z_1;
    wire shift_srl_109Z0Z_2;
    wire shift_srl_109Z0Z_3;
    wire shift_srl_109Z0Z_4;
    wire shift_srl_109Z0Z_5;
    wire shift_srl_109Z0Z_6;
    wire shift_srl_109Z0Z_7;
    wire clk_en_109;
    wire rco_c_105;
    wire shift_srl_105Z0Z_0;
    wire shift_srl_105Z0Z_1;
    wire shift_srl_105Z0Z_2;
    wire shift_srl_105Z0Z_3;
    wire shift_srl_105Z0Z_4;
    wire shift_srl_105Z0Z_10;
    wire shift_srl_105Z0Z_11;
    wire shift_srl_105Z0Z_12;
    wire shift_srl_105Z0Z_13;
    wire shift_srl_105Z0Z_14;
    wire shift_srl_105Z0Z_9;
    wire shift_srl_105Z0Z_7;
    wire shift_srl_105Z0Z_8;
    wire clk_en_105;
    wire shift_srl_104Z0Z_0;
    wire shift_srl_104Z0Z_1;
    wire shift_srl_104Z0Z_2;
    wire shift_srl_104Z0Z_3;
    wire shift_srl_104Z0Z_4;
    wire shift_srl_104Z0Z_5;
    wire shift_srl_104Z0Z_6;
    wire shift_srl_101Z0Z_10;
    wire shift_srl_101Z0Z_11;
    wire shift_srl_101Z0Z_12;
    wire shift_srl_101Z0Z_13;
    wire shift_srl_101Z0Z_9;
    wire shift_srl_101Z0Z_8;
    wire shift_srl_101Z0Z_7;
    wire rco_c_101;
    wire shift_srl_101Z0Z_0;
    wire shift_srl_101Z0Z_1;
    wire shift_srl_101Z0Z_2;
    wire shift_srl_101Z0Z_3;
    wire shift_srl_101Z0Z_4;
    wire shift_srl_101Z0Z_5;
    wire shift_srl_101Z0Z_6;
    wire shift_srl_149_RNIU42SZ0Z_15;
    wire rco_c_149;
    wire shift_srl_148Z0Z_6;
    wire shift_srl_148Z0Z_7;
    wire shift_srl_148Z0Z_2;
    wire shift_srl_148Z0Z_3;
    wire shift_srl_148Z0Z_4;
    wire shift_srl_148Z0Z_5;
    wire clk_en_148;
    wire shift_srl_25Z0Z_3;
    wire shift_srl_25Z0Z_0;
    wire shift_srl_25Z0Z_1;
    wire shift_srl_25Z0Z_2;
    wire rco_c_24;
    wire shift_srl_157Z0Z_0;
    wire shift_srl_157Z0Z_1;
    wire shift_srl_157Z0Z_2;
    wire shift_srl_157Z0Z_3;
    wire shift_srl_157Z0Z_4;
    wire shift_srl_157Z0Z_12;
    wire shift_srl_157Z0Z_13;
    wire shift_srl_157Z0Z_14;
    wire shift_srl_157Z0Z_6;
    wire shift_srl_157Z0Z_7;
    wire clk_en_157;
    wire shift_srl_155Z0Z_0;
    wire shift_srl_155Z0Z_1;
    wire shift_srl_155Z0Z_6;
    wire shift_srl_155Z0Z_9;
    wire shift_srl_155Z0Z_5;
    wire shift_srl_155Z0Z_4;
    wire shift_srl_155Z0Z_7;
    wire shift_srl_155Z0Z_8;
    wire shift_srl_155Z0Z_12;
    wire shift_srl_155Z0Z_13;
    wire shift_srl_155Z0Z_14;
    wire shift_srl_155Z0Z_2;
    wire shift_srl_155Z0Z_3;
    wire shift_srl_155Z0Z_10;
    wire shift_srl_155Z0Z_11;
    wire clk_en_155;
    wire shift_srl_124Z0Z_0;
    wire shift_srl_124Z0Z_1;
    wire shift_srl_124Z0Z_2;
    wire shift_srl_124Z0Z_3;
    wire shift_srl_124Z0Z_4;
    wire shift_srl_124Z0Z_5;
    wire shift_srl_124Z0Z_6;
    wire shift_srl_124Z0Z_7;
    wire shift_srl_144Z0Z_0;
    wire shift_srl_144Z0Z_1;
    wire shift_srl_144Z0Z_2;
    wire shift_srl_144Z0Z_3;
    wire shift_srl_144Z0Z_4;
    wire shift_srl_144Z0Z_5;
    wire shift_srl_144Z0Z_6;
    wire shift_srl_144Z0Z_10;
    wire shift_srl_144Z0Z_11;
    wire shift_srl_144Z0Z_12;
    wire shift_srl_144Z0Z_13;
    wire shift_srl_144Z0Z_14;
    wire shift_srl_144Z0Z_9;
    wire shift_srl_144Z0Z_7;
    wire shift_srl_144Z0Z_8;
    wire shift_srl_116Z0Z_15;
    wire rco_int_0_a2_1_a2_1_118_cascade_;
    wire rco_c_118_cascade_;
    wire rco_int_0_a2_1_a2_1_123;
    wire clk_en_124;
    wire shift_srl_117Z0Z_14;
    wire shift_srl_117Z0Z_13;
    wire shift_srl_117Z0Z_12;
    wire shift_srl_117Z0Z_11;
    wire shift_srl_117Z0Z_10;
    wire shift_srl_114Z0Z_10;
    wire shift_srl_114Z0Z_11;
    wire shift_srl_114Z0Z_12;
    wire shift_srl_114Z0Z_13;
    wire shift_srl_114Z0Z_14;
    wire shift_srl_114Z0Z_9;
    wire shift_srl_114Z0Z_8;
    wire shift_srl_114Z0Z_15;
    wire shift_srl_114Z0Z_0;
    wire shift_srl_114Z0Z_1;
    wire shift_srl_114Z0Z_2;
    wire shift_srl_114Z0Z_3;
    wire shift_srl_114Z0Z_4;
    wire shift_srl_114Z0Z_5;
    wire shift_srl_114Z0Z_6;
    wire shift_srl_114Z0Z_7;
    wire shift_srl_118Z0Z_0;
    wire shift_srl_118Z0Z_1;
    wire shift_srl_118Z0Z_2;
    wire shift_srl_118Z0Z_3;
    wire shift_srl_118Z0Z_4;
    wire shift_srl_118Z0Z_5;
    wire shift_srl_118Z0Z_6;
    wire shift_srl_118Z0Z_7;
    wire shift_srl_100Z0Z_0;
    wire shift_srl_100Z0Z_1;
    wire shift_srl_100Z0Z_2;
    wire shift_srl_100Z0Z_3;
    wire shift_srl_100Z0Z_4;
    wire shift_srl_100Z0Z_5;
    wire shift_srl_104Z0Z_10;
    wire shift_srl_104Z0Z_11;
    wire shift_srl_104Z0Z_12;
    wire shift_srl_104Z0Z_13;
    wire shift_srl_104Z0Z_14;
    wire shift_srl_104Z0Z_9;
    wire shift_srl_104Z0Z_7;
    wire shift_srl_104Z0Z_8;
    wire shift_srl_102_RNIN8GNZ0Z_15_cascade_;
    wire clk_en_104;
    wire shift_srl_101Z0Z_14;
    wire shift_srl_105Z0Z_15;
    wire shift_srl_106Z0Z_15;
    wire clk_en_101;
    wire clk_en_0_a3_0_a2_sx_103_cascade_;
    wire rco_c_102;
    wire rco_c_103;
    wire shift_srl_103Z0Z_0;
    wire shift_srl_103Z0Z_1;
    wire shift_srl_103Z0Z_2;
    wire shift_srl_103Z0Z_3;
    wire shift_srl_103Z0Z_4;
    wire shift_srl_103Z0Z_5;
    wire shift_srl_100Z0Z_9;
    wire shift_srl_100Z0Z_8;
    wire shift_srl_100Z0Z_6;
    wire shift_srl_100Z0Z_7;
    wire shift_srl_103Z0Z_6;
    wire rco_c_165;
    wire shift_srl_90Z0Z_9;
    wire shift_srl_90Z0Z_8;
    wire shift_srl_90Z0Z_6;
    wire shift_srl_90Z0Z_7;
    wire shift_srl_91Z0Z_10;
    wire shift_srl_91Z0Z_11;
    wire shift_srl_91Z0Z_12;
    wire shift_srl_91Z0Z_13;
    wire shift_srl_91Z0Z_14;
    wire shift_srl_91Z0Z_9;
    wire shift_srl_91Z0Z_8;
    wire shift_srl_91Z0Z_0;
    wire shift_srl_91Z0Z_1;
    wire shift_srl_91Z0Z_2;
    wire shift_srl_91Z0Z_3;
    wire shift_srl_91Z0Z_4;
    wire shift_srl_91Z0Z_5;
    wire shift_srl_91Z0Z_6;
    wire shift_srl_91Z0Z_7;
    wire shift_srl_25Z0Z_4;
    wire shift_srl_25Z0Z_5;
    wire shift_srl_25Z0Z_6;
    wire shift_srl_25Z0Z_10;
    wire shift_srl_25Z0Z_11;
    wire shift_srl_25Z0Z_12;
    wire shift_srl_25Z0Z_13;
    wire shift_srl_25Z0Z_14;
    wire shift_srl_25Z0Z_9;
    wire shift_srl_25Z0Z_7;
    wire shift_srl_25Z0Z_8;
    wire clk_en_25;
    wire shift_srl_89Z0Z_0;
    wire shift_srl_89Z0Z_1;
    wire shift_srl_89Z0Z_2;
    wire shift_srl_89Z0Z_3;
    wire shift_srl_89Z0Z_4;
    wire shift_srl_89Z0Z_5;
    wire shift_srl_89Z0Z_6;
    wire shift_srl_89Z0Z_10;
    wire shift_srl_89Z0Z_11;
    wire shift_srl_89Z0Z_12;
    wire shift_srl_89Z0Z_13;
    wire shift_srl_89Z0Z_9;
    wire shift_srl_89Z0Z_7;
    wire shift_srl_89Z0Z_8;
    wire shift_srl_24Z0Z_0;
    wire shift_srl_24Z0Z_1;
    wire shift_srl_24Z0Z_2;
    wire shift_srl_143Z0Z_0;
    wire shift_srl_143Z0Z_1;
    wire shift_srl_143Z0Z_2;
    wire shift_srl_143Z0Z_3;
    wire shift_srl_143Z0Z_4;
    wire shift_srl_143Z0Z_5;
    wire shift_srl_143Z0Z_6;
    wire shift_srl_26Z0Z_0;
    wire shift_srl_26Z0Z_1;
    wire shift_srl_26Z0Z_2;
    wire shift_srl_26Z0Z_3;
    wire shift_srl_26Z0Z_4;
    wire shift_srl_26Z0Z_5;
    wire shift_srl_26Z0Z_6;
    wire shift_srl_121Z0Z_0;
    wire shift_srl_121Z0Z_1;
    wire shift_srl_121Z0Z_2;
    wire shift_srl_121Z0Z_3;
    wire shift_srl_121Z0Z_4;
    wire shift_srl_121Z0Z_5;
    wire shift_srl_121Z0Z_6;
    wire shift_srl_121Z0Z_7;
    wire clk_en_121;
    wire shift_srl_143Z0Z_10;
    wire shift_srl_143Z0Z_11;
    wire shift_srl_143Z0Z_12;
    wire shift_srl_143Z0Z_13;
    wire shift_srl_143Z0Z_14;
    wire shift_srl_143Z0Z_9;
    wire shift_srl_143Z0Z_7;
    wire shift_srl_143Z0Z_8;
    wire shift_srl_117Z0Z_0;
    wire shift_srl_117Z0Z_1;
    wire shift_srl_117Z0Z_2;
    wire shift_srl_117Z0Z_3;
    wire shift_srl_117Z0Z_4;
    wire shift_srl_117Z0Z_5;
    wire shift_srl_117Z0Z_6;
    wire rco_c_143;
    wire rco_c_142;
    wire clk_en_0_a3_0_a2_sx_144_cascade_;
    wire clk_en_144;
    wire clk_en_0_a3_0_a2_sx_143_cascade_;
    wire clk_en_143;
    wire rco_c_99_cascade_;
    wire shift_srl_122Z0Z_15;
    wire shift_srl_122Z0Z_0;
    wire shift_srl_122Z0Z_1;
    wire shift_srl_122Z0Z_2;
    wire shift_srl_122Z0Z_3;
    wire shift_srl_122Z0Z_4;
    wire shift_srl_122Z0Z_5;
    wire shift_srl_122Z0Z_6;
    wire shift_srl_122Z0Z_7;
    wire clk_en_122;
    wire shift_srl_142Z0Z_10;
    wire shift_srl_142Z0Z_11;
    wire shift_srl_142Z0Z_12;
    wire shift_srl_142Z0Z_13;
    wire shift_srl_142Z0Z_14;
    wire shift_srl_142Z0Z_9;
    wire shift_srl_142Z0Z_8;
    wire clk_en_112;
    wire N_91;
    wire shift_srl_118Z0Z_15;
    wire shift_srl_111Z0Z_14;
    wire shift_srl_111Z0Z_13;
    wire shift_srl_111Z0Z_0;
    wire shift_srl_111Z0Z_1;
    wire shift_srl_111Z0Z_2;
    wire shift_srl_111Z0Z_3;
    wire shift_srl_111Z0Z_4;
    wire shift_srl_111Z0Z_5;
    wire shift_srl_111Z0Z_6;
    wire shift_srl_112Z0Z_15;
    wire shift_srl_113Z0Z_15;
    wire shift_srl_112_RNIV16I3Z0Z_15_cascade_;
    wire clk_en_114;
    wire clk_en_118;
    wire shift_srl_111Z0Z_15;
    wire rco_c_111;
    wire rco_int_0_a2_1_a2_1_120;
    wire rco_c_199;
    wire shift_srl_199Z0Z_0;
    wire shift_srl_199Z0Z_1;
    wire shift_srl_199Z0Z_2;
    wire shift_srl_199Z0Z_3;
    wire shift_srl_199Z0Z_4;
    wire shift_srl_199Z0Z_5;
    wire shift_srl_199Z0Z_6;
    wire shift_srl_102Z0Z_10;
    wire shift_srl_102Z0Z_11;
    wire shift_srl_102Z0Z_12;
    wire shift_srl_102Z0Z_13;
    wire shift_srl_102Z0Z_14;
    wire shift_srl_102Z0Z_7;
    wire shift_srl_104Z0Z_15;
    wire shift_srl_101Z0Z_15;
    wire rco_int_0_a3_0_a2_s_0_sx_104;
    wire shift_srl_100Z0Z_14;
    wire shift_srl_100Z0Z_13;
    wire shift_srl_100Z0Z_12;
    wire shift_srl_100Z0Z_10;
    wire shift_srl_100Z0Z_11;
    wire clk_en_100;
    wire shift_srl_103Z0Z_10;
    wire shift_srl_103Z0Z_11;
    wire shift_srl_103Z0Z_12;
    wire shift_srl_103Z0Z_13;
    wire shift_srl_103Z0Z_14;
    wire shift_srl_103Z0Z_15;
    wire shift_srl_103Z0Z_9;
    wire shift_srl_103Z0Z_7;
    wire shift_srl_103Z0Z_8;
    wire clk_en_103;
    wire rco_c_87;
    wire rco_c_86;
    wire shift_srl_90Z0Z_0;
    wire shift_srl_90Z0Z_1;
    wire shift_srl_90Z0Z_2;
    wire shift_srl_90Z0Z_3;
    wire shift_srl_90Z0Z_4;
    wire shift_srl_90Z0Z_5;
    wire clk_en_91;
    wire shift_srl_90Z0Z_14;
    wire shift_srl_90Z0Z_13;
    wire shift_srl_90Z0Z_12;
    wire shift_srl_90Z0Z_10;
    wire shift_srl_90Z0Z_11;
    wire clk_en_90;
    wire shift_srl_87Z0Z_10;
    wire shift_srl_87Z0Z_11;
    wire shift_srl_87Z0Z_12;
    wire shift_srl_87Z0Z_13;
    wire shift_srl_87Z0Z_14;
    wire shift_srl_87Z0Z_9;
    wire shift_srl_87Z0Z_8;
    wire shift_srl_86Z0Z_0;
    wire shift_srl_86Z0Z_1;
    wire shift_srl_86Z0Z_2;
    wire shift_srl_86Z0Z_3;
    wire shift_srl_86Z0Z_4;
    wire shift_srl_86Z0Z_11;
    wire shift_srl_84Z0Z_0;
    wire shift_srl_84Z0Z_1;
    wire shift_srl_84Z0Z_2;
    wire shift_srl_84Z0Z_3;
    wire shift_srl_84Z0Z_4;
    wire shift_srl_84Z0Z_5;
    wire shift_srl_84Z0Z_6;
    wire shift_srl_84Z0Z_10;
    wire shift_srl_84Z0Z_11;
    wire shift_srl_84Z0Z_12;
    wire shift_srl_84Z0Z_13;
    wire shift_srl_84Z0Z_14;
    wire shift_srl_84Z0Z_9;
    wire shift_srl_84Z0Z_7;
    wire shift_srl_84Z0Z_8;
    wire rco_int_0_a2_0_a2_0_sx_91_cascade_;
    wire shift_srl_91_RNI20EN1Z0Z_15_cascade_;
    wire shift_srl_83_RNIKTI68Z0Z_15_cascade_;
    wire clk_en_84;
    wire clk_en_84_cascade_;
    wire shift_srl_89Z0Z_14;
    wire clk_en_89;
    wire shift_srl_24Z0Z_3;
    wire shift_srl_24Z0Z_4;
    wire shift_srl_24Z0Z_7;
    wire shift_srl_24Z0Z_5;
    wire shift_srl_24Z0Z_6;
    wire shift_srl_152Z0Z_10;
    wire shift_srl_152Z0Z_11;
    wire shift_srl_152Z0Z_12;
    wire shift_srl_152Z0Z_13;
    wire shift_srl_152Z0Z_14;
    wire shift_srl_152Z0Z_9;
    wire shift_srl_152Z0Z_8;
    wire shift_srl_153Z0Z_10;
    wire shift_srl_153Z0Z_11;
    wire shift_srl_153Z0Z_12;
    wire shift_srl_153Z0Z_13;
    wire shift_srl_153Z0Z_14;
    wire shift_srl_153Z0Z_9;
    wire shift_srl_153Z0Z_8;
    wire shift_srl_153Z0Z_15;
    wire shift_srl_153Z0Z_0;
    wire shift_srl_153Z0Z_1;
    wire shift_srl_153Z0Z_2;
    wire shift_srl_153Z0Z_3;
    wire shift_srl_153Z0Z_4;
    wire shift_srl_153Z0Z_5;
    wire shift_srl_153Z0Z_6;
    wire shift_srl_153Z0Z_7;
    wire shift_srl_141Z0Z_10;
    wire shift_srl_141Z0Z_11;
    wire shift_srl_141Z0Z_12;
    wire shift_srl_141Z0Z_9;
    wire shift_srl_141Z0Z_7;
    wire shift_srl_141Z0Z_8;
    wire shift_srl_141Z0Z_4;
    wire shift_srl_141Z0Z_5;
    wire shift_srl_141Z0Z_6;
    wire shift_srl_141Z0Z_3;
    wire shift_srl_141Z0Z_13;
    wire shift_srl_144Z0Z_15;
    wire rco_int_0_a2_0_a2_0_sx_144_cascade_;
    wire shift_srl_143Z0Z_15;
    wire shift_srl_141Z0Z_14;
    wire shift_srl_141Z0Z_15;
    wire shift_srl_141Z0Z_0;
    wire shift_srl_141Z0Z_1;
    wire shift_srl_141Z0Z_2;
    wire shift_srl_145Z0Z_10;
    wire shift_srl_145Z0Z_11;
    wire shift_srl_145Z0Z_12;
    wire shift_srl_145Z0Z_13;
    wire shift_srl_145Z0Z_14;
    wire shift_srl_145Z0Z_9;
    wire shift_srl_145Z0Z_8;
    wire rco_int_0_a3_0_a2_138_m6_0_a2_7_4_cascade_;
    wire rco_int_0_a3_0_a2_138_m6_0_a2_7_cascade_;
    wire N_122_i;
    wire rco_c_110;
    wire rco_int_0_a3_0_a2_138_m6_0_a2_7_4_1;
    wire rco_int_0_a3_0_a2_138_m6_0_a2_7_0;
    wire shift_srl_120_RNIG17D2Z0Z_15;
    wire shift_srl_139Z0Z_0;
    wire shift_srl_139Z0Z_1;
    wire shift_srl_139Z0Z_2;
    wire shift_srl_139Z0Z_3;
    wire shift_srl_139Z0Z_4;
    wire shift_srl_139Z0Z_5;
    wire shift_srl_139Z0Z_6;
    wire rco_int_0_a2_0_a2_s_0_1_110_cascade_;
    wire rco_int_0_a2_0_a2_out_5_cascade_;
    wire shift_srl_110Z0Z_14;
    wire clk_en_110;
    wire shift_srl_110Z0Z_15;
    wire shift_srl_109Z0Z_15;
    wire shift_srl_107Z0Z_15;
    wire shift_srl_108Z0Z_15;
    wire rco_int_0_a3_0_a2_s_0_1_104;
    wire shift_srl_110_RNI91581Z0Z_15_cascade_;
    wire rco_int_0_a2_0_a2_s_0_sx_110;
    wire rco_int_0_a3_0_a2_138_m6_0_a2_7_4;
    wire shift_srl_110_RNI4QDG2Z0Z_15_cascade_;
    wire g0_4;
    wire g0_0;
    wire rco_int_0_a3_0_a2_0_132;
    wire g0_9_cascade_;
    wire g0_16_cascade_;
    wire rco_int_0_a3_0_a2_0_138;
    wire g0_12;
    wire rco_int_0_a2_1_a2_out_0;
    wire g0_8;
    wire shift_srl_199Z0Z_10;
    wire shift_srl_199Z0Z_11;
    wire shift_srl_199Z0Z_12;
    wire shift_srl_199Z0Z_13;
    wire shift_srl_199Z0Z_14;
    wire shift_srl_199Z0Z_15;
    wire shift_srl_199Z0Z_9;
    wire shift_srl_199Z0Z_7;
    wire shift_srl_199Z0Z_8;
    wire clk_en_199;
    wire shift_srl_102Z0Z_15;
    wire shift_srl_102Z0Z_0;
    wire shift_srl_102Z0Z_1;
    wire shift_srl_102Z0Z_2;
    wire shift_srl_102Z0Z_3;
    wire shift_srl_102Z0Z_4;
    wire shift_srl_102Z0Z_5;
    wire shift_srl_102Z0Z_6;
    wire shift_srl_102Z0Z_8;
    wire shift_srl_102Z0Z_9;
    wire clk_en_102;
    wire shift_srl_139Z0Z_7;
    wire shift_srl_139Z0Z_8;
    wire shift_srl_139Z0Z_9;
    wire shift_srl_139Z0Z_10;
    wire shift_srl_85Z0Z_10;
    wire shift_srl_85Z0Z_11;
    wire shift_srl_85Z0Z_12;
    wire shift_srl_85Z0Z_13;
    wire shift_srl_85Z0Z_14;
    wire shift_srl_85Z0Z_9;
    wire shift_srl_85Z0Z_8;
    wire shift_srl_88Z0Z_10;
    wire shift_srl_88Z0Z_11;
    wire shift_srl_88Z0Z_12;
    wire shift_srl_88Z0Z_13;
    wire shift_srl_88Z0Z_14;
    wire shift_srl_88Z0Z_9;
    wire shift_srl_88Z0Z_8;
    wire rco_c_88;
    wire rco_c_83_cascade_;
    wire shift_srl_86_RNI8K1LZ0Z_15;
    wire shift_srl_86Z0Z_10;
    wire shift_srl_86Z0Z_5;
    wire shift_srl_86Z0Z_6;
    wire shift_srl_86Z0Z_12;
    wire shift_srl_86Z0Z_13;
    wire shift_srl_86Z0Z_9;
    wire shift_srl_86Z0Z_7;
    wire shift_srl_86Z0Z_8;
    wire shift_srl_43Z0Z_11;
    wire shift_srl_43Z0Z_10;
    wire shift_srl_43Z0Z_12;
    wire shift_srl_43Z0Z_13;
    wire shift_srl_43Z0Z_14;
    wire shift_srl_43Z0Z_9;
    wire shift_srl_43Z0Z_8;
    wire shift_srl_43Z0Z_2;
    wire shift_srl_43Z0Z_3;
    wire shift_srl_43Z0Z_4;
    wire shift_srl_43Z0Z_5;
    wire shift_srl_43Z0Z_0;
    wire shift_srl_43Z0Z_1;
    wire shift_srl_43Z0Z_6;
    wire shift_srl_43Z0Z_7;
    wire shift_srl_24Z0Z_10;
    wire shift_srl_24Z0Z_11;
    wire shift_srl_24Z0Z_12;
    wire shift_srl_24Z0Z_13;
    wire shift_srl_24Z0Z_14;
    wire shift_srl_24Z0Z_8;
    wire shift_srl_24Z0Z_9;
    wire clk_en_24;
    wire shift_srl_152Z0Z_0;
    wire shift_srl_152Z0Z_1;
    wire shift_srl_152Z0Z_2;
    wire shift_srl_152Z0Z_3;
    wire shift_srl_152Z0Z_4;
    wire shift_srl_152Z0Z_5;
    wire shift_srl_152Z0Z_6;
    wire shift_srl_152Z0Z_7;
    wire shift_srl_152Z0Z_15;
    wire clk_en_0_a3_0_a2_sx_153_cascade_;
    wire clk_en_153;
    wire shift_srl_91_RNIUH4HPZ0Z_15_cascade_;
    wire rco_c_145_cascade_;
    wire clk_en_152;
    wire shift_srl_151Z0Z_0;
    wire shift_srl_151Z0Z_1;
    wire shift_srl_151Z0Z_2;
    wire shift_srl_151Z0Z_3;
    wire shift_srl_151Z0Z_4;
    wire shift_srl_151Z0Z_5;
    wire shift_srl_151Z0Z_6;
    wire shift_srl_151Z0Z_10;
    wire shift_srl_151Z0Z_11;
    wire shift_srl_151Z0Z_12;
    wire shift_srl_151Z0Z_13;
    wire shift_srl_151Z0Z_14;
    wire shift_srl_151Z0Z_15;
    wire shift_srl_151Z0Z_9;
    wire shift_srl_151Z0Z_7;
    wire shift_srl_151Z0Z_8;
    wire clk_en_151;
    wire shift_srl_140Z0Z_10;
    wire shift_srl_140Z0Z_11;
    wire shift_srl_140Z0Z_12;
    wire shift_srl_140Z0Z_13;
    wire shift_srl_140Z0Z_14;
    wire shift_srl_140Z0Z_9;
    wire shift_srl_140Z0Z_8;
    wire shift_srl_140Z0Z_0;
    wire shift_srl_140Z0Z_1;
    wire shift_srl_140Z0Z_2;
    wire shift_srl_140Z0Z_3;
    wire shift_srl_140Z0Z_4;
    wire shift_srl_140Z0Z_5;
    wire shift_srl_140Z0Z_6;
    wire shift_srl_140Z0Z_7;
    wire N_124_i;
    wire shift_srl_145Z0Z_15;
    wire shift_srl_145Z0Z_0;
    wire shift_srl_145Z0Z_1;
    wire shift_srl_145Z0Z_2;
    wire shift_srl_145Z0Z_3;
    wire shift_srl_145Z0Z_4;
    wire shift_srl_145Z0Z_5;
    wire shift_srl_145Z0Z_6;
    wire shift_srl_145Z0Z_7;
    wire clk_en_145;
    wire shift_srl_142Z0Z_15;
    wire shift_srl_142Z0Z_0;
    wire shift_srl_142Z0Z_1;
    wire shift_srl_142Z0Z_2;
    wire shift_srl_142Z0Z_3;
    wire shift_srl_142Z0Z_4;
    wire shift_srl_142Z0Z_5;
    wire shift_srl_142Z0Z_6;
    wire shift_srl_142Z0Z_7;
    wire clk_en_142;
    wire shift_srl_120Z0Z_10;
    wire shift_srl_120Z0Z_11;
    wire shift_srl_120Z0Z_12;
    wire shift_srl_120Z0Z_13;
    wire shift_srl_120Z0Z_14;
    wire shift_srl_120Z0Z_9;
    wire shift_srl_120Z0Z_8;
    wire N_162;
    wire rco_c_115;
    wire shift_srl_115Z0Z_15;
    wire shift_srl_115Z0Z_0;
    wire shift_srl_115Z0Z_1;
    wire shift_srl_115Z0Z_2;
    wire shift_srl_115Z0Z_3;
    wire shift_srl_115Z0Z_4;
    wire shift_srl_115Z0Z_5;
    wire shift_srl_115Z0Z_10;
    wire shift_srl_115Z0Z_11;
    wire shift_srl_115Z0Z_12;
    wire shift_srl_115Z0Z_13;
    wire shift_srl_115Z0Z_14;
    wire shift_srl_115Z0Z_9;
    wire shift_srl_115Z0Z_8;
    wire shift_srl_115Z0Z_6;
    wire shift_srl_115Z0Z_7;
    wire clk_en_115;
    wire rco_c_194;
    wire rco_c_193;
    wire rco_c_184;
    wire rco_c_187;
    wire rco_c_191;
    wire rco_c_195;
    wire shift_srl_194Z0Z_0;
    wire shift_srl_139Z0Z_11;
    wire rco_c_90;
    wire rco_c_91;
    wire shift_srl_85Z0Z_0;
    wire shift_srl_85Z0Z_1;
    wire shift_srl_85Z0Z_2;
    wire shift_srl_85Z0Z_3;
    wire shift_srl_85Z0Z_4;
    wire shift_srl_85Z0Z_5;
    wire shift_srl_85Z0Z_6;
    wire shift_srl_85Z0Z_7;
    wire clk_en_85;
    wire shift_srl_88Z0Z_0;
    wire shift_srl_88Z0Z_1;
    wire shift_srl_88Z0Z_2;
    wire shift_srl_88Z0Z_3;
    wire shift_srl_88Z0Z_4;
    wire shift_srl_88Z0Z_5;
    wire shift_srl_88Z0Z_6;
    wire shift_srl_88Z0Z_7;
    wire clk_en_88;
    wire shift_srl_87Z0Z_0;
    wire shift_srl_87Z0Z_1;
    wire shift_srl_87Z0Z_2;
    wire shift_srl_87Z0Z_3;
    wire shift_srl_87Z0Z_4;
    wire shift_srl_87Z0Z_5;
    wire shift_srl_87Z0Z_6;
    wire shift_srl_87Z0Z_7;
    wire clk_en_87;
    wire shift_srl_99Z0Z_10;
    wire shift_srl_99Z0Z_11;
    wire shift_srl_99Z0Z_12;
    wire shift_srl_99Z0Z_13;
    wire shift_srl_99Z0Z_9;
    wire shift_srl_99Z0Z_8;
    wire shift_srl_99Z0Z_6;
    wire shift_srl_99Z0Z_7;
    wire shift_srl_42Z0Z_6;
    wire shift_srl_42Z0Z_5;
    wire shift_srl_42Z0Z_10;
    wire shift_srl_42Z0Z_11;
    wire shift_srl_42Z0Z_12;
    wire shift_srl_42Z0Z_13;
    wire shift_srl_42Z0Z_14;
    wire shift_srl_42Z0Z_9;
    wire shift_srl_42Z0Z_7;
    wire shift_srl_42Z0Z_8;
    wire rco_c_43;
    wire rco_c_42;
    wire shift_srl_42Z0Z_0;
    wire shift_srl_42Z0Z_1;
    wire shift_srl_42Z0Z_2;
    wire shift_srl_42Z0Z_3;
    wire shift_srl_42Z0Z_4;
    wire shift_srl_26Z0Z_10;
    wire shift_srl_26Z0Z_11;
    wire shift_srl_26Z0Z_12;
    wire shift_srl_26Z0Z_13;
    wire shift_srl_26Z0Z_14;
    wire shift_srl_26Z0Z_9;
    wire shift_srl_26Z0Z_7;
    wire shift_srl_26Z0Z_8;
    wire clk_en_26;
    wire shift_srl_28Z0Z_0;
    wire shift_srl_28Z0Z_10;
    wire shift_srl_28Z0Z_9;
    wire shift_srl_28Z0Z_1;
    wire shift_srl_28Z0Z_2;
    wire shift_srl_28Z0Z_3;
    wire shift_srl_28Z0Z_11;
    wire shift_srl_28Z0Z_8;
    wire shift_srl_28Z0Z_12;
    wire shift_srl_28Z0Z_13;
    wire shift_srl_28Z0Z_14;
    wire shift_srl_28Z0Z_4;
    wire shift_srl_28Z0Z_5;
    wire shift_srl_28Z0Z_6;
    wire shift_srl_28Z0Z_7;
    wire shift_srl_117Z0Z_7;
    wire shift_srl_117Z0Z_8;
    wire shift_srl_117Z0Z_9;
    wire clk_en_117;
    wire rco_int_0_a3_0_a2_138_m6_0_a2_7;
    wire rco_int_0_a2_0_a2_out_5;
    wire shift_srl_140Z0Z_15;
    wire shift_srl_139Z0Z_14;
    wire shift_srl_139Z0Z_12;
    wire shift_srl_139Z0Z_13;
    wire clk_en_139;
    wire shift_srl_162Z0Z_10;
    wire shift_srl_162Z0Z_6;
    wire shift_srl_162Z0Z_14;
    wire shift_srl_162Z0Z_9;
    wire shift_srl_162Z0Z_7;
    wire shift_srl_162Z0Z_8;
    wire shift_srl_120Z0Z_6;
    wire shift_srl_120Z0Z_7;
    wire shift_srl_120Z0Z_5;
    wire shift_srl_120Z0Z_3;
    wire shift_srl_120Z0Z_4;
    wire rco_c_119;
    wire shift_srl_120Z0Z_0;
    wire shift_srl_120Z0Z_1;
    wire shift_srl_120Z0Z_2;
    wire clk_en_120;
    wire shift_srl_127Z0Z_10;
    wire shift_srl_127Z0Z_11;
    wire shift_srl_127Z0Z_12;
    wire shift_srl_127Z0Z_13;
    wire shift_srl_127Z0Z_14;
    wire shift_srl_127Z0Z_9;
    wire shift_srl_127Z0Z_8;
    wire rco_int_0_a2_1_a2_0_127;
    wire shift_srl_120Z0Z_15;
    wire rco_int_0_a2_1_a2_0_120;
    wire shift_srl_124Z0Z_15;
    wire rco_int_0_a2_1_a2_0_120_cascade_;
    wire rco_int_0_a2_1_a2_0_123;
    wire shift_srl_126Z0Z_15;
    wire shift_srl_125Z0Z_15;
    wire clk_en_0_a3_0_a2_1_127_cascade_;
    wire rco_c_118;
    wire shift_srl_119Z0Z_14;
    wire clk_en_0_a3_0_a2_sx_119;
    wire rco_int_0_a2_1_a2_0_0_116;
    wire shift_srl_119Z0Z_15;
    wire shift_srl_119Z0Z_0;
    wire shift_srl_119Z0Z_1;
    wire shift_srl_119Z0Z_2;
    wire shift_srl_119Z0Z_3;
    wire shift_srl_119Z0Z_10;
    wire shift_srl_119Z0Z_13;
    wire shift_srl_119Z0Z_9;
    wire shift_srl_119Z0Z_8;
    wire shift_srl_119Z0Z_4;
    wire shift_srl_40Z0Z_8;
    wire shift_srl_40Z0Z_7;
    wire rco_c_116;
    wire shift_srl_117Z0Z_15;
    wire rco_c_117;
    wire rco_c_132;
    wire shift_srl_133Z0Z_15;
    wire rco_c_133;
    wire rco_c_58;
    wire rco_c_85;
    wire shift_srl_92Z0Z_10;
    wire shift_srl_92Z0Z_11;
    wire shift_srl_92Z0Z_12;
    wire shift_srl_92Z0Z_13;
    wire shift_srl_92Z0Z_14;
    wire shift_srl_92Z0Z_9;
    wire shift_srl_94Z0Z_8;
    wire shift_srl_94Z0Z_9;
    wire shift_srl_94Z0Z_7;
    wire shift_srl_94Z0Z_6;
    wire shift_srl_94Z0Z_5;
    wire shift_srl_141_RNI9SAMZ0Z_15;
    wire rco_c_141;
    wire shift_srl_144_RNIIPPI1Z0Z_15;
    wire rco_c_144;
    wire shift_srl_146_RNIVSUTZ0Z_15;
    wire rco_c_150;
    wire rco_c_173;
    wire rco_c_176;
    wire rco_c_179;
    wire rco_c_182;
    wire shift_srl_95Z0Z_10;
    wire shift_srl_95Z0Z_11;
    wire shift_srl_95Z0Z_12;
    wire shift_srl_95Z0Z_9;
    wire shift_srl_95Z0Z_8;
    wire shift_srl_95Z0Z_0;
    wire shift_srl_95Z0Z_1;
    wire shift_srl_95Z0Z_2;
    wire shift_srl_95Z0Z_3;
    wire shift_srl_95Z0Z_4;
    wire shift_srl_95Z0Z_5;
    wire shift_srl_95Z0Z_6;
    wire shift_srl_95Z0Z_7;
    wire shift_srl_86Z0Z_14;
    wire clk_en_86;
    wire shift_srl_86Z0Z_15;
    wire shift_srl_87Z0Z_15;
    wire shift_srl_85Z0Z_15;
    wire shift_srl_89Z0Z_15;
    wire rco_int_0_a2_0_a2_0_sx_89_cascade_;
    wire shift_srl_88Z0Z_15;
    wire shift_srl_91Z0Z_15;
    wire shift_srl_90Z0Z_15;
    wire shift_srl_89_RNIPCQF1Z0Z_15_cascade_;
    wire shift_srl_91_RNIOVG12Z0Z_15_cascade_;
    wire rco_c_93_cascade_;
    wire rco_c_40;
    wire clk_en_42;
    wire rco_c_39_cascade_;
    wire clk_en_40;
    wire rco_c_39;
    wire clk_en_0_a3_0_a2_sx_98_cascade_;
    wire rco_c_97;
    wire shift_srl_45Z0Z_0;
    wire shift_srl_45Z0Z_1;
    wire shift_srl_45Z0Z_2;
    wire shift_srl_45Z0Z_3;
    wire shift_srl_45Z0Z_4;
    wire shift_srl_45Z0Z_5;
    wire shift_srl_45Z0Z_6;
    wire rco_int_0_a2_0_a2_83_m6_0_a2_sx;
    wire shift_srl_59Z0Z_14;
    wire shift_srl_59Z0Z_13;
    wire shift_srl_59Z0Z_12;
    wire shift_srl_59Z0Z_11;
    wire shift_srl_59Z0Z_10;
    wire shift_srl_59Z0Z_8;
    wire shift_srl_59Z0Z_9;
    wire shift_srl_98Z0Z_0;
    wire shift_srl_98Z0Z_1;
    wire shift_srl_98Z0Z_2;
    wire shift_srl_98Z0Z_3;
    wire shift_srl_98Z0Z_4;
    wire shift_srl_98Z0Z_5;
    wire shift_srl_98Z0Z_6;
    wire shift_srl_98Z0Z_10;
    wire shift_srl_98Z0Z_11;
    wire shift_srl_98Z0Z_12;
    wire shift_srl_98Z0Z_13;
    wire shift_srl_98Z0Z_14;
    wire shift_srl_98Z0Z_9;
    wire shift_srl_98Z0Z_7;
    wire shift_srl_98Z0Z_8;
    wire clk_en_98;
    wire shift_srl_99Z0Z_14;
    wire shift_srl_99Z0Z_15;
    wire shift_srl_99Z0Z_0;
    wire shift_srl_99Z0Z_1;
    wire shift_srl_99Z0Z_2;
    wire shift_srl_99Z0Z_3;
    wire shift_srl_99Z0Z_4;
    wire shift_srl_99Z0Z_5;
    wire clk_en_99;
    wire shift_srl_29Z0Z_2;
    wire shift_srl_29Z0Z_3;
    wire shift_srl_29Z0Z_4;
    wire shift_srl_29Z0Z_5;
    wire shift_srl_29Z0Z_6;
    wire shift_srl_29Z0Z_7;
    wire shift_srl_29Z0Z_8;
    wire rco_c_27;
    wire rco_c_27_cascade_;
    wire clk_en_28;
    wire rco_int_0_a2_0_a2_out_1;
    wire rco_c_28;
    wire rco_c_28_cascade_;
    wire shift_srl_27_RNIP5TNZ0Z_15_cascade_;
    wire rco_int_0_a2_0_a2_out_2_cascade_;
    wire shift_srl_29Z0Z_9;
    wire shift_srl_29Z0Z_10;
    wire shift_srl_29Z0Z_11;
    wire shift_srl_29Z0Z_12;
    wire shift_srl_29Z0Z_1;
    wire shift_srl_29Z0Z_0;
    wire shift_srl_29Z0Z_13;
    wire shift_srl_29Z0Z_14;
    wire clk_en_29;
    wire shift_srl_38Z0Z_13;
    wire shift_srl_158Z0Z_0;
    wire shift_srl_158Z0Z_1;
    wire shift_srl_158Z0Z_2;
    wire shift_srl_158Z0Z_3;
    wire shift_srl_158Z0Z_4;
    wire shift_srl_158Z0Z_5;
    wire shift_srl_158Z0Z_6;
    wire shift_srl_162Z0Z_0;
    wire shift_srl_162Z0Z_1;
    wire shift_srl_162Z0Z_2;
    wire shift_srl_162Z0Z_3;
    wire shift_srl_162Z0Z_4;
    wire shift_srl_162Z0Z_5;
    wire shift_srl_162Z0Z_11;
    wire shift_srl_162Z0Z_12;
    wire shift_srl_162Z0Z_13;
    wire shift_srl_156Z0Z_0;
    wire shift_srl_156Z0Z_1;
    wire shift_srl_156Z0Z_2;
    wire shift_srl_156Z0Z_3;
    wire shift_srl_156Z0Z_4;
    wire shift_srl_156Z0Z_5;
    wire shift_srl_156Z0Z_6;
    wire shift_srl_187Z0Z_0;
    wire shift_srl_187Z0Z_1;
    wire shift_srl_187Z0Z_2;
    wire shift_srl_187Z0Z_3;
    wire shift_srl_187Z0Z_4;
    wire shift_srl_187Z0Z_5;
    wire shift_srl_187Z0Z_6;
    wire shift_srl_111Z0Z_10;
    wire shift_srl_111Z0Z_11;
    wire shift_srl_111Z0Z_12;
    wire shift_srl_111Z0Z_9;
    wire shift_srl_111Z0Z_7;
    wire shift_srl_111Z0Z_8;
    wire clk_en_111;
    wire shift_srl_127Z0Z_15;
    wire shift_srl_127Z0Z_0;
    wire shift_srl_127Z0Z_1;
    wire shift_srl_127Z0Z_2;
    wire shift_srl_127Z0Z_3;
    wire shift_srl_127Z0Z_4;
    wire shift_srl_127Z0Z_5;
    wire shift_srl_127Z0Z_6;
    wire shift_srl_127Z0Z_7;
    wire clk_en_127;
    wire shift_srl_173Z0Z_0;
    wire shift_srl_173Z0Z_1;
    wire shift_srl_173Z0Z_2;
    wire shift_srl_173Z0Z_3;
    wire shift_srl_173Z0Z_4;
    wire shift_srl_173Z0Z_5;
    wire shift_srl_173Z0Z_6;
    wire shift_srl_119Z0Z_7;
    wire shift_srl_119Z0Z_5;
    wire shift_srl_119Z0Z_6;
    wire shift_srl_119Z0Z_11;
    wire shift_srl_119Z0Z_12;
    wire clk_en_119;
    wire shift_srl_40Z0Z_0;
    wire shift_srl_40Z0Z_1;
    wire shift_srl_40Z0Z_2;
    wire shift_srl_40Z0Z_3;
    wire shift_srl_40Z0Z_4;
    wire shift_srl_40Z0Z_5;
    wire shift_srl_40Z0Z_6;
    wire rco_c_54;
    wire shift_srl_198Z0Z_6;
    wire shift_srl_93Z0Z_0;
    wire shift_srl_93Z0Z_1;
    wire shift_srl_93Z0Z_2;
    wire shift_srl_93Z0Z_3;
    wire shift_srl_93Z0Z_4;
    wire shift_srl_93Z0Z_5;
    wire shift_srl_84Z0Z_15;
    wire rco_c_84;
    wire shift_srl_89_RNIPCQF1Z0Z_15;
    wire rco_c_89;
    wire shift_srl_91_RNIOVG12Z0Z_15;
    wire rco_c_83;
    wire rco_c_92;
    wire shift_srl_92Z0Z_15;
    wire shift_srl_93Z0Z_10;
    wire shift_srl_93Z0Z_11;
    wire shift_srl_93Z0Z_12;
    wire shift_srl_93Z0Z_13;
    wire shift_srl_93Z0Z_14;
    wire shift_srl_93Z0Z_9;
    wire shift_srl_46Z0Z_0;
    wire shift_srl_46Z0Z_3;
    wire shift_srl_46Z0Z_8;
    wire shift_srl_46Z0Z_9;
    wire shift_srl_46Z0Z_1;
    wire shift_srl_46Z0Z_2;
    wire shift_srl_97Z0Z_10;
    wire shift_srl_97Z0Z_11;
    wire shift_srl_97Z0Z_12;
    wire shift_srl_97Z0Z_13;
    wire shift_srl_97Z0Z_14;
    wire shift_srl_97Z0Z_9;
    wire shift_srl_97Z0Z_8;
    wire shift_srl_95_RNIHJ49Z0Z_15_cascade_;
    wire rco_c_96;
    wire shift_srl_94Z0Z_14;
    wire shift_srl_94Z0Z_13;
    wire shift_srl_94Z0Z_12;
    wire shift_srl_94Z0Z_10;
    wire shift_srl_94Z0Z_11;
    wire shift_srl_96Z0Z_1;
    wire shift_srl_96Z0Z_2;
    wire shift_srl_96Z0Z_3;
    wire shift_srl_96Z0Z_0;
    wire shift_srl_96Z0Z_10;
    wire shift_srl_96Z0Z_11;
    wire shift_srl_96Z0Z_6;
    wire shift_srl_96Z0Z_4;
    wire shift_srl_96Z0Z_5;
    wire shift_srl_96Z0Z_12;
    wire shift_srl_96Z0Z_13;
    wire shift_srl_96Z0Z_14;
    wire shift_srl_96Z0Z_9;
    wire shift_srl_96Z0Z_7;
    wire shift_srl_96Z0Z_8;
    wire clk_en_96;
    wire shift_srl_45Z0Z_10;
    wire shift_srl_45Z0Z_11;
    wire shift_srl_45Z0Z_12;
    wire shift_srl_45Z0Z_13;
    wire shift_srl_45Z0Z_14;
    wire shift_srl_45Z0Z_9;
    wire shift_srl_45Z0Z_7;
    wire shift_srl_45Z0Z_8;
    wire clk_en_43;
    wire N_4016_i_0_a2_1;
    wire rco_int_0_a2_21_m6_0_a2_s_7;
    wire rco_int_0_a2_21_m6_0_a2_s_8;
    wire shift_srl_23_RNI0DK37Z0Z_15_cascade_;
    wire rco_c_9;
    wire rco_c_41_cascade_;
    wire rco_c_41;
    wire clk_en_45;
    wire shift_srl_44Z0Z_0;
    wire shift_srl_44Z0Z_1;
    wire shift_srl_44Z0Z_2;
    wire shift_srl_44Z0Z_3;
    wire shift_srl_44Z0Z_4;
    wire shift_srl_44Z0Z_5;
    wire shift_srl_44Z0Z_6;
    wire shift_srl_48Z0Z_0;
    wire shift_srl_48Z0Z_1;
    wire shift_srl_48Z0Z_2;
    wire shift_srl_48Z0Z_3;
    wire shift_srl_48Z0Z_4;
    wire shift_srl_48Z0Z_5;
    wire shift_srl_94_RNI2F961Z0Z_15_cascade_;
    wire shift_srl_96Z0Z_15;
    wire shift_srl_98Z0Z_15;
    wire shift_srl_98_RNIA7Q31Z0Z_15;
    wire rco_int_0_a2_0_a2_99_m6_0_a2_1;
    wire rco_int_0_a2_0_a2_99_m6_0_a2_9_1_cascade_;
    wire rco_int_0_a2_0_a2_99_m6_0_a2_9_sx;
    wire shift_srl_95Z0Z_15;
    wire rco_c_34;
    wire shift_srl_95Z0Z_13;
    wire shift_srl_95Z0Z_14;
    wire clk_en_95;
    wire shift_srl_93Z0Z_15;
    wire shift_srl_40_fastZ0Z_15;
    wire shift_srl_40Z0Z_14;
    wire shift_srl_40Z0Z_13;
    wire shift_srl_40Z0Z_12;
    wire shift_srl_40Z0Z_11;
    wire shift_srl_40Z0Z_9;
    wire shift_srl_40Z0Z_10;
    wire clk_en_g_40;
    wire rco_int_0_a2_0_a2_out_2;
    wire rco_c_30;
    wire shift_srl_30Z0Z_0;
    wire shift_srl_30Z0Z_1;
    wire shift_srl_30Z0Z_2;
    wire shift_srl_30Z0Z_3;
    wire shift_srl_30Z0Z_4;
    wire shift_srl_30Z0Z_5;
    wire shift_srl_38Z0Z_0;
    wire shift_srl_38Z0Z_1;
    wire shift_srl_38Z0Z_2;
    wire shift_srl_38Z0Z_3;
    wire shift_srl_38Z0Z_4;
    wire shift_srl_38Z0Z_5;
    wire shift_srl_38Z0Z_6;
    wire shift_srl_38Z0Z_10;
    wire shift_srl_38Z0Z_11;
    wire shift_srl_38Z0Z_12;
    wire shift_srl_38Z0Z_14;
    wire shift_srl_38Z0Z_9;
    wire shift_srl_38Z0Z_7;
    wire shift_srl_38Z0Z_8;
    wire clk_en_38;
    wire shift_srl_158Z0Z_10;
    wire shift_srl_158Z0Z_11;
    wire shift_srl_158Z0Z_12;
    wire shift_srl_158Z0Z_13;
    wire shift_srl_158Z0Z_14;
    wire shift_srl_158Z0Z_9;
    wire shift_srl_158Z0Z_7;
    wire shift_srl_158Z0Z_8;
    wire rco_c_158;
    wire rco_c_157;
    wire rco_int_0_a2_0_a2_sx_1_153;
    wire rco_c_153_cascade_;
    wire clk_en_162;
    wire shift_srl_160_RNIFA2R1Z0Z_15;
    wire clk_en_158;
    wire shift_srl_156Z0Z_10;
    wire shift_srl_156Z0Z_11;
    wire shift_srl_156Z0Z_12;
    wire shift_srl_156Z0Z_13;
    wire shift_srl_156Z0Z_14;
    wire shift_srl_156Z0Z_9;
    wire shift_srl_156Z0Z_7;
    wire shift_srl_156Z0Z_8;
    wire clk_en_156;
    wire g0_15;
    wire rco_int_0_a3_0_a2_0_183_cascade_;
    wire clk_en_0_a2_0_a2_1_187_cascade_;
    wire clk_en_0_a2_0_a2_sx_187;
    wire shift_srl_183Z0Z_15;
    wire shift_srl_183Z0Z_0;
    wire shift_srl_187Z0Z_10;
    wire shift_srl_187Z0Z_11;
    wire shift_srl_187Z0Z_12;
    wire shift_srl_187Z0Z_13;
    wire shift_srl_187Z0Z_14;
    wire shift_srl_187Z0Z_9;
    wire shift_srl_187Z0Z_7;
    wire shift_srl_187Z0Z_8;
    wire clk_en_187;
    wire shift_srl_194Z0Z_10;
    wire shift_srl_194Z0Z_11;
    wire shift_srl_194Z0Z_12;
    wire shift_srl_194Z0Z_13;
    wire shift_srl_194Z0Z_14;
    wire shift_srl_194Z0Z_9;
    wire shift_srl_194Z0Z_1;
    wire shift_srl_194Z0Z_2;
    wire shift_srl_194Z0Z_3;
    wire shift_srl_194Z0Z_4;
    wire shift_srl_194Z0Z_5;
    wire shift_srl_194Z0Z_6;
    wire shift_srl_194Z0Z_7;
    wire shift_srl_194Z0Z_8;
    wire shift_srl_175Z0Z_0;
    wire shift_srl_175Z0Z_1;
    wire shift_srl_175Z0Z_2;
    wire shift_srl_175Z0Z_3;
    wire shift_srl_175Z0Z_4;
    wire shift_srl_175Z0Z_5;
    wire shift_srl_175Z0Z_6;
    wire shift_srl_198Z0Z_10;
    wire shift_srl_198Z0Z_11;
    wire shift_srl_198Z0Z_12;
    wire shift_srl_198Z0Z_13;
    wire shift_srl_198Z0Z_14;
    wire shift_srl_198Z0Z_9;
    wire shift_srl_198Z0Z_7;
    wire shift_srl_198Z0Z_8;
    wire rco_c_197;
    wire rco_c_197_cascade_;
    wire rco_c_198;
    wire shift_srl_198Z0Z_15;
    wire shift_srl_198Z0Z_0;
    wire shift_srl_198Z0Z_1;
    wire shift_srl_198Z0Z_2;
    wire shift_srl_198Z0Z_3;
    wire shift_srl_198Z0Z_4;
    wire shift_srl_198Z0Z_5;
    wire shift_srl_197Z0Z_2;
    wire shift_srl_197Z0Z_3;
    wire shift_srl_197Z0Z_4;
    wire shift_srl_197Z0Z_5;
    wire shift_srl_197Z0Z_6;
    wire shift_srl_197Z0Z_0;
    wire shift_srl_197Z0Z_1;
    wire shift_srl_197Z0Z_10;
    wire shift_srl_197Z0Z_11;
    wire shift_srl_197Z0Z_12;
    wire shift_srl_197Z0Z_13;
    wire shift_srl_197Z0Z_14;
    wire shift_srl_197Z0Z_15;
    wire shift_srl_197Z0Z_9;
    wire shift_srl_197Z0Z_7;
    wire shift_srl_197Z0Z_8;
    wire shift_srl_93Z0Z_8;
    wire shift_srl_93Z0Z_6;
    wire shift_srl_93Z0Z_7;
    wire clk_en_93;
    wire shift_srl_92Z0Z_0;
    wire shift_srl_92Z0Z_1;
    wire shift_srl_92Z0Z_2;
    wire shift_srl_92Z0Z_3;
    wire shift_srl_92Z0Z_4;
    wire shift_srl_92Z0Z_5;
    wire shift_srl_92Z0Z_6;
    wire shift_srl_92Z0Z_7;
    wire shift_srl_92Z0Z_8;
    wire clk_en_92;
    wire shift_srl_146Z0Z_15;
    wire rco_c_146;
    wire shift_srl_46Z0Z_7;
    wire shift_srl_46Z0Z_10;
    wire shift_srl_46Z0Z_11;
    wire shift_srl_46Z0Z_12;
    wire shift_srl_46Z0Z_13;
    wire shift_srl_46Z0Z_14;
    wire shift_srl_46Z0Z_6;
    wire shift_srl_46Z0Z_4;
    wire shift_srl_46Z0Z_5;
    wire clk_en_46;
    wire shift_srl_97Z0Z_15;
    wire shift_srl_97Z0Z_0;
    wire shift_srl_97Z0Z_1;
    wire shift_srl_97Z0Z_2;
    wire shift_srl_97Z0Z_3;
    wire shift_srl_97Z0Z_4;
    wire shift_srl_97Z0Z_5;
    wire shift_srl_97Z0Z_6;
    wire shift_srl_97Z0Z_7;
    wire clk_en_97;
    wire shift_srl_51Z0Z_10;
    wire shift_srl_51Z0Z_11;
    wire shift_srl_51Z0Z_12;
    wire shift_srl_51Z0Z_13;
    wire shift_srl_51Z0Z_14;
    wire shift_srl_51Z0Z_6;
    wire shift_srl_53Z0Z_0;
    wire shift_srl_53Z0Z_1;
    wire shift_srl_53Z0Z_2;
    wire shift_srl_53Z0Z_3;
    wire shift_srl_53Z0Z_4;
    wire shift_srl_53Z0Z_5;
    wire shift_srl_53Z0Z_6;
    wire shift_srl_53Z0Z_10;
    wire shift_srl_53Z0Z_11;
    wire shift_srl_53Z0Z_12;
    wire shift_srl_53Z0Z_13;
    wire shift_srl_53Z0Z_14;
    wire shift_srl_53Z0Z_9;
    wire shift_srl_53Z0Z_7;
    wire shift_srl_53Z0Z_8;
    wire shift_srl_41Z0Z_10;
    wire shift_srl_41Z0Z_11;
    wire shift_srl_41Z0Z_12;
    wire shift_srl_41Z0Z_13;
    wire shift_srl_41Z0Z_14;
    wire shift_srl_41Z0Z_9;
    wire shift_srl_41Z0Z_8;
    wire shift_srl_59Z0Z_0;
    wire shift_srl_59Z0Z_1;
    wire shift_srl_59Z0Z_2;
    wire shift_srl_59Z0Z_3;
    wire shift_srl_59Z0Z_4;
    wire shift_srl_59Z0Z_5;
    wire shift_srl_59Z0Z_6;
    wire shift_srl_59Z0Z_7;
    wire shift_srl_44Z0Z_10;
    wire shift_srl_44Z0Z_11;
    wire shift_srl_44Z0Z_12;
    wire shift_srl_44Z0Z_13;
    wire shift_srl_44Z0Z_14;
    wire shift_srl_44Z0Z_9;
    wire shift_srl_44Z0Z_7;
    wire shift_srl_44Z0Z_8;
    wire clk_en_44;
    wire shift_srl_48Z0Z_10;
    wire shift_srl_48Z0Z_9;
    wire shift_srl_48Z0Z_8;
    wire shift_srl_48Z0Z_6;
    wire shift_srl_48Z0Z_7;
    wire shift_srl_39_RNIG4I71Z0Z_15;
    wire shift_srl_39Z0Z_14;
    wire shift_srl_39Z0Z_13;
    wire shift_srl_39Z0Z_12;
    wire shift_srl_39Z0Z_11;
    wire shift_srl_39Z0Z_10;
    wire shift_srl_39Z0Z_9;
    wire shift_srl_61Z0Z_1;
    wire shift_srl_61Z0Z_2;
    wire shift_srl_61Z0Z_3;
    wire shift_srl_61Z0Z_4;
    wire shift_srl_61Z0Z_5;
    wire shift_srl_61Z0Z_6;
    wire shift_srl_61Z0Z_7;
    wire rco_int_0_a2_0_a2_s_0_0_35_cascade_;
    wire shift_srl_31_RNI84161_0Z0Z_15;
    wire shift_srl_37_RNI973EZ0Z_15;
    wire rco_int_0_a2_0_a2_99_m6_0_a2_2;
    wire shift_srl_26Z0Z_15;
    wire shift_srl_25Z0Z_15;
    wire shift_srl_27Z0Z_15;
    wire shift_srl_27_RNIAA521_0Z0Z_15;
    wire rco_int_0_a2_0_a2_99_m6_0_a2_3;
    wire shift_srl_62Z0Z_0;
    wire shift_srl_62Z0Z_1;
    wire shift_srl_62Z0Z_2;
    wire shift_srl_62Z0Z_3;
    wire shift_srl_62Z0Z_4;
    wire shift_srl_62Z0Z_5;
    wire shift_srl_62Z0Z_6;
    wire shift_srl_174Z0Z_0;
    wire shift_srl_174Z0Z_1;
    wire shift_srl_174Z0Z_2;
    wire shift_srl_174Z0Z_3;
    wire shift_srl_174Z0Z_4;
    wire shift_srl_174Z0Z_5;
    wire shift_srl_174Z0Z_6;
    wire rco_c_166;
    wire shift_srl_159_RNIDDRE1Z0Z_15;
    wire rco_c_162_cascade_;
    wire shift_srl_184Z0Z_0;
    wire shift_srl_184Z0Z_1;
    wire shift_srl_184Z0Z_2;
    wire shift_srl_184Z0Z_3;
    wire shift_srl_184Z0Z_4;
    wire shift_srl_184Z0Z_5;
    wire shift_srl_184Z0Z_6;
    wire shift_srl_183Z0Z_10;
    wire shift_srl_183Z0Z_11;
    wire shift_srl_183Z0Z_12;
    wire shift_srl_183Z0Z_13;
    wire shift_srl_183Z0Z_14;
    wire shift_srl_183Z0Z_9;
    wire shift_srl_183Z0Z_8;
    wire shift_srl_183Z0Z_7;
    wire shift_srl_183Z0Z_1;
    wire shift_srl_183Z0Z_2;
    wire shift_srl_183Z0Z_3;
    wire shift_srl_183Z0Z_4;
    wire shift_srl_183Z0Z_5;
    wire shift_srl_183Z0Z_6;
    wire clk_en_183;
    wire rco_c_181;
    wire rco_c_180;
    wire clk_en_0_a3_0_a2_sx_182_cascade_;
    wire shift_srl_91_RNI20EN1Z0Z_15;
    wire rco_int_0_a2_0_a2_99_m6_0_a2_9;
    wire shift_srl_145_RNIN9307Z0Z_15;
    wire rco_int_0_a2_0_a2_1_1_145;
    wire rco_int_0_a3_0_a2_sx_183_cascade_;
    wire shift_srl_195Z0Z_10;
    wire shift_srl_195Z0Z_11;
    wire shift_srl_195Z0Z_12;
    wire shift_srl_195Z0Z_13;
    wire shift_srl_195Z0Z_14;
    wire shift_srl_195Z0Z_9;
    wire shift_srl_195Z0Z_8;
    wire shift_srl_185Z0Z_0;
    wire shift_srl_185Z0Z_1;
    wire shift_srl_185Z0Z_2;
    wire shift_srl_185Z0Z_3;
    wire shift_srl_185Z0Z_4;
    wire shift_srl_185Z0Z_5;
    wire shift_srl_185Z0Z_6;
    wire clk_en_194;
    wire N_4183;
    wire clk_en_198;
    wire rco_c_172_cascade_;
    wire shift_srl_196Z0Z_0;
    wire shift_srl_196Z0Z_1;
    wire shift_srl_196Z0Z_2;
    wire shift_srl_196Z0Z_3;
    wire shift_srl_196Z0Z_4;
    wire shift_srl_196Z0Z_5;
    wire shift_srl_196Z0Z_6;
    wire shift_srl_196Z0Z_7;
    wire shift_srl_196Z0Z_8;
    wire shift_srl_196Z0Z_9;
    wire clk_en_197;
    wire shift_srl_196Z0Z_15;
    wire rco_c_196;
    wire shift_srl_196Z0Z_14;
    wire shift_srl_196Z0Z_13;
    wire shift_srl_196Z0Z_12;
    wire shift_srl_196Z0Z_10;
    wire shift_srl_196Z0Z_11;
    wire clk_en_196;
    wire shift_srl_182Z0Z_10;
    wire shift_srl_182Z0Z_11;
    wire shift_srl_182Z0Z_12;
    wire shift_srl_182Z0Z_13;
    wire shift_srl_182Z0Z_14;
    wire shift_srl_182Z0Z_9;
    wire shift_srl_182Z0Z_8;
    wire shift_srl_182Z0Z_0;
    wire shift_srl_182Z0Z_1;
    wire shift_srl_182Z0Z_2;
    wire shift_srl_182Z0Z_3;
    wire shift_srl_182Z0Z_4;
    wire shift_srl_182Z0Z_5;
    wire shift_srl_182Z0Z_6;
    wire shift_srl_182Z0Z_7;
    wire clk_en_182;
    wire rco_c_94;
    wire shift_srl_95_RNIHJ49Z0Z_15;
    wire rco_c_95;
    wire shift_srl_94_RNI2F961Z0Z_15;
    wire rco_c_93;
    wire rco_c_98;
    wire shift_srl_94Z0Z_15;
    wire shift_srl_94Z0Z_0;
    wire shift_srl_94Z0Z_1;
    wire shift_srl_94Z0Z_2;
    wire shift_srl_94Z0Z_3;
    wire shift_srl_94Z0Z_4;
    wire clk_en_94;
    wire shift_srl_49Z0Z_9;
    wire shift_srl_49Z0Z_8;
    wire shift_srl_49Z0Z_7;
    wire shift_srl_51Z0Z_0;
    wire shift_srl_51Z0Z_1;
    wire shift_srl_51Z0Z_2;
    wire shift_srl_51Z0Z_3;
    wire shift_srl_51Z0Z_4;
    wire shift_srl_51Z0Z_5;
    wire shift_srl_51Z0Z_7;
    wire shift_srl_51Z0Z_8;
    wire shift_srl_51Z0Z_9;
    wire clk_en_53;
    wire shift_srl_50_RNI869CZ0Z_15_cascade_;
    wire clk_en_51;
    wire shift_srl_49Z0Z_14;
    wire shift_srl_49Z0Z_13;
    wire shift_srl_49Z0Z_12;
    wire shift_srl_49Z0Z_10;
    wire shift_srl_49Z0Z_11;
    wire rco_int_0_a2_0_a2_0_39_cascade_;
    wire rco_int_0_a2_0_a2_83_m6_0_a2_3_sx_cascade_;
    wire rco_int_0_a2_0_a2_83_m6_0_a2_3;
    wire shift_srl_53Z0Z_15;
    wire shift_srl_53_RNI66TQZ0Z_15_cascade_;
    wire shift_srl_56Z0Z_10;
    wire shift_srl_56Z0Z_11;
    wire shift_srl_56Z0Z_12;
    wire shift_srl_56Z0Z_13;
    wire shift_srl_56Z0Z_14;
    wire shift_srl_56Z0Z_9;
    wire shift_srl_58_RNIQMNUZ0Z_15_cascade_;
    wire shift_srl_54_RNIEAU71Z0Z_15_cascade_;
    wire clk_en_59;
    wire shift_srl_55Z0Z_14;
    wire shift_srl_55Z0Z_13;
    wire shift_srl_55Z0Z_12;
    wire shift_srl_55Z0Z_11;
    wire shift_srl_55Z0Z_0;
    wire shift_srl_55Z0Z_1;
    wire shift_srl_55Z0Z_2;
    wire shift_srl_55Z0Z_3;
    wire shift_srl_55Z0Z_4;
    wire shift_srl_55Z0Z_5;
    wire shift_srl_55Z0Z_6;
    wire shift_srl_44Z0Z_15;
    wire shift_srl_43Z0Z_15;
    wire shift_srl_42Z0Z_15;
    wire rco_int_0_a2_1_a2_0_44_cascade_;
    wire shift_srl_48Z0Z_14;
    wire shift_srl_48Z0Z_13;
    wire shift_srl_48Z0Z_11;
    wire shift_srl_48Z0Z_12;
    wire clk_en_48;
    wire shift_srl_55Z0Z_10;
    wire shift_srl_55Z0Z_9;
    wire shift_srl_55Z0Z_7;
    wire shift_srl_55Z0Z_8;
    wire shift_srl_61Z0Z_0;
    wire shift_srl_61Z0Z_12;
    wire shift_srl_61Z0Z_13;
    wire shift_srl_61Z0Z_14;
    wire shift_srl_61Z0Z_10;
    wire shift_srl_61Z0Z_11;
    wire shift_srl_61Z0Z_8;
    wire shift_srl_61Z0Z_9;
    wire shift_srl_61_RNI3LM9Z0Z_15_cascade_;
    wire shift_srl_61Z0Z_15;
    wire shift_srl_62_RNIM5RKZ0Z_15_cascade_;
    wire clk_en_61;
    wire shift_srl_62Z0Z_10;
    wire shift_srl_62Z0Z_11;
    wire shift_srl_62Z0Z_12;
    wire shift_srl_62Z0Z_13;
    wire shift_srl_62Z0Z_14;
    wire shift_srl_62Z0Z_15;
    wire shift_srl_62Z0Z_9;
    wire shift_srl_62Z0Z_7;
    wire shift_srl_62Z0Z_8;
    wire clk_en_62;
    wire shift_srl_174Z0Z_10;
    wire shift_srl_174Z0Z_11;
    wire shift_srl_174Z0Z_12;
    wire shift_srl_174Z0Z_13;
    wire shift_srl_174Z0Z_14;
    wire shift_srl_174Z0Z_9;
    wire shift_srl_174Z0Z_7;
    wire shift_srl_174Z0Z_8;
    wire clk_en_174;
    wire shift_srl_166Z0Z_1;
    wire shift_srl_166Z0Z_2;
    wire shift_srl_166Z0Z_3;
    wire shift_srl_166Z0Z_4;
    wire shift_srl_166Z0Z_5;
    wire shift_srl_166Z0Z_6;
    wire shift_srl_166Z0Z_7;
    wire shift_srl_166Z0Z_10;
    wire shift_srl_166Z0Z_11;
    wire shift_srl_166Z0Z_12;
    wire shift_srl_166Z0Z_13;
    wire shift_srl_166Z0Z_14;
    wire shift_srl_166Z0Z_8;
    wire shift_srl_166Z0Z_9;
    wire shift_srl_166Z0Z_0;
    wire clk_en_166;
    wire shift_srl_184Z0Z_10;
    wire shift_srl_184Z0Z_11;
    wire shift_srl_184Z0Z_12;
    wire shift_srl_184Z0Z_13;
    wire shift_srl_184Z0Z_9;
    wire shift_srl_184Z0Z_7;
    wire shift_srl_184Z0Z_8;
    wire shift_srl_186Z0Z_0;
    wire shift_srl_186Z0Z_1;
    wire shift_srl_186Z0Z_2;
    wire shift_srl_186Z0Z_3;
    wire shift_srl_186Z0Z_4;
    wire shift_srl_186Z0Z_5;
    wire shift_srl_186Z0Z_6;
    wire shift_srl_184Z0Z_14;
    wire clk_en_184;
    wire clk_en_0_a2_0_a2_0_sx_192_cascade_;
    wire N_4179_cascade_;
    wire shift_srl_194Z0Z_15;
    wire N_4179;
    wire N_4181;
    wire clk_en_0_a2_0_a2_0_sx_192;
    wire shift_srl_195Z0Z_15;
    wire shift_srl_195Z0Z_0;
    wire shift_srl_195Z0Z_1;
    wire shift_srl_195Z0Z_2;
    wire shift_srl_195Z0Z_3;
    wire shift_srl_195Z0Z_4;
    wire shift_srl_195Z0Z_5;
    wire shift_srl_195Z0Z_6;
    wire shift_srl_195Z0Z_7;
    wire clk_en_195;
    wire shift_srl_185Z0Z_10;
    wire shift_srl_185Z0Z_11;
    wire shift_srl_185Z0Z_12;
    wire shift_srl_185Z0Z_13;
    wire shift_srl_185Z0Z_14;
    wire shift_srl_185Z0Z_9;
    wire shift_srl_185Z0Z_7;
    wire shift_srl_185Z0Z_8;
    wire clk_en_185;
    wire shift_srl_175Z0Z_10;
    wire shift_srl_175Z0Z_11;
    wire shift_srl_175Z0Z_12;
    wire shift_srl_175Z0Z_13;
    wire shift_srl_175Z0Z_14;
    wire shift_srl_175Z0Z_9;
    wire shift_srl_175Z0Z_7;
    wire shift_srl_175Z0Z_8;
    wire clk_en_175;
    wire shift_srl_192Z0Z_0;
    wire shift_srl_192Z0Z_1;
    wire shift_srl_192Z0Z_2;
    wire shift_srl_192Z0Z_3;
    wire shift_srl_192Z0Z_4;
    wire shift_srl_192Z0Z_5;
    wire shift_srl_192Z0Z_6;
    wire N_4177;
    wire shift_srl_192Z0Z_15;
    wire rco_c_192;
    wire shift_srl_192Z0Z_14;
    wire shift_srl_192Z0Z_13;
    wire shift_srl_192Z0Z_12;
    wire shift_srl_192Z0Z_11;
    wire shift_srl_192Z0Z_10;
    wire rco_c_46;
    wire shift_srl_49Z0Z_0;
    wire shift_srl_49Z0Z_1;
    wire shift_srl_49Z0Z_2;
    wire shift_srl_49Z0Z_3;
    wire shift_srl_49Z0Z_4;
    wire shift_srl_49Z0Z_5;
    wire shift_srl_49Z0Z_6;
    wire rco_c_44_cascade_;
    wire rco_int_0_a2_0_a2_0_0_37;
    wire clk_en_0_a3_0_a2_sx_49_cascade_;
    wire clk_en_49;
    wire shift_srl_46Z0Z_15;
    wire shift_srl_47_RNIV3QLZ0Z_15_cascade_;
    wire rco_c_47;
    wire shift_srl_50Z0Z_14;
    wire shift_srl_50Z0Z_11;
    wire shift_srl_50Z0Z_12;
    wire shift_srl_50Z0Z_13;
    wire shift_srl_52Z0Z_10;
    wire shift_srl_52Z0Z_11;
    wire shift_srl_52Z0Z_12;
    wire shift_srl_52Z0Z_13;
    wire shift_srl_52Z0Z_14;
    wire shift_srl_52Z0Z_9;
    wire shift_srl_52Z0Z_8;
    wire rco_c_52;
    wire rco_c_51;
    wire rco_int_0_a2_0_a2_0_39;
    wire shift_srl_40Z0Z_15;
    wire shift_srl_51Z0Z_15;
    wire rco_c_48_cascade_;
    wire clk_en_55;
    wire shift_srl_55Z0Z_15;
    wire shift_srl_54Z0Z_14;
    wire shift_srl_54Z0Z_13;
    wire shift_srl_54Z0Z_12;
    wire shift_srl_54Z0Z_11;
    wire shift_srl_54Z0Z_10;
    wire shift_srl_57Z0Z_10;
    wire shift_srl_57Z0Z_11;
    wire shift_srl_57Z0Z_12;
    wire shift_srl_57Z0Z_13;
    wire shift_srl_57Z0Z_14;
    wire shift_srl_57Z0Z_9;
    wire shift_srl_57Z0Z_8;
    wire shift_srl_60Z0Z_10;
    wire shift_srl_60Z0Z_11;
    wire shift_srl_60Z0Z_12;
    wire shift_srl_60Z0Z_13;
    wire shift_srl_60Z0Z_9;
    wire shift_srl_60Z0Z_8;
    wire shift_srl_60Z0Z_14;
    wire shift_srl_60Z0Z_4;
    wire shift_srl_60Z0Z_5;
    wire shift_srl_60Z0Z_6;
    wire shift_srl_60Z0Z_7;
    wire rco_int_0_a2_0_a2_sx_153;
    wire clk_en_0_a3_0_a2_sx_179_cascade_;
    wire rco_int_0_a2_0_a2_93_m6_0_a2_4_7_0;
    wire rco_int_0_a2_1_a2_0_44;
    wire rco_int_0_a2_0_a2_93_m6_0_a2_4_7_4_sx_cascade_;
    wire rco_int_0_a2_0_a2_93_m6_0_a2_4_7_4_cascade_;
    wire rco_int_0_a2_0_a2_93_m6_0_a2_4_7;
    wire rco_int_0_a3_0_a2_0_0_66;
    wire shift_srl_63Z0Z_0;
    wire shift_srl_63Z0Z_1;
    wire shift_srl_63Z0Z_2;
    wire shift_srl_63Z0Z_3;
    wire shift_srl_63Z0Z_4;
    wire shift_srl_63Z0Z_5;
    wire shift_srl_63Z0Z_6;
    wire rco_c_60;
    wire shift_srl_61_RNI3LM9Z0Z_15;
    wire rco_c_61;
    wire rco_c_62;
    wire rco_c_65;
    wire shift_srl_60Z0Z_15;
    wire shift_srl_60Z0Z_0;
    wire shift_srl_60Z0Z_1;
    wire shift_srl_60Z0Z_2;
    wire shift_srl_60Z0Z_3;
    wire shift_srl_159Z0Z_10;
    wire shift_srl_159Z0Z_9;
    wire shift_srl_159Z0Z_11;
    wire shift_srl_159Z0Z_12;
    wire shift_srl_159Z0Z_5;
    wire shift_srl_159Z0Z_13;
    wire shift_srl_159Z0Z_0;
    wire shift_srl_159Z0Z_6;
    wire shift_srl_159Z0Z_3;
    wire shift_srl_159Z0Z_4;
    wire shift_srl_159Z0Z_7;
    wire shift_srl_159Z0Z_8;
    wire shift_srl_159Z0Z_1;
    wire shift_srl_159Z0Z_2;
    wire shift_srl_171Z0Z_2;
    wire shift_srl_171Z0Z_3;
    wire shift_srl_171Z0Z_4;
    wire shift_srl_171Z0Z_5;
    wire shift_srl_171Z0Z_6;
    wire shift_srl_171Z0Z_7;
    wire shift_srl_179Z0Z_0;
    wire shift_srl_179Z0Z_1;
    wire shift_srl_179Z0Z_2;
    wire shift_srl_179Z0Z_3;
    wire shift_srl_179Z0Z_4;
    wire shift_srl_179Z0Z_5;
    wire shift_srl_179Z0Z_6;
    wire shift_srl_186Z0Z_10;
    wire shift_srl_186Z0Z_11;
    wire shift_srl_186Z0Z_12;
    wire shift_srl_186Z0Z_13;
    wire shift_srl_186Z0Z_14;
    wire shift_srl_186Z0Z_9;
    wire shift_srl_186Z0Z_7;
    wire shift_srl_186Z0Z_8;
    wire clk_en_186;
    wire shift_srl_178Z0Z_0;
    wire shift_srl_178Z0Z_1;
    wire shift_srl_178Z0Z_2;
    wire shift_srl_178Z0Z_3;
    wire shift_srl_178Z0Z_4;
    wire shift_srl_178Z0Z_9;
    wire shift_srl_181Z0Z_1;
    wire shift_srl_181Z0Z_2;
    wire shift_srl_181Z0Z_3;
    wire shift_srl_181Z0Z_4;
    wire shift_srl_181Z0Z_5;
    wire shift_srl_181Z0Z_0;
    wire shift_srl_176Z0Z_10;
    wire shift_srl_176Z0Z_11;
    wire shift_srl_176Z0Z_12;
    wire shift_srl_176Z0Z_13;
    wire shift_srl_176Z0Z_14;
    wire shift_srl_176Z0Z_9;
    wire shift_srl_176Z0Z_8;
    wire rco_c_175;
    wire rco_c_174;
    wire clk_en_0_a3_0_a2cf1_176_cascade_;
    wire shift_srl_175Z0Z_15;
    wire shift_srl_174Z0Z_15;
    wire shift_srl_173Z0Z_15;
    wire shift_srl_182Z0Z_15;
    wire shift_srl_181Z0Z_15;
    wire shift_srl_176_RNIUGI51Z0Z_15_cascade_;
    wire shift_srl_182_RNIEPSC2Z0Z_15;
    wire shift_srl_193Z0Z_10;
    wire shift_srl_193Z0Z_11;
    wire shift_srl_193Z0Z_12;
    wire shift_srl_193Z0Z_13;
    wire shift_srl_193Z0Z_14;
    wire shift_srl_193Z0Z_9;
    wire shift_srl_193Z0Z_8;
    wire shift_srl_193Z0Z_15;
    wire shift_srl_193Z0Z_0;
    wire shift_srl_193Z0Z_1;
    wire shift_srl_193Z0Z_2;
    wire shift_srl_193Z0Z_3;
    wire shift_srl_193Z0Z_4;
    wire shift_srl_193Z0Z_5;
    wire shift_srl_193Z0Z_6;
    wire shift_srl_193Z0Z_7;
    wire clk_en_193;
    wire shift_srl_45Z0Z_15;
    wire rco_c_45;
    wire shift_srl_47Z0Z_0;
    wire shift_srl_47Z0Z_1;
    wire shift_srl_47Z0Z_2;
    wire shift_srl_47Z0Z_3;
    wire shift_srl_47Z0Z_4;
    wire shift_srl_47Z0Z_5;
    wire shift_srl_47Z0Z_15;
    wire shift_srl_47Z0Z_10;
    wire shift_srl_47Z0Z_11;
    wire shift_srl_47Z0Z_12;
    wire shift_srl_47Z0Z_13;
    wire shift_srl_47Z0Z_14;
    wire shift_srl_47Z0Z_6;
    wire shift_srl_47Z0Z_9;
    wire shift_srl_47Z0Z_7;
    wire shift_srl_47Z0Z_8;
    wire clk_en_47;
    wire shift_srl_50Z0Z_10;
    wire shift_srl_50Z0Z_5;
    wire shift_srl_50Z0Z_6;
    wire shift_srl_50Z0Z_9;
    wire shift_srl_50Z0Z_7;
    wire shift_srl_50Z0Z_8;
    wire shift_srl_50Z0Z_15;
    wire shift_srl_50Z0Z_0;
    wire shift_srl_50Z0Z_1;
    wire shift_srl_50Z0Z_2;
    wire shift_srl_50Z0Z_3;
    wire shift_srl_50Z0Z_4;
    wire clk_en_50;
    wire shift_srl_52Z0Z_15;
    wire shift_srl_52Z0Z_0;
    wire shift_srl_52Z0Z_1;
    wire shift_srl_52Z0Z_2;
    wire shift_srl_52Z0Z_3;
    wire shift_srl_52Z0Z_4;
    wire shift_srl_52Z0Z_5;
    wire shift_srl_52Z0Z_6;
    wire shift_srl_52Z0Z_7;
    wire clk_en_52;
    wire rco_c_57;
    wire rco_c_56;
    wire clk_en_54_cascade_;
    wire rco_c_55;
    wire shift_srl_48Z0Z_15;
    wire shift_srl_56Z0Z_15;
    wire shift_srl_55_RNI9BJMZ0Z_15;
    wire rco_c_44;
    wire clk_en_0_a3_0_a2_sx_57_cascade_;
    wire shift_srl_47_RNIV3QLZ0Z_15;
    wire shift_srl_57Z0Z_15;
    wire shift_srl_57Z0Z_0;
    wire shift_srl_57Z0Z_1;
    wire shift_srl_57Z0Z_2;
    wire shift_srl_57Z0Z_3;
    wire shift_srl_57Z0Z_4;
    wire shift_srl_57Z0Z_5;
    wire shift_srl_57Z0Z_6;
    wire shift_srl_57Z0Z_7;
    wire clk_en_57;
    wire rco_int_0_a2_1_a2_sx_53;
    wire rco_c_53;
    wire shift_srl_54Z0Z_15;
    wire shift_srl_54Z0Z_0;
    wire shift_srl_54Z0Z_1;
    wire shift_srl_54Z0Z_2;
    wire shift_srl_54Z0Z_3;
    wire shift_srl_64Z0Z_10;
    wire shift_srl_64Z0Z_11;
    wire shift_srl_64Z0Z_12;
    wire shift_srl_64Z0Z_13;
    wire shift_srl_64Z0Z_14;
    wire shift_srl_64Z0Z_9;
    wire shift_srl_64Z0Z_8;
    wire shift_srl_65Z0Z_10;
    wire shift_srl_65Z0Z_11;
    wire shift_srl_65Z0Z_12;
    wire shift_srl_65Z0Z_13;
    wire shift_srl_65Z0Z_14;
    wire shift_srl_65Z0Z_9;
    wire shift_srl_65Z0Z_8;
    wire shift_srl_63Z0Z_7;
    wire shift_srl_63Z0Z_8;
    wire shift_srl_31Z0Z_0;
    wire shift_srl_31Z0Z_1;
    wire shift_srl_31Z0Z_2;
    wire shift_srl_31Z0Z_3;
    wire shift_srl_31Z0Z_4;
    wire shift_srl_31Z0Z_5;
    wire shift_srl_31Z0Z_6;
    wire shift_srl_31Z0Z_10;
    wire shift_srl_31Z0Z_11;
    wire shift_srl_31Z0Z_12;
    wire shift_srl_31Z0Z_13;
    wire shift_srl_31Z0Z_14;
    wire shift_srl_31Z0Z_9;
    wire shift_srl_31Z0Z_7;
    wire shift_srl_31Z0Z_8;
    wire shift_srl_160Z0Z_15;
    wire shift_srl_162Z0Z_15;
    wire shift_srl_161Z0Z_15;
    wire rco_int_0_a3_0_a2_0_sx_162_cascade_;
    wire rco_int_0_a3_0_a2_0_162_cascade_;
    wire shift_srl_159Z0Z_14;
    wire shift_srl_159Z0Z_15;
    wire shift_srl_158Z0Z_15;
    wire shift_srl_157Z0Z_15;
    wire rco_int_0_a2_0_a2_1_145;
    wire clk_en_0_a3_0_a2_sx_159_cascade_;
    wire clk_en_159;
    wire shift_srl_156Z0Z_15;
    wire shift_srl_155Z0Z_15;
    wire shift_srl_154Z0Z_15;
    wire shift_srl_156_RNII4IKZ0Z_15;
    wire shift_srl_171Z0Z_10;
    wire shift_srl_171Z0Z_11;
    wire shift_srl_171Z0Z_12;
    wire shift_srl_171Z0Z_13;
    wire shift_srl_171Z0Z_14;
    wire shift_srl_171Z0Z_8;
    wire shift_srl_171Z0Z_9;
    wire shift_srl_171Z0Z_0;
    wire shift_srl_171Z0Z_1;
    wire clk_en_171;
    wire shift_srl_179Z0Z_10;
    wire shift_srl_179Z0Z_11;
    wire shift_srl_179Z0Z_12;
    wire shift_srl_179Z0Z_13;
    wire shift_srl_179Z0Z_14;
    wire shift_srl_179Z0Z_9;
    wire shift_srl_179Z0Z_7;
    wire shift_srl_179Z0Z_8;
    wire clk_en_179;
    wire shift_srl_178Z0Z_5;
    wire shift_srl_178Z0Z_10;
    wire shift_srl_178Z0Z_11;
    wire shift_srl_178Z0Z_12;
    wire shift_srl_178Z0Z_6;
    wire shift_srl_178Z0Z_13;
    wire shift_srl_178Z0Z_14;
    wire shift_srl_178Z0Z_7;
    wire shift_srl_178Z0Z_8;
    wire rco_int_0_a2_1_a2_0_sx_179;
    wire shift_srl_179_RNIVNOT1Z0Z_15_cascade_;
    wire shift_srl_179_RNIVNOT1Z0Z_15;
    wire shift_srl_179Z0Z_15;
    wire rco_int_0_a2_1_a2_0_sx_182;
    wire clk_en_178;
    wire shift_srl_177Z0Z_14;
    wire shift_srl_181Z0Z_10;
    wire shift_srl_181Z0Z_11;
    wire shift_srl_181Z0Z_12;
    wire shift_srl_181Z0Z_6;
    wire shift_srl_181Z0Z_13;
    wire shift_srl_181Z0Z_14;
    wire shift_srl_181Z0Z_9;
    wire shift_srl_181Z0Z_7;
    wire shift_srl_181Z0Z_8;
    wire clk_en_181;
    wire shift_srl_189Z0Z_10;
    wire shift_srl_189Z0Z_11;
    wire shift_srl_189Z0Z_12;
    wire shift_srl_189Z0Z_13;
    wire shift_srl_189Z0Z_14;
    wire shift_srl_189Z0Z_9;
    wire shift_srl_189Z0Z_8;
    wire shift_srl_188Z0Z_0;
    wire shift_srl_188Z0Z_1;
    wire shift_srl_188Z0Z_2;
    wire shift_srl_188Z0Z_3;
    wire shift_srl_188Z0Z_4;
    wire shift_srl_188Z0Z_5;
    wire shift_srl_188Z0Z_6;
    wire shift_srl_176Z0Z_15;
    wire shift_srl_176Z0Z_0;
    wire shift_srl_176Z0Z_1;
    wire shift_srl_176Z0Z_2;
    wire shift_srl_176Z0Z_3;
    wire shift_srl_176Z0Z_4;
    wire shift_srl_176Z0Z_5;
    wire shift_srl_176Z0Z_6;
    wire shift_srl_176Z0Z_7;
    wire clk_en_176;
    wire rco_c_120;
    wire shift_srl_121Z0Z_15;
    wire rco_c_121;
    wire rco_c_177;
    wire shift_srl_83Z0Z_12;
    wire shift_srl_83Z0Z_13;
    wire shift_srl_83Z0Z_14;
    wire shift_srl_83Z0Z_11;
    wire shift_srl_83Z0Z_0;
    wire shift_srl_83Z0Z_1;
    wire shift_srl_83Z0Z_2;
    wire shift_srl_83Z0Z_3;
    wire shift_srl_83Z0Z_7;
    wire shift_srl_83Z0Z_4;
    wire shift_srl_83Z0Z_5;
    wire shift_srl_83Z0Z_6;
    wire shift_srl_82Z0Z_0;
    wire shift_srl_82Z0Z_1;
    wire shift_srl_82Z0Z_2;
    wire shift_srl_82Z0Z_3;
    wire shift_srl_82Z0Z_4;
    wire shift_srl_82Z0Z_5;
    wire shift_srl_82Z0Z_6;
    wire shift_srl_41Z0Z_15;
    wire shift_srl_41Z0Z_0;
    wire shift_srl_41Z0Z_1;
    wire shift_srl_41Z0Z_2;
    wire shift_srl_41Z0Z_3;
    wire shift_srl_41Z0Z_4;
    wire shift_srl_41Z0Z_5;
    wire shift_srl_41Z0Z_6;
    wire shift_srl_41Z0Z_7;
    wire clk_en_41;
    wire shift_srl_56Z0Z_0;
    wire shift_srl_56Z0Z_1;
    wire shift_srl_56Z0Z_6;
    wire shift_srl_56Z0Z_2;
    wire shift_srl_56Z0Z_5;
    wire shift_srl_56Z0Z_3;
    wire shift_srl_56Z0Z_4;
    wire shift_srl_56Z0Z_7;
    wire shift_srl_56Z0Z_8;
    wire clk_en_56;
    wire shift_srl_58Z0Z_0;
    wire shift_srl_58Z0Z_1;
    wire shift_srl_58Z0Z_2;
    wire shift_srl_58Z0Z_3;
    wire shift_srl_58Z0Z_4;
    wire shift_srl_58Z0Z_5;
    wire shift_srl_58Z0Z_6;
    wire shift_srl_58Z0Z_10;
    wire shift_srl_58Z0Z_11;
    wire shift_srl_58Z0Z_12;
    wire shift_srl_58Z0Z_13;
    wire shift_srl_58Z0Z_14;
    wire shift_srl_58Z0Z_15;
    wire shift_srl_58Z0Z_9;
    wire shift_srl_58Z0Z_7;
    wire shift_srl_58Z0Z_8;
    wire clk_en_58;
    wire shift_srl_64Z0Z_0;
    wire shift_srl_64Z0Z_1;
    wire shift_srl_64Z0Z_2;
    wire shift_srl_64Z0Z_3;
    wire shift_srl_64Z0Z_4;
    wire shift_srl_64Z0Z_5;
    wire shift_srl_64Z0Z_6;
    wire shift_srl_64Z0Z_7;
    wire clk_en_64;
    wire clk_en_60;
    wire shift_srl_63Z0Z_14;
    wire shift_srl_63Z0Z_13;
    wire shift_srl_63Z0Z_12;
    wire shift_srl_63Z0Z_11;
    wire shift_srl_63Z0Z_9;
    wire shift_srl_63Z0Z_10;
    wire clk_en_63;
    wire shift_srl_65Z0Z_0;
    wire shift_srl_65Z0Z_1;
    wire shift_srl_65Z0Z_2;
    wire shift_srl_65Z0Z_3;
    wire shift_srl_65Z0Z_4;
    wire shift_srl_65Z0Z_5;
    wire shift_srl_65Z0Z_6;
    wire shift_srl_65Z0Z_7;
    wire clk_en_65;
    wire shift_srl_30Z0Z_6;
    wire shift_srl_38Z0Z_15;
    wire rco_c_38;
    wire rco_c_38_cascade_;
    wire shift_srl_30Z0Z_7;
    wire shift_srl_100Z0Z_15;
    wire rco_c_100;
    wire rco_int_0_a3_0_a2_out_0;
    wire rco_c_99;
    wire rco_c_104;
    wire rco_c_29;
    wire clk_en_31;
    wire shift_srl_30Z0Z_14;
    wire shift_srl_30Z0Z_13;
    wire shift_srl_30Z0Z_12;
    wire shift_srl_30Z0Z_11;
    wire shift_srl_30Z0Z_10;
    wire shift_srl_30Z0Z_8;
    wire shift_srl_30Z0Z_9;
    wire clk_en_30;
    wire shift_srl_165Z0Z_10;
    wire shift_srl_165Z0Z_11;
    wire shift_srl_165Z0Z_12;
    wire shift_srl_165Z0Z_13;
    wire shift_srl_165Z0Z_14;
    wire shift_srl_165Z0Z_9;
    wire shift_srl_165Z0Z_8;
    wire shift_srl_165Z0Z_0;
    wire shift_srl_165Z0Z_1;
    wire shift_srl_165Z0Z_2;
    wire shift_srl_165Z0Z_3;
    wire shift_srl_165Z0Z_4;
    wire shift_srl_165Z0Z_5;
    wire shift_srl_165Z0Z_6;
    wire shift_srl_165Z0Z_7;
    wire clk_en_165;
    wire shift_srl_167Z0Z_10;
    wire shift_srl_167Z0Z_11;
    wire shift_srl_167Z0Z_12;
    wire shift_srl_167Z0Z_13;
    wire shift_srl_167Z0Z_14;
    wire shift_srl_167Z0Z_9;
    wire shift_srl_167Z0Z_8;
    wire shift_srl_167Z0Z_0;
    wire shift_srl_167Z0Z_1;
    wire shift_srl_167Z0Z_2;
    wire shift_srl_167Z0Z_3;
    wire shift_srl_167Z0Z_4;
    wire shift_srl_167Z0Z_5;
    wire shift_srl_167Z0Z_6;
    wire shift_srl_167Z0Z_7;
    wire shift_srl_170Z0Z_0;
    wire shift_srl_170Z0Z_1;
    wire shift_srl_170Z0Z_2;
    wire shift_srl_170Z0Z_3;
    wire shift_srl_170Z0Z_4;
    wire shift_srl_170Z0Z_5;
    wire shift_srl_170Z0Z_6;
    wire shift_srl_177Z0Z_0;
    wire shift_srl_177Z0Z_1;
    wire shift_srl_177Z0Z_2;
    wire shift_srl_177Z0Z_3;
    wire shift_srl_177Z0Z_4;
    wire shift_srl_177Z0Z_5;
    wire shift_srl_177Z0Z_13;
    wire shift_srl_180Z0Z_0;
    wire shift_srl_180Z0Z_1;
    wire shift_srl_180Z0Z_2;
    wire shift_srl_180Z0Z_3;
    wire shift_srl_180Z0Z_7;
    wire shift_srl_180Z0Z_6;
    wire N_4173;
    wire rco_c_188;
    wire shift_srl_188Z0Z_14;
    wire shift_srl_188Z0Z_13;
    wire shift_srl_188Z0Z_12;
    wire shift_srl_188Z0Z_11;
    wire shift_srl_188Z0Z_10;
    wire shift_srl_192Z0Z_7;
    wire shift_srl_192Z0Z_8;
    wire shift_srl_192Z0Z_9;
    wire clk_en_192;
    wire shift_srl_173Z0Z_10;
    wire shift_srl_173Z0Z_11;
    wire shift_srl_173Z0Z_12;
    wire shift_srl_173Z0Z_13;
    wire shift_srl_173Z0Z_14;
    wire shift_srl_173Z0Z_9;
    wire shift_srl_173Z0Z_7;
    wire shift_srl_173Z0Z_8;
    wire clk_en_173;
    wire shift_srl_176_RNIUGI51Z0Z_15;
    wire shift_srl_177Z0Z_15;
    wire shift_srl_178Z0Z_15;
    wire rco_c_178;
    wire shift_srl_83Z0Z_10;
    wire shift_srl_83Z0Z_8;
    wire shift_srl_83Z0Z_9;
    wire shift_srl_82Z0Z_10;
    wire shift_srl_82Z0Z_11;
    wire shift_srl_82Z0Z_12;
    wire shift_srl_82Z0Z_13;
    wire shift_srl_82Z0Z_14;
    wire shift_srl_82Z0Z_9;
    wire shift_srl_82Z0Z_7;
    wire shift_srl_82Z0Z_8;
    wire N_3998_i;
    wire shift_srl_80_RNIG3FB1Z0Z_15_cascade_;
    wire clk_en_0_a3_0_a2_0_83_cascade_;
    wire clk_en_83;
    wire N_787;
    wire shift_srl_82Z0Z_15;
    wire shift_srl_83Z0Z_15;
    wire rco_int_0_a2_0_a2_0_83;
    wire shift_srl_76Z0Z_10;
    wire shift_srl_76Z0Z_11;
    wire shift_srl_76Z0Z_12;
    wire shift_srl_76Z0Z_13;
    wire shift_srl_76Z0Z_14;
    wire shift_srl_76Z0Z_9;
    wire shift_srl_76Z0Z_8;
    wire shift_srl_76Z0Z_0;
    wire shift_srl_76Z0Z_1;
    wire shift_srl_76Z0Z_2;
    wire shift_srl_76Z0Z_3;
    wire shift_srl_76Z0Z_4;
    wire shift_srl_76Z0Z_5;
    wire shift_srl_76Z0Z_6;
    wire shift_srl_76Z0Z_7;
    wire rco_c_64;
    wire rco_c_63;
    wire shift_srl_63Z0Z_15;
    wire shift_srl_64Z0Z_15;
    wire shift_srl_62_RNIM5RKZ0Z_15;
    wire shift_srl_65Z0Z_15;
    wire shift_srl_65_RNILFDF1Z0Z_15;
    wire shift_srl_65_RNILFDF1Z0Z_15_cascade_;
    wire shift_srl_59Z0Z_15;
    wire rco_int_0_a2_1_a2_0_53;
    wire shift_srl_54_RNIEAU71Z0Z_15;
    wire rco_int_0_a2_1_a2_0_0_59;
    wire rco_int_0_a3_0_a2cf1_1_66;
    wire rco_int_0_a2_1_a2_1_48;
    wire rco_int_0_a2_1_a2_0_0_59_cascade_;
    wire rco_int_0_a3_0_a2cf1_66_cascade_;
    wire rco_c_37;
    wire rco_c_66_cascade_;
    wire clk_en_76;
    wire shift_srl_66Z0Z_0;
    wire shift_srl_66Z0Z_1;
    wire shift_srl_66Z0Z_2;
    wire shift_srl_66Z0Z_3;
    wire shift_srl_66Z0Z_4;
    wire shift_srl_66Z0Z_5;
    wire shift_srl_66Z0Z_6;
    wire shift_srl_66Z0Z_10;
    wire shift_srl_66Z0Z_11;
    wire shift_srl_66Z0Z_12;
    wire shift_srl_66Z0Z_13;
    wire shift_srl_66Z0Z_14;
    wire shift_srl_66Z0Z_15;
    wire shift_srl_66Z0Z_9;
    wire shift_srl_66Z0Z_7;
    wire shift_srl_66Z0Z_8;
    wire clk_en_66;
    wire shift_srl_35Z0Z_10;
    wire shift_srl_35Z0Z_11;
    wire shift_srl_35Z0Z_12;
    wire shift_srl_35Z0Z_13;
    wire shift_srl_35Z0Z_14;
    wire shift_srl_35Z0Z_9;
    wire shift_srl_35Z0Z_8;
    wire shift_srl_34Z0Z_14;
    wire shift_srl_34Z0Z_13;
    wire shift_srl_34Z0Z_12;
    wire shift_srl_34Z0Z_11;
    wire shift_srl_34Z0Z_10;
    wire shift_srl_34Z0Z_9;
    wire shift_srl_35Z0Z_15;
    wire shift_srl_35Z0Z_0;
    wire shift_srl_35Z0Z_1;
    wire shift_srl_35Z0Z_2;
    wire shift_srl_35Z0Z_3;
    wire shift_srl_35Z0Z_4;
    wire shift_srl_35Z0Z_5;
    wire shift_srl_35Z0Z_6;
    wire shift_srl_35Z0Z_7;
    wire clk_en_35;
    wire shift_srl_39Z0Z_15;
    wire shift_srl_39Z0Z_0;
    wire shift_srl_39Z0Z_1;
    wire shift_srl_39Z0Z_2;
    wire shift_srl_39Z0Z_3;
    wire shift_srl_39Z0Z_4;
    wire shift_srl_39Z0Z_5;
    wire shift_srl_39Z0Z_6;
    wire shift_srl_169Z0Z_4;
    wire shift_srl_169Z0Z_5;
    wire shift_srl_169Z0Z_6;
    wire shift_srl_39Z0Z_7;
    wire shift_srl_39Z0Z_8;
    wire clk_en_39;
    wire shift_srl_169Z0Z_10;
    wire shift_srl_169Z0Z_11;
    wire shift_srl_169Z0Z_2;
    wire shift_srl_169Z0Z_3;
    wire shift_srl_169Z0Z_12;
    wire shift_srl_169Z0Z_13;
    wire shift_srl_169Z0Z_14;
    wire shift_srl_169Z0Z_9;
    wire shift_srl_169Z0Z_7;
    wire shift_srl_169Z0Z_8;
    wire shift_srl_164_RNIBMOLZ0Z_15;
    wire clk_en_167;
    wire rco_int_0_a2_0_a2_0_153;
    wire rco_c_145;
    wire clk_en_163_cascade_;
    wire shift_srl_169Z0Z_0;
    wire shift_srl_169Z0Z_1;
    wire clk_en_169;
    wire shift_srl_170Z0Z_10;
    wire shift_srl_170Z0Z_11;
    wire shift_srl_170Z0Z_12;
    wire shift_srl_170Z0Z_13;
    wire shift_srl_170Z0Z_14;
    wire shift_srl_170Z0Z_9;
    wire shift_srl_170Z0Z_7;
    wire shift_srl_170Z0Z_8;
    wire clk_en_170;
    wire shift_srl_177Z0Z_10;
    wire shift_srl_177Z0Z_11;
    wire shift_srl_177Z0Z_12;
    wire shift_srl_177Z0Z_6;
    wire shift_srl_177Z0Z_9;
    wire shift_srl_177Z0Z_7;
    wire shift_srl_177Z0Z_8;
    wire clk_en_177;
    wire shift_srl_180Z0Z_10;
    wire shift_srl_180Z0Z_4;
    wire shift_srl_180Z0Z_5;
    wire shift_srl_180Z0Z_13;
    wire shift_srl_180Z0Z_14;
    wire shift_srl_180Z0Z_15;
    wire shift_srl_180Z0Z_11;
    wire shift_srl_180Z0Z_12;
    wire shift_srl_180Z0Z_8;
    wire shift_srl_180Z0Z_9;
    wire clk_en_180;
    wire shift_srl_189Z0Z_0;
    wire shift_srl_189Z0Z_1;
    wire shift_srl_189Z0Z_2;
    wire shift_srl_189Z0Z_3;
    wire shift_srl_189Z0Z_4;
    wire shift_srl_189Z0Z_5;
    wire shift_srl_189Z0Z_6;
    wire shift_srl_189Z0Z_7;
    wire clk_en_189;
    wire shift_srl_188Z0Z_7;
    wire shift_srl_188Z0Z_8;
    wire shift_srl_188Z0Z_9;
    wire clk_en_188;
    wire shift_srl_80Z0Z_0;
    wire shift_srl_80Z0Z_1;
    wire shift_srl_80Z0Z_2;
    wire shift_srl_80Z0Z_3;
    wire shift_srl_80Z0Z_4;
    wire shift_srl_80Z0Z_5;
    wire shift_srl_80Z0Z_6;
    wire shift_srl_80Z0Z_7;
    wire shift_srl_78Z0Z_10;
    wire shift_srl_78Z0Z_11;
    wire shift_srl_78Z0Z_12;
    wire shift_srl_78Z0Z_13;
    wire shift_srl_78Z0Z_14;
    wire shift_srl_78Z0Z_9;
    wire shift_srl_78Z0Z_8;
    wire shift_srl_78Z0Z_0;
    wire shift_srl_78Z0Z_1;
    wire shift_srl_78Z0Z_2;
    wire shift_srl_78Z0Z_3;
    wire shift_srl_78Z0Z_4;
    wire shift_srl_78Z0Z_5;
    wire shift_srl_78Z0Z_6;
    wire shift_srl_78Z0Z_7;
    wire shift_srl_69Z0Z_0;
    wire shift_srl_69Z0Z_1;
    wire shift_srl_69Z0Z_2;
    wire shift_srl_69Z0Z_3;
    wire shift_srl_69Z0Z_4;
    wire shift_srl_69Z0Z_5;
    wire shift_srl_67Z0Z_9;
    wire shift_srl_67Z0Z_8;
    wire shift_srl_67Z0Z_7;
    wire shift_srl_67Z0Z_6;
    wire shift_srl_67Z0Z_5;
    wire rco_c_67;
    wire rco_c_68;
    wire rco_c_69;
    wire shift_srl_67Z0Z_0;
    wire shift_srl_67Z0Z_1;
    wire shift_srl_67Z0Z_2;
    wire shift_srl_67Z0Z_3;
    wire shift_srl_67Z0Z_4;
    wire shift_srl_71Z0Z_10;
    wire shift_srl_71Z0Z_3;
    wire shift_srl_71Z0Z_9;
    wire shift_srl_71Z0Z_0;
    wire shift_srl_71Z0Z_1;
    wire shift_srl_71Z0Z_2;
    wire shift_srl_68_RNIHDC4Z0Z_15_cascade_;
    wire shift_srl_69_RNIBQRCZ0Z_15;
    wire shift_srl_69_RNIBQRCZ0Z_15_cascade_;
    wire shift_srl_67Z0Z_14;
    wire shift_srl_67Z0Z_13;
    wire shift_srl_67Z0Z_12;
    wire shift_srl_67Z0Z_10;
    wire shift_srl_67Z0Z_11;
    wire shift_srl_70Z0Z_1;
    wire shift_srl_70Z0Z_2;
    wire shift_srl_70Z0Z_3;
    wire shift_srl_70Z0Z_4;
    wire shift_srl_70Z0Z_5;
    wire shift_srl_70Z0Z_6;
    wire shift_srl_70Z0Z_7;
    wire shift_srl_34Z0Z_15;
    wire shift_srl_34Z0Z_0;
    wire shift_srl_34Z0Z_1;
    wire shift_srl_34Z0Z_2;
    wire shift_srl_34Z0Z_3;
    wire shift_srl_37Z0Z_14;
    wire shift_srl_37Z0Z_15;
    wire shift_srl_37Z0Z_0;
    wire shift_srl_37Z0Z_1;
    wire shift_srl_37Z0Z_2;
    wire shift_srl_37Z0Z_3;
    wire shift_srl_37Z0Z_4;
    wire rco_c_32;
    wire rco_c_32_cascade_;
    wire shift_srl_29Z0Z_15;
    wire shift_srl_28Z0Z_15;
    wire shift_srl_24Z0Z_15;
    wire shift_srl_30Z0Z_15;
    wire shift_srl_27_RNIP5TNZ0Z_15;
    wire shift_srl_29_RNISHF41Z0Z_15_cascade_;
    wire shift_srl_31Z0Z_15;
    wire rco_int_0_a2_0_a2_out_4_cascade_;
    wire rco_c_33;
    wire rco_int_0_a2_0_a2_out_4;
    wire rco_int_0_a2_0_a2_s_0_0_35;
    wire rco_c_36;
    wire rco_c_35;
    wire shift_srl_36Z0Z_15;
    wire shift_srl_36Z0Z_0;
    wire shift_srl_36Z0Z_1;
    wire shift_srl_36Z0Z_2;
    wire shift_srl_36Z0Z_3;
    wire shift_srl_36Z0Z_4;
    wire rco_c_169;
    wire rco_c_168;
    wire shift_srl_166Z0Z_15;
    wire shift_srl_165Z0Z_15;
    wire shift_srl_167Z0Z_15;
    wire shift_srl_167_RNIUC2TZ0Z_15_cascade_;
    wire shift_srl_170Z0Z_15;
    wire shift_srl_169Z0Z_15;
    wire shift_srl_163_RNI3MR51Z0Z_15_cascade_;
    wire shift_srl_170_RNIRM2S1Z0Z_15_cascade_;
    wire rco_int_0_a3_0_a2_0_172;
    wire rco_int_0_a3_0_a2_0_172_cascade_;
    wire clk_en_0_a3_0_a2cf1_1_176;
    wire shift_srl_163Z0Z_10;
    wire shift_srl_163Z0Z_11;
    wire shift_srl_163Z0Z_12;
    wire shift_srl_163Z0Z_13;
    wire shift_srl_163Z0Z_14;
    wire shift_srl_163Z0Z_9;
    wire shift_srl_163Z0Z_8;
    wire shift_srl_36Z0Z_10;
    wire shift_srl_36Z0Z_11;
    wire shift_srl_36Z0Z_12;
    wire shift_srl_36Z0Z_9;
    wire shift_srl_36Z0Z_8;
    wire shift_srl_36Z0Z_7;
    wire shift_srl_191Z0Z_10;
    wire shift_srl_191Z0Z_11;
    wire shift_srl_191Z0Z_12;
    wire shift_srl_191Z0Z_13;
    wire shift_srl_191Z0Z_14;
    wire shift_srl_191Z0Z_9;
    wire shift_srl_191Z0Z_8;
    wire shift_srl_36Z0Z_5;
    wire shift_srl_36Z0Z_6;
    wire rco_c_79;
    wire N_785;
    wire shift_srl_81Z0Z_0;
    wire shift_srl_81Z0Z_1;
    wire shift_srl_81Z0Z_2;
    wire shift_srl_81Z0Z_3;
    wire shift_srl_81Z0Z_4;
    wire shift_srl_81Z0Z_5;
    wire shift_srl_81Z0Z_6;
    wire shift_srl_79_RNITG241Z0Z_15;
    wire shift_srl_79_RNITG241Z0Z_15_cascade_;
    wire rco_c_78;
    wire shift_srl_79Z0Z_0;
    wire shift_srl_78Z0Z_15;
    wire rco_int_0_a2_0_a2_0_1_83;
    wire shift_srl_80Z0Z_15;
    wire shift_srl_80Z0Z_14;
    wire shift_srl_80Z0Z_13;
    wire shift_srl_80Z0Z_12;
    wire shift_srl_80Z0Z_11;
    wire shift_srl_80Z0Z_10;
    wire shift_srl_80Z0Z_8;
    wire shift_srl_80Z0Z_9;
    wire clk_en_80;
    wire shift_srl_76Z0Z_15;
    wire shift_srl_76_RNIF788Z0Z_15_cascade_;
    wire clk_en_78;
    wire shift_srl_75Z0Z_14;
    wire shift_srl_75Z0Z_13;
    wire shift_srl_75Z0Z_12;
    wire shift_srl_75Z0Z_11;
    wire shift_srl_68Z0Z_0;
    wire shift_srl_68Z0Z_1;
    wire shift_srl_68Z0Z_2;
    wire shift_srl_68Z0Z_3;
    wire shift_srl_68Z0Z_4;
    wire shift_srl_68Z0Z_5;
    wire shift_srl_68Z0Z_6;
    wire rco_c_70;
    wire shift_srl_71_RNIGP6RZ0Z_15_cascade_;
    wire rco_int_0_a2_1_a2_sx_59;
    wire rco_int_0_a2_1_a2_sx_44;
    wire N_4016_i;
    wire rco_c_59_cascade_;
    wire rco_int_0_a3_0_a2_0_66;
    wire rco_c_59;
    wire shift_srl_68_RNIHDC4Z0Z_15;
    wire shift_srl_69Z0Z_14;
    wire shift_srl_69Z0Z_13;
    wire shift_srl_69Z0Z_12;
    wire shift_srl_69Z0Z_11;
    wire shift_srl_69Z0Z_10;
    wire shift_srl_71Z0Z_4;
    wire shift_srl_71Z0Z_5;
    wire shift_srl_71Z0Z_6;
    wire shift_srl_71Z0Z_13;
    wire shift_srl_71Z0Z_14;
    wire shift_srl_71Z0Z_11;
    wire shift_srl_71Z0Z_12;
    wire shift_srl_71Z0Z_7;
    wire shift_srl_71Z0Z_8;
    wire clk_en_71;
    wire shift_srl_69Z0Z_6;
    wire shift_srl_69Z0Z_7;
    wire shift_srl_69Z0Z_8;
    wire shift_srl_69Z0Z_9;
    wire clk_en_69;
    wire shift_srl_70Z0Z_10;
    wire shift_srl_70Z0Z_11;
    wire shift_srl_70Z0Z_12;
    wire shift_srl_70Z0Z_13;
    wire shift_srl_70Z0Z_14;
    wire shift_srl_70Z0Z_8;
    wire shift_srl_70Z0Z_9;
    wire shift_srl_70Z0Z_0;
    wire clk_en_70;
    wire shift_srl_34Z0Z_4;
    wire shift_srl_34Z0Z_5;
    wire shift_srl_37Z0Z_12;
    wire shift_srl_37Z0Z_13;
    wire shift_srl_37Z0Z_5;
    wire shift_srl_37Z0Z_6;
    wire shift_srl_37Z0Z_9;
    wire shift_srl_37Z0Z_7;
    wire shift_srl_37Z0Z_8;
    wire shift_srl_33Z0Z_0;
    wire shift_srl_33Z0Z_1;
    wire shift_srl_33Z0Z_2;
    wire shift_srl_33Z0Z_3;
    wire shift_srl_33Z0Z_13;
    wire shift_srl_33Z0Z_14;
    wire shift_srl_33Z0Z_15;
    wire shift_srl_33Z0Z_10;
    wire shift_srl_33Z0Z_11;
    wire shift_srl_33Z0Z_12;
    wire shift_srl_33Z0Z_4;
    wire shift_srl_33Z0Z_5;
    wire shift_srl_33Z0Z_6;
    wire shift_srl_33Z0Z_9;
    wire shift_srl_33Z0Z_7;
    wire shift_srl_33Z0Z_8;
    wire clk_en_33;
    wire shift_srl_164Z0Z_10;
    wire shift_srl_164Z0Z_13;
    wire shift_srl_164Z0Z_14;
    wire shift_srl_164Z0Z_8;
    wire shift_srl_164Z0Z_9;
    wire shift_srl_164Z0Z_6;
    wire shift_srl_164Z0Z_7;
    wire shift_srl_163Z0Z_0;
    wire shift_srl_163Z0Z_1;
    wire shift_srl_163Z0Z_2;
    wire shift_srl_163Z0Z_3;
    wire shift_srl_163Z0Z_4;
    wire shift_srl_163Z0Z_5;
    wire shift_srl_163Z0Z_6;
    wire shift_srl_163Z0Z_7;
    wire clk_en_163;
    wire shift_srl_191Z0Z_15;
    wire shift_srl_191Z0Z_0;
    wire shift_srl_191Z0Z_1;
    wire shift_srl_191Z0Z_2;
    wire shift_srl_191Z0Z_3;
    wire shift_srl_191Z0Z_4;
    wire shift_srl_191Z0Z_5;
    wire shift_srl_191Z0Z_6;
    wire shift_srl_191Z0Z_7;
    wire shift_srl_187Z0Z_15;
    wire shift_srl_189Z0Z_15;
    wire clk_en_0_a3_0_a2_0_sx_190_cascade_;
    wire shift_srl_188Z0Z_15;
    wire N_4175_cascade_;
    wire clk_en_191;
    wire rco_int_0_a3_0_a2_0_183;
    wire rco_c_172;
    wire shift_srl_79Z0Z_1;
    wire shift_srl_79Z0Z_2;
    wire shift_srl_79Z0Z_3;
    wire shift_srl_79Z0Z_4;
    wire shift_srl_79Z0Z_5;
    wire shift_srl_79Z0Z_6;
    wire shift_srl_81Z0Z_10;
    wire shift_srl_81Z0Z_11;
    wire shift_srl_81Z0Z_12;
    wire shift_srl_81Z0Z_13;
    wire shift_srl_81Z0Z_14;
    wire shift_srl_81Z0Z_15;
    wire shift_srl_81Z0Z_9;
    wire shift_srl_81Z0Z_7;
    wire shift_srl_81Z0Z_8;
    wire N_786;
    wire shift_srl_79Z0Z_10;
    wire shift_srl_79Z0Z_11;
    wire shift_srl_79Z0Z_12;
    wire shift_srl_79Z0Z_13;
    wire shift_srl_79Z0Z_14;
    wire shift_srl_79Z0Z_15;
    wire shift_srl_79Z0Z_9;
    wire shift_srl_79Z0Z_7;
    wire shift_srl_79Z0Z_8;
    wire clk_en_79;
    wire shift_srl_77Z0Z_10;
    wire shift_srl_77Z0Z_11;
    wire shift_srl_77Z0Z_12;
    wire shift_srl_77Z0Z_13;
    wire shift_srl_77Z0Z_14;
    wire shift_srl_77Z0Z_9;
    wire shift_srl_77Z0Z_8;
    wire shift_srl_68Z0Z_10;
    wire shift_srl_68Z0Z_11;
    wire shift_srl_68Z0Z_12;
    wire shift_srl_68Z0Z_13;
    wire shift_srl_68Z0Z_14;
    wire shift_srl_68Z0Z_9;
    wire shift_srl_68Z0Z_7;
    wire shift_srl_68Z0Z_8;
    wire clk_en_68;
    wire shift_srl_72Z0Z_0;
    wire shift_srl_72Z0Z_1;
    wire shift_srl_72Z0Z_2;
    wire shift_srl_72Z0Z_3;
    wire shift_srl_72Z0Z_4;
    wire shift_srl_72Z0Z_5;
    wire shift_srl_72Z0Z_6;
    wire clk_en_67;
    wire shift_srl_68Z0Z_15;
    wire shift_srl_67Z0Z_15;
    wire shift_srl_74_RNIS4SRZ0Z_15_cascade_;
    wire rco_int_0_a3_0_a2_0_74;
    wire shift_srl_71Z0Z_15;
    wire shift_srl_70Z0Z_15;
    wire shift_srl_69Z0Z_15;
    wire rco_int_0_a3_0_a2_0_1_74;
    wire shift_srl_72Z0Z_10;
    wire shift_srl_72Z0Z_11;
    wire shift_srl_72Z0Z_12;
    wire shift_srl_72Z0Z_13;
    wire shift_srl_72Z0Z_14;
    wire shift_srl_72Z0Z_9;
    wire shift_srl_72Z0Z_7;
    wire shift_srl_72Z0Z_8;
    wire clk_en_72;
    wire shift_srl_34Z0Z_6;
    wire shift_srl_54Z0Z_4;
    wire shift_srl_54Z0Z_5;
    wire shift_srl_54Z0Z_6;
    wire shift_srl_54Z0Z_7;
    wire shift_srl_54Z0Z_8;
    wire shift_srl_54Z0Z_9;
    wire clk_en_54;
    wire shift_srl_34Z0Z_7;
    wire shift_srl_34Z0Z_8;
    wire clk_en_34;
    wire shift_srl_32Z0Z_10;
    wire shift_srl_32Z0Z_11;
    wire shift_srl_32Z0Z_12;
    wire shift_srl_32Z0Z_13;
    wire shift_srl_32Z0Z_14;
    wire shift_srl_32Z0Z_9;
    wire shift_srl_32Z0Z_8;
    wire rco_c_31;
    wire shift_srl_32Z0Z_15;
    wire shift_srl_32Z0Z_0;
    wire shift_srl_32Z0Z_1;
    wire shift_srl_164Z0Z_15;
    wire shift_srl_164Z0Z_0;
    wire shift_srl_164Z0Z_1;
    wire shift_srl_164Z0Z_2;
    wire shift_srl_164Z0Z_3;
    wire shift_srl_164Z0Z_4;
    wire shift_srl_164Z0Z_5;
    wire shift_srl_164Z0Z_11;
    wire shift_srl_164Z0Z_12;
    wire rco_c_171;
    wire shift_srl_171Z0Z_15;
    wire shift_srl_171_RNIVSP62Z0Z_15;
    wire shift_srl_171_RNIVSP62Z0Z_15_cascade_;
    wire shift_srl_170_RNIRM2S1Z0Z_15;
    wire rco_c_170;
    wire shift_srl_163_RNI3MR51Z0Z_15;
    wire rco_c_167;
    wire rco_int_0_a3_0_a2_0_162;
    wire rco_c_153;
    wire clk_en_164;
    wire shift_srl_163Z0Z_15;
    wire rco_c_162;
    wire rco_c_163;
    wire shift_srl_168Z0Z_0;
    wire shift_srl_168Z0Z_1;
    wire shift_srl_168Z0Z_2;
    wire shift_srl_168Z0Z_3;
    wire shift_srl_168Z0Z_4;
    wire shift_srl_168Z0Z_5;
    wire shift_srl_168Z0Z_6;
    wire shift_srl_190Z0Z_9;
    wire shift_srl_190Z0Z_3;
    wire shift_srl_190Z0Z_4;
    wire shift_srl_190Z0Z_10;
    wire shift_srl_190Z0Z_5;
    wire shift_srl_190Z0Z_11;
    wire shift_srl_190Z0Z_8;
    wire shift_srl_190Z0Z_6;
    wire shift_srl_190Z0Z_7;
    wire shift_srl_190Z0Z_12;
    wire shift_srl_190Z0Z_13;
    wire shift_srl_190Z0Z_14;
    wire shift_srl_190Z0Z_2;
    wire shift_srl_190Z0Z_0;
    wire shift_srl_190Z0Z_1;
    wire clk_en_190;
    wire shift_srl_139Z0Z_15;
    wire rco_c_139;
    wire shift_srl_50_RNI869CZ0Z_15;
    wire rco_c_50;
    wire shift_srl_77Z0Z_15;
    wire shift_srl_77Z0Z_0;
    wire shift_srl_77Z0Z_1;
    wire shift_srl_77Z0Z_2;
    wire shift_srl_77Z0Z_3;
    wire shift_srl_77Z0Z_4;
    wire shift_srl_77Z0Z_5;
    wire shift_srl_77Z0Z_6;
    wire shift_srl_77Z0Z_7;
    wire clk_en_77;
    wire rco_c_75;
    wire shift_srl_76_RNIF788Z0Z_15;
    wire rco_c_76;
    wire shift_srl_77_RNI8HLIZ0Z_15;
    wire rco_c_77;
    wire rco_c_74;
    wire shift_srl_80_RNIG3FB1Z0Z_15;
    wire rco_c_80;
    wire shift_srl_75Z0Z_15;
    wire shift_srl_75Z0Z_0;
    wire shift_srl_75Z0Z_1;
    wire shift_srl_75Z0Z_2;
    wire shift_srl_75Z0Z_10;
    wire shift_srl_75Z0Z_9;
    wire shift_srl_75Z0Z_8;
    wire shift_srl_75Z0Z_7;
    wire shift_srl_75Z0Z_6;
    wire shift_srl_75Z0Z_5;
    wire shift_srl_75Z0Z_3;
    wire shift_srl_75Z0Z_4;
    wire clk_en_75;
    wire shift_srl_74Z0Z_0;
    wire shift_srl_74Z0Z_1;
    wire shift_srl_74Z0Z_2;
    wire shift_srl_74Z0Z_3;
    wire shift_srl_74Z0Z_4;
    wire shift_srl_74Z0Z_5;
    wire shift_srl_74Z0Z_6;
    wire shift_srl_74Z0Z_10;
    wire shift_srl_74Z0Z_11;
    wire shift_srl_74Z0Z_12;
    wire shift_srl_74Z0Z_13;
    wire shift_srl_74Z0Z_14;
    wire shift_srl_74Z0Z_15;
    wire shift_srl_74Z0Z_9;
    wire shift_srl_74Z0Z_7;
    wire shift_srl_74Z0Z_8;
    wire clk_en_74;
    wire shift_srl_32Z0Z_7;
    wire shift_srl_32Z0Z_6;
    wire shift_srl_32Z0Z_4;
    wire shift_srl_32Z0Z_5;
    wire shift_srl_32Z0Z_2;
    wire shift_srl_32Z0Z_3;
    wire clk_en_32;
    wire shift_srl_172Z0Z_10;
    wire shift_srl_172Z0Z_11;
    wire shift_srl_172Z0Z_12;
    wire shift_srl_172Z0Z_13;
    wire shift_srl_172Z0Z_14;
    wire shift_srl_172Z0Z_9;
    wire shift_srl_172Z0Z_8;
    wire shift_srl_172Z0Z_15;
    wire shift_srl_172Z0Z_0;
    wire shift_srl_172Z0Z_1;
    wire shift_srl_172Z0Z_2;
    wire shift_srl_172Z0Z_3;
    wire shift_srl_172Z0Z_4;
    wire shift_srl_172Z0Z_5;
    wire shift_srl_172Z0Z_6;
    wire shift_srl_172Z0Z_7;
    wire clk_en_172;
    wire shift_srl_168Z0Z_13;
    wire shift_srl_168Z0Z_14;
    wire shift_srl_168Z0Z_15;
    wire shift_srl_168Z0Z_12;
    wire shift_srl_168Z0Z_7;
    wire shift_srl_168Z0Z_8;
    wire shift_srl_168Z0Z_9;
    wire shift_srl_168Z0Z_10;
    wire shift_srl_168Z0Z_11;
    wire clk_en_168;
    wire rco_c_72;
    wire shift_srl_73Z0Z_10;
    wire shift_srl_73Z0Z_11;
    wire shift_srl_73Z0Z_12;
    wire shift_srl_73Z0Z_13;
    wire shift_srl_73Z0Z_14;
    wire shift_srl_73Z0Z_9;
    wire shift_srl_73Z0Z_8;
    wire rco_c_0;
    wire shift_srl_73Z0Z_0;
    wire shift_srl_73Z0Z_1;
    wire shift_srl_73Z0Z_2;
    wire shift_srl_73Z0Z_3;
    wire shift_srl_73Z0Z_4;
    wire shift_srl_73Z0Z_5;
    wire shift_srl_73Z0Z_6;
    wire shift_srl_73Z0Z_7;
    wire clk_en_73;
    wire shift_srl_36Z0Z_13;
    wire shift_srl_36Z0Z_14;
    wire clk_en_36;
    wire shift_srl_73Z0Z_15;
    wire shift_srl_72Z0Z_15;
    wire rco_c_73;
    wire shift_srl_71_RNIGP6RZ0Z_15;
    wire rco_c_66;
    wire rco_c_71;
    wire shift_srl_37Z0Z_10;
    wire shift_srl_37Z0Z_11;
    wire clk_c_g;
    wire clk_en_37;
    wire shift_srl_186Z0Z_15;
    wire rco_c_186;
    wire shift_srl_185Z0Z_15;
    wire shift_srl_184Z0Z_15;
    wire rco_c_185;
    wire shift_srl_190Z0Z_15;
    wire rco_c_190;
    wire N_4175;
    wire rco_c_183;
    wire rco_c_189;
    wire shift_srl_129_RNIDM4DZ0Z_15;
    wire rco_c_129;
    wire rco_c_127;
    wire shift_srl_128Z0Z_15;
    wire rco_c_128;
    wire shift_srl_140_RNI85IAZ0Z_15;
    wire rco_c_138;
    wire N_125_i;
    wire rco_c_48;
    wire shift_srl_49Z0Z_15;
    wire rco_c_49;
    wire _gnd_net_;

    PRE_IO_GBUF clk_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__95450),
            .GLOBALBUFFEROUTPUT(clk_c_g));
    IO_PAD clk_ibuf_gb_io_iopad (
            .OE(N__95452),
            .DIN(N__95451),
            .DOUT(N__95450),
            .PACKAGEPIN(clk));
    defparam clk_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam clk_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_ibuf_gb_io_preio (
            .PADOEN(N__95452),
            .PADOUT(N__95451),
            .PADIN(N__95450),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD en_in_ibuf_iopad (
            .OE(N__95441),
            .DIN(N__95440),
            .DOUT(N__95439),
            .PACKAGEPIN(en_in));
    defparam en_in_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam en_in_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO en_in_ibuf_preio (
            .PADOEN(N__95441),
            .PADOUT(N__95440),
            .PADIN(N__95439),
            .CLOCKENABLE(),
            .DIN0(en_in_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_0_iopad (
            .OE(N__95432),
            .DIN(N__95431),
            .DOUT(N__95430),
            .PACKAGEPIN(rco[0]));
    defparam rco_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_0_preio (
            .PADOEN(N__95432),
            .PADOUT(N__95431),
            .PADIN(N__95430),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__90307),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_1_iopad (
            .OE(N__95423),
            .DIN(N__95422),
            .DOUT(N__95421),
            .PACKAGEPIN(rco[1]));
    defparam rco_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_1_preio (
            .PADOEN(N__95423),
            .PADOUT(N__95422),
            .PADIN(N__95421),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__57133),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_10_iopad (
            .OE(N__95414),
            .DIN(N__95413),
            .DOUT(N__95412),
            .PACKAGEPIN(rco[10]));
    defparam rco_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_10_preio (
            .PADOEN(N__95414),
            .PADOUT(N__95413),
            .PADIN(N__95412),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__52327),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_100_iopad (
            .OE(N__95405),
            .DIN(N__95404),
            .DOUT(N__95403),
            .PACKAGEPIN(rco[100]));
    defparam rco_obuf_100_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_100_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_100_preio (
            .PADOEN(N__95405),
            .PADOUT(N__95404),
            .PADIN(N__95403),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__79638),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_101_iopad (
            .OE(N__95396),
            .DIN(N__95395),
            .DOUT(N__95394),
            .PACKAGEPIN(rco[101]));
    defparam rco_obuf_101_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_101_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_101_preio (
            .PADOEN(N__95396),
            .PADOUT(N__95395),
            .PADIN(N__95394),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__58186),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_102_iopad (
            .OE(N__95387),
            .DIN(N__95386),
            .DOUT(N__95385),
            .PACKAGEPIN(rco[102]));
    defparam rco_obuf_102_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_102_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_102_preio (
            .PADOEN(N__95387),
            .PADOUT(N__95386),
            .PADIN(N__95385),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__59167),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_103_iopad (
            .OE(N__95378),
            .DIN(N__95377),
            .DOUT(N__95376),
            .PACKAGEPIN(rco[103]));
    defparam rco_obuf_103_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_103_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_103_preio (
            .PADOEN(N__95378),
            .PADOUT(N__95377),
            .PADIN(N__95376),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__59140),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_104_iopad (
            .OE(N__95369),
            .DIN(N__95368),
            .DOUT(N__95367),
            .PACKAGEPIN(rco[104]));
    defparam rco_obuf_104_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_104_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_104_preio (
            .PADOEN(N__95369),
            .PADOUT(N__95368),
            .PADIN(N__95367),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__79248),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_105_iopad (
            .OE(N__95360),
            .DIN(N__95359),
            .DOUT(N__95358),
            .PACKAGEPIN(rco[105]));
    defparam rco_obuf_105_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_105_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_105_preio (
            .PADOEN(N__95360),
            .PADOUT(N__95359),
            .PADIN(N__95358),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__57982),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_106_iopad (
            .OE(N__95351),
            .DIN(N__95350),
            .DOUT(N__95349),
            .PACKAGEPIN(rco[106]));
    defparam rco_obuf_106_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_106_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_106_preio (
            .PADOEN(N__95351),
            .PADOUT(N__95350),
            .PADIN(N__95349),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__56647),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_107_iopad (
            .OE(N__95342),
            .DIN(N__95341),
            .DOUT(N__95340),
            .PACKAGEPIN(rco[107]));
    defparam rco_obuf_107_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_107_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_107_preio (
            .PADOEN(N__95342),
            .PADOUT(N__95341),
            .PADIN(N__95340),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__55519),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_108_iopad (
            .OE(N__95333),
            .DIN(N__95332),
            .DOUT(N__95331),
            .PACKAGEPIN(rco[108]));
    defparam rco_obuf_108_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_108_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_108_preio (
            .PADOEN(N__95333),
            .PADOUT(N__95332),
            .PADIN(N__95331),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__55546),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_109_iopad (
            .OE(N__95324),
            .DIN(N__95323),
            .DOUT(N__95322),
            .PACKAGEPIN(rco[109]));
    defparam rco_obuf_109_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_109_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_109_preio (
            .PADOEN(N__95324),
            .PADOUT(N__95323),
            .PADIN(N__95322),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__55531),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_11_iopad (
            .OE(N__95315),
            .DIN(N__95314),
            .DOUT(N__95313),
            .PACKAGEPIN(rco[11]));
    defparam rco_obuf_11_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_11_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_11_preio (
            .PADOEN(N__95315),
            .PADOUT(N__95314),
            .PADIN(N__95313),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__50377),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_110_iopad (
            .OE(N__95306),
            .DIN(N__95305),
            .DOUT(N__95304),
            .PACKAGEPIN(rco[110]));
    defparam rco_obuf_110_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_110_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_110_preio (
            .PADOEN(N__95306),
            .PADOUT(N__95305),
            .PADIN(N__95304),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__62011),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_111_iopad (
            .OE(N__95297),
            .DIN(N__95296),
            .DOUT(N__95295),
            .PACKAGEPIN(rco[111]));
    defparam rco_obuf_111_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_111_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_111_preio (
            .PADOEN(N__95297),
            .PADOUT(N__95296),
            .PADIN(N__95295),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__60670),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_112_iopad (
            .OE(N__95288),
            .DIN(N__95287),
            .DOUT(N__95286),
            .PACKAGEPIN(rco[112]));
    defparam rco_obuf_112_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_112_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_112_preio (
            .PADOEN(N__95288),
            .PADOUT(N__95287),
            .PADIN(N__95286),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__60364),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_113_iopad (
            .OE(N__95279),
            .DIN(N__95278),
            .DOUT(N__95277),
            .PACKAGEPIN(rco[113]));
    defparam rco_obuf_113_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_113_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_113_preio (
            .PADOEN(N__95279),
            .PADOUT(N__95278),
            .PADIN(N__95277),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__53260),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_114_iopad (
            .OE(N__95270),
            .DIN(N__95269),
            .DOUT(N__95268),
            .PACKAGEPIN(rco[114]));
    defparam rco_obuf_114_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_114_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_114_preio (
            .PADOEN(N__95270),
            .PADOUT(N__95269),
            .PADIN(N__95268),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__63880),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_115_iopad (
            .OE(N__95261),
            .DIN(N__95260),
            .DOUT(N__95259),
            .PACKAGEPIN(rco[115]));
    defparam rco_obuf_115_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_115_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_115_preio (
            .PADOEN(N__95261),
            .PADOUT(N__95260),
            .PADIN(N__95259),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__63856),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_116_iopad (
            .OE(N__95252),
            .DIN(N__95251),
            .DOUT(N__95250),
            .PACKAGEPIN(rco[116]));
    defparam rco_obuf_116_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_116_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_116_preio (
            .PADOEN(N__95252),
            .PADOUT(N__95251),
            .PADIN(N__95250),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__66496),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_117_iopad (
            .OE(N__95243),
            .DIN(N__95242),
            .DOUT(N__95241),
            .PACKAGEPIN(rco[117]));
    defparam rco_obuf_117_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_117_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_117_preio (
            .PADOEN(N__95243),
            .PADOUT(N__95242),
            .PADIN(N__95241),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__66334),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_118_iopad (
            .OE(N__95234),
            .DIN(N__95233),
            .DOUT(N__95232),
            .PACKAGEPIN(rco[118]));
    defparam rco_obuf_118_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_118_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_118_preio (
            .PADOEN(N__95234),
            .PADOUT(N__95233),
            .PADIN(N__95232),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__65977),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_119_iopad (
            .OE(N__95225),
            .DIN(N__95224),
            .DOUT(N__95223),
            .PACKAGEPIN(rco[119]));
    defparam rco_obuf_119_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_119_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_119_preio (
            .PADOEN(N__95225),
            .PADOUT(N__95224),
            .PADIN(N__95223),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__65227),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_12_iopad (
            .OE(N__95216),
            .DIN(N__95215),
            .DOUT(N__95214),
            .PACKAGEPIN(rco[12]));
    defparam rco_obuf_12_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_12_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_12_preio (
            .PADOEN(N__95216),
            .PADOUT(N__95215),
            .PADIN(N__95214),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__49528),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_120_iopad (
            .OE(N__95207),
            .DIN(N__95206),
            .DOUT(N__95205),
            .PACKAGEPIN(rco[120]));
    defparam rco_obuf_120_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_120_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_120_preio (
            .PADOEN(N__95207),
            .PADOUT(N__95206),
            .PADIN(N__95205),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__78519),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_121_iopad (
            .OE(N__95198),
            .DIN(N__95197),
            .DOUT(N__95196),
            .PACKAGEPIN(rco[121]));
    defparam rco_obuf_121_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_121_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_121_preio (
            .PADOEN(N__95198),
            .PADOUT(N__95197),
            .PADIN(N__95196),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__78415),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_122_iopad (
            .OE(N__95189),
            .DIN(N__95188),
            .DOUT(N__95187),
            .PACKAGEPIN(rco[122]));
    defparam rco_obuf_122_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_122_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_122_preio (
            .PADOEN(N__95189),
            .PADOUT(N__95188),
            .PADIN(N__95187),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__55318),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_123_iopad (
            .OE(N__95180),
            .DIN(N__95179),
            .DOUT(N__95178),
            .PACKAGEPIN(rco[123]));
    defparam rco_obuf_123_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_123_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_123_preio (
            .PADOEN(N__95180),
            .PADOUT(N__95179),
            .PADIN(N__95178),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__57625),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_124_iopad (
            .OE(N__95171),
            .DIN(N__95170),
            .DOUT(N__95169),
            .PACKAGEPIN(rco[124]));
    defparam rco_obuf_124_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_124_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_124_preio (
            .PADOEN(N__95171),
            .PADOUT(N__95170),
            .PADIN(N__95169),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__50179),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_125_iopad (
            .OE(N__95162),
            .DIN(N__95161),
            .DOUT(N__95160),
            .PACKAGEPIN(rco[125]));
    defparam rco_obuf_125_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_125_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_125_preio (
            .PADOEN(N__95162),
            .PADOUT(N__95161),
            .PADIN(N__95160),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__51181),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_126_iopad (
            .OE(N__95153),
            .DIN(N__95152),
            .DOUT(N__95151),
            .PACKAGEPIN(rco[126]));
    defparam rco_obuf_126_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_126_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_126_preio (
            .PADOEN(N__95153),
            .PADOUT(N__95152),
            .PADIN(N__95151),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__57646),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_127_iopad (
            .OE(N__95144),
            .DIN(N__95143),
            .DOUT(N__95142),
            .PACKAGEPIN(rco[127]));
    defparam rco_obuf_127_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_127_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_127_preio (
            .PADOEN(N__95144),
            .PADOUT(N__95143),
            .PADIN(N__95142),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__91334),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_128_iopad (
            .OE(N__95135),
            .DIN(N__95134),
            .DOUT(N__95133),
            .PACKAGEPIN(rco[128]));
    defparam rco_obuf_128_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_128_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_128_preio (
            .PADOEN(N__95135),
            .PADOUT(N__95134),
            .PADIN(N__95133),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__91174),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_129_iopad (
            .OE(N__95126),
            .DIN(N__95125),
            .DOUT(N__95124),
            .PACKAGEPIN(rco[129]));
    defparam rco_obuf_129_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_129_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_129_preio (
            .PADOEN(N__95126),
            .PADOUT(N__95125),
            .PADIN(N__95124),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__91351),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_13_iopad (
            .OE(N__95117),
            .DIN(N__95116),
            .DOUT(N__95115),
            .PACKAGEPIN(rco[13]));
    defparam rco_obuf_13_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_13_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_13_preio (
            .PADOEN(N__95117),
            .PADOUT(N__95116),
            .PADIN(N__95115),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__49276),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_130_iopad (
            .OE(N__95108),
            .DIN(N__95107),
            .DOUT(N__95106),
            .PACKAGEPIN(rco[130]));
    defparam rco_obuf_130_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_130_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_130_preio (
            .PADOEN(N__95108),
            .PADOUT(N__95107),
            .PADIN(N__95106),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__51007),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_131_iopad (
            .OE(N__95099),
            .DIN(N__95098),
            .DOUT(N__95097),
            .PACKAGEPIN(rco[131]));
    defparam rco_obuf_131_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_131_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_131_preio (
            .PADOEN(N__95099),
            .PADOUT(N__95098),
            .PADIN(N__95097),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__51025),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_132_iopad (
            .OE(N__95090),
            .DIN(N__95089),
            .DOUT(N__95088),
            .PACKAGEPIN(rco[132]));
    defparam rco_obuf_132_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_132_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_132_preio (
            .PADOEN(N__95090),
            .PADOUT(N__95089),
            .PADIN(N__95088),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__66316),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_133_iopad (
            .OE(N__95081),
            .DIN(N__95080),
            .DOUT(N__95079),
            .PACKAGEPIN(rco[133]));
    defparam rco_obuf_133_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_133_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_133_preio (
            .PADOEN(N__95081),
            .PADOUT(N__95080),
            .PADIN(N__95079),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__66184),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_134_iopad (
            .OE(N__95072),
            .DIN(N__95071),
            .DOUT(N__95070),
            .PACKAGEPIN(rco[134]));
    defparam rco_obuf_134_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_134_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_134_preio (
            .PADOEN(N__95072),
            .PADOUT(N__95071),
            .PADIN(N__95070),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__51235),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_135_iopad (
            .OE(N__95063),
            .DIN(N__95062),
            .DOUT(N__95061),
            .PACKAGEPIN(rco[135]));
    defparam rco_obuf_135_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_135_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_135_preio (
            .PADOEN(N__95063),
            .PADOUT(N__95062),
            .PADIN(N__95061),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__51199),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_136_iopad (
            .OE(N__95054),
            .DIN(N__95053),
            .DOUT(N__95052),
            .PACKAGEPIN(rco[136]));
    defparam rco_obuf_136_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_136_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_136_preio (
            .PADOEN(N__95054),
            .PADOUT(N__95053),
            .PADIN(N__95052),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__51307),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_137_iopad (
            .OE(N__95045),
            .DIN(N__95044),
            .DOUT(N__95043),
            .PACKAGEPIN(rco[137]));
    defparam rco_obuf_137_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_137_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_137_preio (
            .PADOEN(N__95045),
            .PADOUT(N__95044),
            .PADIN(N__95043),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__51124),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_138_iopad (
            .OE(N__95036),
            .DIN(N__95035),
            .DOUT(N__95034),
            .PACKAGEPIN(rco[138]));
    defparam rco_obuf_138_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_138_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_138_preio (
            .PADOEN(N__95036),
            .PADOUT(N__95035),
            .PADIN(N__95034),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__91126),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_139_iopad (
            .OE(N__95027),
            .DIN(N__95026),
            .DOUT(N__95025),
            .PACKAGEPIN(rco[139]));
    defparam rco_obuf_139_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_139_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_139_preio (
            .PADOEN(N__95027),
            .PADOUT(N__95026),
            .PADIN(N__95025),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__88069),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_14_iopad (
            .OE(N__95018),
            .DIN(N__95017),
            .DOUT(N__95016),
            .PACKAGEPIN(rco[14]));
    defparam rco_obuf_14_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_14_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_14_preio (
            .PADOEN(N__95018),
            .PADOUT(N__95017),
            .PADIN(N__95016),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__50599),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_140_iopad (
            .OE(N__95009),
            .DIN(N__95008),
            .DOUT(N__95007),
            .PACKAGEPIN(rco[140]));
    defparam rco_obuf_140_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_140_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_140_preio (
            .PADOEN(N__95009),
            .PADOUT(N__95008),
            .PADIN(N__95007),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__91048),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_141_iopad (
            .OE(N__95000),
            .DIN(N__94999),
            .DOUT(N__94998),
            .PACKAGEPIN(rco[141]));
    defparam rco_obuf_141_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_141_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_141_preio (
            .PADOEN(N__95000),
            .PADOUT(N__94999),
            .PADIN(N__94998),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__66562),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_142_iopad (
            .OE(N__94991),
            .DIN(N__94990),
            .DOUT(N__94989),
            .PACKAGEPIN(rco[142]));
    defparam rco_obuf_142_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_142_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_142_preio (
            .PADOEN(N__94991),
            .PADOUT(N__94990),
            .PADIN(N__94989),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__60013),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_143_iopad (
            .OE(N__94982),
            .DIN(N__94981),
            .DOUT(N__94980),
            .PACKAGEPIN(rco[143]));
    defparam rco_obuf_143_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_143_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_143_preio (
            .PADOEN(N__94982),
            .PADOUT(N__94981),
            .PADIN(N__94980),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__60025),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_144_iopad (
            .OE(N__94973),
            .DIN(N__94972),
            .DOUT(N__94971),
            .PACKAGEPIN(rco[144]));
    defparam rco_obuf_144_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_144_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_144_preio (
            .PADOEN(N__94973),
            .PADOUT(N__94972),
            .PADIN(N__94971),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__66511),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_145_iopad (
            .OE(N__94964),
            .DIN(N__94963),
            .DOUT(N__94962),
            .PACKAGEPIN(rco[145]));
    defparam rco_obuf_145_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_145_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_145_preio (
            .PADOEN(N__94964),
            .PADOUT(N__94963),
            .PADIN(N__94962),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__82221),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_146_iopad (
            .OE(N__94955),
            .DIN(N__94954),
            .DOUT(N__94953),
            .PACKAGEPIN(rco[146]));
    defparam rco_obuf_146_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_146_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_146_preio (
            .PADOEN(N__94955),
            .PADOUT(N__94954),
            .PADIN(N__94953),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__70669),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_147_iopad (
            .OE(N__94946),
            .DIN(N__94945),
            .DOUT(N__94944),
            .PACKAGEPIN(rco[147]));
    defparam rco_obuf_147_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_147_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_147_preio (
            .PADOEN(N__94946),
            .PADOUT(N__94945),
            .PADIN(N__94944),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__56002),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_148_iopad (
            .OE(N__94937),
            .DIN(N__94936),
            .DOUT(N__94935),
            .PACKAGEPIN(rco[148]));
    defparam rco_obuf_148_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_148_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_148_preio (
            .PADOEN(N__94937),
            .PADOUT(N__94936),
            .PADIN(N__94935),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__56026),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_149_iopad (
            .OE(N__94928),
            .DIN(N__94927),
            .DOUT(N__94926),
            .PACKAGEPIN(rco[149]));
    defparam rco_obuf_149_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_149_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_149_preio (
            .PADOEN(N__94928),
            .PADOUT(N__94927),
            .PADIN(N__94926),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__58294),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_15_iopad (
            .OE(N__94919),
            .DIN(N__94918),
            .DOUT(N__94917),
            .PACKAGEPIN(rco[15]));
    defparam rco_obuf_15_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_15_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_15_preio (
            .PADOEN(N__94919),
            .PADOUT(N__94918),
            .PADIN(N__94917),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__50461),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_150_iopad (
            .OE(N__94910),
            .DIN(N__94909),
            .DOUT(N__94908),
            .PACKAGEPIN(rco[150]));
    defparam rco_obuf_150_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_150_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_150_preio (
            .PADOEN(N__94910),
            .PADOUT(N__94909),
            .PADIN(N__94908),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__66751),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_151_iopad (
            .OE(N__94901),
            .DIN(N__94900),
            .DOUT(N__94899),
            .PACKAGEPIN(rco[151]));
    defparam rco_obuf_151_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_151_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_151_preio (
            .PADOEN(N__94901),
            .PADOUT(N__94900),
            .PADIN(N__94899),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__54712),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_152_iopad (
            .OE(N__94892),
            .DIN(N__94891),
            .DOUT(N__94890),
            .PACKAGEPIN(rco[152]));
    defparam rco_obuf_152_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_152_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_152_preio (
            .PADOEN(N__94892),
            .PADOUT(N__94891),
            .PADIN(N__94890),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__55573),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_153_iopad (
            .OE(N__94883),
            .DIN(N__94882),
            .DOUT(N__94881),
            .PACKAGEPIN(rco[153]));
    defparam rco_obuf_153_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_153_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_153_preio (
            .PADOEN(N__94883),
            .PADOUT(N__94882),
            .PADIN(N__94881),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__87916),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_154_iopad (
            .OE(N__94874),
            .DIN(N__94873),
            .DOUT(N__94872),
            .PACKAGEPIN(rco[154]));
    defparam rco_obuf_154_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_154_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_154_preio (
            .PADOEN(N__94874),
            .PADOUT(N__94873),
            .PADIN(N__94872),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__53545),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_155_iopad (
            .OE(N__94865),
            .DIN(N__94864),
            .DOUT(N__94863),
            .PACKAGEPIN(rco[155]));
    defparam rco_obuf_155_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_155_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_155_preio (
            .PADOEN(N__94865),
            .PADOUT(N__94864),
            .PADIN(N__94863),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__53563),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_156_iopad (
            .OE(N__94856),
            .DIN(N__94855),
            .DOUT(N__94854),
            .PACKAGEPIN(rco[156]));
    defparam rco_obuf_156_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_156_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_156_preio (
            .PADOEN(N__94856),
            .PADOUT(N__94855),
            .PADIN(N__94854),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__53527),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_157_iopad (
            .OE(N__94847),
            .DIN(N__94846),
            .DOUT(N__94845),
            .PACKAGEPIN(rco[157]));
    defparam rco_obuf_157_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_157_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_157_preio (
            .PADOEN(N__94847),
            .PADOUT(N__94846),
            .PADIN(N__94845),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__69931),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_158_iopad (
            .OE(N__94838),
            .DIN(N__94837),
            .DOUT(N__94836),
            .PACKAGEPIN(rco[158]));
    defparam rco_obuf_158_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_158_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_158_preio (
            .PADOEN(N__94838),
            .PADOUT(N__94837),
            .PADIN(N__94836),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__69955),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_159_iopad (
            .OE(N__94829),
            .DIN(N__94828),
            .DOUT(N__94827),
            .PACKAGEPIN(rco[159]));
    defparam rco_obuf_159_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_159_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_159_preio (
            .PADOEN(N__94829),
            .PADOUT(N__94828),
            .PADIN(N__94827),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__53509),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_16_iopad (
            .OE(N__94820),
            .DIN(N__94819),
            .DOUT(N__94818),
            .PACKAGEPIN(rco[16]));
    defparam rco_obuf_16_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_16_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_16_preio (
            .PADOEN(N__94820),
            .PADOUT(N__94819),
            .PADIN(N__94818),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__49603),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_160_iopad (
            .OE(N__94811),
            .DIN(N__94810),
            .DOUT(N__94809),
            .PACKAGEPIN(rco[160]));
    defparam rco_obuf_160_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_160_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_160_preio (
            .PADOEN(N__94811),
            .PADOUT(N__94810),
            .PADIN(N__94809),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__53491),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_161_iopad (
            .OE(N__94802),
            .DIN(N__94801),
            .DOUT(N__94800),
            .PACKAGEPIN(rco[161]));
    defparam rco_obuf_161_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_161_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_161_preio (
            .PADOEN(N__94802),
            .PADOUT(N__94801),
            .PADIN(N__94800),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__53473),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_162_iopad (
            .OE(N__94793),
            .DIN(N__94792),
            .DOUT(N__94791),
            .PACKAGEPIN(rco[162]));
    defparam rco_obuf_162_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_162_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_162_preio (
            .PADOEN(N__94793),
            .PADOUT(N__94792),
            .PADIN(N__94791),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__87720),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_163_iopad (
            .OE(N__94784),
            .DIN(N__94783),
            .DOUT(N__94782),
            .PACKAGEPIN(rco[163]));
    defparam rco_obuf_163_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_163_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_163_preio (
            .PADOEN(N__94784),
            .PADOUT(N__94783),
            .PADIN(N__94782),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__87586),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_164_iopad (
            .OE(N__94775),
            .DIN(N__94774),
            .DOUT(N__94773),
            .PACKAGEPIN(rco[164]));
    defparam rco_obuf_164_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_164_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_164_preio (
            .PADOEN(N__94775),
            .PADOUT(N__94774),
            .PADIN(N__94773),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__53236),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_165_iopad (
            .OE(N__94766),
            .DIN(N__94765),
            .DOUT(N__94764),
            .PACKAGEPIN(rco[165]));
    defparam rco_obuf_165_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_165_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_165_preio (
            .PADOEN(N__94766),
            .PADOUT(N__94765),
            .PADIN(N__94764),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__59413),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_166_iopad (
            .OE(N__94757),
            .DIN(N__94756),
            .DOUT(N__94755),
            .PACKAGEPIN(rco[166]));
    defparam rco_obuf_166_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_166_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_166_preio (
            .PADOEN(N__94757),
            .PADOUT(N__94756),
            .PADIN(N__94755),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__71683),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_167_iopad (
            .OE(N__94748),
            .DIN(N__94747),
            .DOUT(N__94746),
            .PACKAGEPIN(rco[167]));
    defparam rco_obuf_167_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_167_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_167_preio (
            .PADOEN(N__94748),
            .PADOUT(N__94747),
            .PADIN(N__94746),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__87388),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_168_iopad (
            .OE(N__94739),
            .DIN(N__94738),
            .DOUT(N__94737),
            .PACKAGEPIN(rco[168]));
    defparam rco_obuf_168_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_168_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_168_preio (
            .PADOEN(N__94739),
            .PADOUT(N__94738),
            .PADIN(N__94737),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__84037),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_169_iopad (
            .OE(N__94730),
            .DIN(N__94729),
            .DOUT(N__94728),
            .PACKAGEPIN(rco[169]));
    defparam rco_obuf_169_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_169_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_169_preio (
            .PADOEN(N__94730),
            .PADOUT(N__94729),
            .PADIN(N__94728),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__84058),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_17_iopad (
            .OE(N__94721),
            .DIN(N__94720),
            .DOUT(N__94719),
            .PACKAGEPIN(rco[17]));
    defparam rco_obuf_17_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_17_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_17_preio (
            .PADOEN(N__94721),
            .PADOUT(N__94720),
            .PADIN(N__94719),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__50317),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_170_iopad (
            .OE(N__94712),
            .DIN(N__94711),
            .DOUT(N__94710),
            .PACKAGEPIN(rco[170]));
    defparam rco_obuf_170_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_170_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_170_preio (
            .PADOEN(N__94712),
            .PADOUT(N__94711),
            .PADIN(N__94710),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__87442),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_171_iopad (
            .OE(N__94703),
            .DIN(N__94702),
            .DOUT(N__94701),
            .PACKAGEPIN(rco[171]));
    defparam rco_obuf_171_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_171_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_171_preio (
            .PADOEN(N__94703),
            .PADOUT(N__94702),
            .PADIN(N__94701),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__87508),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_172_iopad (
            .OE(N__94694),
            .DIN(N__94693),
            .DOUT(N__94692),
            .PACKAGEPIN(rco[172]));
    defparam rco_obuf_172_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_172_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_172_preio (
            .PADOEN(N__94694),
            .PADOUT(N__94693),
            .PADIN(N__94692),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__85993),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_173_iopad (
            .OE(N__94685),
            .DIN(N__94684),
            .DOUT(N__94683),
            .PACKAGEPIN(rco[173]));
    defparam rco_obuf_173_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_173_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_173_preio (
            .PADOEN(N__94685),
            .PADOUT(N__94684),
            .PADIN(N__94683),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__66739),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_174_iopad (
            .OE(N__94676),
            .DIN(N__94675),
            .DOUT(N__94674),
            .PACKAGEPIN(rco[174]));
    defparam rco_obuf_174_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_174_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_174_preio (
            .PADOEN(N__94676),
            .PADOUT(N__94675),
            .PADIN(N__94674),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__75733),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_175_iopad (
            .OE(N__94667),
            .DIN(N__94666),
            .DOUT(N__94665),
            .PACKAGEPIN(rco[175]));
    defparam rco_obuf_175_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_175_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_175_preio (
            .PADOEN(N__94667),
            .PADOUT(N__94666),
            .PADIN(N__94665),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__75748),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_176_iopad (
            .OE(N__94658),
            .DIN(N__94657),
            .DOUT(N__94656),
            .PACKAGEPIN(rco[176]));
    defparam rco_obuf_176_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_176_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_176_preio (
            .PADOEN(N__94658),
            .PADOUT(N__94657),
            .PADIN(N__94656),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__66724),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_177_iopad (
            .OE(N__94649),
            .DIN(N__94648),
            .DOUT(N__94647),
            .PACKAGEPIN(rco[177]));
    defparam rco_obuf_177_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_177_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_177_preio (
            .PADOEN(N__94649),
            .PADOUT(N__94648),
            .PADIN(N__94647),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__78403),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_178_iopad (
            .OE(N__94640),
            .DIN(N__94639),
            .DOUT(N__94638),
            .PACKAGEPIN(rco[178]));
    defparam rco_obuf_178_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_178_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_178_preio (
            .PADOEN(N__94640),
            .PADOUT(N__94639),
            .PADIN(N__94638),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__80377),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_179_iopad (
            .OE(N__94631),
            .DIN(N__94630),
            .DOUT(N__94629),
            .PACKAGEPIN(rco[179]));
    defparam rco_obuf_179_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_179_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_179_preio (
            .PADOEN(N__94631),
            .PADOUT(N__94630),
            .PADIN(N__94629),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__66712),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_18_iopad (
            .OE(N__94622),
            .DIN(N__94621),
            .DOUT(N__94620),
            .PACKAGEPIN(rco[18]));
    defparam rco_obuf_18_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_18_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_18_preio (
            .PADOEN(N__94622),
            .PADOUT(N__94621),
            .PADIN(N__94620),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__50578),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_180_iopad (
            .OE(N__94613),
            .DIN(N__94612),
            .DOUT(N__94611),
            .PACKAGEPIN(rco[180]));
    defparam rco_obuf_180_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_180_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_180_preio (
            .PADOEN(N__94613),
            .PADOUT(N__94612),
            .PADIN(N__94611),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__71821),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_181_iopad (
            .OE(N__94604),
            .DIN(N__94603),
            .DOUT(N__94602),
            .PACKAGEPIN(rco[181]));
    defparam rco_obuf_181_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_181_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_181_preio (
            .PADOEN(N__94604),
            .PADOUT(N__94603),
            .PADIN(N__94602),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__71839),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_182_iopad (
            .OE(N__94595),
            .DIN(N__94594),
            .DOUT(N__94593),
            .PACKAGEPIN(rco[182]));
    defparam rco_obuf_182_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_182_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_182_preio (
            .PADOEN(N__94595),
            .PADOUT(N__94594),
            .PADIN(N__94593),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__66700),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_183_iopad (
            .OE(N__94586),
            .DIN(N__94585),
            .DOUT(N__94584),
            .PACKAGEPIN(rco[183]));
    defparam rco_obuf_183_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_183_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_183_preio (
            .PADOEN(N__94586),
            .PADOUT(N__94585),
            .PADIN(N__94584),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__91540),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_184_iopad (
            .OE(N__94577),
            .DIN(N__94576),
            .DOUT(N__94575),
            .PACKAGEPIN(rco[184]));
    defparam rco_obuf_184_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_184_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_184_preio (
            .PADOEN(N__94577),
            .PADOUT(N__94576),
            .PADIN(N__94575),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__64006),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_185_iopad (
            .OE(N__94568),
            .DIN(N__94567),
            .DOUT(N__94566),
            .PACKAGEPIN(rco[185]));
    defparam rco_obuf_185_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_185_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_185_preio (
            .PADOEN(N__94568),
            .PADOUT(N__94567),
            .PADIN(N__94566),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__91621),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_186_iopad (
            .OE(N__94559),
            .DIN(N__94558),
            .DOUT(N__94557),
            .PACKAGEPIN(rco[186]));
    defparam rco_obuf_186_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_186_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_186_preio (
            .PADOEN(N__94559),
            .PADOUT(N__94558),
            .PADIN(N__94557),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__91777),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_187_iopad (
            .OE(N__94550),
            .DIN(N__94549),
            .DOUT(N__94548),
            .PACKAGEPIN(rco[187]));
    defparam rco_obuf_187_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_187_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_187_preio (
            .PADOEN(N__94550),
            .PADOUT(N__94549),
            .PADIN(N__94548),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__63988),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_188_iopad (
            .OE(N__94541),
            .DIN(N__94540),
            .DOUT(N__94539),
            .PACKAGEPIN(rco[188]));
    defparam rco_obuf_188_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_188_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_188_preio (
            .PADOEN(N__94541),
            .PADOUT(N__94540),
            .PADIN(N__94539),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__80314),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_189_iopad (
            .OE(N__94532),
            .DIN(N__94531),
            .DOUT(N__94530),
            .PACKAGEPIN(rco[189]));
    defparam rco_obuf_189_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_189_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_189_preio (
            .PADOEN(N__94532),
            .PADOUT(N__94531),
            .PADIN(N__94530),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__91399),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_19_iopad (
            .OE(N__94523),
            .DIN(N__94522),
            .DOUT(N__94521),
            .PACKAGEPIN(rco[19]));
    defparam rco_obuf_19_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_19_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_19_preio (
            .PADOEN(N__94523),
            .PADOUT(N__94522),
            .PADIN(N__94521),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__49585),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_190_iopad (
            .OE(N__94514),
            .DIN(N__94513),
            .DOUT(N__94512),
            .PACKAGEPIN(rco[190]));
    defparam rco_obuf_190_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_190_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_190_preio (
            .PADOEN(N__94514),
            .PADOUT(N__94513),
            .PADIN(N__94512),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__91582),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_191_iopad (
            .OE(N__94505),
            .DIN(N__94504),
            .DOUT(N__94503),
            .PACKAGEPIN(rco[191]));
    defparam rco_obuf_191_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_191_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_191_preio (
            .PADOEN(N__94505),
            .PADOUT(N__94504),
            .PADIN(N__94503),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__64216),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_192_iopad (
            .OE(N__94496),
            .DIN(N__94495),
            .DOUT(N__94494),
            .PACKAGEPIN(rco[192]));
    defparam rco_obuf_192_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_192_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_192_preio (
            .PADOEN(N__94496),
            .PADOUT(N__94495),
            .PADIN(N__94494),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__74194),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_193_iopad (
            .OE(N__94487),
            .DIN(N__94486),
            .DOUT(N__94485),
            .PACKAGEPIN(rco[193]));
    defparam rco_obuf_193_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_193_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_193_preio (
            .PADOEN(N__94487),
            .PADOUT(N__94486),
            .PADIN(N__94485),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__64027),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_194_iopad (
            .OE(N__94478),
            .DIN(N__94477),
            .DOUT(N__94476),
            .PACKAGEPIN(rco[194]));
    defparam rco_obuf_194_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_194_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_194_preio (
            .PADOEN(N__94478),
            .PADOUT(N__94477),
            .PADIN(N__94476),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__64048),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_195_iopad (
            .OE(N__94469),
            .DIN(N__94468),
            .DOUT(N__94467),
            .PACKAGEPIN(rco[195]));
    defparam rco_obuf_195_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_195_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_195_preio (
            .PADOEN(N__94469),
            .PADOUT(N__94468),
            .PADIN(N__94467),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__64192),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_196_iopad (
            .OE(N__94460),
            .DIN(N__94459),
            .DOUT(N__94458),
            .PACKAGEPIN(rco[196]));
    defparam rco_obuf_196_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_196_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_196_preio (
            .PADOEN(N__94460),
            .PADOUT(N__94459),
            .PADIN(N__94458),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__72352),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_197_iopad (
            .OE(N__94451),
            .DIN(N__94450),
            .DOUT(N__94449),
            .PACKAGEPIN(rco[197]));
    defparam rco_obuf_197_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_197_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_197_preio (
            .PADOEN(N__94451),
            .PADOUT(N__94450),
            .PADIN(N__94449),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__70483),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_198_iopad (
            .OE(N__94442),
            .DIN(N__94441),
            .DOUT(N__94440),
            .PACKAGEPIN(rco[198]));
    defparam rco_obuf_198_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_198_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_198_preio (
            .PADOEN(N__94442),
            .PADOUT(N__94441),
            .PADIN(N__94440),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__70459),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_199_iopad (
            .OE(N__94433),
            .DIN(N__94432),
            .DOUT(N__94431),
            .PACKAGEPIN(rco[199]));
    defparam rco_obuf_199_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_199_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_199_preio (
            .PADOEN(N__94433),
            .PADOUT(N__94432),
            .PADIN(N__94431),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__60616),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_2_iopad (
            .OE(N__94424),
            .DIN(N__94423),
            .DOUT(N__94422),
            .PACKAGEPIN(rco[2]));
    defparam rco_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_2_preio (
            .PADOEN(N__94424),
            .PADOUT(N__94423),
            .PADIN(N__94422),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__52285),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_20_iopad (
            .OE(N__94415),
            .DIN(N__94414),
            .DOUT(N__94413),
            .PACKAGEPIN(rco[20]));
    defparam rco_obuf_20_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_20_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_20_preio (
            .PADOEN(N__94415),
            .PADOUT(N__94414),
            .PADIN(N__94413),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__50338),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_21_iopad (
            .OE(N__94406),
            .DIN(N__94405),
            .DOUT(N__94404),
            .PACKAGEPIN(rco[21]));
    defparam rco_obuf_21_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_21_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_21_preio (
            .PADOEN(N__94406),
            .PADOUT(N__94405),
            .PADIN(N__94404),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__52147),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_22_iopad (
            .OE(N__94397),
            .DIN(N__94396),
            .DOUT(N__94395),
            .PACKAGEPIN(rco[22]));
    defparam rco_obuf_22_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_22_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_22_preio (
            .PADOEN(N__94397),
            .PADOUT(N__94396),
            .PADIN(N__94395),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__48157),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_23_iopad (
            .OE(N__94388),
            .DIN(N__94387),
            .DOUT(N__94386),
            .PACKAGEPIN(rco[23]));
    defparam rco_obuf_23_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_23_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_23_preio (
            .PADOEN(N__94388),
            .PADOUT(N__94387),
            .PADIN(N__94386),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__85231),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_24_iopad (
            .OE(N__94379),
            .DIN(N__94378),
            .DOUT(N__94377),
            .PACKAGEPIN(rco[24]));
    defparam rco_obuf_24_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_24_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_24_preio (
            .PADOEN(N__94379),
            .PADOUT(N__94378),
            .PADIN(N__94377),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__58366),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_25_iopad (
            .OE(N__94370),
            .DIN(N__94369),
            .DOUT(N__94368),
            .PACKAGEPIN(rco[25]));
    defparam rco_obuf_25_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_25_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_25_preio (
            .PADOEN(N__94370),
            .PADOUT(N__94369),
            .PADIN(N__94368),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__53950),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_26_iopad (
            .OE(N__94361),
            .DIN(N__94360),
            .DOUT(N__94359),
            .PACKAGEPIN(rco[26]));
    defparam rco_obuf_26_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_26_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_26_preio (
            .PADOEN(N__94361),
            .PADOUT(N__94360),
            .PADIN(N__94359),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__53848),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_27_iopad (
            .OE(N__94352),
            .DIN(N__94351),
            .DOUT(N__94350),
            .PACKAGEPIN(rco[27]));
    defparam rco_obuf_27_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_27_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_27_preio (
            .PADOEN(N__94352),
            .PADOUT(N__94351),
            .PADIN(N__94350),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__67732),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_28_iopad (
            .OE(N__94343),
            .DIN(N__94342),
            .DOUT(N__94341),
            .PACKAGEPIN(rco[28]));
    defparam rco_obuf_28_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_28_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_28_preio (
            .PADOEN(N__94343),
            .PADOUT(N__94342),
            .PADIN(N__94341),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__67696),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_29_iopad (
            .OE(N__94334),
            .DIN(N__94333),
            .DOUT(N__94332),
            .PACKAGEPIN(rco[29]));
    defparam rco_obuf_29_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_29_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_29_preio (
            .PADOEN(N__94334),
            .PADOUT(N__94333),
            .PADIN(N__94332),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__79936),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_3_iopad (
            .OE(N__94325),
            .DIN(N__94324),
            .DOUT(N__94323),
            .PACKAGEPIN(rco[3]));
    defparam rco_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_3_preio (
            .PADOEN(N__94325),
            .PADOUT(N__94324),
            .PADIN(N__94323),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__48274),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_30_iopad (
            .OE(N__94316),
            .DIN(N__94315),
            .DOUT(N__94314),
            .PACKAGEPIN(rco[30]));
    defparam rco_obuf_30_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_30_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_30_preio (
            .PADOEN(N__94316),
            .PADOUT(N__94315),
            .PADIN(N__94314),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__69652),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_31_iopad (
            .OE(N__94307),
            .DIN(N__94306),
            .DOUT(N__94305),
            .PACKAGEPIN(rco[31]));
    defparam rco_obuf_31_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_31_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_31_preio (
            .PADOEN(N__94307),
            .PADOUT(N__94306),
            .PADIN(N__94305),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__87367),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_32_iopad (
            .OE(N__94298),
            .DIN(N__94297),
            .DOUT(N__94296),
            .PACKAGEPIN(rco[32]));
    defparam rco_obuf_32_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_32_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_32_preio (
            .PADOEN(N__94298),
            .PADOUT(N__94297),
            .PADIN(N__94296),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__83389),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_33_iopad (
            .OE(N__94289),
            .DIN(N__94288),
            .DOUT(N__94287),
            .PACKAGEPIN(rco[33]));
    defparam rco_obuf_33_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_33_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_33_preio (
            .PADOEN(N__94289),
            .PADOUT(N__94288),
            .PADIN(N__94287),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__83626),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_34_iopad (
            .OE(N__94280),
            .DIN(N__94279),
            .DOUT(N__94278),
            .PACKAGEPIN(rco[34]));
    defparam rco_obuf_34_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_34_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_34_preio (
            .PADOEN(N__94280),
            .PADOUT(N__94279),
            .PADIN(N__94278),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__69595),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_35_iopad (
            .OE(N__94271),
            .DIN(N__94270),
            .DOUT(N__94269),
            .PACKAGEPIN(rco[35]));
    defparam rco_obuf_35_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_35_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_35_preio (
            .PADOEN(N__94271),
            .PADOUT(N__94270),
            .PADIN(N__94269),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__83515),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_36_iopad (
            .OE(N__94262),
            .DIN(N__94261),
            .DOUT(N__94260),
            .PACKAGEPIN(rco[36]));
    defparam rco_obuf_36_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_36_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_36_preio (
            .PADOEN(N__94262),
            .PADOUT(N__94261),
            .PADIN(N__94260),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__83542),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_37_iopad (
            .OE(N__94253),
            .DIN(N__94252),
            .DOUT(N__94251),
            .PACKAGEPIN(rco[37]));
    defparam rco_obuf_37_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_37_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_37_preio (
            .PADOEN(N__94253),
            .PADOUT(N__94252),
            .PADIN(N__94251),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__81340),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_38_iopad (
            .OE(N__94244),
            .DIN(N__94243),
            .DOUT(N__94242),
            .PACKAGEPIN(rco[38]));
    defparam rco_obuf_38_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_38_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_38_preio (
            .PADOEN(N__94244),
            .PADOUT(N__94243),
            .PADIN(N__94242),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__79714),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_39_iopad (
            .OE(N__94235),
            .DIN(N__94234),
            .DOUT(N__94233),
            .PACKAGEPIN(rco[39]));
    defparam rco_obuf_39_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_39_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_39_preio (
            .PADOEN(N__94235),
            .PADOUT(N__94234),
            .PADIN(N__94233),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__67252),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_4_iopad (
            .OE(N__94226),
            .DIN(N__94225),
            .DOUT(N__94224),
            .PACKAGEPIN(rco[4]));
    defparam rco_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_4_preio (
            .PADOEN(N__94226),
            .PADOUT(N__94225),
            .PADIN(N__94224),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__48406),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_40_iopad (
            .OE(N__94217),
            .DIN(N__94216),
            .DOUT(N__94215),
            .PACKAGEPIN(rco[40]));
    defparam rco_obuf_40_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_40_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_40_preio (
            .PADOEN(N__94217),
            .PADOUT(N__94216),
            .PADIN(N__94215),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__67324),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_41_iopad (
            .OE(N__94208),
            .DIN(N__94207),
            .DOUT(N__94206),
            .PACKAGEPIN(rco[41]));
    defparam rco_obuf_41_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_41_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_41_preio (
            .PADOEN(N__94208),
            .PADOUT(N__94207),
            .PADIN(N__94206),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__69130),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_42_iopad (
            .OE(N__94199),
            .DIN(N__94198),
            .DOUT(N__94197),
            .PACKAGEPIN(rco[42]));
    defparam rco_obuf_42_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_42_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_42_preio (
            .PADOEN(N__94199),
            .PADOUT(N__94198),
            .PADIN(N__94197),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__64528),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_43_iopad (
            .OE(N__94190),
            .DIN(N__94189),
            .DOUT(N__94188),
            .PACKAGEPIN(rco[43]));
    defparam rco_obuf_43_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_43_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_43_preio (
            .PADOEN(N__94190),
            .PADOUT(N__94189),
            .PADIN(N__94188),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__64549),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_44_iopad (
            .OE(N__94181),
            .DIN(N__94180),
            .DOUT(N__94179),
            .PACKAGEPIN(rco[44]));
    defparam rco_obuf_44_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_44_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_44_preio (
            .PADOEN(N__94181),
            .PADOUT(N__94180),
            .PADIN(N__94179),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__76912),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_45_iopad (
            .OE(N__94172),
            .DIN(N__94171),
            .DOUT(N__94170),
            .PACKAGEPIN(rco[45]));
    defparam rco_obuf_45_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_45_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_45_preio (
            .PADOEN(N__94172),
            .PADOUT(N__94171),
            .PADIN(N__94170),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__76168),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_46_iopad (
            .OE(N__94163),
            .DIN(N__94162),
            .DOUT(N__94161),
            .PACKAGEPIN(rco[46]));
    defparam rco_obuf_46_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_46_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_46_preio (
            .PADOEN(N__94163),
            .PADOUT(N__94162),
            .PADIN(N__94161),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__74326),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_47_iopad (
            .OE(N__94154),
            .DIN(N__94153),
            .DOUT(N__94152),
            .PACKAGEPIN(rco[47]));
    defparam rco_obuf_47_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_47_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_47_preio (
            .PADOEN(N__94154),
            .PADOUT(N__94153),
            .PADIN(N__94152),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__74599),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_48_iopad (
            .OE(N__94145),
            .DIN(N__94144),
            .DOUT(N__94143),
            .PACKAGEPIN(rco[48]));
    defparam rco_obuf_48_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_48_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_48_preio (
            .PADOEN(N__94145),
            .PADOUT(N__94144),
            .PADIN(N__94143),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__93622),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_49_iopad (
            .OE(N__94136),
            .DIN(N__94135),
            .DOUT(N__94134),
            .PACKAGEPIN(rco[49]));
    defparam rco_obuf_49_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_49_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_49_preio (
            .PADOEN(N__94136),
            .PADOUT(N__94135),
            .PADIN(N__94134),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__93451),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_5_iopad (
            .OE(N__94127),
            .DIN(N__94126),
            .DOUT(N__94125),
            .PACKAGEPIN(rco[5]));
    defparam rco_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_5_preio (
            .PADOEN(N__94127),
            .PADOUT(N__94126),
            .PADIN(N__94125),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__48424),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_50_iopad (
            .OE(N__94118),
            .DIN(N__94117),
            .DOUT(N__94116),
            .PACKAGEPIN(rco[50]));
    defparam rco_obuf_50_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_50_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_50_preio (
            .PADOEN(N__94118),
            .PADOUT(N__94117),
            .PADIN(N__94116),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__88291),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_51_iopad (
            .OE(N__94109),
            .DIN(N__94108),
            .DOUT(N__94107),
            .PACKAGEPIN(rco[51]));
    defparam rco_obuf_51_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_51_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_51_preio (
            .PADOEN(N__94109),
            .PADOUT(N__94108),
            .PADIN(N__94107),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__74788),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_52_iopad (
            .OE(N__94100),
            .DIN(N__94099),
            .DOUT(N__94098),
            .PACKAGEPIN(rco[52]));
    defparam rco_obuf_52_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_52_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_52_preio (
            .PADOEN(N__94100),
            .PADOUT(N__94099),
            .PADIN(N__94098),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__74806),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_53_iopad (
            .OE(N__94091),
            .DIN(N__94090),
            .DOUT(N__94089),
            .PACKAGEPIN(rco[53]));
    defparam rco_obuf_53_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_53_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_53_preio (
            .PADOEN(N__94091),
            .PADOUT(N__94090),
            .PADIN(N__94089),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__77089),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_54_iopad (
            .OE(N__94082),
            .DIN(N__94081),
            .DOUT(N__94080),
            .PACKAGEPIN(rco[54]));
    defparam rco_obuf_54_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_54_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_54_preio (
            .PADOEN(N__94082),
            .PADOUT(N__94081),
            .PADIN(N__94080),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__68380),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_55_iopad (
            .OE(N__94073),
            .DIN(N__94072),
            .DOUT(N__94071),
            .PACKAGEPIN(rco[55]));
    defparam rco_obuf_55_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_55_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_55_preio (
            .PADOEN(N__94073),
            .PADOUT(N__94072),
            .PADIN(N__94071),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__76639),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_56_iopad (
            .OE(N__94064),
            .DIN(N__94063),
            .DOUT(N__94062),
            .PACKAGEPIN(rco[56]));
    defparam rco_obuf_56_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_56_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_56_preio (
            .PADOEN(N__94064),
            .PADOUT(N__94063),
            .PADIN(N__94062),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__76660),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_57_iopad (
            .OE(N__94055),
            .DIN(N__94054),
            .DOUT(N__94053),
            .PACKAGEPIN(rco[57]));
    defparam rco_obuf_57_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_57_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_57_preio (
            .PADOEN(N__94055),
            .PADOUT(N__94054),
            .PADIN(N__94053),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__76678),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_58_iopad (
            .OE(N__94046),
            .DIN(N__94045),
            .DOUT(N__94044),
            .PACKAGEPIN(rco[58]));
    defparam rco_obuf_58_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_58_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_58_preio (
            .PADOEN(N__94046),
            .PADOUT(N__94045),
            .PADIN(N__94044),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__66169),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_59_iopad (
            .OE(N__94037),
            .DIN(N__94036),
            .DOUT(N__94035),
            .PACKAGEPIN(rco[59]));
    defparam rco_obuf_59_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_59_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_59_preio (
            .PADOEN(N__94037),
            .PADOUT(N__94036),
            .PADIN(N__94035),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__84921),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_6_iopad (
            .OE(N__94028),
            .DIN(N__94027),
            .DOUT(N__94026),
            .PACKAGEPIN(rco[6]));
    defparam rco_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_6_preio (
            .PADOEN(N__94028),
            .PADOUT(N__94027),
            .PADIN(N__94026),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__48790),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_60_iopad (
            .OE(N__94019),
            .DIN(N__94018),
            .DOUT(N__94017),
            .PACKAGEPIN(rco[60]));
    defparam rco_obuf_60_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_60_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_60_preio (
            .PADOEN(N__94019),
            .PADOUT(N__94018),
            .PADIN(N__94017),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__75235),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_61_iopad (
            .OE(N__94010),
            .DIN(N__94009),
            .DOUT(N__94008),
            .PACKAGEPIN(rco[61]));
    defparam rco_obuf_61_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_61_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_61_preio (
            .PADOEN(N__94010),
            .PADOUT(N__94009),
            .PADIN(N__94008),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__75394),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_62_iopad (
            .OE(N__94001),
            .DIN(N__94000),
            .DOUT(N__93999),
            .PACKAGEPIN(rco[62]));
    defparam rco_obuf_62_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_62_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_62_preio (
            .PADOEN(N__94001),
            .PADOUT(N__94000),
            .PADIN(N__93999),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__75379),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_63_iopad (
            .OE(N__93992),
            .DIN(N__93991),
            .DOUT(N__93990),
            .PACKAGEPIN(rco[63]));
    defparam rco_obuf_63_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_63_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_63_preio (
            .PADOEN(N__93992),
            .PADOUT(N__93991),
            .PADIN(N__93990),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__81157),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_64_iopad (
            .OE(N__93983),
            .DIN(N__93982),
            .DOUT(N__93981),
            .PACKAGEPIN(rco[64]));
    defparam rco_obuf_64_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_64_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_64_preio (
            .PADOEN(N__93983),
            .PADOUT(N__93982),
            .PADIN(N__93981),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__81175),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_65_iopad (
            .OE(N__93974),
            .DIN(N__93973),
            .DOUT(N__93972),
            .PACKAGEPIN(rco[65]));
    defparam rco_obuf_65_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_65_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_65_preio (
            .PADOEN(N__93974),
            .PADOUT(N__93973),
            .PADIN(N__93972),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__75358),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_66_iopad (
            .OE(N__93965),
            .DIN(N__93964),
            .DOUT(N__93963),
            .PACKAGEPIN(rco[66]));
    defparam rco_obuf_66_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_66_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_66_preio (
            .PADOEN(N__93965),
            .PADOUT(N__93964),
            .PADIN(N__93963),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__90727),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_67_iopad (
            .OE(N__93956),
            .DIN(N__93955),
            .DOUT(N__93954),
            .PACKAGEPIN(rco[67]));
    defparam rco_obuf_67_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_67_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_67_preio (
            .PADOEN(N__93956),
            .PADOUT(N__93955),
            .PADIN(N__93954),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__83083),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_68_iopad (
            .OE(N__93947),
            .DIN(N__93946),
            .DOUT(N__93945),
            .PACKAGEPIN(rco[68]));
    defparam rco_obuf_68_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_68_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_68_preio (
            .PADOEN(N__93947),
            .PADOUT(N__93946),
            .PADIN(N__93945),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__83059),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_69_iopad (
            .OE(N__93938),
            .DIN(N__93937),
            .DOUT(N__93936),
            .PACKAGEPIN(rco[69]));
    defparam rco_obuf_69_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_69_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_69_preio (
            .PADOEN(N__93938),
            .PADOUT(N__93937),
            .PADIN(N__93936),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__83179),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_7_iopad (
            .OE(N__93929),
            .DIN(N__93928),
            .DOUT(N__93927),
            .PACKAGEPIN(rco[7]));
    defparam rco_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_7_preio (
            .PADOEN(N__93929),
            .PADOUT(N__93928),
            .PADIN(N__93927),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__51690),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_70_iopad (
            .OE(N__93920),
            .DIN(N__93919),
            .DOUT(N__93918),
            .PACKAGEPIN(rco[70]));
    defparam rco_obuf_70_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_70_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_70_preio (
            .PADOEN(N__93920),
            .PADOUT(N__93919),
            .PADIN(N__93918),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__84745),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_71_iopad (
            .OE(N__93911),
            .DIN(N__93910),
            .DOUT(N__93909),
            .PACKAGEPIN(rco[71]));
    defparam rco_obuf_71_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_71_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_71_preio (
            .PADOEN(N__93911),
            .PADOUT(N__93910),
            .PADIN(N__93909),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__90631),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_72_iopad (
            .OE(N__93902),
            .DIN(N__93901),
            .DOUT(N__93900),
            .PACKAGEPIN(rco[72]));
    defparam rco_obuf_72_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_72_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_72_preio (
            .PADOEN(N__93902),
            .PADOUT(N__93901),
            .PADIN(N__93900),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__89068),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_73_iopad (
            .OE(N__93893),
            .DIN(N__93892),
            .DOUT(N__93891),
            .PACKAGEPIN(rco[73]));
    defparam rco_obuf_73_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_73_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_73_preio (
            .PADOEN(N__93893),
            .PADOUT(N__93892),
            .PADIN(N__93891),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__90799),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_74_iopad (
            .OE(N__93884),
            .DIN(N__93883),
            .DOUT(N__93882),
            .PACKAGEPIN(rco[74]));
    defparam rco_obuf_74_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_74_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_74_preio (
            .PADOEN(N__93884),
            .PADOUT(N__93883),
            .PADIN(N__93882),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__88523),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_75_iopad (
            .OE(N__93875),
            .DIN(N__93874),
            .DOUT(N__93873),
            .PACKAGEPIN(rco[75]));
    defparam rco_obuf_75_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_75_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_75_preio (
            .PADOEN(N__93875),
            .PADOUT(N__93874),
            .PADIN(N__93873),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__88654),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_76_iopad (
            .OE(N__93866),
            .DIN(N__93865),
            .DOUT(N__93864),
            .PACKAGEPIN(rco[76]));
    defparam rco_obuf_76_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_76_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_76_preio (
            .PADOEN(N__93866),
            .PADOUT(N__93865),
            .PADIN(N__93864),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__88627),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_77_iopad (
            .OE(N__93857),
            .DIN(N__93856),
            .DOUT(N__93855),
            .PACKAGEPIN(rco[77]));
    defparam rco_obuf_77_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_77_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_77_preio (
            .PADOEN(N__93857),
            .PADOUT(N__93856),
            .PADIN(N__93855),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__88561),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_78_iopad (
            .OE(N__93848),
            .DIN(N__93847),
            .DOUT(N__93846),
            .PACKAGEPIN(rco[78]));
    defparam rco_obuf_78_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_78_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_78_preio (
            .PADOEN(N__93848),
            .PADOUT(N__93847),
            .PADIN(N__93846),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__84529),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_79_iopad (
            .OE(N__93839),
            .DIN(N__93838),
            .DOUT(N__93837),
            .PACKAGEPIN(rco[79]));
    defparam rco_obuf_79_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_79_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_79_preio (
            .PADOEN(N__93839),
            .PADOUT(N__93838),
            .PADIN(N__93837),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__84445),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_8_iopad (
            .OE(N__93830),
            .DIN(N__93829),
            .DOUT(N__93828),
            .PACKAGEPIN(rco[8]));
    defparam rco_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_8_preio (
            .PADOEN(N__93830),
            .PADOUT(N__93829),
            .PADIN(N__93828),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__52641),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_80_iopad (
            .OE(N__93821),
            .DIN(N__93820),
            .DOUT(N__93819),
            .PACKAGEPIN(rco[80]));
    defparam rco_obuf_80_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_80_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_80_preio (
            .PADOEN(N__93821),
            .PADOUT(N__93820),
            .PADIN(N__93819),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__88417),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_81_iopad (
            .OE(N__93812),
            .DIN(N__93811),
            .DOUT(N__93810),
            .PACKAGEPIN(rco[81]));
    defparam rco_obuf_81_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_81_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_81_preio (
            .PADOEN(N__93812),
            .PADOUT(N__93811),
            .PADIN(N__93810),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__84433),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_82_iopad (
            .OE(N__93803),
            .DIN(N__93802),
            .DOUT(N__93801),
            .PACKAGEPIN(rco[82]));
    defparam rco_obuf_82_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_82_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_82_preio (
            .PADOEN(N__93803),
            .PADOUT(N__93802),
            .PADIN(N__93801),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__80893),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_83_iopad (
            .OE(N__93794),
            .DIN(N__93793),
            .DOUT(N__93792),
            .PACKAGEPIN(rco[83]));
    defparam rco_obuf_83_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_83_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_83_preio (
            .PADOEN(N__93794),
            .PADOUT(N__93793),
            .PADIN(N__93792),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__68533),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_84_iopad (
            .OE(N__93785),
            .DIN(N__93784),
            .DOUT(N__93783),
            .PACKAGEPIN(rco[84]));
    defparam rco_obuf_84_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_84_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_84_preio (
            .PADOEN(N__93785),
            .PADOUT(N__93784),
            .PADIN(N__93783),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__68626),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_85_iopad (
            .OE(N__93776),
            .DIN(N__93775),
            .DOUT(N__93774),
            .PACKAGEPIN(rco[85]));
    defparam rco_obuf_85_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_85_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_85_preio (
            .PADOEN(N__93776),
            .PADOUT(N__93775),
            .PADIN(N__93774),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__66157),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_86_iopad (
            .OE(N__93767),
            .DIN(N__93766),
            .DOUT(N__93765),
            .PACKAGEPIN(rco[86]));
    defparam rco_obuf_86_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_86_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_86_preio (
            .PADOEN(N__93767),
            .PADOUT(N__93766),
            .PADIN(N__93765),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__61012),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_87_iopad (
            .OE(N__93758),
            .DIN(N__93757),
            .DOUT(N__93756),
            .PACKAGEPIN(rco[87]));
    defparam rco_obuf_87_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_87_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_87_preio (
            .PADOEN(N__93758),
            .PADOUT(N__93757),
            .PADIN(N__93756),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__61024),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_88_iopad (
            .OE(N__93749),
            .DIN(N__93748),
            .DOUT(N__93747),
            .PACKAGEPIN(rco[88]));
    defparam rco_obuf_88_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_88_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_88_preio (
            .PADOEN(N__93749),
            .PADOUT(N__93748),
            .PADIN(N__93747),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__62908),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_89_iopad (
            .OE(N__93740),
            .DIN(N__93739),
            .DOUT(N__93738),
            .PACKAGEPIN(rco[89]));
    defparam rco_obuf_89_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_89_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_89_preio (
            .PADOEN(N__93740),
            .PADOUT(N__93739),
            .PADIN(N__93738),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__68572),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_9_iopad (
            .OE(N__93731),
            .DIN(N__93730),
            .DOUT(N__93729),
            .PACKAGEPIN(rco[9]));
    defparam rco_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_9_preio (
            .PADOEN(N__93731),
            .PADOUT(N__93730),
            .PADIN(N__93729),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__69193),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_90_iopad (
            .OE(N__93722),
            .DIN(N__93721),
            .DOUT(N__93720),
            .PACKAGEPIN(rco[90]));
    defparam rco_obuf_90_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_90_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_90_preio (
            .PADOEN(N__93722),
            .PADOUT(N__93721),
            .PADIN(N__93720),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__64162),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_91_iopad (
            .OE(N__93713),
            .DIN(N__93712),
            .DOUT(N__93711),
            .PACKAGEPIN(rco[91]));
    defparam rco_obuf_91_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_91_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_91_preio (
            .PADOEN(N__93713),
            .PADOUT(N__93712),
            .PADIN(N__93711),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__64150),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_92_iopad (
            .OE(N__93704),
            .DIN(N__93703),
            .DOUT(N__93702),
            .PACKAGEPIN(rco[92]));
    defparam rco_obuf_92_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_92_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_92_preio (
            .PADOEN(N__93704),
            .PADOUT(N__93703),
            .PADIN(N__93702),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__68431),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_93_iopad (
            .OE(N__93695),
            .DIN(N__93694),
            .DOUT(N__93693),
            .PACKAGEPIN(rco[93]));
    defparam rco_obuf_93_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_93_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_93_preio (
            .PADOEN(N__93695),
            .PADOUT(N__93694),
            .PADIN(N__93693),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__72796),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_94_iopad (
            .OE(N__93686),
            .DIN(N__93685),
            .DOUT(N__93684),
            .PACKAGEPIN(rco[94]));
    defparam rco_obuf_94_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_94_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_94_preio (
            .PADOEN(N__93686),
            .PADOUT(N__93685),
            .PADIN(N__93684),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__72532),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_95_iopad (
            .OE(N__93677),
            .DIN(N__93676),
            .DOUT(N__93675),
            .PACKAGEPIN(rco[95]));
    defparam rco_obuf_95_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_95_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_95_preio (
            .PADOEN(N__93677),
            .PADOUT(N__93676),
            .PADIN(N__93675),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__72841),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_96_iopad (
            .OE(N__93668),
            .DIN(N__93667),
            .DOUT(N__93666),
            .PACKAGEPIN(rco[96]));
    defparam rco_obuf_96_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_96_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_96_preio (
            .PADOEN(N__93668),
            .PADOUT(N__93667),
            .PADIN(N__93666),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__68815),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_97_iopad (
            .OE(N__93659),
            .DIN(N__93658),
            .DOUT(N__93657),
            .PACKAGEPIN(rco[97]));
    defparam rco_obuf_97_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_97_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_97_preio (
            .PADOEN(N__93659),
            .PADOUT(N__93658),
            .PADIN(N__93657),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__67216),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_98_iopad (
            .OE(N__93650),
            .DIN(N__93649),
            .DOUT(N__93648),
            .PACKAGEPIN(rco[98]));
    defparam rco_obuf_98_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_98_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_98_preio (
            .PADOEN(N__93650),
            .PADOUT(N__93649),
            .PADIN(N__93648),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__72736),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rco_obuf_99_iopad (
            .OE(N__93641),
            .DIN(N__93640),
            .DOUT(N__93639),
            .PACKAGEPIN(rco[99]));
    defparam rco_obuf_99_preio.NEG_TRIGGER=1'b0;
    defparam rco_obuf_99_preio.PIN_TYPE=6'b011001;
    PRE_IO rco_obuf_99_preio (
            .PADOEN(N__93641),
            .PADOUT(N__93640),
            .PADIN(N__93639),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__79567),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IoInMux I__19184 (
            .O(N__93622),
            .I(N__93619));
    LocalMux I__19183 (
            .O(N__93619),
            .I(N__93616));
    IoSpan4Mux I__19182 (
            .O(N__93616),
            .I(N__93612));
    InMux I__19181 (
            .O(N__93615),
            .I(N__93609));
    Span4Mux_s0_h I__19180 (
            .O(N__93612),
            .I(N__93604));
    LocalMux I__19179 (
            .O(N__93609),
            .I(N__93604));
    Span4Mux_h I__19178 (
            .O(N__93604),
            .I(N__93600));
    InMux I__19177 (
            .O(N__93603),
            .I(N__93597));
    Span4Mux_v I__19176 (
            .O(N__93600),
            .I(N__93588));
    LocalMux I__19175 (
            .O(N__93597),
            .I(N__93588));
    InMux I__19174 (
            .O(N__93596),
            .I(N__93584));
    InMux I__19173 (
            .O(N__93595),
            .I(N__93577));
    InMux I__19172 (
            .O(N__93594),
            .I(N__93577));
    InMux I__19171 (
            .O(N__93593),
            .I(N__93577));
    Span4Mux_v I__19170 (
            .O(N__93588),
            .I(N__93573));
    InMux I__19169 (
            .O(N__93587),
            .I(N__93570));
    LocalMux I__19168 (
            .O(N__93584),
            .I(N__93567));
    LocalMux I__19167 (
            .O(N__93577),
            .I(N__93561));
    CascadeMux I__19166 (
            .O(N__93576),
            .I(N__93558));
    Sp12to4 I__19165 (
            .O(N__93573),
            .I(N__93549));
    LocalMux I__19164 (
            .O(N__93570),
            .I(N__93544));
    Span4Mux_h I__19163 (
            .O(N__93567),
            .I(N__93544));
    InMux I__19162 (
            .O(N__93566),
            .I(N__93541));
    InMux I__19161 (
            .O(N__93565),
            .I(N__93538));
    InMux I__19160 (
            .O(N__93564),
            .I(N__93535));
    Span4Mux_v I__19159 (
            .O(N__93561),
            .I(N__93532));
    InMux I__19158 (
            .O(N__93558),
            .I(N__93521));
    InMux I__19157 (
            .O(N__93557),
            .I(N__93521));
    InMux I__19156 (
            .O(N__93556),
            .I(N__93521));
    InMux I__19155 (
            .O(N__93555),
            .I(N__93521));
    InMux I__19154 (
            .O(N__93554),
            .I(N__93521));
    InMux I__19153 (
            .O(N__93553),
            .I(N__93516));
    InMux I__19152 (
            .O(N__93552),
            .I(N__93516));
    Odrv12 I__19151 (
            .O(N__93549),
            .I(rco_c_48));
    Odrv4 I__19150 (
            .O(N__93544),
            .I(rco_c_48));
    LocalMux I__19149 (
            .O(N__93541),
            .I(rco_c_48));
    LocalMux I__19148 (
            .O(N__93538),
            .I(rco_c_48));
    LocalMux I__19147 (
            .O(N__93535),
            .I(rco_c_48));
    Odrv4 I__19146 (
            .O(N__93532),
            .I(rco_c_48));
    LocalMux I__19145 (
            .O(N__93521),
            .I(rco_c_48));
    LocalMux I__19144 (
            .O(N__93516),
            .I(rco_c_48));
    InMux I__19143 (
            .O(N__93499),
            .I(N__93496));
    LocalMux I__19142 (
            .O(N__93496),
            .I(N__93492));
    InMux I__19141 (
            .O(N__93495),
            .I(N__93488));
    Span12Mux_v I__19140 (
            .O(N__93492),
            .I(N__93485));
    InMux I__19139 (
            .O(N__93491),
            .I(N__93482));
    LocalMux I__19138 (
            .O(N__93488),
            .I(N__93479));
    Span12Mux_h I__19137 (
            .O(N__93485),
            .I(N__93474));
    LocalMux I__19136 (
            .O(N__93482),
            .I(N__93471));
    Span4Mux_h I__19135 (
            .O(N__93479),
            .I(N__93468));
    InMux I__19134 (
            .O(N__93478),
            .I(N__93465));
    InMux I__19133 (
            .O(N__93477),
            .I(N__93462));
    Odrv12 I__19132 (
            .O(N__93474),
            .I(shift_srl_49Z0Z_15));
    Odrv4 I__19131 (
            .O(N__93471),
            .I(shift_srl_49Z0Z_15));
    Odrv4 I__19130 (
            .O(N__93468),
            .I(shift_srl_49Z0Z_15));
    LocalMux I__19129 (
            .O(N__93465),
            .I(shift_srl_49Z0Z_15));
    LocalMux I__19128 (
            .O(N__93462),
            .I(shift_srl_49Z0Z_15));
    IoInMux I__19127 (
            .O(N__93451),
            .I(N__93448));
    LocalMux I__19126 (
            .O(N__93448),
            .I(rco_c_49));
    InMux I__19125 (
            .O(N__93445),
            .I(N__93442));
    LocalMux I__19124 (
            .O(N__93442),
            .I(N__93439));
    Odrv12 I__19123 (
            .O(N__93439),
            .I(shift_srl_37Z0Z_10));
    InMux I__19122 (
            .O(N__93436),
            .I(N__93433));
    LocalMux I__19121 (
            .O(N__93433),
            .I(N__93430));
    Odrv12 I__19120 (
            .O(N__93430),
            .I(shift_srl_37Z0Z_11));
    ClkMux I__19119 (
            .O(N__93427),
            .I(N__91864));
    ClkMux I__19118 (
            .O(N__93426),
            .I(N__91864));
    ClkMux I__19117 (
            .O(N__93425),
            .I(N__91864));
    ClkMux I__19116 (
            .O(N__93424),
            .I(N__91864));
    ClkMux I__19115 (
            .O(N__93423),
            .I(N__91864));
    ClkMux I__19114 (
            .O(N__93422),
            .I(N__91864));
    ClkMux I__19113 (
            .O(N__93421),
            .I(N__91864));
    ClkMux I__19112 (
            .O(N__93420),
            .I(N__91864));
    ClkMux I__19111 (
            .O(N__93419),
            .I(N__91864));
    ClkMux I__19110 (
            .O(N__93418),
            .I(N__91864));
    ClkMux I__19109 (
            .O(N__93417),
            .I(N__91864));
    ClkMux I__19108 (
            .O(N__93416),
            .I(N__91864));
    ClkMux I__19107 (
            .O(N__93415),
            .I(N__91864));
    ClkMux I__19106 (
            .O(N__93414),
            .I(N__91864));
    ClkMux I__19105 (
            .O(N__93413),
            .I(N__91864));
    ClkMux I__19104 (
            .O(N__93412),
            .I(N__91864));
    ClkMux I__19103 (
            .O(N__93411),
            .I(N__91864));
    ClkMux I__19102 (
            .O(N__93410),
            .I(N__91864));
    ClkMux I__19101 (
            .O(N__93409),
            .I(N__91864));
    ClkMux I__19100 (
            .O(N__93408),
            .I(N__91864));
    ClkMux I__19099 (
            .O(N__93407),
            .I(N__91864));
    ClkMux I__19098 (
            .O(N__93406),
            .I(N__91864));
    ClkMux I__19097 (
            .O(N__93405),
            .I(N__91864));
    ClkMux I__19096 (
            .O(N__93404),
            .I(N__91864));
    ClkMux I__19095 (
            .O(N__93403),
            .I(N__91864));
    ClkMux I__19094 (
            .O(N__93402),
            .I(N__91864));
    ClkMux I__19093 (
            .O(N__93401),
            .I(N__91864));
    ClkMux I__19092 (
            .O(N__93400),
            .I(N__91864));
    ClkMux I__19091 (
            .O(N__93399),
            .I(N__91864));
    ClkMux I__19090 (
            .O(N__93398),
            .I(N__91864));
    ClkMux I__19089 (
            .O(N__93397),
            .I(N__91864));
    ClkMux I__19088 (
            .O(N__93396),
            .I(N__91864));
    ClkMux I__19087 (
            .O(N__93395),
            .I(N__91864));
    ClkMux I__19086 (
            .O(N__93394),
            .I(N__91864));
    ClkMux I__19085 (
            .O(N__93393),
            .I(N__91864));
    ClkMux I__19084 (
            .O(N__93392),
            .I(N__91864));
    ClkMux I__19083 (
            .O(N__93391),
            .I(N__91864));
    ClkMux I__19082 (
            .O(N__93390),
            .I(N__91864));
    ClkMux I__19081 (
            .O(N__93389),
            .I(N__91864));
    ClkMux I__19080 (
            .O(N__93388),
            .I(N__91864));
    ClkMux I__19079 (
            .O(N__93387),
            .I(N__91864));
    ClkMux I__19078 (
            .O(N__93386),
            .I(N__91864));
    ClkMux I__19077 (
            .O(N__93385),
            .I(N__91864));
    ClkMux I__19076 (
            .O(N__93384),
            .I(N__91864));
    ClkMux I__19075 (
            .O(N__93383),
            .I(N__91864));
    ClkMux I__19074 (
            .O(N__93382),
            .I(N__91864));
    ClkMux I__19073 (
            .O(N__93381),
            .I(N__91864));
    ClkMux I__19072 (
            .O(N__93380),
            .I(N__91864));
    ClkMux I__19071 (
            .O(N__93379),
            .I(N__91864));
    ClkMux I__19070 (
            .O(N__93378),
            .I(N__91864));
    ClkMux I__19069 (
            .O(N__93377),
            .I(N__91864));
    ClkMux I__19068 (
            .O(N__93376),
            .I(N__91864));
    ClkMux I__19067 (
            .O(N__93375),
            .I(N__91864));
    ClkMux I__19066 (
            .O(N__93374),
            .I(N__91864));
    ClkMux I__19065 (
            .O(N__93373),
            .I(N__91864));
    ClkMux I__19064 (
            .O(N__93372),
            .I(N__91864));
    ClkMux I__19063 (
            .O(N__93371),
            .I(N__91864));
    ClkMux I__19062 (
            .O(N__93370),
            .I(N__91864));
    ClkMux I__19061 (
            .O(N__93369),
            .I(N__91864));
    ClkMux I__19060 (
            .O(N__93368),
            .I(N__91864));
    ClkMux I__19059 (
            .O(N__93367),
            .I(N__91864));
    ClkMux I__19058 (
            .O(N__93366),
            .I(N__91864));
    ClkMux I__19057 (
            .O(N__93365),
            .I(N__91864));
    ClkMux I__19056 (
            .O(N__93364),
            .I(N__91864));
    ClkMux I__19055 (
            .O(N__93363),
            .I(N__91864));
    ClkMux I__19054 (
            .O(N__93362),
            .I(N__91864));
    ClkMux I__19053 (
            .O(N__93361),
            .I(N__91864));
    ClkMux I__19052 (
            .O(N__93360),
            .I(N__91864));
    ClkMux I__19051 (
            .O(N__93359),
            .I(N__91864));
    ClkMux I__19050 (
            .O(N__93358),
            .I(N__91864));
    ClkMux I__19049 (
            .O(N__93357),
            .I(N__91864));
    ClkMux I__19048 (
            .O(N__93356),
            .I(N__91864));
    ClkMux I__19047 (
            .O(N__93355),
            .I(N__91864));
    ClkMux I__19046 (
            .O(N__93354),
            .I(N__91864));
    ClkMux I__19045 (
            .O(N__93353),
            .I(N__91864));
    ClkMux I__19044 (
            .O(N__93352),
            .I(N__91864));
    ClkMux I__19043 (
            .O(N__93351),
            .I(N__91864));
    ClkMux I__19042 (
            .O(N__93350),
            .I(N__91864));
    ClkMux I__19041 (
            .O(N__93349),
            .I(N__91864));
    ClkMux I__19040 (
            .O(N__93348),
            .I(N__91864));
    ClkMux I__19039 (
            .O(N__93347),
            .I(N__91864));
    ClkMux I__19038 (
            .O(N__93346),
            .I(N__91864));
    ClkMux I__19037 (
            .O(N__93345),
            .I(N__91864));
    ClkMux I__19036 (
            .O(N__93344),
            .I(N__91864));
    ClkMux I__19035 (
            .O(N__93343),
            .I(N__91864));
    ClkMux I__19034 (
            .O(N__93342),
            .I(N__91864));
    ClkMux I__19033 (
            .O(N__93341),
            .I(N__91864));
    ClkMux I__19032 (
            .O(N__93340),
            .I(N__91864));
    ClkMux I__19031 (
            .O(N__93339),
            .I(N__91864));
    ClkMux I__19030 (
            .O(N__93338),
            .I(N__91864));
    ClkMux I__19029 (
            .O(N__93337),
            .I(N__91864));
    ClkMux I__19028 (
            .O(N__93336),
            .I(N__91864));
    ClkMux I__19027 (
            .O(N__93335),
            .I(N__91864));
    ClkMux I__19026 (
            .O(N__93334),
            .I(N__91864));
    ClkMux I__19025 (
            .O(N__93333),
            .I(N__91864));
    ClkMux I__19024 (
            .O(N__93332),
            .I(N__91864));
    ClkMux I__19023 (
            .O(N__93331),
            .I(N__91864));
    ClkMux I__19022 (
            .O(N__93330),
            .I(N__91864));
    ClkMux I__19021 (
            .O(N__93329),
            .I(N__91864));
    ClkMux I__19020 (
            .O(N__93328),
            .I(N__91864));
    ClkMux I__19019 (
            .O(N__93327),
            .I(N__91864));
    ClkMux I__19018 (
            .O(N__93326),
            .I(N__91864));
    ClkMux I__19017 (
            .O(N__93325),
            .I(N__91864));
    ClkMux I__19016 (
            .O(N__93324),
            .I(N__91864));
    ClkMux I__19015 (
            .O(N__93323),
            .I(N__91864));
    ClkMux I__19014 (
            .O(N__93322),
            .I(N__91864));
    ClkMux I__19013 (
            .O(N__93321),
            .I(N__91864));
    ClkMux I__19012 (
            .O(N__93320),
            .I(N__91864));
    ClkMux I__19011 (
            .O(N__93319),
            .I(N__91864));
    ClkMux I__19010 (
            .O(N__93318),
            .I(N__91864));
    ClkMux I__19009 (
            .O(N__93317),
            .I(N__91864));
    ClkMux I__19008 (
            .O(N__93316),
            .I(N__91864));
    ClkMux I__19007 (
            .O(N__93315),
            .I(N__91864));
    ClkMux I__19006 (
            .O(N__93314),
            .I(N__91864));
    ClkMux I__19005 (
            .O(N__93313),
            .I(N__91864));
    ClkMux I__19004 (
            .O(N__93312),
            .I(N__91864));
    ClkMux I__19003 (
            .O(N__93311),
            .I(N__91864));
    ClkMux I__19002 (
            .O(N__93310),
            .I(N__91864));
    ClkMux I__19001 (
            .O(N__93309),
            .I(N__91864));
    ClkMux I__19000 (
            .O(N__93308),
            .I(N__91864));
    ClkMux I__18999 (
            .O(N__93307),
            .I(N__91864));
    ClkMux I__18998 (
            .O(N__93306),
            .I(N__91864));
    ClkMux I__18997 (
            .O(N__93305),
            .I(N__91864));
    ClkMux I__18996 (
            .O(N__93304),
            .I(N__91864));
    ClkMux I__18995 (
            .O(N__93303),
            .I(N__91864));
    ClkMux I__18994 (
            .O(N__93302),
            .I(N__91864));
    ClkMux I__18993 (
            .O(N__93301),
            .I(N__91864));
    ClkMux I__18992 (
            .O(N__93300),
            .I(N__91864));
    ClkMux I__18991 (
            .O(N__93299),
            .I(N__91864));
    ClkMux I__18990 (
            .O(N__93298),
            .I(N__91864));
    ClkMux I__18989 (
            .O(N__93297),
            .I(N__91864));
    ClkMux I__18988 (
            .O(N__93296),
            .I(N__91864));
    ClkMux I__18987 (
            .O(N__93295),
            .I(N__91864));
    ClkMux I__18986 (
            .O(N__93294),
            .I(N__91864));
    ClkMux I__18985 (
            .O(N__93293),
            .I(N__91864));
    ClkMux I__18984 (
            .O(N__93292),
            .I(N__91864));
    ClkMux I__18983 (
            .O(N__93291),
            .I(N__91864));
    ClkMux I__18982 (
            .O(N__93290),
            .I(N__91864));
    ClkMux I__18981 (
            .O(N__93289),
            .I(N__91864));
    ClkMux I__18980 (
            .O(N__93288),
            .I(N__91864));
    ClkMux I__18979 (
            .O(N__93287),
            .I(N__91864));
    ClkMux I__18978 (
            .O(N__93286),
            .I(N__91864));
    ClkMux I__18977 (
            .O(N__93285),
            .I(N__91864));
    ClkMux I__18976 (
            .O(N__93284),
            .I(N__91864));
    ClkMux I__18975 (
            .O(N__93283),
            .I(N__91864));
    ClkMux I__18974 (
            .O(N__93282),
            .I(N__91864));
    ClkMux I__18973 (
            .O(N__93281),
            .I(N__91864));
    ClkMux I__18972 (
            .O(N__93280),
            .I(N__91864));
    ClkMux I__18971 (
            .O(N__93279),
            .I(N__91864));
    ClkMux I__18970 (
            .O(N__93278),
            .I(N__91864));
    ClkMux I__18969 (
            .O(N__93277),
            .I(N__91864));
    ClkMux I__18968 (
            .O(N__93276),
            .I(N__91864));
    ClkMux I__18967 (
            .O(N__93275),
            .I(N__91864));
    ClkMux I__18966 (
            .O(N__93274),
            .I(N__91864));
    ClkMux I__18965 (
            .O(N__93273),
            .I(N__91864));
    ClkMux I__18964 (
            .O(N__93272),
            .I(N__91864));
    ClkMux I__18963 (
            .O(N__93271),
            .I(N__91864));
    ClkMux I__18962 (
            .O(N__93270),
            .I(N__91864));
    ClkMux I__18961 (
            .O(N__93269),
            .I(N__91864));
    ClkMux I__18960 (
            .O(N__93268),
            .I(N__91864));
    ClkMux I__18959 (
            .O(N__93267),
            .I(N__91864));
    ClkMux I__18958 (
            .O(N__93266),
            .I(N__91864));
    ClkMux I__18957 (
            .O(N__93265),
            .I(N__91864));
    ClkMux I__18956 (
            .O(N__93264),
            .I(N__91864));
    ClkMux I__18955 (
            .O(N__93263),
            .I(N__91864));
    ClkMux I__18954 (
            .O(N__93262),
            .I(N__91864));
    ClkMux I__18953 (
            .O(N__93261),
            .I(N__91864));
    ClkMux I__18952 (
            .O(N__93260),
            .I(N__91864));
    ClkMux I__18951 (
            .O(N__93259),
            .I(N__91864));
    ClkMux I__18950 (
            .O(N__93258),
            .I(N__91864));
    ClkMux I__18949 (
            .O(N__93257),
            .I(N__91864));
    ClkMux I__18948 (
            .O(N__93256),
            .I(N__91864));
    ClkMux I__18947 (
            .O(N__93255),
            .I(N__91864));
    ClkMux I__18946 (
            .O(N__93254),
            .I(N__91864));
    ClkMux I__18945 (
            .O(N__93253),
            .I(N__91864));
    ClkMux I__18944 (
            .O(N__93252),
            .I(N__91864));
    ClkMux I__18943 (
            .O(N__93251),
            .I(N__91864));
    ClkMux I__18942 (
            .O(N__93250),
            .I(N__91864));
    ClkMux I__18941 (
            .O(N__93249),
            .I(N__91864));
    ClkMux I__18940 (
            .O(N__93248),
            .I(N__91864));
    ClkMux I__18939 (
            .O(N__93247),
            .I(N__91864));
    ClkMux I__18938 (
            .O(N__93246),
            .I(N__91864));
    ClkMux I__18937 (
            .O(N__93245),
            .I(N__91864));
    ClkMux I__18936 (
            .O(N__93244),
            .I(N__91864));
    ClkMux I__18935 (
            .O(N__93243),
            .I(N__91864));
    ClkMux I__18934 (
            .O(N__93242),
            .I(N__91864));
    ClkMux I__18933 (
            .O(N__93241),
            .I(N__91864));
    ClkMux I__18932 (
            .O(N__93240),
            .I(N__91864));
    ClkMux I__18931 (
            .O(N__93239),
            .I(N__91864));
    ClkMux I__18930 (
            .O(N__93238),
            .I(N__91864));
    ClkMux I__18929 (
            .O(N__93237),
            .I(N__91864));
    ClkMux I__18928 (
            .O(N__93236),
            .I(N__91864));
    ClkMux I__18927 (
            .O(N__93235),
            .I(N__91864));
    ClkMux I__18926 (
            .O(N__93234),
            .I(N__91864));
    ClkMux I__18925 (
            .O(N__93233),
            .I(N__91864));
    ClkMux I__18924 (
            .O(N__93232),
            .I(N__91864));
    ClkMux I__18923 (
            .O(N__93231),
            .I(N__91864));
    ClkMux I__18922 (
            .O(N__93230),
            .I(N__91864));
    ClkMux I__18921 (
            .O(N__93229),
            .I(N__91864));
    ClkMux I__18920 (
            .O(N__93228),
            .I(N__91864));
    ClkMux I__18919 (
            .O(N__93227),
            .I(N__91864));
    ClkMux I__18918 (
            .O(N__93226),
            .I(N__91864));
    ClkMux I__18917 (
            .O(N__93225),
            .I(N__91864));
    ClkMux I__18916 (
            .O(N__93224),
            .I(N__91864));
    ClkMux I__18915 (
            .O(N__93223),
            .I(N__91864));
    ClkMux I__18914 (
            .O(N__93222),
            .I(N__91864));
    ClkMux I__18913 (
            .O(N__93221),
            .I(N__91864));
    ClkMux I__18912 (
            .O(N__93220),
            .I(N__91864));
    ClkMux I__18911 (
            .O(N__93219),
            .I(N__91864));
    ClkMux I__18910 (
            .O(N__93218),
            .I(N__91864));
    ClkMux I__18909 (
            .O(N__93217),
            .I(N__91864));
    ClkMux I__18908 (
            .O(N__93216),
            .I(N__91864));
    ClkMux I__18907 (
            .O(N__93215),
            .I(N__91864));
    ClkMux I__18906 (
            .O(N__93214),
            .I(N__91864));
    ClkMux I__18905 (
            .O(N__93213),
            .I(N__91864));
    ClkMux I__18904 (
            .O(N__93212),
            .I(N__91864));
    ClkMux I__18903 (
            .O(N__93211),
            .I(N__91864));
    ClkMux I__18902 (
            .O(N__93210),
            .I(N__91864));
    ClkMux I__18901 (
            .O(N__93209),
            .I(N__91864));
    ClkMux I__18900 (
            .O(N__93208),
            .I(N__91864));
    ClkMux I__18899 (
            .O(N__93207),
            .I(N__91864));
    ClkMux I__18898 (
            .O(N__93206),
            .I(N__91864));
    ClkMux I__18897 (
            .O(N__93205),
            .I(N__91864));
    ClkMux I__18896 (
            .O(N__93204),
            .I(N__91864));
    ClkMux I__18895 (
            .O(N__93203),
            .I(N__91864));
    ClkMux I__18894 (
            .O(N__93202),
            .I(N__91864));
    ClkMux I__18893 (
            .O(N__93201),
            .I(N__91864));
    ClkMux I__18892 (
            .O(N__93200),
            .I(N__91864));
    ClkMux I__18891 (
            .O(N__93199),
            .I(N__91864));
    ClkMux I__18890 (
            .O(N__93198),
            .I(N__91864));
    ClkMux I__18889 (
            .O(N__93197),
            .I(N__91864));
    ClkMux I__18888 (
            .O(N__93196),
            .I(N__91864));
    ClkMux I__18887 (
            .O(N__93195),
            .I(N__91864));
    ClkMux I__18886 (
            .O(N__93194),
            .I(N__91864));
    ClkMux I__18885 (
            .O(N__93193),
            .I(N__91864));
    ClkMux I__18884 (
            .O(N__93192),
            .I(N__91864));
    ClkMux I__18883 (
            .O(N__93191),
            .I(N__91864));
    ClkMux I__18882 (
            .O(N__93190),
            .I(N__91864));
    ClkMux I__18881 (
            .O(N__93189),
            .I(N__91864));
    ClkMux I__18880 (
            .O(N__93188),
            .I(N__91864));
    ClkMux I__18879 (
            .O(N__93187),
            .I(N__91864));
    ClkMux I__18878 (
            .O(N__93186),
            .I(N__91864));
    ClkMux I__18877 (
            .O(N__93185),
            .I(N__91864));
    ClkMux I__18876 (
            .O(N__93184),
            .I(N__91864));
    ClkMux I__18875 (
            .O(N__93183),
            .I(N__91864));
    ClkMux I__18874 (
            .O(N__93182),
            .I(N__91864));
    ClkMux I__18873 (
            .O(N__93181),
            .I(N__91864));
    ClkMux I__18872 (
            .O(N__93180),
            .I(N__91864));
    ClkMux I__18871 (
            .O(N__93179),
            .I(N__91864));
    ClkMux I__18870 (
            .O(N__93178),
            .I(N__91864));
    ClkMux I__18869 (
            .O(N__93177),
            .I(N__91864));
    ClkMux I__18868 (
            .O(N__93176),
            .I(N__91864));
    ClkMux I__18867 (
            .O(N__93175),
            .I(N__91864));
    ClkMux I__18866 (
            .O(N__93174),
            .I(N__91864));
    ClkMux I__18865 (
            .O(N__93173),
            .I(N__91864));
    ClkMux I__18864 (
            .O(N__93172),
            .I(N__91864));
    ClkMux I__18863 (
            .O(N__93171),
            .I(N__91864));
    ClkMux I__18862 (
            .O(N__93170),
            .I(N__91864));
    ClkMux I__18861 (
            .O(N__93169),
            .I(N__91864));
    ClkMux I__18860 (
            .O(N__93168),
            .I(N__91864));
    ClkMux I__18859 (
            .O(N__93167),
            .I(N__91864));
    ClkMux I__18858 (
            .O(N__93166),
            .I(N__91864));
    ClkMux I__18857 (
            .O(N__93165),
            .I(N__91864));
    ClkMux I__18856 (
            .O(N__93164),
            .I(N__91864));
    ClkMux I__18855 (
            .O(N__93163),
            .I(N__91864));
    ClkMux I__18854 (
            .O(N__93162),
            .I(N__91864));
    ClkMux I__18853 (
            .O(N__93161),
            .I(N__91864));
    ClkMux I__18852 (
            .O(N__93160),
            .I(N__91864));
    ClkMux I__18851 (
            .O(N__93159),
            .I(N__91864));
    ClkMux I__18850 (
            .O(N__93158),
            .I(N__91864));
    ClkMux I__18849 (
            .O(N__93157),
            .I(N__91864));
    ClkMux I__18848 (
            .O(N__93156),
            .I(N__91864));
    ClkMux I__18847 (
            .O(N__93155),
            .I(N__91864));
    ClkMux I__18846 (
            .O(N__93154),
            .I(N__91864));
    ClkMux I__18845 (
            .O(N__93153),
            .I(N__91864));
    ClkMux I__18844 (
            .O(N__93152),
            .I(N__91864));
    ClkMux I__18843 (
            .O(N__93151),
            .I(N__91864));
    ClkMux I__18842 (
            .O(N__93150),
            .I(N__91864));
    ClkMux I__18841 (
            .O(N__93149),
            .I(N__91864));
    ClkMux I__18840 (
            .O(N__93148),
            .I(N__91864));
    ClkMux I__18839 (
            .O(N__93147),
            .I(N__91864));
    ClkMux I__18838 (
            .O(N__93146),
            .I(N__91864));
    ClkMux I__18837 (
            .O(N__93145),
            .I(N__91864));
    ClkMux I__18836 (
            .O(N__93144),
            .I(N__91864));
    ClkMux I__18835 (
            .O(N__93143),
            .I(N__91864));
    ClkMux I__18834 (
            .O(N__93142),
            .I(N__91864));
    ClkMux I__18833 (
            .O(N__93141),
            .I(N__91864));
    ClkMux I__18832 (
            .O(N__93140),
            .I(N__91864));
    ClkMux I__18831 (
            .O(N__93139),
            .I(N__91864));
    ClkMux I__18830 (
            .O(N__93138),
            .I(N__91864));
    ClkMux I__18829 (
            .O(N__93137),
            .I(N__91864));
    ClkMux I__18828 (
            .O(N__93136),
            .I(N__91864));
    ClkMux I__18827 (
            .O(N__93135),
            .I(N__91864));
    ClkMux I__18826 (
            .O(N__93134),
            .I(N__91864));
    ClkMux I__18825 (
            .O(N__93133),
            .I(N__91864));
    ClkMux I__18824 (
            .O(N__93132),
            .I(N__91864));
    ClkMux I__18823 (
            .O(N__93131),
            .I(N__91864));
    ClkMux I__18822 (
            .O(N__93130),
            .I(N__91864));
    ClkMux I__18821 (
            .O(N__93129),
            .I(N__91864));
    ClkMux I__18820 (
            .O(N__93128),
            .I(N__91864));
    ClkMux I__18819 (
            .O(N__93127),
            .I(N__91864));
    ClkMux I__18818 (
            .O(N__93126),
            .I(N__91864));
    ClkMux I__18817 (
            .O(N__93125),
            .I(N__91864));
    ClkMux I__18816 (
            .O(N__93124),
            .I(N__91864));
    ClkMux I__18815 (
            .O(N__93123),
            .I(N__91864));
    ClkMux I__18814 (
            .O(N__93122),
            .I(N__91864));
    ClkMux I__18813 (
            .O(N__93121),
            .I(N__91864));
    ClkMux I__18812 (
            .O(N__93120),
            .I(N__91864));
    ClkMux I__18811 (
            .O(N__93119),
            .I(N__91864));
    ClkMux I__18810 (
            .O(N__93118),
            .I(N__91864));
    ClkMux I__18809 (
            .O(N__93117),
            .I(N__91864));
    ClkMux I__18808 (
            .O(N__93116),
            .I(N__91864));
    ClkMux I__18807 (
            .O(N__93115),
            .I(N__91864));
    ClkMux I__18806 (
            .O(N__93114),
            .I(N__91864));
    ClkMux I__18805 (
            .O(N__93113),
            .I(N__91864));
    ClkMux I__18804 (
            .O(N__93112),
            .I(N__91864));
    ClkMux I__18803 (
            .O(N__93111),
            .I(N__91864));
    ClkMux I__18802 (
            .O(N__93110),
            .I(N__91864));
    ClkMux I__18801 (
            .O(N__93109),
            .I(N__91864));
    ClkMux I__18800 (
            .O(N__93108),
            .I(N__91864));
    ClkMux I__18799 (
            .O(N__93107),
            .I(N__91864));
    ClkMux I__18798 (
            .O(N__93106),
            .I(N__91864));
    ClkMux I__18797 (
            .O(N__93105),
            .I(N__91864));
    ClkMux I__18796 (
            .O(N__93104),
            .I(N__91864));
    ClkMux I__18795 (
            .O(N__93103),
            .I(N__91864));
    ClkMux I__18794 (
            .O(N__93102),
            .I(N__91864));
    ClkMux I__18793 (
            .O(N__93101),
            .I(N__91864));
    ClkMux I__18792 (
            .O(N__93100),
            .I(N__91864));
    ClkMux I__18791 (
            .O(N__93099),
            .I(N__91864));
    ClkMux I__18790 (
            .O(N__93098),
            .I(N__91864));
    ClkMux I__18789 (
            .O(N__93097),
            .I(N__91864));
    ClkMux I__18788 (
            .O(N__93096),
            .I(N__91864));
    ClkMux I__18787 (
            .O(N__93095),
            .I(N__91864));
    ClkMux I__18786 (
            .O(N__93094),
            .I(N__91864));
    ClkMux I__18785 (
            .O(N__93093),
            .I(N__91864));
    ClkMux I__18784 (
            .O(N__93092),
            .I(N__91864));
    ClkMux I__18783 (
            .O(N__93091),
            .I(N__91864));
    ClkMux I__18782 (
            .O(N__93090),
            .I(N__91864));
    ClkMux I__18781 (
            .O(N__93089),
            .I(N__91864));
    ClkMux I__18780 (
            .O(N__93088),
            .I(N__91864));
    ClkMux I__18779 (
            .O(N__93087),
            .I(N__91864));
    ClkMux I__18778 (
            .O(N__93086),
            .I(N__91864));
    ClkMux I__18777 (
            .O(N__93085),
            .I(N__91864));
    ClkMux I__18776 (
            .O(N__93084),
            .I(N__91864));
    ClkMux I__18775 (
            .O(N__93083),
            .I(N__91864));
    ClkMux I__18774 (
            .O(N__93082),
            .I(N__91864));
    ClkMux I__18773 (
            .O(N__93081),
            .I(N__91864));
    ClkMux I__18772 (
            .O(N__93080),
            .I(N__91864));
    ClkMux I__18771 (
            .O(N__93079),
            .I(N__91864));
    ClkMux I__18770 (
            .O(N__93078),
            .I(N__91864));
    ClkMux I__18769 (
            .O(N__93077),
            .I(N__91864));
    ClkMux I__18768 (
            .O(N__93076),
            .I(N__91864));
    ClkMux I__18767 (
            .O(N__93075),
            .I(N__91864));
    ClkMux I__18766 (
            .O(N__93074),
            .I(N__91864));
    ClkMux I__18765 (
            .O(N__93073),
            .I(N__91864));
    ClkMux I__18764 (
            .O(N__93072),
            .I(N__91864));
    ClkMux I__18763 (
            .O(N__93071),
            .I(N__91864));
    ClkMux I__18762 (
            .O(N__93070),
            .I(N__91864));
    ClkMux I__18761 (
            .O(N__93069),
            .I(N__91864));
    ClkMux I__18760 (
            .O(N__93068),
            .I(N__91864));
    ClkMux I__18759 (
            .O(N__93067),
            .I(N__91864));
    ClkMux I__18758 (
            .O(N__93066),
            .I(N__91864));
    ClkMux I__18757 (
            .O(N__93065),
            .I(N__91864));
    ClkMux I__18756 (
            .O(N__93064),
            .I(N__91864));
    ClkMux I__18755 (
            .O(N__93063),
            .I(N__91864));
    ClkMux I__18754 (
            .O(N__93062),
            .I(N__91864));
    ClkMux I__18753 (
            .O(N__93061),
            .I(N__91864));
    ClkMux I__18752 (
            .O(N__93060),
            .I(N__91864));
    ClkMux I__18751 (
            .O(N__93059),
            .I(N__91864));
    ClkMux I__18750 (
            .O(N__93058),
            .I(N__91864));
    ClkMux I__18749 (
            .O(N__93057),
            .I(N__91864));
    ClkMux I__18748 (
            .O(N__93056),
            .I(N__91864));
    ClkMux I__18747 (
            .O(N__93055),
            .I(N__91864));
    ClkMux I__18746 (
            .O(N__93054),
            .I(N__91864));
    ClkMux I__18745 (
            .O(N__93053),
            .I(N__91864));
    ClkMux I__18744 (
            .O(N__93052),
            .I(N__91864));
    ClkMux I__18743 (
            .O(N__93051),
            .I(N__91864));
    ClkMux I__18742 (
            .O(N__93050),
            .I(N__91864));
    ClkMux I__18741 (
            .O(N__93049),
            .I(N__91864));
    ClkMux I__18740 (
            .O(N__93048),
            .I(N__91864));
    ClkMux I__18739 (
            .O(N__93047),
            .I(N__91864));
    ClkMux I__18738 (
            .O(N__93046),
            .I(N__91864));
    ClkMux I__18737 (
            .O(N__93045),
            .I(N__91864));
    ClkMux I__18736 (
            .O(N__93044),
            .I(N__91864));
    ClkMux I__18735 (
            .O(N__93043),
            .I(N__91864));
    ClkMux I__18734 (
            .O(N__93042),
            .I(N__91864));
    ClkMux I__18733 (
            .O(N__93041),
            .I(N__91864));
    ClkMux I__18732 (
            .O(N__93040),
            .I(N__91864));
    ClkMux I__18731 (
            .O(N__93039),
            .I(N__91864));
    ClkMux I__18730 (
            .O(N__93038),
            .I(N__91864));
    ClkMux I__18729 (
            .O(N__93037),
            .I(N__91864));
    ClkMux I__18728 (
            .O(N__93036),
            .I(N__91864));
    ClkMux I__18727 (
            .O(N__93035),
            .I(N__91864));
    ClkMux I__18726 (
            .O(N__93034),
            .I(N__91864));
    ClkMux I__18725 (
            .O(N__93033),
            .I(N__91864));
    ClkMux I__18724 (
            .O(N__93032),
            .I(N__91864));
    ClkMux I__18723 (
            .O(N__93031),
            .I(N__91864));
    ClkMux I__18722 (
            .O(N__93030),
            .I(N__91864));
    ClkMux I__18721 (
            .O(N__93029),
            .I(N__91864));
    ClkMux I__18720 (
            .O(N__93028),
            .I(N__91864));
    ClkMux I__18719 (
            .O(N__93027),
            .I(N__91864));
    ClkMux I__18718 (
            .O(N__93026),
            .I(N__91864));
    ClkMux I__18717 (
            .O(N__93025),
            .I(N__91864));
    ClkMux I__18716 (
            .O(N__93024),
            .I(N__91864));
    ClkMux I__18715 (
            .O(N__93023),
            .I(N__91864));
    ClkMux I__18714 (
            .O(N__93022),
            .I(N__91864));
    ClkMux I__18713 (
            .O(N__93021),
            .I(N__91864));
    ClkMux I__18712 (
            .O(N__93020),
            .I(N__91864));
    ClkMux I__18711 (
            .O(N__93019),
            .I(N__91864));
    ClkMux I__18710 (
            .O(N__93018),
            .I(N__91864));
    ClkMux I__18709 (
            .O(N__93017),
            .I(N__91864));
    ClkMux I__18708 (
            .O(N__93016),
            .I(N__91864));
    ClkMux I__18707 (
            .O(N__93015),
            .I(N__91864));
    ClkMux I__18706 (
            .O(N__93014),
            .I(N__91864));
    ClkMux I__18705 (
            .O(N__93013),
            .I(N__91864));
    ClkMux I__18704 (
            .O(N__93012),
            .I(N__91864));
    ClkMux I__18703 (
            .O(N__93011),
            .I(N__91864));
    ClkMux I__18702 (
            .O(N__93010),
            .I(N__91864));
    ClkMux I__18701 (
            .O(N__93009),
            .I(N__91864));
    ClkMux I__18700 (
            .O(N__93008),
            .I(N__91864));
    ClkMux I__18699 (
            .O(N__93007),
            .I(N__91864));
    ClkMux I__18698 (
            .O(N__93006),
            .I(N__91864));
    ClkMux I__18697 (
            .O(N__93005),
            .I(N__91864));
    ClkMux I__18696 (
            .O(N__93004),
            .I(N__91864));
    ClkMux I__18695 (
            .O(N__93003),
            .I(N__91864));
    ClkMux I__18694 (
            .O(N__93002),
            .I(N__91864));
    ClkMux I__18693 (
            .O(N__93001),
            .I(N__91864));
    ClkMux I__18692 (
            .O(N__93000),
            .I(N__91864));
    ClkMux I__18691 (
            .O(N__92999),
            .I(N__91864));
    ClkMux I__18690 (
            .O(N__92998),
            .I(N__91864));
    ClkMux I__18689 (
            .O(N__92997),
            .I(N__91864));
    ClkMux I__18688 (
            .O(N__92996),
            .I(N__91864));
    ClkMux I__18687 (
            .O(N__92995),
            .I(N__91864));
    ClkMux I__18686 (
            .O(N__92994),
            .I(N__91864));
    ClkMux I__18685 (
            .O(N__92993),
            .I(N__91864));
    ClkMux I__18684 (
            .O(N__92992),
            .I(N__91864));
    ClkMux I__18683 (
            .O(N__92991),
            .I(N__91864));
    ClkMux I__18682 (
            .O(N__92990),
            .I(N__91864));
    ClkMux I__18681 (
            .O(N__92989),
            .I(N__91864));
    ClkMux I__18680 (
            .O(N__92988),
            .I(N__91864));
    ClkMux I__18679 (
            .O(N__92987),
            .I(N__91864));
    ClkMux I__18678 (
            .O(N__92986),
            .I(N__91864));
    ClkMux I__18677 (
            .O(N__92985),
            .I(N__91864));
    ClkMux I__18676 (
            .O(N__92984),
            .I(N__91864));
    ClkMux I__18675 (
            .O(N__92983),
            .I(N__91864));
    ClkMux I__18674 (
            .O(N__92982),
            .I(N__91864));
    ClkMux I__18673 (
            .O(N__92981),
            .I(N__91864));
    ClkMux I__18672 (
            .O(N__92980),
            .I(N__91864));
    ClkMux I__18671 (
            .O(N__92979),
            .I(N__91864));
    ClkMux I__18670 (
            .O(N__92978),
            .I(N__91864));
    ClkMux I__18669 (
            .O(N__92977),
            .I(N__91864));
    ClkMux I__18668 (
            .O(N__92976),
            .I(N__91864));
    ClkMux I__18667 (
            .O(N__92975),
            .I(N__91864));
    ClkMux I__18666 (
            .O(N__92974),
            .I(N__91864));
    ClkMux I__18665 (
            .O(N__92973),
            .I(N__91864));
    ClkMux I__18664 (
            .O(N__92972),
            .I(N__91864));
    ClkMux I__18663 (
            .O(N__92971),
            .I(N__91864));
    ClkMux I__18662 (
            .O(N__92970),
            .I(N__91864));
    ClkMux I__18661 (
            .O(N__92969),
            .I(N__91864));
    ClkMux I__18660 (
            .O(N__92968),
            .I(N__91864));
    ClkMux I__18659 (
            .O(N__92967),
            .I(N__91864));
    ClkMux I__18658 (
            .O(N__92966),
            .I(N__91864));
    ClkMux I__18657 (
            .O(N__92965),
            .I(N__91864));
    ClkMux I__18656 (
            .O(N__92964),
            .I(N__91864));
    ClkMux I__18655 (
            .O(N__92963),
            .I(N__91864));
    ClkMux I__18654 (
            .O(N__92962),
            .I(N__91864));
    ClkMux I__18653 (
            .O(N__92961),
            .I(N__91864));
    ClkMux I__18652 (
            .O(N__92960),
            .I(N__91864));
    ClkMux I__18651 (
            .O(N__92959),
            .I(N__91864));
    ClkMux I__18650 (
            .O(N__92958),
            .I(N__91864));
    ClkMux I__18649 (
            .O(N__92957),
            .I(N__91864));
    ClkMux I__18648 (
            .O(N__92956),
            .I(N__91864));
    ClkMux I__18647 (
            .O(N__92955),
            .I(N__91864));
    ClkMux I__18646 (
            .O(N__92954),
            .I(N__91864));
    ClkMux I__18645 (
            .O(N__92953),
            .I(N__91864));
    ClkMux I__18644 (
            .O(N__92952),
            .I(N__91864));
    ClkMux I__18643 (
            .O(N__92951),
            .I(N__91864));
    ClkMux I__18642 (
            .O(N__92950),
            .I(N__91864));
    ClkMux I__18641 (
            .O(N__92949),
            .I(N__91864));
    ClkMux I__18640 (
            .O(N__92948),
            .I(N__91864));
    ClkMux I__18639 (
            .O(N__92947),
            .I(N__91864));
    ClkMux I__18638 (
            .O(N__92946),
            .I(N__91864));
    ClkMux I__18637 (
            .O(N__92945),
            .I(N__91864));
    ClkMux I__18636 (
            .O(N__92944),
            .I(N__91864));
    ClkMux I__18635 (
            .O(N__92943),
            .I(N__91864));
    ClkMux I__18634 (
            .O(N__92942),
            .I(N__91864));
    ClkMux I__18633 (
            .O(N__92941),
            .I(N__91864));
    ClkMux I__18632 (
            .O(N__92940),
            .I(N__91864));
    ClkMux I__18631 (
            .O(N__92939),
            .I(N__91864));
    ClkMux I__18630 (
            .O(N__92938),
            .I(N__91864));
    ClkMux I__18629 (
            .O(N__92937),
            .I(N__91864));
    ClkMux I__18628 (
            .O(N__92936),
            .I(N__91864));
    ClkMux I__18627 (
            .O(N__92935),
            .I(N__91864));
    ClkMux I__18626 (
            .O(N__92934),
            .I(N__91864));
    ClkMux I__18625 (
            .O(N__92933),
            .I(N__91864));
    ClkMux I__18624 (
            .O(N__92932),
            .I(N__91864));
    ClkMux I__18623 (
            .O(N__92931),
            .I(N__91864));
    ClkMux I__18622 (
            .O(N__92930),
            .I(N__91864));
    ClkMux I__18621 (
            .O(N__92929),
            .I(N__91864));
    ClkMux I__18620 (
            .O(N__92928),
            .I(N__91864));
    ClkMux I__18619 (
            .O(N__92927),
            .I(N__91864));
    ClkMux I__18618 (
            .O(N__92926),
            .I(N__91864));
    ClkMux I__18617 (
            .O(N__92925),
            .I(N__91864));
    ClkMux I__18616 (
            .O(N__92924),
            .I(N__91864));
    ClkMux I__18615 (
            .O(N__92923),
            .I(N__91864));
    ClkMux I__18614 (
            .O(N__92922),
            .I(N__91864));
    ClkMux I__18613 (
            .O(N__92921),
            .I(N__91864));
    ClkMux I__18612 (
            .O(N__92920),
            .I(N__91864));
    ClkMux I__18611 (
            .O(N__92919),
            .I(N__91864));
    ClkMux I__18610 (
            .O(N__92918),
            .I(N__91864));
    ClkMux I__18609 (
            .O(N__92917),
            .I(N__91864));
    ClkMux I__18608 (
            .O(N__92916),
            .I(N__91864));
    ClkMux I__18607 (
            .O(N__92915),
            .I(N__91864));
    ClkMux I__18606 (
            .O(N__92914),
            .I(N__91864));
    ClkMux I__18605 (
            .O(N__92913),
            .I(N__91864));
    ClkMux I__18604 (
            .O(N__92912),
            .I(N__91864));
    ClkMux I__18603 (
            .O(N__92911),
            .I(N__91864));
    ClkMux I__18602 (
            .O(N__92910),
            .I(N__91864));
    ClkMux I__18601 (
            .O(N__92909),
            .I(N__91864));
    ClkMux I__18600 (
            .O(N__92908),
            .I(N__91864));
    ClkMux I__18599 (
            .O(N__92907),
            .I(N__91864));
    GlobalMux I__18598 (
            .O(N__91864),
            .I(N__91861));
    gio2CtrlBuf I__18597 (
            .O(N__91861),
            .I(clk_c_g));
    CEMux I__18596 (
            .O(N__91858),
            .I(N__91852));
    CEMux I__18595 (
            .O(N__91857),
            .I(N__91849));
    CEMux I__18594 (
            .O(N__91856),
            .I(N__91846));
    CEMux I__18593 (
            .O(N__91855),
            .I(N__91843));
    LocalMux I__18592 (
            .O(N__91852),
            .I(N__91838));
    LocalMux I__18591 (
            .O(N__91849),
            .I(N__91838));
    LocalMux I__18590 (
            .O(N__91846),
            .I(N__91835));
    LocalMux I__18589 (
            .O(N__91843),
            .I(N__91832));
    Odrv12 I__18588 (
            .O(N__91838),
            .I(clk_en_37));
    Odrv12 I__18587 (
            .O(N__91835),
            .I(clk_en_37));
    Odrv4 I__18586 (
            .O(N__91832),
            .I(clk_en_37));
    InMux I__18585 (
            .O(N__91825),
            .I(N__91822));
    LocalMux I__18584 (
            .O(N__91822),
            .I(N__91818));
    InMux I__18583 (
            .O(N__91821),
            .I(N__91815));
    Span4Mux_v I__18582 (
            .O(N__91818),
            .I(N__91811));
    LocalMux I__18581 (
            .O(N__91815),
            .I(N__91808));
    InMux I__18580 (
            .O(N__91814),
            .I(N__91804));
    Span4Mux_h I__18579 (
            .O(N__91811),
            .I(N__91799));
    Span4Mux_v I__18578 (
            .O(N__91808),
            .I(N__91799));
    InMux I__18577 (
            .O(N__91807),
            .I(N__91795));
    LocalMux I__18576 (
            .O(N__91804),
            .I(N__91792));
    Span4Mux_h I__18575 (
            .O(N__91799),
            .I(N__91789));
    InMux I__18574 (
            .O(N__91798),
            .I(N__91786));
    LocalMux I__18573 (
            .O(N__91795),
            .I(shift_srl_186Z0Z_15));
    Odrv4 I__18572 (
            .O(N__91792),
            .I(shift_srl_186Z0Z_15));
    Odrv4 I__18571 (
            .O(N__91789),
            .I(shift_srl_186Z0Z_15));
    LocalMux I__18570 (
            .O(N__91786),
            .I(shift_srl_186Z0Z_15));
    IoInMux I__18569 (
            .O(N__91777),
            .I(N__91774));
    LocalMux I__18568 (
            .O(N__91774),
            .I(N__91771));
    Odrv12 I__18567 (
            .O(N__91771),
            .I(rco_c_186));
    CascadeMux I__18566 (
            .O(N__91768),
            .I(N__91764));
    InMux I__18565 (
            .O(N__91767),
            .I(N__91758));
    InMux I__18564 (
            .O(N__91764),
            .I(N__91755));
    InMux I__18563 (
            .O(N__91763),
            .I(N__91752));
    InMux I__18562 (
            .O(N__91762),
            .I(N__91749));
    InMux I__18561 (
            .O(N__91761),
            .I(N__91746));
    LocalMux I__18560 (
            .O(N__91758),
            .I(N__91743));
    LocalMux I__18559 (
            .O(N__91755),
            .I(N__91737));
    LocalMux I__18558 (
            .O(N__91752),
            .I(N__91737));
    LocalMux I__18557 (
            .O(N__91749),
            .I(N__91733));
    LocalMux I__18556 (
            .O(N__91746),
            .I(N__91728));
    Span4Mux_h I__18555 (
            .O(N__91743),
            .I(N__91728));
    InMux I__18554 (
            .O(N__91742),
            .I(N__91725));
    Span12Mux_v I__18553 (
            .O(N__91737),
            .I(N__91722));
    InMux I__18552 (
            .O(N__91736),
            .I(N__91719));
    Span4Mux_v I__18551 (
            .O(N__91733),
            .I(N__91716));
    Span4Mux_h I__18550 (
            .O(N__91728),
            .I(N__91713));
    LocalMux I__18549 (
            .O(N__91725),
            .I(N__91710));
    Odrv12 I__18548 (
            .O(N__91722),
            .I(shift_srl_185Z0Z_15));
    LocalMux I__18547 (
            .O(N__91719),
            .I(shift_srl_185Z0Z_15));
    Odrv4 I__18546 (
            .O(N__91716),
            .I(shift_srl_185Z0Z_15));
    Odrv4 I__18545 (
            .O(N__91713),
            .I(shift_srl_185Z0Z_15));
    Odrv4 I__18544 (
            .O(N__91710),
            .I(shift_srl_185Z0Z_15));
    InMux I__18543 (
            .O(N__91699),
            .I(N__91695));
    InMux I__18542 (
            .O(N__91698),
            .I(N__91692));
    LocalMux I__18541 (
            .O(N__91695),
            .I(N__91683));
    LocalMux I__18540 (
            .O(N__91692),
            .I(N__91683));
    InMux I__18539 (
            .O(N__91691),
            .I(N__91679));
    InMux I__18538 (
            .O(N__91690),
            .I(N__91676));
    InMux I__18537 (
            .O(N__91689),
            .I(N__91673));
    InMux I__18536 (
            .O(N__91688),
            .I(N__91670));
    Span4Mux_v I__18535 (
            .O(N__91683),
            .I(N__91667));
    InMux I__18534 (
            .O(N__91682),
            .I(N__91664));
    LocalMux I__18533 (
            .O(N__91679),
            .I(N__91661));
    LocalMux I__18532 (
            .O(N__91676),
            .I(N__91658));
    LocalMux I__18531 (
            .O(N__91673),
            .I(N__91653));
    LocalMux I__18530 (
            .O(N__91670),
            .I(N__91653));
    Span4Mux_h I__18529 (
            .O(N__91667),
            .I(N__91648));
    LocalMux I__18528 (
            .O(N__91664),
            .I(N__91648));
    Span12Mux_s9_v I__18527 (
            .O(N__91661),
            .I(N__91643));
    Span4Mux_v I__18526 (
            .O(N__91658),
            .I(N__91638));
    Span4Mux_v I__18525 (
            .O(N__91653),
            .I(N__91638));
    Span4Mux_h I__18524 (
            .O(N__91648),
            .I(N__91635));
    InMux I__18523 (
            .O(N__91647),
            .I(N__91630));
    InMux I__18522 (
            .O(N__91646),
            .I(N__91630));
    Odrv12 I__18521 (
            .O(N__91643),
            .I(shift_srl_184Z0Z_15));
    Odrv4 I__18520 (
            .O(N__91638),
            .I(shift_srl_184Z0Z_15));
    Odrv4 I__18519 (
            .O(N__91635),
            .I(shift_srl_184Z0Z_15));
    LocalMux I__18518 (
            .O(N__91630),
            .I(shift_srl_184Z0Z_15));
    IoInMux I__18517 (
            .O(N__91621),
            .I(N__91618));
    LocalMux I__18516 (
            .O(N__91618),
            .I(N__91615));
    Odrv12 I__18515 (
            .O(N__91615),
            .I(rco_c_185));
    InMux I__18514 (
            .O(N__91612),
            .I(N__91609));
    LocalMux I__18513 (
            .O(N__91609),
            .I(N__91603));
    InMux I__18512 (
            .O(N__91608),
            .I(N__91600));
    InMux I__18511 (
            .O(N__91607),
            .I(N__91597));
    InMux I__18510 (
            .O(N__91606),
            .I(N__91594));
    Span12Mux_v I__18509 (
            .O(N__91603),
            .I(N__91589));
    LocalMux I__18508 (
            .O(N__91600),
            .I(N__91589));
    LocalMux I__18507 (
            .O(N__91597),
            .I(shift_srl_190Z0Z_15));
    LocalMux I__18506 (
            .O(N__91594),
            .I(shift_srl_190Z0Z_15));
    Odrv12 I__18505 (
            .O(N__91589),
            .I(shift_srl_190Z0Z_15));
    IoInMux I__18504 (
            .O(N__91582),
            .I(N__91579));
    LocalMux I__18503 (
            .O(N__91579),
            .I(N__91576));
    Span4Mux_s1_h I__18502 (
            .O(N__91576),
            .I(N__91573));
    Odrv4 I__18501 (
            .O(N__91573),
            .I(rco_c_190));
    InMux I__18500 (
            .O(N__91570),
            .I(N__91567));
    LocalMux I__18499 (
            .O(N__91567),
            .I(N__91562));
    InMux I__18498 (
            .O(N__91566),
            .I(N__91559));
    CascadeMux I__18497 (
            .O(N__91565),
            .I(N__91556));
    Span4Mux_v I__18496 (
            .O(N__91562),
            .I(N__91553));
    LocalMux I__18495 (
            .O(N__91559),
            .I(N__91550));
    InMux I__18494 (
            .O(N__91556),
            .I(N__91547));
    Odrv4 I__18493 (
            .O(N__91553),
            .I(N_4175));
    Odrv12 I__18492 (
            .O(N__91550),
            .I(N_4175));
    LocalMux I__18491 (
            .O(N__91547),
            .I(N_4175));
    IoInMux I__18490 (
            .O(N__91540),
            .I(N__91534));
    InMux I__18489 (
            .O(N__91539),
            .I(N__91522));
    InMux I__18488 (
            .O(N__91538),
            .I(N__91517));
    InMux I__18487 (
            .O(N__91537),
            .I(N__91517));
    LocalMux I__18486 (
            .O(N__91534),
            .I(N__91513));
    InMux I__18485 (
            .O(N__91533),
            .I(N__91506));
    InMux I__18484 (
            .O(N__91532),
            .I(N__91506));
    InMux I__18483 (
            .O(N__91531),
            .I(N__91497));
    InMux I__18482 (
            .O(N__91530),
            .I(N__91497));
    InMux I__18481 (
            .O(N__91529),
            .I(N__91497));
    InMux I__18480 (
            .O(N__91528),
            .I(N__91497));
    InMux I__18479 (
            .O(N__91527),
            .I(N__91494));
    InMux I__18478 (
            .O(N__91526),
            .I(N__91488));
    InMux I__18477 (
            .O(N__91525),
            .I(N__91488));
    LocalMux I__18476 (
            .O(N__91522),
            .I(N__91483));
    LocalMux I__18475 (
            .O(N__91517),
            .I(N__91483));
    InMux I__18474 (
            .O(N__91516),
            .I(N__91480));
    IoSpan4Mux I__18473 (
            .O(N__91513),
            .I(N__91475));
    InMux I__18472 (
            .O(N__91512),
            .I(N__91470));
    InMux I__18471 (
            .O(N__91511),
            .I(N__91470));
    LocalMux I__18470 (
            .O(N__91506),
            .I(N__91465));
    LocalMux I__18469 (
            .O(N__91497),
            .I(N__91465));
    LocalMux I__18468 (
            .O(N__91494),
            .I(N__91462));
    InMux I__18467 (
            .O(N__91493),
            .I(N__91459));
    LocalMux I__18466 (
            .O(N__91488),
            .I(N__91454));
    Span12Mux_v I__18465 (
            .O(N__91483),
            .I(N__91451));
    LocalMux I__18464 (
            .O(N__91480),
            .I(N__91448));
    InMux I__18463 (
            .O(N__91479),
            .I(N__91443));
    InMux I__18462 (
            .O(N__91478),
            .I(N__91443));
    Span4Mux_s2_v I__18461 (
            .O(N__91475),
            .I(N__91438));
    LocalMux I__18460 (
            .O(N__91470),
            .I(N__91438));
    Span4Mux_v I__18459 (
            .O(N__91465),
            .I(N__91435));
    Span12Mux_s3_h I__18458 (
            .O(N__91462),
            .I(N__91430));
    LocalMux I__18457 (
            .O(N__91459),
            .I(N__91430));
    InMux I__18456 (
            .O(N__91458),
            .I(N__91425));
    InMux I__18455 (
            .O(N__91457),
            .I(N__91425));
    Span4Mux_h I__18454 (
            .O(N__91454),
            .I(N__91422));
    Span12Mux_h I__18453 (
            .O(N__91451),
            .I(N__91415));
    Sp12to4 I__18452 (
            .O(N__91448),
            .I(N__91415));
    LocalMux I__18451 (
            .O(N__91443),
            .I(N__91415));
    Span4Mux_v I__18450 (
            .O(N__91438),
            .I(N__91412));
    Odrv4 I__18449 (
            .O(N__91435),
            .I(rco_c_183));
    Odrv12 I__18448 (
            .O(N__91430),
            .I(rco_c_183));
    LocalMux I__18447 (
            .O(N__91425),
            .I(rco_c_183));
    Odrv4 I__18446 (
            .O(N__91422),
            .I(rco_c_183));
    Odrv12 I__18445 (
            .O(N__91415),
            .I(rco_c_183));
    Odrv4 I__18444 (
            .O(N__91412),
            .I(rco_c_183));
    IoInMux I__18443 (
            .O(N__91399),
            .I(N__91396));
    LocalMux I__18442 (
            .O(N__91396),
            .I(N__91393));
    Span4Mux_s1_h I__18441 (
            .O(N__91393),
            .I(N__91390));
    Odrv4 I__18440 (
            .O(N__91390),
            .I(rco_c_189));
    InMux I__18439 (
            .O(N__91387),
            .I(N__91384));
    LocalMux I__18438 (
            .O(N__91384),
            .I(N__91381));
    Span4Mux_v I__18437 (
            .O(N__91381),
            .I(N__91378));
    Span4Mux_v I__18436 (
            .O(N__91378),
            .I(N__91375));
    Sp12to4 I__18435 (
            .O(N__91375),
            .I(N__91371));
    CascadeMux I__18434 (
            .O(N__91374),
            .I(N__91368));
    Span12Mux_s11_h I__18433 (
            .O(N__91371),
            .I(N__91365));
    InMux I__18432 (
            .O(N__91368),
            .I(N__91362));
    Span12Mux_h I__18431 (
            .O(N__91365),
            .I(N__91359));
    LocalMux I__18430 (
            .O(N__91362),
            .I(N__91356));
    Odrv12 I__18429 (
            .O(N__91359),
            .I(shift_srl_129_RNIDM4DZ0Z_15));
    Odrv4 I__18428 (
            .O(N__91356),
            .I(shift_srl_129_RNIDM4DZ0Z_15));
    IoInMux I__18427 (
            .O(N__91351),
            .I(N__91348));
    LocalMux I__18426 (
            .O(N__91348),
            .I(N__91345));
    Span4Mux_s1_h I__18425 (
            .O(N__91345),
            .I(N__91342));
    Sp12to4 I__18424 (
            .O(N__91342),
            .I(N__91339));
    Odrv12 I__18423 (
            .O(N__91339),
            .I(rco_c_129));
    InMux I__18422 (
            .O(N__91336),
            .I(N__91329));
    InMux I__18421 (
            .O(N__91335),
            .I(N__91329));
    IoInMux I__18420 (
            .O(N__91334),
            .I(N__91326));
    LocalMux I__18419 (
            .O(N__91329),
            .I(N__91322));
    LocalMux I__18418 (
            .O(N__91326),
            .I(N__91319));
    InMux I__18417 (
            .O(N__91325),
            .I(N__91316));
    Span4Mux_v I__18416 (
            .O(N__91322),
            .I(N__91313));
    IoSpan4Mux I__18415 (
            .O(N__91319),
            .I(N__91310));
    LocalMux I__18414 (
            .O(N__91316),
            .I(N__91307));
    Span4Mux_v I__18413 (
            .O(N__91313),
            .I(N__91303));
    Span4Mux_s3_h I__18412 (
            .O(N__91310),
            .I(N__91300));
    Span4Mux_v I__18411 (
            .O(N__91307),
            .I(N__91297));
    InMux I__18410 (
            .O(N__91306),
            .I(N__91294));
    Sp12to4 I__18409 (
            .O(N__91303),
            .I(N__91291));
    Sp12to4 I__18408 (
            .O(N__91300),
            .I(N__91284));
    Sp12to4 I__18407 (
            .O(N__91297),
            .I(N__91284));
    LocalMux I__18406 (
            .O(N__91294),
            .I(N__91284));
    Span12Mux_s11_h I__18405 (
            .O(N__91291),
            .I(N__91279));
    Span12Mux_s8_h I__18404 (
            .O(N__91284),
            .I(N__91279));
    Odrv12 I__18403 (
            .O(N__91279),
            .I(rco_c_127));
    InMux I__18402 (
            .O(N__91276),
            .I(N__91273));
    LocalMux I__18401 (
            .O(N__91273),
            .I(N__91270));
    Span12Mux_v I__18400 (
            .O(N__91270),
            .I(N__91263));
    InMux I__18399 (
            .O(N__91269),
            .I(N__91260));
    CascadeMux I__18398 (
            .O(N__91268),
            .I(N__91257));
    InMux I__18397 (
            .O(N__91267),
            .I(N__91251));
    InMux I__18396 (
            .O(N__91266),
            .I(N__91251));
    Span12Mux_h I__18395 (
            .O(N__91263),
            .I(N__91242));
    LocalMux I__18394 (
            .O(N__91260),
            .I(N__91239));
    InMux I__18393 (
            .O(N__91257),
            .I(N__91236));
    InMux I__18392 (
            .O(N__91256),
            .I(N__91233));
    LocalMux I__18391 (
            .O(N__91251),
            .I(N__91230));
    InMux I__18390 (
            .O(N__91250),
            .I(N__91221));
    InMux I__18389 (
            .O(N__91249),
            .I(N__91221));
    InMux I__18388 (
            .O(N__91248),
            .I(N__91221));
    InMux I__18387 (
            .O(N__91247),
            .I(N__91221));
    InMux I__18386 (
            .O(N__91246),
            .I(N__91218));
    CascadeMux I__18385 (
            .O(N__91245),
            .I(N__91215));
    Span12Mux_h I__18384 (
            .O(N__91242),
            .I(N__91210));
    Span4Mux_h I__18383 (
            .O(N__91239),
            .I(N__91205));
    LocalMux I__18382 (
            .O(N__91236),
            .I(N__91205));
    LocalMux I__18381 (
            .O(N__91233),
            .I(N__91200));
    Span4Mux_h I__18380 (
            .O(N__91230),
            .I(N__91200));
    LocalMux I__18379 (
            .O(N__91221),
            .I(N__91195));
    LocalMux I__18378 (
            .O(N__91218),
            .I(N__91195));
    InMux I__18377 (
            .O(N__91215),
            .I(N__91192));
    InMux I__18376 (
            .O(N__91214),
            .I(N__91187));
    InMux I__18375 (
            .O(N__91213),
            .I(N__91187));
    Odrv12 I__18374 (
            .O(N__91210),
            .I(shift_srl_128Z0Z_15));
    Odrv4 I__18373 (
            .O(N__91205),
            .I(shift_srl_128Z0Z_15));
    Odrv4 I__18372 (
            .O(N__91200),
            .I(shift_srl_128Z0Z_15));
    Odrv12 I__18371 (
            .O(N__91195),
            .I(shift_srl_128Z0Z_15));
    LocalMux I__18370 (
            .O(N__91192),
            .I(shift_srl_128Z0Z_15));
    LocalMux I__18369 (
            .O(N__91187),
            .I(shift_srl_128Z0Z_15));
    IoInMux I__18368 (
            .O(N__91174),
            .I(N__91171));
    LocalMux I__18367 (
            .O(N__91171),
            .I(N__91168));
    IoSpan4Mux I__18366 (
            .O(N__91168),
            .I(N__91165));
    Odrv4 I__18365 (
            .O(N__91165),
            .I(rco_c_128));
    InMux I__18364 (
            .O(N__91162),
            .I(N__91159));
    LocalMux I__18363 (
            .O(N__91159),
            .I(N__91156));
    Span4Mux_h I__18362 (
            .O(N__91156),
            .I(N__91152));
    CascadeMux I__18361 (
            .O(N__91155),
            .I(N__91149));
    Sp12to4 I__18360 (
            .O(N__91152),
            .I(N__91146));
    InMux I__18359 (
            .O(N__91149),
            .I(N__91143));
    Span12Mux_v I__18358 (
            .O(N__91146),
            .I(N__91140));
    LocalMux I__18357 (
            .O(N__91143),
            .I(N__91137));
    Span12Mux_h I__18356 (
            .O(N__91140),
            .I(N__91134));
    Span4Mux_v I__18355 (
            .O(N__91137),
            .I(N__91131));
    Odrv12 I__18354 (
            .O(N__91134),
            .I(shift_srl_140_RNI85IAZ0Z_15));
    Odrv4 I__18353 (
            .O(N__91131),
            .I(shift_srl_140_RNI85IAZ0Z_15));
    IoInMux I__18352 (
            .O(N__91126),
            .I(N__91123));
    LocalMux I__18351 (
            .O(N__91123),
            .I(N__91120));
    IoSpan4Mux I__18350 (
            .O(N__91120),
            .I(N__91117));
    IoSpan4Mux I__18349 (
            .O(N__91117),
            .I(N__91114));
    Span4Mux_s1_v I__18348 (
            .O(N__91114),
            .I(N__91107));
    InMux I__18347 (
            .O(N__91113),
            .I(N__91104));
    InMux I__18346 (
            .O(N__91112),
            .I(N__91101));
    InMux I__18345 (
            .O(N__91111),
            .I(N__91096));
    InMux I__18344 (
            .O(N__91110),
            .I(N__91096));
    Span4Mux_v I__18343 (
            .O(N__91107),
            .I(N__91093));
    LocalMux I__18342 (
            .O(N__91104),
            .I(N__91090));
    LocalMux I__18341 (
            .O(N__91101),
            .I(N__91087));
    LocalMux I__18340 (
            .O(N__91096),
            .I(N__91084));
    Sp12to4 I__18339 (
            .O(N__91093),
            .I(N__91077));
    Span12Mux_s4_h I__18338 (
            .O(N__91090),
            .I(N__91077));
    Span12Mux_v I__18337 (
            .O(N__91087),
            .I(N__91074));
    Span4Mux_h I__18336 (
            .O(N__91084),
            .I(N__91071));
    InMux I__18335 (
            .O(N__91083),
            .I(N__91066));
    InMux I__18334 (
            .O(N__91082),
            .I(N__91066));
    Span12Mux_h I__18333 (
            .O(N__91077),
            .I(N__91061));
    Span12Mux_h I__18332 (
            .O(N__91074),
            .I(N__91061));
    Sp12to4 I__18331 (
            .O(N__91071),
            .I(N__91058));
    LocalMux I__18330 (
            .O(N__91066),
            .I(N__91055));
    Odrv12 I__18329 (
            .O(N__91061),
            .I(rco_c_138));
    Odrv12 I__18328 (
            .O(N__91058),
            .I(rco_c_138));
    Odrv12 I__18327 (
            .O(N__91055),
            .I(rco_c_138));
    IoInMux I__18326 (
            .O(N__91048),
            .I(N__91045));
    LocalMux I__18325 (
            .O(N__91045),
            .I(N__91042));
    IoSpan4Mux I__18324 (
            .O(N__91042),
            .I(N__91039));
    Odrv4 I__18323 (
            .O(N__91039),
            .I(N_125_i));
    InMux I__18322 (
            .O(N__91036),
            .I(N__91033));
    LocalMux I__18321 (
            .O(N__91033),
            .I(shift_srl_73Z0Z_2));
    InMux I__18320 (
            .O(N__91030),
            .I(N__91027));
    LocalMux I__18319 (
            .O(N__91027),
            .I(shift_srl_73Z0Z_3));
    InMux I__18318 (
            .O(N__91024),
            .I(N__91021));
    LocalMux I__18317 (
            .O(N__91021),
            .I(shift_srl_73Z0Z_4));
    InMux I__18316 (
            .O(N__91018),
            .I(N__91015));
    LocalMux I__18315 (
            .O(N__91015),
            .I(shift_srl_73Z0Z_5));
    InMux I__18314 (
            .O(N__91012),
            .I(N__91009));
    LocalMux I__18313 (
            .O(N__91009),
            .I(shift_srl_73Z0Z_6));
    InMux I__18312 (
            .O(N__91006),
            .I(N__91003));
    LocalMux I__18311 (
            .O(N__91003),
            .I(N__91000));
    Odrv4 I__18310 (
            .O(N__91000),
            .I(shift_srl_73Z0Z_7));
    CEMux I__18309 (
            .O(N__90997),
            .I(N__90993));
    CEMux I__18308 (
            .O(N__90996),
            .I(N__90990));
    LocalMux I__18307 (
            .O(N__90993),
            .I(N__90987));
    LocalMux I__18306 (
            .O(N__90990),
            .I(N__90984));
    Span4Mux_s2_h I__18305 (
            .O(N__90987),
            .I(N__90981));
    Odrv12 I__18304 (
            .O(N__90984),
            .I(clk_en_73));
    Odrv4 I__18303 (
            .O(N__90981),
            .I(clk_en_73));
    InMux I__18302 (
            .O(N__90976),
            .I(N__90973));
    LocalMux I__18301 (
            .O(N__90973),
            .I(N__90970));
    Span4Mux_h I__18300 (
            .O(N__90970),
            .I(N__90967));
    Odrv4 I__18299 (
            .O(N__90967),
            .I(shift_srl_36Z0Z_13));
    InMux I__18298 (
            .O(N__90964),
            .I(N__90961));
    LocalMux I__18297 (
            .O(N__90961),
            .I(N__90958));
    Span4Mux_h I__18296 (
            .O(N__90958),
            .I(N__90955));
    Span4Mux_v I__18295 (
            .O(N__90955),
            .I(N__90952));
    Span4Mux_h I__18294 (
            .O(N__90952),
            .I(N__90949));
    Span4Mux_h I__18293 (
            .O(N__90949),
            .I(N__90946));
    Odrv4 I__18292 (
            .O(N__90946),
            .I(shift_srl_36Z0Z_14));
    CEMux I__18291 (
            .O(N__90943),
            .I(N__90939));
    CEMux I__18290 (
            .O(N__90942),
            .I(N__90935));
    LocalMux I__18289 (
            .O(N__90939),
            .I(N__90932));
    CEMux I__18288 (
            .O(N__90938),
            .I(N__90929));
    LocalMux I__18287 (
            .O(N__90935),
            .I(N__90926));
    Span4Mux_v I__18286 (
            .O(N__90932),
            .I(N__90923));
    LocalMux I__18285 (
            .O(N__90929),
            .I(N__90920));
    Span4Mux_h I__18284 (
            .O(N__90926),
            .I(N__90915));
    Span4Mux_h I__18283 (
            .O(N__90923),
            .I(N__90910));
    Span4Mux_h I__18282 (
            .O(N__90920),
            .I(N__90910));
    CEMux I__18281 (
            .O(N__90919),
            .I(N__90907));
    CEMux I__18280 (
            .O(N__90918),
            .I(N__90904));
    Span4Mux_h I__18279 (
            .O(N__90915),
            .I(N__90901));
    Span4Mux_v I__18278 (
            .O(N__90910),
            .I(N__90898));
    LocalMux I__18277 (
            .O(N__90907),
            .I(N__90895));
    LocalMux I__18276 (
            .O(N__90904),
            .I(N__90892));
    Odrv4 I__18275 (
            .O(N__90901),
            .I(clk_en_36));
    Odrv4 I__18274 (
            .O(N__90898),
            .I(clk_en_36));
    Odrv12 I__18273 (
            .O(N__90895),
            .I(clk_en_36));
    Odrv4 I__18272 (
            .O(N__90892),
            .I(clk_en_36));
    InMux I__18271 (
            .O(N__90883),
            .I(N__90879));
    InMux I__18270 (
            .O(N__90882),
            .I(N__90876));
    LocalMux I__18269 (
            .O(N__90879),
            .I(N__90870));
    LocalMux I__18268 (
            .O(N__90876),
            .I(N__90870));
    InMux I__18267 (
            .O(N__90875),
            .I(N__90866));
    Span4Mux_v I__18266 (
            .O(N__90870),
            .I(N__90863));
    InMux I__18265 (
            .O(N__90869),
            .I(N__90860));
    LocalMux I__18264 (
            .O(N__90866),
            .I(N__90857));
    Span4Mux_h I__18263 (
            .O(N__90863),
            .I(N__90854));
    LocalMux I__18262 (
            .O(N__90860),
            .I(shift_srl_73Z0Z_15));
    Odrv4 I__18261 (
            .O(N__90857),
            .I(shift_srl_73Z0Z_15));
    Odrv4 I__18260 (
            .O(N__90854),
            .I(shift_srl_73Z0Z_15));
    InMux I__18259 (
            .O(N__90847),
            .I(N__90843));
    InMux I__18258 (
            .O(N__90846),
            .I(N__90840));
    LocalMux I__18257 (
            .O(N__90843),
            .I(N__90835));
    LocalMux I__18256 (
            .O(N__90840),
            .I(N__90831));
    InMux I__18255 (
            .O(N__90839),
            .I(N__90828));
    CascadeMux I__18254 (
            .O(N__90838),
            .I(N__90824));
    Span4Mux_v I__18253 (
            .O(N__90835),
            .I(N__90821));
    InMux I__18252 (
            .O(N__90834),
            .I(N__90818));
    Span4Mux_v I__18251 (
            .O(N__90831),
            .I(N__90813));
    LocalMux I__18250 (
            .O(N__90828),
            .I(N__90813));
    InMux I__18249 (
            .O(N__90827),
            .I(N__90808));
    InMux I__18248 (
            .O(N__90824),
            .I(N__90808));
    Odrv4 I__18247 (
            .O(N__90821),
            .I(shift_srl_72Z0Z_15));
    LocalMux I__18246 (
            .O(N__90818),
            .I(shift_srl_72Z0Z_15));
    Odrv4 I__18245 (
            .O(N__90813),
            .I(shift_srl_72Z0Z_15));
    LocalMux I__18244 (
            .O(N__90808),
            .I(shift_srl_72Z0Z_15));
    IoInMux I__18243 (
            .O(N__90799),
            .I(N__90796));
    LocalMux I__18242 (
            .O(N__90796),
            .I(N__90793));
    IoSpan4Mux I__18241 (
            .O(N__90793),
            .I(N__90790));
    Odrv4 I__18240 (
            .O(N__90790),
            .I(rco_c_73));
    InMux I__18239 (
            .O(N__90787),
            .I(N__90782));
    InMux I__18238 (
            .O(N__90786),
            .I(N__90779));
    CascadeMux I__18237 (
            .O(N__90785),
            .I(N__90776));
    LocalMux I__18236 (
            .O(N__90782),
            .I(N__90770));
    LocalMux I__18235 (
            .O(N__90779),
            .I(N__90770));
    InMux I__18234 (
            .O(N__90776),
            .I(N__90767));
    InMux I__18233 (
            .O(N__90775),
            .I(N__90763));
    Span4Mux_v I__18232 (
            .O(N__90770),
            .I(N__90758));
    LocalMux I__18231 (
            .O(N__90767),
            .I(N__90758));
    CascadeMux I__18230 (
            .O(N__90766),
            .I(N__90755));
    LocalMux I__18229 (
            .O(N__90763),
            .I(N__90752));
    Span4Mux_h I__18228 (
            .O(N__90758),
            .I(N__90749));
    InMux I__18227 (
            .O(N__90755),
            .I(N__90746));
    Odrv12 I__18226 (
            .O(N__90752),
            .I(shift_srl_71_RNIGP6RZ0Z_15));
    Odrv4 I__18225 (
            .O(N__90749),
            .I(shift_srl_71_RNIGP6RZ0Z_15));
    LocalMux I__18224 (
            .O(N__90746),
            .I(shift_srl_71_RNIGP6RZ0Z_15));
    CascadeMux I__18223 (
            .O(N__90739),
            .I(N__90735));
    CascadeMux I__18222 (
            .O(N__90738),
            .I(N__90730));
    InMux I__18221 (
            .O(N__90735),
            .I(N__90724));
    InMux I__18220 (
            .O(N__90734),
            .I(N__90721));
    InMux I__18219 (
            .O(N__90733),
            .I(N__90718));
    InMux I__18218 (
            .O(N__90730),
            .I(N__90715));
    InMux I__18217 (
            .O(N__90729),
            .I(N__90710));
    InMux I__18216 (
            .O(N__90728),
            .I(N__90707));
    IoInMux I__18215 (
            .O(N__90727),
            .I(N__90704));
    LocalMux I__18214 (
            .O(N__90724),
            .I(N__90697));
    LocalMux I__18213 (
            .O(N__90721),
            .I(N__90697));
    LocalMux I__18212 (
            .O(N__90718),
            .I(N__90697));
    LocalMux I__18211 (
            .O(N__90715),
            .I(N__90690));
    InMux I__18210 (
            .O(N__90714),
            .I(N__90685));
    InMux I__18209 (
            .O(N__90713),
            .I(N__90685));
    LocalMux I__18208 (
            .O(N__90710),
            .I(N__90680));
    LocalMux I__18207 (
            .O(N__90707),
            .I(N__90680));
    LocalMux I__18206 (
            .O(N__90704),
            .I(N__90677));
    Span4Mux_v I__18205 (
            .O(N__90697),
            .I(N__90674));
    InMux I__18204 (
            .O(N__90696),
            .I(N__90667));
    InMux I__18203 (
            .O(N__90695),
            .I(N__90667));
    InMux I__18202 (
            .O(N__90694),
            .I(N__90667));
    InMux I__18201 (
            .O(N__90693),
            .I(N__90664));
    Span4Mux_v I__18200 (
            .O(N__90690),
            .I(N__90659));
    LocalMux I__18199 (
            .O(N__90685),
            .I(N__90659));
    Span4Mux_h I__18198 (
            .O(N__90680),
            .I(N__90656));
    Span12Mux_s8_h I__18197 (
            .O(N__90677),
            .I(N__90653));
    Sp12to4 I__18196 (
            .O(N__90674),
            .I(N__90646));
    LocalMux I__18195 (
            .O(N__90667),
            .I(N__90646));
    LocalMux I__18194 (
            .O(N__90664),
            .I(N__90646));
    Span4Mux_h I__18193 (
            .O(N__90659),
            .I(N__90643));
    Span4Mux_v I__18192 (
            .O(N__90656),
            .I(N__90640));
    Odrv12 I__18191 (
            .O(N__90653),
            .I(rco_c_66));
    Odrv12 I__18190 (
            .O(N__90646),
            .I(rco_c_66));
    Odrv4 I__18189 (
            .O(N__90643),
            .I(rco_c_66));
    Odrv4 I__18188 (
            .O(N__90640),
            .I(rco_c_66));
    IoInMux I__18187 (
            .O(N__90631),
            .I(N__90628));
    LocalMux I__18186 (
            .O(N__90628),
            .I(N__90625));
    Odrv4 I__18185 (
            .O(N__90625),
            .I(rco_c_71));
    InMux I__18184 (
            .O(N__90622),
            .I(N__90619));
    LocalMux I__18183 (
            .O(N__90619),
            .I(shift_srl_73Z0Z_11));
    InMux I__18182 (
            .O(N__90616),
            .I(N__90613));
    LocalMux I__18181 (
            .O(N__90613),
            .I(shift_srl_73Z0Z_12));
    InMux I__18180 (
            .O(N__90610),
            .I(N__90607));
    LocalMux I__18179 (
            .O(N__90607),
            .I(shift_srl_73Z0Z_13));
    InMux I__18178 (
            .O(N__90604),
            .I(N__90601));
    LocalMux I__18177 (
            .O(N__90601),
            .I(shift_srl_73Z0Z_14));
    InMux I__18176 (
            .O(N__90598),
            .I(N__90595));
    LocalMux I__18175 (
            .O(N__90595),
            .I(shift_srl_73Z0Z_9));
    InMux I__18174 (
            .O(N__90592),
            .I(N__90589));
    LocalMux I__18173 (
            .O(N__90589),
            .I(shift_srl_73Z0Z_8));
    CascadeMux I__18172 (
            .O(N__90586),
            .I(N__90581));
    InMux I__18171 (
            .O(N__90585),
            .I(N__90572));
    InMux I__18170 (
            .O(N__90584),
            .I(N__90572));
    InMux I__18169 (
            .O(N__90581),
            .I(N__90572));
    CascadeMux I__18168 (
            .O(N__90580),
            .I(N__90566));
    CascadeMux I__18167 (
            .O(N__90579),
            .I(N__90547));
    LocalMux I__18166 (
            .O(N__90572),
            .I(N__90543));
    InMux I__18165 (
            .O(N__90571),
            .I(N__90534));
    InMux I__18164 (
            .O(N__90570),
            .I(N__90534));
    InMux I__18163 (
            .O(N__90569),
            .I(N__90534));
    InMux I__18162 (
            .O(N__90566),
            .I(N__90534));
    InMux I__18161 (
            .O(N__90565),
            .I(N__90523));
    InMux I__18160 (
            .O(N__90564),
            .I(N__90523));
    InMux I__18159 (
            .O(N__90563),
            .I(N__90523));
    CascadeMux I__18158 (
            .O(N__90562),
            .I(N__90520));
    InMux I__18157 (
            .O(N__90561),
            .I(N__90514));
    CascadeMux I__18156 (
            .O(N__90560),
            .I(N__90510));
    InMux I__18155 (
            .O(N__90559),
            .I(N__90501));
    InMux I__18154 (
            .O(N__90558),
            .I(N__90501));
    InMux I__18153 (
            .O(N__90557),
            .I(N__90501));
    InMux I__18152 (
            .O(N__90556),
            .I(N__90501));
    CascadeMux I__18151 (
            .O(N__90555),
            .I(N__90498));
    CascadeMux I__18150 (
            .O(N__90554),
            .I(N__90495));
    CascadeMux I__18149 (
            .O(N__90553),
            .I(N__90489));
    CascadeMux I__18148 (
            .O(N__90552),
            .I(N__90479));
    CascadeMux I__18147 (
            .O(N__90551),
            .I(N__90476));
    CascadeMux I__18146 (
            .O(N__90550),
            .I(N__90468));
    InMux I__18145 (
            .O(N__90547),
            .I(N__90465));
    CascadeMux I__18144 (
            .O(N__90546),
            .I(N__90455));
    Span4Mux_h I__18143 (
            .O(N__90543),
            .I(N__90444));
    LocalMux I__18142 (
            .O(N__90534),
            .I(N__90444));
    CascadeMux I__18141 (
            .O(N__90533),
            .I(N__90440));
    CascadeMux I__18140 (
            .O(N__90532),
            .I(N__90436));
    CascadeMux I__18139 (
            .O(N__90531),
            .I(N__90417));
    CascadeMux I__18138 (
            .O(N__90530),
            .I(N__90414));
    LocalMux I__18137 (
            .O(N__90523),
            .I(N__90410));
    InMux I__18136 (
            .O(N__90520),
            .I(N__90407));
    CascadeMux I__18135 (
            .O(N__90519),
            .I(N__90400));
    InMux I__18134 (
            .O(N__90518),
            .I(N__90396));
    CascadeMux I__18133 (
            .O(N__90517),
            .I(N__90392));
    LocalMux I__18132 (
            .O(N__90514),
            .I(N__90386));
    InMux I__18131 (
            .O(N__90513),
            .I(N__90381));
    InMux I__18130 (
            .O(N__90510),
            .I(N__90381));
    LocalMux I__18129 (
            .O(N__90501),
            .I(N__90378));
    InMux I__18128 (
            .O(N__90498),
            .I(N__90371));
    InMux I__18127 (
            .O(N__90495),
            .I(N__90371));
    InMux I__18126 (
            .O(N__90494),
            .I(N__90371));
    CascadeMux I__18125 (
            .O(N__90493),
            .I(N__90367));
    CascadeMux I__18124 (
            .O(N__90492),
            .I(N__90364));
    InMux I__18123 (
            .O(N__90489),
            .I(N__90357));
    InMux I__18122 (
            .O(N__90488),
            .I(N__90357));
    InMux I__18121 (
            .O(N__90487),
            .I(N__90357));
    InMux I__18120 (
            .O(N__90486),
            .I(N__90354));
    InMux I__18119 (
            .O(N__90485),
            .I(N__90351));
    CascadeMux I__18118 (
            .O(N__90484),
            .I(N__90346));
    CascadeMux I__18117 (
            .O(N__90483),
            .I(N__90341));
    InMux I__18116 (
            .O(N__90482),
            .I(N__90338));
    InMux I__18115 (
            .O(N__90479),
            .I(N__90335));
    InMux I__18114 (
            .O(N__90476),
            .I(N__90330));
    InMux I__18113 (
            .O(N__90475),
            .I(N__90330));
    CascadeMux I__18112 (
            .O(N__90474),
            .I(N__90325));
    InMux I__18111 (
            .O(N__90473),
            .I(N__90322));
    InMux I__18110 (
            .O(N__90472),
            .I(N__90313));
    InMux I__18109 (
            .O(N__90471),
            .I(N__90313));
    InMux I__18108 (
            .O(N__90468),
            .I(N__90310));
    LocalMux I__18107 (
            .O(N__90465),
            .I(N__90304));
    InMux I__18106 (
            .O(N__90464),
            .I(N__90301));
    InMux I__18105 (
            .O(N__90463),
            .I(N__90298));
    InMux I__18104 (
            .O(N__90462),
            .I(N__90293));
    InMux I__18103 (
            .O(N__90461),
            .I(N__90293));
    InMux I__18102 (
            .O(N__90460),
            .I(N__90289));
    InMux I__18101 (
            .O(N__90459),
            .I(N__90286));
    InMux I__18100 (
            .O(N__90458),
            .I(N__90282));
    InMux I__18099 (
            .O(N__90455),
            .I(N__90279));
    InMux I__18098 (
            .O(N__90454),
            .I(N__90273));
    InMux I__18097 (
            .O(N__90453),
            .I(N__90273));
    InMux I__18096 (
            .O(N__90452),
            .I(N__90266));
    InMux I__18095 (
            .O(N__90451),
            .I(N__90266));
    InMux I__18094 (
            .O(N__90450),
            .I(N__90266));
    InMux I__18093 (
            .O(N__90449),
            .I(N__90260));
    Span4Mux_v I__18092 (
            .O(N__90444),
            .I(N__90257));
    InMux I__18091 (
            .O(N__90443),
            .I(N__90248));
    InMux I__18090 (
            .O(N__90440),
            .I(N__90248));
    InMux I__18089 (
            .O(N__90439),
            .I(N__90248));
    InMux I__18088 (
            .O(N__90436),
            .I(N__90248));
    CascadeMux I__18087 (
            .O(N__90435),
            .I(N__90245));
    CascadeMux I__18086 (
            .O(N__90434),
            .I(N__90239));
    CascadeMux I__18085 (
            .O(N__90433),
            .I(N__90231));
    CascadeMux I__18084 (
            .O(N__90432),
            .I(N__90221));
    InMux I__18083 (
            .O(N__90431),
            .I(N__90218));
    InMux I__18082 (
            .O(N__90430),
            .I(N__90213));
    InMux I__18081 (
            .O(N__90429),
            .I(N__90213));
    CascadeMux I__18080 (
            .O(N__90428),
            .I(N__90207));
    CascadeMux I__18079 (
            .O(N__90427),
            .I(N__90204));
    InMux I__18078 (
            .O(N__90426),
            .I(N__90201));
    InMux I__18077 (
            .O(N__90425),
            .I(N__90198));
    InMux I__18076 (
            .O(N__90424),
            .I(N__90195));
    InMux I__18075 (
            .O(N__90423),
            .I(N__90190));
    InMux I__18074 (
            .O(N__90422),
            .I(N__90190));
    InMux I__18073 (
            .O(N__90421),
            .I(N__90187));
    InMux I__18072 (
            .O(N__90420),
            .I(N__90180));
    InMux I__18071 (
            .O(N__90417),
            .I(N__90175));
    InMux I__18070 (
            .O(N__90414),
            .I(N__90175));
    InMux I__18069 (
            .O(N__90413),
            .I(N__90172));
    Span4Mux_h I__18068 (
            .O(N__90410),
            .I(N__90167));
    LocalMux I__18067 (
            .O(N__90407),
            .I(N__90167));
    CascadeMux I__18066 (
            .O(N__90406),
            .I(N__90164));
    InMux I__18065 (
            .O(N__90405),
            .I(N__90158));
    InMux I__18064 (
            .O(N__90404),
            .I(N__90158));
    InMux I__18063 (
            .O(N__90403),
            .I(N__90153));
    InMux I__18062 (
            .O(N__90400),
            .I(N__90153));
    InMux I__18061 (
            .O(N__90399),
            .I(N__90150));
    LocalMux I__18060 (
            .O(N__90396),
            .I(N__90147));
    InMux I__18059 (
            .O(N__90395),
            .I(N__90142));
    InMux I__18058 (
            .O(N__90392),
            .I(N__90142));
    InMux I__18057 (
            .O(N__90391),
            .I(N__90134));
    InMux I__18056 (
            .O(N__90390),
            .I(N__90134));
    InMux I__18055 (
            .O(N__90389),
            .I(N__90134));
    Span4Mux_v I__18054 (
            .O(N__90386),
            .I(N__90130));
    LocalMux I__18053 (
            .O(N__90381),
            .I(N__90123));
    Span4Mux_h I__18052 (
            .O(N__90378),
            .I(N__90123));
    LocalMux I__18051 (
            .O(N__90371),
            .I(N__90123));
    InMux I__18050 (
            .O(N__90370),
            .I(N__90120));
    InMux I__18049 (
            .O(N__90367),
            .I(N__90117));
    InMux I__18048 (
            .O(N__90364),
            .I(N__90114));
    LocalMux I__18047 (
            .O(N__90357),
            .I(N__90109));
    LocalMux I__18046 (
            .O(N__90354),
            .I(N__90109));
    LocalMux I__18045 (
            .O(N__90351),
            .I(N__90106));
    InMux I__18044 (
            .O(N__90350),
            .I(N__90101));
    InMux I__18043 (
            .O(N__90349),
            .I(N__90101));
    InMux I__18042 (
            .O(N__90346),
            .I(N__90092));
    InMux I__18041 (
            .O(N__90345),
            .I(N__90092));
    InMux I__18040 (
            .O(N__90344),
            .I(N__90092));
    InMux I__18039 (
            .O(N__90341),
            .I(N__90092));
    LocalMux I__18038 (
            .O(N__90338),
            .I(N__90085));
    LocalMux I__18037 (
            .O(N__90335),
            .I(N__90085));
    LocalMux I__18036 (
            .O(N__90330),
            .I(N__90085));
    InMux I__18035 (
            .O(N__90329),
            .I(N__90078));
    InMux I__18034 (
            .O(N__90328),
            .I(N__90078));
    InMux I__18033 (
            .O(N__90325),
            .I(N__90078));
    LocalMux I__18032 (
            .O(N__90322),
            .I(N__90072));
    InMux I__18031 (
            .O(N__90321),
            .I(N__90068));
    InMux I__18030 (
            .O(N__90320),
            .I(N__90065));
    InMux I__18029 (
            .O(N__90319),
            .I(N__90062));
    InMux I__18028 (
            .O(N__90318),
            .I(N__90059));
    LocalMux I__18027 (
            .O(N__90313),
            .I(N__90054));
    LocalMux I__18026 (
            .O(N__90310),
            .I(N__90054));
    InMux I__18025 (
            .O(N__90309),
            .I(N__90051));
    InMux I__18024 (
            .O(N__90308),
            .I(N__90048));
    IoInMux I__18023 (
            .O(N__90307),
            .I(N__90045));
    Span4Mux_v I__18022 (
            .O(N__90304),
            .I(N__90033));
    LocalMux I__18021 (
            .O(N__90301),
            .I(N__90033));
    LocalMux I__18020 (
            .O(N__90298),
            .I(N__90033));
    LocalMux I__18019 (
            .O(N__90293),
            .I(N__90030));
    InMux I__18018 (
            .O(N__90292),
            .I(N__90027));
    LocalMux I__18017 (
            .O(N__90289),
            .I(N__90017));
    LocalMux I__18016 (
            .O(N__90286),
            .I(N__90017));
    CascadeMux I__18015 (
            .O(N__90285),
            .I(N__90014));
    LocalMux I__18014 (
            .O(N__90282),
            .I(N__90010));
    LocalMux I__18013 (
            .O(N__90279),
            .I(N__90007));
    InMux I__18012 (
            .O(N__90278),
            .I(N__90004));
    LocalMux I__18011 (
            .O(N__90273),
            .I(N__90001));
    LocalMux I__18010 (
            .O(N__90266),
            .I(N__89998));
    InMux I__18009 (
            .O(N__90265),
            .I(N__89993));
    InMux I__18008 (
            .O(N__90264),
            .I(N__89993));
    InMux I__18007 (
            .O(N__90263),
            .I(N__89990));
    LocalMux I__18006 (
            .O(N__90260),
            .I(N__89987));
    Span4Mux_h I__18005 (
            .O(N__90257),
            .I(N__89982));
    LocalMux I__18004 (
            .O(N__90248),
            .I(N__89982));
    InMux I__18003 (
            .O(N__90245),
            .I(N__89979));
    CascadeMux I__18002 (
            .O(N__90244),
            .I(N__89975));
    CascadeMux I__18001 (
            .O(N__90243),
            .I(N__89969));
    CascadeMux I__18000 (
            .O(N__90242),
            .I(N__89964));
    InMux I__17999 (
            .O(N__90239),
            .I(N__89959));
    InMux I__17998 (
            .O(N__90238),
            .I(N__89959));
    InMux I__17997 (
            .O(N__90237),
            .I(N__89952));
    InMux I__17996 (
            .O(N__90236),
            .I(N__89952));
    InMux I__17995 (
            .O(N__90235),
            .I(N__89952));
    InMux I__17994 (
            .O(N__90234),
            .I(N__89947));
    InMux I__17993 (
            .O(N__90231),
            .I(N__89940));
    InMux I__17992 (
            .O(N__90230),
            .I(N__89935));
    InMux I__17991 (
            .O(N__90229),
            .I(N__89935));
    CascadeMux I__17990 (
            .O(N__90228),
            .I(N__89932));
    InMux I__17989 (
            .O(N__90227),
            .I(N__89927));
    InMux I__17988 (
            .O(N__90226),
            .I(N__89922));
    InMux I__17987 (
            .O(N__90225),
            .I(N__89922));
    InMux I__17986 (
            .O(N__90224),
            .I(N__89917));
    InMux I__17985 (
            .O(N__90221),
            .I(N__89917));
    LocalMux I__17984 (
            .O(N__90218),
            .I(N__89911));
    LocalMux I__17983 (
            .O(N__90213),
            .I(N__89911));
    CascadeMux I__17982 (
            .O(N__90212),
            .I(N__89908));
    InMux I__17981 (
            .O(N__90211),
            .I(N__89903));
    InMux I__17980 (
            .O(N__90210),
            .I(N__89903));
    InMux I__17979 (
            .O(N__90207),
            .I(N__89897));
    InMux I__17978 (
            .O(N__90204),
            .I(N__89897));
    LocalMux I__17977 (
            .O(N__90201),
            .I(N__89892));
    LocalMux I__17976 (
            .O(N__90198),
            .I(N__89892));
    LocalMux I__17975 (
            .O(N__90195),
            .I(N__89887));
    LocalMux I__17974 (
            .O(N__90190),
            .I(N__89887));
    LocalMux I__17973 (
            .O(N__90187),
            .I(N__89884));
    InMux I__17972 (
            .O(N__90186),
            .I(N__89881));
    InMux I__17971 (
            .O(N__90185),
            .I(N__89876));
    InMux I__17970 (
            .O(N__90184),
            .I(N__89876));
    InMux I__17969 (
            .O(N__90183),
            .I(N__89873));
    LocalMux I__17968 (
            .O(N__90180),
            .I(N__89866));
    LocalMux I__17967 (
            .O(N__90175),
            .I(N__89866));
    LocalMux I__17966 (
            .O(N__90172),
            .I(N__89866));
    Span4Mux_v I__17965 (
            .O(N__90167),
            .I(N__89863));
    InMux I__17964 (
            .O(N__90164),
            .I(N__89858));
    InMux I__17963 (
            .O(N__90163),
            .I(N__89858));
    LocalMux I__17962 (
            .O(N__90158),
            .I(N__89853));
    LocalMux I__17961 (
            .O(N__90153),
            .I(N__89853));
    LocalMux I__17960 (
            .O(N__90150),
            .I(N__89850));
    Span4Mux_h I__17959 (
            .O(N__90147),
            .I(N__89845));
    LocalMux I__17958 (
            .O(N__90142),
            .I(N__89845));
    InMux I__17957 (
            .O(N__90141),
            .I(N__89842));
    LocalMux I__17956 (
            .O(N__90134),
            .I(N__89839));
    InMux I__17955 (
            .O(N__90133),
            .I(N__89836));
    Span4Mux_v I__17954 (
            .O(N__90130),
            .I(N__89831));
    Span4Mux_v I__17953 (
            .O(N__90123),
            .I(N__89831));
    LocalMux I__17952 (
            .O(N__90120),
            .I(N__89826));
    LocalMux I__17951 (
            .O(N__90117),
            .I(N__89826));
    LocalMux I__17950 (
            .O(N__90114),
            .I(N__89823));
    Span4Mux_v I__17949 (
            .O(N__90109),
            .I(N__89820));
    Span4Mux_h I__17948 (
            .O(N__90106),
            .I(N__89809));
    LocalMux I__17947 (
            .O(N__90101),
            .I(N__89809));
    LocalMux I__17946 (
            .O(N__90092),
            .I(N__89809));
    Span4Mux_v I__17945 (
            .O(N__90085),
            .I(N__89809));
    LocalMux I__17944 (
            .O(N__90078),
            .I(N__89809));
    CascadeMux I__17943 (
            .O(N__90077),
            .I(N__89806));
    CascadeMux I__17942 (
            .O(N__90076),
            .I(N__89803));
    CascadeMux I__17941 (
            .O(N__90075),
            .I(N__89800));
    Span4Mux_v I__17940 (
            .O(N__90072),
            .I(N__89795));
    CascadeMux I__17939 (
            .O(N__90071),
            .I(N__89789));
    LocalMux I__17938 (
            .O(N__90068),
            .I(N__89777));
    LocalMux I__17937 (
            .O(N__90065),
            .I(N__89777));
    LocalMux I__17936 (
            .O(N__90062),
            .I(N__89777));
    LocalMux I__17935 (
            .O(N__90059),
            .I(N__89777));
    Span4Mux_v I__17934 (
            .O(N__90054),
            .I(N__89774));
    LocalMux I__17933 (
            .O(N__90051),
            .I(N__89769));
    LocalMux I__17932 (
            .O(N__90048),
            .I(N__89769));
    LocalMux I__17931 (
            .O(N__90045),
            .I(N__89766));
    InMux I__17930 (
            .O(N__90044),
            .I(N__89762));
    CascadeMux I__17929 (
            .O(N__90043),
            .I(N__89756));
    CascadeMux I__17928 (
            .O(N__90042),
            .I(N__89753));
    InMux I__17927 (
            .O(N__90041),
            .I(N__89748));
    InMux I__17926 (
            .O(N__90040),
            .I(N__89748));
    Span4Mux_h I__17925 (
            .O(N__90033),
            .I(N__89743));
    Span4Mux_h I__17924 (
            .O(N__90030),
            .I(N__89743));
    LocalMux I__17923 (
            .O(N__90027),
            .I(N__89740));
    InMux I__17922 (
            .O(N__90026),
            .I(N__89729));
    InMux I__17921 (
            .O(N__90025),
            .I(N__89729));
    InMux I__17920 (
            .O(N__90024),
            .I(N__89729));
    InMux I__17919 (
            .O(N__90023),
            .I(N__89729));
    InMux I__17918 (
            .O(N__90022),
            .I(N__89729));
    Span4Mux_h I__17917 (
            .O(N__90017),
            .I(N__89726));
    InMux I__17916 (
            .O(N__90014),
            .I(N__89723));
    InMux I__17915 (
            .O(N__90013),
            .I(N__89720));
    Span4Mux_v I__17914 (
            .O(N__90010),
            .I(N__89717));
    Span12Mux_s9_v I__17913 (
            .O(N__90007),
            .I(N__89704));
    LocalMux I__17912 (
            .O(N__90004),
            .I(N__89704));
    Span12Mux_s9_h I__17911 (
            .O(N__90001),
            .I(N__89704));
    Sp12to4 I__17910 (
            .O(N__89998),
            .I(N__89704));
    LocalMux I__17909 (
            .O(N__89993),
            .I(N__89704));
    LocalMux I__17908 (
            .O(N__89990),
            .I(N__89704));
    Span4Mux_h I__17907 (
            .O(N__89987),
            .I(N__89701));
    Span4Mux_h I__17906 (
            .O(N__89982),
            .I(N__89696));
    LocalMux I__17905 (
            .O(N__89979),
            .I(N__89696));
    InMux I__17904 (
            .O(N__89978),
            .I(N__89687));
    InMux I__17903 (
            .O(N__89975),
            .I(N__89687));
    InMux I__17902 (
            .O(N__89974),
            .I(N__89687));
    InMux I__17901 (
            .O(N__89973),
            .I(N__89687));
    InMux I__17900 (
            .O(N__89972),
            .I(N__89684));
    InMux I__17899 (
            .O(N__89969),
            .I(N__89681));
    InMux I__17898 (
            .O(N__89968),
            .I(N__89674));
    InMux I__17897 (
            .O(N__89967),
            .I(N__89674));
    InMux I__17896 (
            .O(N__89964),
            .I(N__89674));
    LocalMux I__17895 (
            .O(N__89959),
            .I(N__89671));
    LocalMux I__17894 (
            .O(N__89952),
            .I(N__89668));
    InMux I__17893 (
            .O(N__89951),
            .I(N__89663));
    InMux I__17892 (
            .O(N__89950),
            .I(N__89663));
    LocalMux I__17891 (
            .O(N__89947),
            .I(N__89660));
    CascadeMux I__17890 (
            .O(N__89946),
            .I(N__89655));
    InMux I__17889 (
            .O(N__89945),
            .I(N__89648));
    InMux I__17888 (
            .O(N__89944),
            .I(N__89648));
    InMux I__17887 (
            .O(N__89943),
            .I(N__89648));
    LocalMux I__17886 (
            .O(N__89940),
            .I(N__89645));
    LocalMux I__17885 (
            .O(N__89935),
            .I(N__89642));
    InMux I__17884 (
            .O(N__89932),
            .I(N__89635));
    InMux I__17883 (
            .O(N__89931),
            .I(N__89635));
    InMux I__17882 (
            .O(N__89930),
            .I(N__89635));
    LocalMux I__17881 (
            .O(N__89927),
            .I(N__89628));
    LocalMux I__17880 (
            .O(N__89922),
            .I(N__89628));
    LocalMux I__17879 (
            .O(N__89917),
            .I(N__89628));
    InMux I__17878 (
            .O(N__89916),
            .I(N__89625));
    Span4Mux_v I__17877 (
            .O(N__89911),
            .I(N__89622));
    InMux I__17876 (
            .O(N__89908),
            .I(N__89619));
    LocalMux I__17875 (
            .O(N__89903),
            .I(N__89610));
    InMux I__17874 (
            .O(N__89902),
            .I(N__89607));
    LocalMux I__17873 (
            .O(N__89897),
            .I(N__89600));
    Span4Mux_v I__17872 (
            .O(N__89892),
            .I(N__89600));
    Span4Mux_h I__17871 (
            .O(N__89887),
            .I(N__89600));
    Span4Mux_h I__17870 (
            .O(N__89884),
            .I(N__89593));
    LocalMux I__17869 (
            .O(N__89881),
            .I(N__89593));
    LocalMux I__17868 (
            .O(N__89876),
            .I(N__89593));
    LocalMux I__17867 (
            .O(N__89873),
            .I(N__89590));
    Span4Mux_h I__17866 (
            .O(N__89866),
            .I(N__89587));
    Span4Mux_h I__17865 (
            .O(N__89863),
            .I(N__89582));
    LocalMux I__17864 (
            .O(N__89858),
            .I(N__89582));
    Span4Mux_h I__17863 (
            .O(N__89853),
            .I(N__89579));
    Span4Mux_h I__17862 (
            .O(N__89850),
            .I(N__89574));
    Span4Mux_v I__17861 (
            .O(N__89845),
            .I(N__89574));
    LocalMux I__17860 (
            .O(N__89842),
            .I(N__89571));
    Span4Mux_v I__17859 (
            .O(N__89839),
            .I(N__89568));
    LocalMux I__17858 (
            .O(N__89836),
            .I(N__89565));
    Span4Mux_v I__17857 (
            .O(N__89831),
            .I(N__89562));
    Span4Mux_v I__17856 (
            .O(N__89826),
            .I(N__89559));
    Span4Mux_v I__17855 (
            .O(N__89823),
            .I(N__89552));
    Span4Mux_h I__17854 (
            .O(N__89820),
            .I(N__89552));
    Span4Mux_v I__17853 (
            .O(N__89809),
            .I(N__89552));
    InMux I__17852 (
            .O(N__89806),
            .I(N__89549));
    InMux I__17851 (
            .O(N__89803),
            .I(N__89546));
    InMux I__17850 (
            .O(N__89800),
            .I(N__89539));
    InMux I__17849 (
            .O(N__89799),
            .I(N__89539));
    InMux I__17848 (
            .O(N__89798),
            .I(N__89539));
    Sp12to4 I__17847 (
            .O(N__89795),
            .I(N__89536));
    InMux I__17846 (
            .O(N__89794),
            .I(N__89531));
    InMux I__17845 (
            .O(N__89793),
            .I(N__89531));
    InMux I__17844 (
            .O(N__89792),
            .I(N__89526));
    InMux I__17843 (
            .O(N__89789),
            .I(N__89526));
    InMux I__17842 (
            .O(N__89788),
            .I(N__89519));
    InMux I__17841 (
            .O(N__89787),
            .I(N__89519));
    InMux I__17840 (
            .O(N__89786),
            .I(N__89516));
    Span12Mux_v I__17839 (
            .O(N__89777),
            .I(N__89509));
    Sp12to4 I__17838 (
            .O(N__89774),
            .I(N__89509));
    Span12Mux_v I__17837 (
            .O(N__89769),
            .I(N__89509));
    Span4Mux_s1_v I__17836 (
            .O(N__89766),
            .I(N__89506));
    InMux I__17835 (
            .O(N__89765),
            .I(N__89503));
    LocalMux I__17834 (
            .O(N__89762),
            .I(N__89500));
    InMux I__17833 (
            .O(N__89761),
            .I(N__89497));
    CascadeMux I__17832 (
            .O(N__89760),
            .I(N__89494));
    InMux I__17831 (
            .O(N__89759),
            .I(N__89491));
    InMux I__17830 (
            .O(N__89756),
            .I(N__89486));
    InMux I__17829 (
            .O(N__89753),
            .I(N__89486));
    LocalMux I__17828 (
            .O(N__89748),
            .I(N__89483));
    Span4Mux_h I__17827 (
            .O(N__89743),
            .I(N__89480));
    Span12Mux_s9_h I__17826 (
            .O(N__89740),
            .I(N__89465));
    LocalMux I__17825 (
            .O(N__89729),
            .I(N__89465));
    Sp12to4 I__17824 (
            .O(N__89726),
            .I(N__89465));
    LocalMux I__17823 (
            .O(N__89723),
            .I(N__89465));
    LocalMux I__17822 (
            .O(N__89720),
            .I(N__89465));
    Sp12to4 I__17821 (
            .O(N__89717),
            .I(N__89465));
    Span12Mux_v I__17820 (
            .O(N__89704),
            .I(N__89465));
    Span4Mux_h I__17819 (
            .O(N__89701),
            .I(N__89460));
    Span4Mux_h I__17818 (
            .O(N__89696),
            .I(N__89460));
    LocalMux I__17817 (
            .O(N__89687),
            .I(N__89455));
    LocalMux I__17816 (
            .O(N__89684),
            .I(N__89450));
    LocalMux I__17815 (
            .O(N__89681),
            .I(N__89450));
    LocalMux I__17814 (
            .O(N__89674),
            .I(N__89447));
    Span4Mux_v I__17813 (
            .O(N__89671),
            .I(N__89444));
    Span4Mux_h I__17812 (
            .O(N__89668),
            .I(N__89437));
    LocalMux I__17811 (
            .O(N__89663),
            .I(N__89437));
    Span4Mux_h I__17810 (
            .O(N__89660),
            .I(N__89437));
    InMux I__17809 (
            .O(N__89659),
            .I(N__89430));
    InMux I__17808 (
            .O(N__89658),
            .I(N__89430));
    InMux I__17807 (
            .O(N__89655),
            .I(N__89430));
    LocalMux I__17806 (
            .O(N__89648),
            .I(N__89421));
    Span4Mux_h I__17805 (
            .O(N__89645),
            .I(N__89421));
    Span4Mux_v I__17804 (
            .O(N__89642),
            .I(N__89421));
    LocalMux I__17803 (
            .O(N__89635),
            .I(N__89421));
    Span4Mux_v I__17802 (
            .O(N__89628),
            .I(N__89418));
    LocalMux I__17801 (
            .O(N__89625),
            .I(N__89411));
    Span4Mux_v I__17800 (
            .O(N__89622),
            .I(N__89411));
    LocalMux I__17799 (
            .O(N__89619),
            .I(N__89411));
    InMux I__17798 (
            .O(N__89618),
            .I(N__89408));
    InMux I__17797 (
            .O(N__89617),
            .I(N__89405));
    InMux I__17796 (
            .O(N__89616),
            .I(N__89402));
    InMux I__17795 (
            .O(N__89615),
            .I(N__89395));
    InMux I__17794 (
            .O(N__89614),
            .I(N__89395));
    InMux I__17793 (
            .O(N__89613),
            .I(N__89395));
    Span4Mux_h I__17792 (
            .O(N__89610),
            .I(N__89390));
    LocalMux I__17791 (
            .O(N__89607),
            .I(N__89390));
    Span4Mux_h I__17790 (
            .O(N__89600),
            .I(N__89385));
    Span4Mux_h I__17789 (
            .O(N__89593),
            .I(N__89385));
    Span4Mux_h I__17788 (
            .O(N__89590),
            .I(N__89378));
    Span4Mux_h I__17787 (
            .O(N__89587),
            .I(N__89378));
    Span4Mux_v I__17786 (
            .O(N__89582),
            .I(N__89378));
    Span4Mux_h I__17785 (
            .O(N__89579),
            .I(N__89373));
    Span4Mux_h I__17784 (
            .O(N__89574),
            .I(N__89373));
    Span12Mux_v I__17783 (
            .O(N__89571),
            .I(N__89360));
    Sp12to4 I__17782 (
            .O(N__89568),
            .I(N__89360));
    Span12Mux_s10_h I__17781 (
            .O(N__89565),
            .I(N__89360));
    Sp12to4 I__17780 (
            .O(N__89562),
            .I(N__89360));
    Sp12to4 I__17779 (
            .O(N__89559),
            .I(N__89360));
    Sp12to4 I__17778 (
            .O(N__89552),
            .I(N__89360));
    LocalMux I__17777 (
            .O(N__89549),
            .I(N__89347));
    LocalMux I__17776 (
            .O(N__89546),
            .I(N__89347));
    LocalMux I__17775 (
            .O(N__89539),
            .I(N__89347));
    Span12Mux_h I__17774 (
            .O(N__89536),
            .I(N__89347));
    LocalMux I__17773 (
            .O(N__89531),
            .I(N__89347));
    LocalMux I__17772 (
            .O(N__89526),
            .I(N__89347));
    InMux I__17771 (
            .O(N__89525),
            .I(N__89344));
    InMux I__17770 (
            .O(N__89524),
            .I(N__89341));
    LocalMux I__17769 (
            .O(N__89519),
            .I(N__89338));
    LocalMux I__17768 (
            .O(N__89516),
            .I(N__89335));
    Span12Mux_h I__17767 (
            .O(N__89509),
            .I(N__89332));
    Span4Mux_v I__17766 (
            .O(N__89506),
            .I(N__89328));
    LocalMux I__17765 (
            .O(N__89503),
            .I(N__89325));
    Span4Mux_h I__17764 (
            .O(N__89500),
            .I(N__89320));
    LocalMux I__17763 (
            .O(N__89497),
            .I(N__89320));
    InMux I__17762 (
            .O(N__89494),
            .I(N__89317));
    LocalMux I__17761 (
            .O(N__89491),
            .I(N__89304));
    LocalMux I__17760 (
            .O(N__89486),
            .I(N__89304));
    Span12Mux_s10_h I__17759 (
            .O(N__89483),
            .I(N__89304));
    Sp12to4 I__17758 (
            .O(N__89480),
            .I(N__89304));
    Span12Mux_h I__17757 (
            .O(N__89465),
            .I(N__89304));
    Sp12to4 I__17756 (
            .O(N__89460),
            .I(N__89304));
    InMux I__17755 (
            .O(N__89459),
            .I(N__89301));
    InMux I__17754 (
            .O(N__89458),
            .I(N__89298));
    Span4Mux_v I__17753 (
            .O(N__89455),
            .I(N__89293));
    Span4Mux_v I__17752 (
            .O(N__89450),
            .I(N__89293));
    Span4Mux_h I__17751 (
            .O(N__89447),
            .I(N__89286));
    Span4Mux_h I__17750 (
            .O(N__89444),
            .I(N__89286));
    Span4Mux_v I__17749 (
            .O(N__89437),
            .I(N__89286));
    LocalMux I__17748 (
            .O(N__89430),
            .I(N__89283));
    Span4Mux_v I__17747 (
            .O(N__89421),
            .I(N__89276));
    Span4Mux_h I__17746 (
            .O(N__89418),
            .I(N__89276));
    Span4Mux_v I__17745 (
            .O(N__89411),
            .I(N__89276));
    LocalMux I__17744 (
            .O(N__89408),
            .I(N__89255));
    LocalMux I__17743 (
            .O(N__89405),
            .I(N__89255));
    LocalMux I__17742 (
            .O(N__89402),
            .I(N__89255));
    LocalMux I__17741 (
            .O(N__89395),
            .I(N__89255));
    Sp12to4 I__17740 (
            .O(N__89390),
            .I(N__89255));
    Sp12to4 I__17739 (
            .O(N__89385),
            .I(N__89255));
    Sp12to4 I__17738 (
            .O(N__89378),
            .I(N__89255));
    Sp12to4 I__17737 (
            .O(N__89373),
            .I(N__89255));
    Span12Mux_h I__17736 (
            .O(N__89360),
            .I(N__89255));
    Span12Mux_v I__17735 (
            .O(N__89347),
            .I(N__89255));
    LocalMux I__17734 (
            .O(N__89344),
            .I(N__89244));
    LocalMux I__17733 (
            .O(N__89341),
            .I(N__89244));
    Sp12to4 I__17732 (
            .O(N__89338),
            .I(N__89244));
    Sp12to4 I__17731 (
            .O(N__89335),
            .I(N__89244));
    Span12Mux_h I__17730 (
            .O(N__89332),
            .I(N__89244));
    InMux I__17729 (
            .O(N__89331),
            .I(N__89241));
    Span4Mux_h I__17728 (
            .O(N__89328),
            .I(N__89234));
    Span4Mux_v I__17727 (
            .O(N__89325),
            .I(N__89234));
    Span4Mux_v I__17726 (
            .O(N__89320),
            .I(N__89234));
    LocalMux I__17725 (
            .O(N__89317),
            .I(N__89229));
    Span12Mux_v I__17724 (
            .O(N__89304),
            .I(N__89229));
    LocalMux I__17723 (
            .O(N__89301),
            .I(N__89214));
    LocalMux I__17722 (
            .O(N__89298),
            .I(N__89214));
    Sp12to4 I__17721 (
            .O(N__89293),
            .I(N__89214));
    Sp12to4 I__17720 (
            .O(N__89286),
            .I(N__89214));
    Span12Mux_v I__17719 (
            .O(N__89283),
            .I(N__89214));
    Sp12to4 I__17718 (
            .O(N__89276),
            .I(N__89214));
    Span12Mux_v I__17717 (
            .O(N__89255),
            .I(N__89214));
    Span12Mux_v I__17716 (
            .O(N__89244),
            .I(N__89211));
    LocalMux I__17715 (
            .O(N__89241),
            .I(rco_c_0));
    Odrv4 I__17714 (
            .O(N__89234),
            .I(rco_c_0));
    Odrv12 I__17713 (
            .O(N__89229),
            .I(rco_c_0));
    Odrv12 I__17712 (
            .O(N__89214),
            .I(rco_c_0));
    Odrv12 I__17711 (
            .O(N__89211),
            .I(rco_c_0));
    InMux I__17710 (
            .O(N__89200),
            .I(N__89197));
    LocalMux I__17709 (
            .O(N__89197),
            .I(shift_srl_73Z0Z_0));
    InMux I__17708 (
            .O(N__89194),
            .I(N__89191));
    LocalMux I__17707 (
            .O(N__89191),
            .I(shift_srl_73Z0Z_1));
    InMux I__17706 (
            .O(N__89188),
            .I(N__89185));
    LocalMux I__17705 (
            .O(N__89185),
            .I(shift_srl_168Z0Z_14));
    InMux I__17704 (
            .O(N__89182),
            .I(N__89171));
    InMux I__17703 (
            .O(N__89181),
            .I(N__89171));
    InMux I__17702 (
            .O(N__89180),
            .I(N__89171));
    InMux I__17701 (
            .O(N__89179),
            .I(N__89165));
    InMux I__17700 (
            .O(N__89178),
            .I(N__89165));
    LocalMux I__17699 (
            .O(N__89171),
            .I(N__89162));
    InMux I__17698 (
            .O(N__89170),
            .I(N__89159));
    LocalMux I__17697 (
            .O(N__89165),
            .I(N__89156));
    Span4Mux_h I__17696 (
            .O(N__89162),
            .I(N__89153));
    LocalMux I__17695 (
            .O(N__89159),
            .I(shift_srl_168Z0Z_15));
    Odrv12 I__17694 (
            .O(N__89156),
            .I(shift_srl_168Z0Z_15));
    Odrv4 I__17693 (
            .O(N__89153),
            .I(shift_srl_168Z0Z_15));
    InMux I__17692 (
            .O(N__89146),
            .I(N__89143));
    LocalMux I__17691 (
            .O(N__89143),
            .I(shift_srl_168Z0Z_12));
    InMux I__17690 (
            .O(N__89140),
            .I(N__89137));
    LocalMux I__17689 (
            .O(N__89137),
            .I(shift_srl_168Z0Z_7));
    InMux I__17688 (
            .O(N__89134),
            .I(N__89131));
    LocalMux I__17687 (
            .O(N__89131),
            .I(shift_srl_168Z0Z_8));
    InMux I__17686 (
            .O(N__89128),
            .I(N__89125));
    LocalMux I__17685 (
            .O(N__89125),
            .I(shift_srl_168Z0Z_9));
    InMux I__17684 (
            .O(N__89122),
            .I(N__89119));
    LocalMux I__17683 (
            .O(N__89119),
            .I(shift_srl_168Z0Z_10));
    InMux I__17682 (
            .O(N__89116),
            .I(N__89113));
    LocalMux I__17681 (
            .O(N__89113),
            .I(N__89110));
    Odrv4 I__17680 (
            .O(N__89110),
            .I(shift_srl_168Z0Z_11));
    CEMux I__17679 (
            .O(N__89107),
            .I(N__89101));
    CEMux I__17678 (
            .O(N__89106),
            .I(N__89098));
    CEMux I__17677 (
            .O(N__89105),
            .I(N__89095));
    CEMux I__17676 (
            .O(N__89104),
            .I(N__89092));
    LocalMux I__17675 (
            .O(N__89101),
            .I(N__89085));
    LocalMux I__17674 (
            .O(N__89098),
            .I(N__89085));
    LocalMux I__17673 (
            .O(N__89095),
            .I(N__89085));
    LocalMux I__17672 (
            .O(N__89092),
            .I(N__89082));
    Span4Mux_v I__17671 (
            .O(N__89085),
            .I(N__89079));
    Span4Mux_h I__17670 (
            .O(N__89082),
            .I(N__89076));
    Span4Mux_s3_h I__17669 (
            .O(N__89079),
            .I(N__89073));
    Odrv4 I__17668 (
            .O(N__89076),
            .I(clk_en_168));
    Odrv4 I__17667 (
            .O(N__89073),
            .I(clk_en_168));
    IoInMux I__17666 (
            .O(N__89068),
            .I(N__89065));
    LocalMux I__17665 (
            .O(N__89065),
            .I(N__89062));
    Odrv4 I__17664 (
            .O(N__89062),
            .I(rco_c_72));
    InMux I__17663 (
            .O(N__89059),
            .I(N__89056));
    LocalMux I__17662 (
            .O(N__89056),
            .I(shift_srl_73Z0Z_10));
    InMux I__17661 (
            .O(N__89053),
            .I(N__89050));
    LocalMux I__17660 (
            .O(N__89050),
            .I(shift_srl_172Z0Z_0));
    InMux I__17659 (
            .O(N__89047),
            .I(N__89044));
    LocalMux I__17658 (
            .O(N__89044),
            .I(shift_srl_172Z0Z_1));
    InMux I__17657 (
            .O(N__89041),
            .I(N__89038));
    LocalMux I__17656 (
            .O(N__89038),
            .I(shift_srl_172Z0Z_2));
    InMux I__17655 (
            .O(N__89035),
            .I(N__89032));
    LocalMux I__17654 (
            .O(N__89032),
            .I(shift_srl_172Z0Z_3));
    InMux I__17653 (
            .O(N__89029),
            .I(N__89026));
    LocalMux I__17652 (
            .O(N__89026),
            .I(shift_srl_172Z0Z_4));
    InMux I__17651 (
            .O(N__89023),
            .I(N__89020));
    LocalMux I__17650 (
            .O(N__89020),
            .I(shift_srl_172Z0Z_5));
    InMux I__17649 (
            .O(N__89017),
            .I(N__89014));
    LocalMux I__17648 (
            .O(N__89014),
            .I(shift_srl_172Z0Z_6));
    InMux I__17647 (
            .O(N__89011),
            .I(N__89008));
    LocalMux I__17646 (
            .O(N__89008),
            .I(shift_srl_172Z0Z_7));
    CEMux I__17645 (
            .O(N__89005),
            .I(N__89001));
    CEMux I__17644 (
            .O(N__89004),
            .I(N__88998));
    LocalMux I__17643 (
            .O(N__89001),
            .I(clk_en_172));
    LocalMux I__17642 (
            .O(N__88998),
            .I(clk_en_172));
    InMux I__17641 (
            .O(N__88993),
            .I(N__88990));
    LocalMux I__17640 (
            .O(N__88990),
            .I(shift_srl_168Z0Z_13));
    InMux I__17639 (
            .O(N__88987),
            .I(N__88984));
    LocalMux I__17638 (
            .O(N__88984),
            .I(shift_srl_172Z0Z_10));
    InMux I__17637 (
            .O(N__88981),
            .I(N__88978));
    LocalMux I__17636 (
            .O(N__88978),
            .I(shift_srl_172Z0Z_11));
    InMux I__17635 (
            .O(N__88975),
            .I(N__88972));
    LocalMux I__17634 (
            .O(N__88972),
            .I(shift_srl_172Z0Z_12));
    InMux I__17633 (
            .O(N__88969),
            .I(N__88966));
    LocalMux I__17632 (
            .O(N__88966),
            .I(shift_srl_172Z0Z_13));
    InMux I__17631 (
            .O(N__88963),
            .I(N__88960));
    LocalMux I__17630 (
            .O(N__88960),
            .I(shift_srl_172Z0Z_14));
    InMux I__17629 (
            .O(N__88957),
            .I(N__88954));
    LocalMux I__17628 (
            .O(N__88954),
            .I(shift_srl_172Z0Z_9));
    InMux I__17627 (
            .O(N__88951),
            .I(N__88948));
    LocalMux I__17626 (
            .O(N__88948),
            .I(shift_srl_172Z0Z_8));
    InMux I__17625 (
            .O(N__88945),
            .I(N__88942));
    LocalMux I__17624 (
            .O(N__88942),
            .I(N__88939));
    Span4Mux_v I__17623 (
            .O(N__88939),
            .I(N__88935));
    InMux I__17622 (
            .O(N__88938),
            .I(N__88932));
    Span4Mux_h I__17621 (
            .O(N__88935),
            .I(N__88929));
    LocalMux I__17620 (
            .O(N__88932),
            .I(shift_srl_172Z0Z_15));
    Odrv4 I__17619 (
            .O(N__88929),
            .I(shift_srl_172Z0Z_15));
    InMux I__17618 (
            .O(N__88924),
            .I(N__88921));
    LocalMux I__17617 (
            .O(N__88921),
            .I(shift_srl_74Z0Z_13));
    InMux I__17616 (
            .O(N__88918),
            .I(N__88915));
    LocalMux I__17615 (
            .O(N__88915),
            .I(shift_srl_74Z0Z_14));
    InMux I__17614 (
            .O(N__88912),
            .I(N__88908));
    InMux I__17613 (
            .O(N__88911),
            .I(N__88905));
    LocalMux I__17612 (
            .O(N__88908),
            .I(shift_srl_74Z0Z_15));
    LocalMux I__17611 (
            .O(N__88905),
            .I(shift_srl_74Z0Z_15));
    InMux I__17610 (
            .O(N__88900),
            .I(N__88897));
    LocalMux I__17609 (
            .O(N__88897),
            .I(shift_srl_74Z0Z_9));
    InMux I__17608 (
            .O(N__88894),
            .I(N__88891));
    LocalMux I__17607 (
            .O(N__88891),
            .I(shift_srl_74Z0Z_7));
    InMux I__17606 (
            .O(N__88888),
            .I(N__88885));
    LocalMux I__17605 (
            .O(N__88885),
            .I(shift_srl_74Z0Z_8));
    CEMux I__17604 (
            .O(N__88882),
            .I(N__88878));
    CEMux I__17603 (
            .O(N__88881),
            .I(N__88875));
    LocalMux I__17602 (
            .O(N__88878),
            .I(clk_en_74));
    LocalMux I__17601 (
            .O(N__88875),
            .I(clk_en_74));
    InMux I__17600 (
            .O(N__88870),
            .I(N__88867));
    LocalMux I__17599 (
            .O(N__88867),
            .I(shift_srl_32Z0Z_7));
    InMux I__17598 (
            .O(N__88864),
            .I(N__88861));
    LocalMux I__17597 (
            .O(N__88861),
            .I(shift_srl_32Z0Z_6));
    InMux I__17596 (
            .O(N__88858),
            .I(N__88855));
    LocalMux I__17595 (
            .O(N__88855),
            .I(shift_srl_32Z0Z_4));
    InMux I__17594 (
            .O(N__88852),
            .I(N__88849));
    LocalMux I__17593 (
            .O(N__88849),
            .I(shift_srl_32Z0Z_5));
    InMux I__17592 (
            .O(N__88846),
            .I(N__88843));
    LocalMux I__17591 (
            .O(N__88843),
            .I(shift_srl_32Z0Z_2));
    InMux I__17590 (
            .O(N__88840),
            .I(N__88837));
    LocalMux I__17589 (
            .O(N__88837),
            .I(shift_srl_32Z0Z_3));
    CEMux I__17588 (
            .O(N__88834),
            .I(N__88829));
    CEMux I__17587 (
            .O(N__88833),
            .I(N__88826));
    CEMux I__17586 (
            .O(N__88832),
            .I(N__88822));
    LocalMux I__17585 (
            .O(N__88829),
            .I(N__88817));
    LocalMux I__17584 (
            .O(N__88826),
            .I(N__88817));
    CEMux I__17583 (
            .O(N__88825),
            .I(N__88814));
    LocalMux I__17582 (
            .O(N__88822),
            .I(N__88811));
    Span4Mux_v I__17581 (
            .O(N__88817),
            .I(N__88808));
    LocalMux I__17580 (
            .O(N__88814),
            .I(N__88805));
    Span4Mux_h I__17579 (
            .O(N__88811),
            .I(N__88802));
    Span4Mux_s3_h I__17578 (
            .O(N__88808),
            .I(N__88799));
    Odrv4 I__17577 (
            .O(N__88805),
            .I(clk_en_32));
    Odrv4 I__17576 (
            .O(N__88802),
            .I(clk_en_32));
    Odrv4 I__17575 (
            .O(N__88799),
            .I(clk_en_32));
    InMux I__17574 (
            .O(N__88792),
            .I(N__88789));
    LocalMux I__17573 (
            .O(N__88789),
            .I(shift_srl_74Z0Z_2));
    InMux I__17572 (
            .O(N__88786),
            .I(N__88783));
    LocalMux I__17571 (
            .O(N__88783),
            .I(shift_srl_74Z0Z_3));
    InMux I__17570 (
            .O(N__88780),
            .I(N__88777));
    LocalMux I__17569 (
            .O(N__88777),
            .I(shift_srl_74Z0Z_4));
    InMux I__17568 (
            .O(N__88774),
            .I(N__88771));
    LocalMux I__17567 (
            .O(N__88771),
            .I(shift_srl_74Z0Z_5));
    InMux I__17566 (
            .O(N__88768),
            .I(N__88765));
    LocalMux I__17565 (
            .O(N__88765),
            .I(shift_srl_74Z0Z_6));
    InMux I__17564 (
            .O(N__88762),
            .I(N__88759));
    LocalMux I__17563 (
            .O(N__88759),
            .I(shift_srl_74Z0Z_10));
    InMux I__17562 (
            .O(N__88756),
            .I(N__88753));
    LocalMux I__17561 (
            .O(N__88753),
            .I(shift_srl_74Z0Z_11));
    InMux I__17560 (
            .O(N__88750),
            .I(N__88747));
    LocalMux I__17559 (
            .O(N__88747),
            .I(shift_srl_74Z0Z_12));
    InMux I__17558 (
            .O(N__88744),
            .I(N__88741));
    LocalMux I__17557 (
            .O(N__88741),
            .I(shift_srl_75Z0Z_9));
    InMux I__17556 (
            .O(N__88738),
            .I(N__88735));
    LocalMux I__17555 (
            .O(N__88735),
            .I(shift_srl_75Z0Z_8));
    InMux I__17554 (
            .O(N__88732),
            .I(N__88729));
    LocalMux I__17553 (
            .O(N__88729),
            .I(shift_srl_75Z0Z_7));
    InMux I__17552 (
            .O(N__88726),
            .I(N__88723));
    LocalMux I__17551 (
            .O(N__88723),
            .I(shift_srl_75Z0Z_6));
    InMux I__17550 (
            .O(N__88720),
            .I(N__88717));
    LocalMux I__17549 (
            .O(N__88717),
            .I(shift_srl_75Z0Z_5));
    InMux I__17548 (
            .O(N__88714),
            .I(N__88711));
    LocalMux I__17547 (
            .O(N__88711),
            .I(shift_srl_75Z0Z_3));
    InMux I__17546 (
            .O(N__88708),
            .I(N__88705));
    LocalMux I__17545 (
            .O(N__88705),
            .I(shift_srl_75Z0Z_4));
    CEMux I__17544 (
            .O(N__88702),
            .I(N__88697));
    CEMux I__17543 (
            .O(N__88701),
            .I(N__88694));
    CEMux I__17542 (
            .O(N__88700),
            .I(N__88691));
    LocalMux I__17541 (
            .O(N__88697),
            .I(N__88688));
    LocalMux I__17540 (
            .O(N__88694),
            .I(N__88685));
    LocalMux I__17539 (
            .O(N__88691),
            .I(N__88682));
    Span4Mux_h I__17538 (
            .O(N__88688),
            .I(N__88679));
    Span4Mux_v I__17537 (
            .O(N__88685),
            .I(N__88676));
    Span4Mux_v I__17536 (
            .O(N__88682),
            .I(N__88673));
    Odrv4 I__17535 (
            .O(N__88679),
            .I(clk_en_75));
    Odrv4 I__17534 (
            .O(N__88676),
            .I(clk_en_75));
    Odrv4 I__17533 (
            .O(N__88673),
            .I(clk_en_75));
    InMux I__17532 (
            .O(N__88666),
            .I(N__88663));
    LocalMux I__17531 (
            .O(N__88663),
            .I(shift_srl_74Z0Z_0));
    InMux I__17530 (
            .O(N__88660),
            .I(N__88657));
    LocalMux I__17529 (
            .O(N__88657),
            .I(shift_srl_74Z0Z_1));
    IoInMux I__17528 (
            .O(N__88654),
            .I(N__88651));
    LocalMux I__17527 (
            .O(N__88651),
            .I(N__88648));
    IoSpan4Mux I__17526 (
            .O(N__88648),
            .I(N__88645));
    Span4Mux_s0_h I__17525 (
            .O(N__88645),
            .I(N__88642));
    Odrv4 I__17524 (
            .O(N__88642),
            .I(rco_c_75));
    InMux I__17523 (
            .O(N__88639),
            .I(N__88636));
    LocalMux I__17522 (
            .O(N__88636),
            .I(N__88633));
    Span4Mux_v I__17521 (
            .O(N__88633),
            .I(N__88630));
    Odrv4 I__17520 (
            .O(N__88630),
            .I(shift_srl_76_RNIF788Z0Z_15));
    IoInMux I__17519 (
            .O(N__88627),
            .I(N__88624));
    LocalMux I__17518 (
            .O(N__88624),
            .I(N__88621));
    Span4Mux_s3_h I__17517 (
            .O(N__88621),
            .I(N__88618));
    Odrv4 I__17516 (
            .O(N__88618),
            .I(rco_c_76));
    InMux I__17515 (
            .O(N__88615),
            .I(N__88612));
    LocalMux I__17514 (
            .O(N__88612),
            .I(N__88606));
    InMux I__17513 (
            .O(N__88611),
            .I(N__88602));
    InMux I__17512 (
            .O(N__88610),
            .I(N__88597));
    InMux I__17511 (
            .O(N__88609),
            .I(N__88597));
    Span4Mux_v I__17510 (
            .O(N__88606),
            .I(N__88594));
    InMux I__17509 (
            .O(N__88605),
            .I(N__88591));
    LocalMux I__17508 (
            .O(N__88602),
            .I(N__88586));
    LocalMux I__17507 (
            .O(N__88597),
            .I(N__88586));
    Sp12to4 I__17506 (
            .O(N__88594),
            .I(N__88581));
    LocalMux I__17505 (
            .O(N__88591),
            .I(N__88578));
    Span4Mux_h I__17504 (
            .O(N__88586),
            .I(N__88575));
    InMux I__17503 (
            .O(N__88585),
            .I(N__88570));
    InMux I__17502 (
            .O(N__88584),
            .I(N__88570));
    Odrv12 I__17501 (
            .O(N__88581),
            .I(shift_srl_77_RNI8HLIZ0Z_15));
    Odrv4 I__17500 (
            .O(N__88578),
            .I(shift_srl_77_RNI8HLIZ0Z_15));
    Odrv4 I__17499 (
            .O(N__88575),
            .I(shift_srl_77_RNI8HLIZ0Z_15));
    LocalMux I__17498 (
            .O(N__88570),
            .I(shift_srl_77_RNI8HLIZ0Z_15));
    IoInMux I__17497 (
            .O(N__88561),
            .I(N__88558));
    LocalMux I__17496 (
            .O(N__88558),
            .I(N__88555));
    Span12Mux_s3_h I__17495 (
            .O(N__88555),
            .I(N__88552));
    Odrv12 I__17494 (
            .O(N__88552),
            .I(rco_c_77));
    InMux I__17493 (
            .O(N__88549),
            .I(N__88546));
    LocalMux I__17492 (
            .O(N__88546),
            .I(N__88538));
    InMux I__17491 (
            .O(N__88545),
            .I(N__88535));
    InMux I__17490 (
            .O(N__88544),
            .I(N__88524));
    InMux I__17489 (
            .O(N__88543),
            .I(N__88524));
    InMux I__17488 (
            .O(N__88542),
            .I(N__88524));
    InMux I__17487 (
            .O(N__88541),
            .I(N__88524));
    Span4Mux_s1_v I__17486 (
            .O(N__88538),
            .I(N__88518));
    LocalMux I__17485 (
            .O(N__88535),
            .I(N__88518));
    InMux I__17484 (
            .O(N__88534),
            .I(N__88513));
    InMux I__17483 (
            .O(N__88533),
            .I(N__88513));
    LocalMux I__17482 (
            .O(N__88524),
            .I(N__88510));
    IoInMux I__17481 (
            .O(N__88523),
            .I(N__88505));
    Span4Mux_v I__17480 (
            .O(N__88518),
            .I(N__88500));
    LocalMux I__17479 (
            .O(N__88513),
            .I(N__88500));
    Span4Mux_v I__17478 (
            .O(N__88510),
            .I(N__88497));
    InMux I__17477 (
            .O(N__88509),
            .I(N__88492));
    InMux I__17476 (
            .O(N__88508),
            .I(N__88492));
    LocalMux I__17475 (
            .O(N__88505),
            .I(N__88489));
    Span4Mux_h I__17474 (
            .O(N__88500),
            .I(N__88486));
    Span4Mux_h I__17473 (
            .O(N__88497),
            .I(N__88481));
    LocalMux I__17472 (
            .O(N__88492),
            .I(N__88481));
    Span12Mux_s9_v I__17471 (
            .O(N__88489),
            .I(N__88478));
    Span4Mux_v I__17470 (
            .O(N__88486),
            .I(N__88475));
    Span4Mux_h I__17469 (
            .O(N__88481),
            .I(N__88472));
    Odrv12 I__17468 (
            .O(N__88478),
            .I(rco_c_74));
    Odrv4 I__17467 (
            .O(N__88475),
            .I(rco_c_74));
    Odrv4 I__17466 (
            .O(N__88472),
            .I(rco_c_74));
    InMux I__17465 (
            .O(N__88465),
            .I(N__88461));
    CascadeMux I__17464 (
            .O(N__88464),
            .I(N__88457));
    LocalMux I__17463 (
            .O(N__88461),
            .I(N__88454));
    InMux I__17462 (
            .O(N__88460),
            .I(N__88451));
    InMux I__17461 (
            .O(N__88457),
            .I(N__88448));
    Span4Mux_v I__17460 (
            .O(N__88454),
            .I(N__88444));
    LocalMux I__17459 (
            .O(N__88451),
            .I(N__88439));
    LocalMux I__17458 (
            .O(N__88448),
            .I(N__88439));
    CascadeMux I__17457 (
            .O(N__88447),
            .I(N__88435));
    Span4Mux_h I__17456 (
            .O(N__88444),
            .I(N__88432));
    Span4Mux_v I__17455 (
            .O(N__88439),
            .I(N__88429));
    InMux I__17454 (
            .O(N__88438),
            .I(N__88424));
    InMux I__17453 (
            .O(N__88435),
            .I(N__88424));
    Odrv4 I__17452 (
            .O(N__88432),
            .I(shift_srl_80_RNIG3FB1Z0Z_15));
    Odrv4 I__17451 (
            .O(N__88429),
            .I(shift_srl_80_RNIG3FB1Z0Z_15));
    LocalMux I__17450 (
            .O(N__88424),
            .I(shift_srl_80_RNIG3FB1Z0Z_15));
    IoInMux I__17449 (
            .O(N__88417),
            .I(N__88414));
    LocalMux I__17448 (
            .O(N__88414),
            .I(N__88411));
    IoSpan4Mux I__17447 (
            .O(N__88411),
            .I(N__88408));
    Odrv4 I__17446 (
            .O(N__88408),
            .I(rco_c_80));
    InMux I__17445 (
            .O(N__88405),
            .I(N__88398));
    InMux I__17444 (
            .O(N__88404),
            .I(N__88398));
    InMux I__17443 (
            .O(N__88403),
            .I(N__88395));
    LocalMux I__17442 (
            .O(N__88398),
            .I(N__88391));
    LocalMux I__17441 (
            .O(N__88395),
            .I(N__88387));
    InMux I__17440 (
            .O(N__88394),
            .I(N__88384));
    Span4Mux_h I__17439 (
            .O(N__88391),
            .I(N__88381));
    InMux I__17438 (
            .O(N__88390),
            .I(N__88378));
    Span4Mux_v I__17437 (
            .O(N__88387),
            .I(N__88373));
    LocalMux I__17436 (
            .O(N__88384),
            .I(N__88373));
    Odrv4 I__17435 (
            .O(N__88381),
            .I(shift_srl_75Z0Z_15));
    LocalMux I__17434 (
            .O(N__88378),
            .I(shift_srl_75Z0Z_15));
    Odrv4 I__17433 (
            .O(N__88373),
            .I(shift_srl_75Z0Z_15));
    InMux I__17432 (
            .O(N__88366),
            .I(N__88363));
    LocalMux I__17431 (
            .O(N__88363),
            .I(shift_srl_75Z0Z_0));
    InMux I__17430 (
            .O(N__88360),
            .I(N__88357));
    LocalMux I__17429 (
            .O(N__88357),
            .I(shift_srl_75Z0Z_1));
    InMux I__17428 (
            .O(N__88354),
            .I(N__88351));
    LocalMux I__17427 (
            .O(N__88351),
            .I(shift_srl_75Z0Z_2));
    InMux I__17426 (
            .O(N__88348),
            .I(N__88345));
    LocalMux I__17425 (
            .O(N__88345),
            .I(N__88342));
    Span4Mux_h I__17424 (
            .O(N__88342),
            .I(N__88339));
    Odrv4 I__17423 (
            .O(N__88339),
            .I(shift_srl_75Z0Z_10));
    InMux I__17422 (
            .O(N__88336),
            .I(N__88333));
    LocalMux I__17421 (
            .O(N__88333),
            .I(N__88330));
    Span4Mux_v I__17420 (
            .O(N__88330),
            .I(N__88326));
    CascadeMux I__17419 (
            .O(N__88329),
            .I(N__88321));
    Span4Mux_h I__17418 (
            .O(N__88326),
            .I(N__88317));
    InMux I__17417 (
            .O(N__88325),
            .I(N__88310));
    InMux I__17416 (
            .O(N__88324),
            .I(N__88310));
    InMux I__17415 (
            .O(N__88321),
            .I(N__88310));
    CascadeMux I__17414 (
            .O(N__88320),
            .I(N__88307));
    Span4Mux_h I__17413 (
            .O(N__88317),
            .I(N__88304));
    LocalMux I__17412 (
            .O(N__88310),
            .I(N__88301));
    InMux I__17411 (
            .O(N__88307),
            .I(N__88298));
    Odrv4 I__17410 (
            .O(N__88304),
            .I(shift_srl_50_RNI869CZ0Z_15));
    Odrv4 I__17409 (
            .O(N__88301),
            .I(shift_srl_50_RNI869CZ0Z_15));
    LocalMux I__17408 (
            .O(N__88298),
            .I(shift_srl_50_RNI869CZ0Z_15));
    IoInMux I__17407 (
            .O(N__88291),
            .I(N__88288));
    LocalMux I__17406 (
            .O(N__88288),
            .I(N__88285));
    IoSpan4Mux I__17405 (
            .O(N__88285),
            .I(N__88282));
    Odrv4 I__17404 (
            .O(N__88282),
            .I(rco_c_50));
    InMux I__17403 (
            .O(N__88279),
            .I(N__88275));
    InMux I__17402 (
            .O(N__88278),
            .I(N__88272));
    LocalMux I__17401 (
            .O(N__88275),
            .I(N__88269));
    LocalMux I__17400 (
            .O(N__88272),
            .I(N__88266));
    Odrv4 I__17399 (
            .O(N__88269),
            .I(shift_srl_77Z0Z_15));
    Odrv12 I__17398 (
            .O(N__88266),
            .I(shift_srl_77Z0Z_15));
    InMux I__17397 (
            .O(N__88261),
            .I(N__88258));
    LocalMux I__17396 (
            .O(N__88258),
            .I(shift_srl_77Z0Z_0));
    InMux I__17395 (
            .O(N__88255),
            .I(N__88252));
    LocalMux I__17394 (
            .O(N__88252),
            .I(shift_srl_77Z0Z_1));
    InMux I__17393 (
            .O(N__88249),
            .I(N__88246));
    LocalMux I__17392 (
            .O(N__88246),
            .I(shift_srl_77Z0Z_2));
    InMux I__17391 (
            .O(N__88243),
            .I(N__88240));
    LocalMux I__17390 (
            .O(N__88240),
            .I(shift_srl_77Z0Z_3));
    InMux I__17389 (
            .O(N__88237),
            .I(N__88234));
    LocalMux I__17388 (
            .O(N__88234),
            .I(shift_srl_77Z0Z_4));
    InMux I__17387 (
            .O(N__88231),
            .I(N__88228));
    LocalMux I__17386 (
            .O(N__88228),
            .I(shift_srl_77Z0Z_5));
    InMux I__17385 (
            .O(N__88225),
            .I(N__88222));
    LocalMux I__17384 (
            .O(N__88222),
            .I(shift_srl_77Z0Z_6));
    InMux I__17383 (
            .O(N__88219),
            .I(N__88216));
    LocalMux I__17382 (
            .O(N__88216),
            .I(N__88213));
    Span4Mux_h I__17381 (
            .O(N__88213),
            .I(N__88210));
    Odrv4 I__17380 (
            .O(N__88210),
            .I(shift_srl_77Z0Z_7));
    CEMux I__17379 (
            .O(N__88207),
            .I(N__88204));
    LocalMux I__17378 (
            .O(N__88204),
            .I(N__88200));
    CEMux I__17377 (
            .O(N__88203),
            .I(N__88197));
    Span4Mux_h I__17376 (
            .O(N__88200),
            .I(N__88194));
    LocalMux I__17375 (
            .O(N__88197),
            .I(N__88191));
    Odrv4 I__17374 (
            .O(N__88194),
            .I(clk_en_77));
    Odrv4 I__17373 (
            .O(N__88191),
            .I(clk_en_77));
    InMux I__17372 (
            .O(N__88186),
            .I(N__88183));
    LocalMux I__17371 (
            .O(N__88183),
            .I(shift_srl_190Z0Z_8));
    InMux I__17370 (
            .O(N__88180),
            .I(N__88177));
    LocalMux I__17369 (
            .O(N__88177),
            .I(shift_srl_190Z0Z_6));
    InMux I__17368 (
            .O(N__88174),
            .I(N__88171));
    LocalMux I__17367 (
            .O(N__88171),
            .I(shift_srl_190Z0Z_7));
    InMux I__17366 (
            .O(N__88168),
            .I(N__88165));
    LocalMux I__17365 (
            .O(N__88165),
            .I(shift_srl_190Z0Z_12));
    InMux I__17364 (
            .O(N__88162),
            .I(N__88159));
    LocalMux I__17363 (
            .O(N__88159),
            .I(shift_srl_190Z0Z_13));
    InMux I__17362 (
            .O(N__88156),
            .I(N__88153));
    LocalMux I__17361 (
            .O(N__88153),
            .I(shift_srl_190Z0Z_14));
    InMux I__17360 (
            .O(N__88150),
            .I(N__88147));
    LocalMux I__17359 (
            .O(N__88147),
            .I(shift_srl_190Z0Z_2));
    InMux I__17358 (
            .O(N__88144),
            .I(N__88141));
    LocalMux I__17357 (
            .O(N__88141),
            .I(shift_srl_190Z0Z_0));
    InMux I__17356 (
            .O(N__88138),
            .I(N__88135));
    LocalMux I__17355 (
            .O(N__88135),
            .I(shift_srl_190Z0Z_1));
    CEMux I__17354 (
            .O(N__88132),
            .I(N__88129));
    LocalMux I__17353 (
            .O(N__88129),
            .I(N__88125));
    CEMux I__17352 (
            .O(N__88128),
            .I(N__88122));
    Span4Mux_h I__17351 (
            .O(N__88125),
            .I(N__88117));
    LocalMux I__17350 (
            .O(N__88122),
            .I(N__88117));
    Odrv4 I__17349 (
            .O(N__88117),
            .I(clk_en_190));
    InMux I__17348 (
            .O(N__88114),
            .I(N__88109));
    InMux I__17347 (
            .O(N__88113),
            .I(N__88106));
    InMux I__17346 (
            .O(N__88112),
            .I(N__88103));
    LocalMux I__17345 (
            .O(N__88109),
            .I(N__88098));
    LocalMux I__17344 (
            .O(N__88106),
            .I(N__88092));
    LocalMux I__17343 (
            .O(N__88103),
            .I(N__88092));
    InMux I__17342 (
            .O(N__88102),
            .I(N__88087));
    InMux I__17341 (
            .O(N__88101),
            .I(N__88087));
    Span12Mux_v I__17340 (
            .O(N__88098),
            .I(N__88084));
    InMux I__17339 (
            .O(N__88097),
            .I(N__88081));
    Span4Mux_v I__17338 (
            .O(N__88092),
            .I(N__88076));
    LocalMux I__17337 (
            .O(N__88087),
            .I(N__88076));
    Odrv12 I__17336 (
            .O(N__88084),
            .I(shift_srl_139Z0Z_15));
    LocalMux I__17335 (
            .O(N__88081),
            .I(shift_srl_139Z0Z_15));
    Odrv4 I__17334 (
            .O(N__88076),
            .I(shift_srl_139Z0Z_15));
    IoInMux I__17333 (
            .O(N__88069),
            .I(N__88066));
    LocalMux I__17332 (
            .O(N__88066),
            .I(N__88063));
    Span4Mux_s1_h I__17331 (
            .O(N__88063),
            .I(N__88060));
    Span4Mux_v I__17330 (
            .O(N__88060),
            .I(N__88057));
    Odrv4 I__17329 (
            .O(N__88057),
            .I(rco_c_139));
    InMux I__17328 (
            .O(N__88054),
            .I(N__88051));
    LocalMux I__17327 (
            .O(N__88051),
            .I(shift_srl_168Z0Z_6));
    InMux I__17326 (
            .O(N__88048),
            .I(N__88045));
    LocalMux I__17325 (
            .O(N__88045),
            .I(shift_srl_190Z0Z_9));
    InMux I__17324 (
            .O(N__88042),
            .I(N__88039));
    LocalMux I__17323 (
            .O(N__88039),
            .I(shift_srl_190Z0Z_3));
    InMux I__17322 (
            .O(N__88036),
            .I(N__88033));
    LocalMux I__17321 (
            .O(N__88033),
            .I(shift_srl_190Z0Z_4));
    InMux I__17320 (
            .O(N__88030),
            .I(N__88027));
    LocalMux I__17319 (
            .O(N__88027),
            .I(shift_srl_190Z0Z_10));
    InMux I__17318 (
            .O(N__88024),
            .I(N__88021));
    LocalMux I__17317 (
            .O(N__88021),
            .I(shift_srl_190Z0Z_5));
    InMux I__17316 (
            .O(N__88018),
            .I(N__88015));
    LocalMux I__17315 (
            .O(N__88015),
            .I(shift_srl_190Z0Z_11));
    CascadeMux I__17314 (
            .O(N__88012),
            .I(N__88006));
    InMux I__17313 (
            .O(N__88011),
            .I(N__87997));
    InMux I__17312 (
            .O(N__88010),
            .I(N__87997));
    InMux I__17311 (
            .O(N__88009),
            .I(N__87997));
    InMux I__17310 (
            .O(N__88006),
            .I(N__87993));
    CascadeMux I__17309 (
            .O(N__88005),
            .I(N__87989));
    CascadeMux I__17308 (
            .O(N__88004),
            .I(N__87985));
    LocalMux I__17307 (
            .O(N__87997),
            .I(N__87981));
    InMux I__17306 (
            .O(N__87996),
            .I(N__87978));
    LocalMux I__17305 (
            .O(N__87993),
            .I(N__87975));
    InMux I__17304 (
            .O(N__87992),
            .I(N__87972));
    InMux I__17303 (
            .O(N__87989),
            .I(N__87967));
    InMux I__17302 (
            .O(N__87988),
            .I(N__87967));
    InMux I__17301 (
            .O(N__87985),
            .I(N__87964));
    InMux I__17300 (
            .O(N__87984),
            .I(N__87961));
    Span4Mux_v I__17299 (
            .O(N__87981),
            .I(N__87957));
    LocalMux I__17298 (
            .O(N__87978),
            .I(N__87954));
    Span4Mux_v I__17297 (
            .O(N__87975),
            .I(N__87947));
    LocalMux I__17296 (
            .O(N__87972),
            .I(N__87947));
    LocalMux I__17295 (
            .O(N__87967),
            .I(N__87947));
    LocalMux I__17294 (
            .O(N__87964),
            .I(N__87944));
    LocalMux I__17293 (
            .O(N__87961),
            .I(N__87941));
    InMux I__17292 (
            .O(N__87960),
            .I(N__87938));
    Span4Mux_h I__17291 (
            .O(N__87957),
            .I(N__87933));
    Span4Mux_v I__17290 (
            .O(N__87954),
            .I(N__87933));
    Span4Mux_v I__17289 (
            .O(N__87947),
            .I(N__87930));
    Span4Mux_h I__17288 (
            .O(N__87944),
            .I(N__87925));
    Span4Mux_v I__17287 (
            .O(N__87941),
            .I(N__87925));
    LocalMux I__17286 (
            .O(N__87938),
            .I(rco_int_0_a3_0_a2_0_162));
    Odrv4 I__17285 (
            .O(N__87933),
            .I(rco_int_0_a3_0_a2_0_162));
    Odrv4 I__17284 (
            .O(N__87930),
            .I(rco_int_0_a3_0_a2_0_162));
    Odrv4 I__17283 (
            .O(N__87925),
            .I(rco_int_0_a3_0_a2_0_162));
    IoInMux I__17282 (
            .O(N__87916),
            .I(N__87913));
    LocalMux I__17281 (
            .O(N__87913),
            .I(N__87910));
    Span4Mux_s1_h I__17280 (
            .O(N__87910),
            .I(N__87901));
    InMux I__17279 (
            .O(N__87909),
            .I(N__87887));
    InMux I__17278 (
            .O(N__87908),
            .I(N__87887));
    InMux I__17277 (
            .O(N__87907),
            .I(N__87887));
    InMux I__17276 (
            .O(N__87906),
            .I(N__87887));
    InMux I__17275 (
            .O(N__87905),
            .I(N__87887));
    InMux I__17274 (
            .O(N__87904),
            .I(N__87887));
    Span4Mux_h I__17273 (
            .O(N__87901),
            .I(N__87884));
    InMux I__17272 (
            .O(N__87900),
            .I(N__87881));
    LocalMux I__17271 (
            .O(N__87887),
            .I(N__87876));
    Sp12to4 I__17270 (
            .O(N__87884),
            .I(N__87870));
    LocalMux I__17269 (
            .O(N__87881),
            .I(N__87866));
    InMux I__17268 (
            .O(N__87880),
            .I(N__87861));
    InMux I__17267 (
            .O(N__87879),
            .I(N__87861));
    Span4Mux_h I__17266 (
            .O(N__87876),
            .I(N__87858));
    InMux I__17265 (
            .O(N__87875),
            .I(N__87851));
    InMux I__17264 (
            .O(N__87874),
            .I(N__87851));
    InMux I__17263 (
            .O(N__87873),
            .I(N__87851));
    Span12Mux_v I__17262 (
            .O(N__87870),
            .I(N__87848));
    CascadeMux I__17261 (
            .O(N__87869),
            .I(N__87845));
    Span4Mux_v I__17260 (
            .O(N__87866),
            .I(N__87839));
    LocalMux I__17259 (
            .O(N__87861),
            .I(N__87836));
    Sp12to4 I__17258 (
            .O(N__87858),
            .I(N__87833));
    LocalMux I__17257 (
            .O(N__87851),
            .I(N__87830));
    Span12Mux_h I__17256 (
            .O(N__87848),
            .I(N__87827));
    InMux I__17255 (
            .O(N__87845),
            .I(N__87818));
    InMux I__17254 (
            .O(N__87844),
            .I(N__87818));
    InMux I__17253 (
            .O(N__87843),
            .I(N__87818));
    InMux I__17252 (
            .O(N__87842),
            .I(N__87818));
    Span4Mux_h I__17251 (
            .O(N__87839),
            .I(N__87815));
    Span4Mux_h I__17250 (
            .O(N__87836),
            .I(N__87812));
    Span12Mux_v I__17249 (
            .O(N__87833),
            .I(N__87807));
    Span12Mux_s9_h I__17248 (
            .O(N__87830),
            .I(N__87807));
    Odrv12 I__17247 (
            .O(N__87827),
            .I(rco_c_153));
    LocalMux I__17246 (
            .O(N__87818),
            .I(rco_c_153));
    Odrv4 I__17245 (
            .O(N__87815),
            .I(rco_c_153));
    Odrv4 I__17244 (
            .O(N__87812),
            .I(rco_c_153));
    Odrv12 I__17243 (
            .O(N__87807),
            .I(rco_c_153));
    CEMux I__17242 (
            .O(N__87796),
            .I(N__87792));
    CEMux I__17241 (
            .O(N__87795),
            .I(N__87789));
    LocalMux I__17240 (
            .O(N__87792),
            .I(N__87786));
    LocalMux I__17239 (
            .O(N__87789),
            .I(N__87782));
    Span4Mux_h I__17238 (
            .O(N__87786),
            .I(N__87779));
    CEMux I__17237 (
            .O(N__87785),
            .I(N__87776));
    Span4Mux_h I__17236 (
            .O(N__87782),
            .I(N__87773));
    Sp12to4 I__17235 (
            .O(N__87779),
            .I(N__87768));
    LocalMux I__17234 (
            .O(N__87776),
            .I(N__87768));
    Odrv4 I__17233 (
            .O(N__87773),
            .I(clk_en_164));
    Odrv12 I__17232 (
            .O(N__87768),
            .I(clk_en_164));
    InMux I__17231 (
            .O(N__87763),
            .I(N__87758));
    InMux I__17230 (
            .O(N__87762),
            .I(N__87753));
    InMux I__17229 (
            .O(N__87761),
            .I(N__87753));
    LocalMux I__17228 (
            .O(N__87758),
            .I(N__87750));
    LocalMux I__17227 (
            .O(N__87753),
            .I(N__87746));
    Span4Mux_h I__17226 (
            .O(N__87750),
            .I(N__87743));
    InMux I__17225 (
            .O(N__87749),
            .I(N__87739));
    Span4Mux_h I__17224 (
            .O(N__87746),
            .I(N__87734));
    Span4Mux_v I__17223 (
            .O(N__87743),
            .I(N__87734));
    InMux I__17222 (
            .O(N__87742),
            .I(N__87731));
    LocalMux I__17221 (
            .O(N__87739),
            .I(shift_srl_163Z0Z_15));
    Odrv4 I__17220 (
            .O(N__87734),
            .I(shift_srl_163Z0Z_15));
    LocalMux I__17219 (
            .O(N__87731),
            .I(shift_srl_163Z0Z_15));
    InMux I__17218 (
            .O(N__87724),
            .I(N__87721));
    LocalMux I__17217 (
            .O(N__87721),
            .I(N__87713));
    IoInMux I__17216 (
            .O(N__87720),
            .I(N__87709));
    InMux I__17215 (
            .O(N__87719),
            .I(N__87699));
    InMux I__17214 (
            .O(N__87718),
            .I(N__87699));
    InMux I__17213 (
            .O(N__87717),
            .I(N__87699));
    InMux I__17212 (
            .O(N__87716),
            .I(N__87699));
    Span4Mux_v I__17211 (
            .O(N__87713),
            .I(N__87695));
    CascadeMux I__17210 (
            .O(N__87712),
            .I(N__87692));
    LocalMux I__17209 (
            .O(N__87709),
            .I(N__87688));
    InMux I__17208 (
            .O(N__87708),
            .I(N__87685));
    LocalMux I__17207 (
            .O(N__87699),
            .I(N__87682));
    InMux I__17206 (
            .O(N__87698),
            .I(N__87679));
    Span4Mux_v I__17205 (
            .O(N__87695),
            .I(N__87676));
    InMux I__17204 (
            .O(N__87692),
            .I(N__87671));
    InMux I__17203 (
            .O(N__87691),
            .I(N__87671));
    Span12Mux_s0_v I__17202 (
            .O(N__87688),
            .I(N__87666));
    LocalMux I__17201 (
            .O(N__87685),
            .I(N__87663));
    Span4Mux_v I__17200 (
            .O(N__87682),
            .I(N__87657));
    LocalMux I__17199 (
            .O(N__87679),
            .I(N__87657));
    Span4Mux_v I__17198 (
            .O(N__87676),
            .I(N__87654));
    LocalMux I__17197 (
            .O(N__87671),
            .I(N__87651));
    InMux I__17196 (
            .O(N__87670),
            .I(N__87648));
    InMux I__17195 (
            .O(N__87669),
            .I(N__87645));
    Span12Mux_h I__17194 (
            .O(N__87666),
            .I(N__87642));
    Span12Mux_v I__17193 (
            .O(N__87663),
            .I(N__87639));
    CascadeMux I__17192 (
            .O(N__87662),
            .I(N__87636));
    Span4Mux_h I__17191 (
            .O(N__87657),
            .I(N__87630));
    Span4Mux_v I__17190 (
            .O(N__87654),
            .I(N__87627));
    Span4Mux_v I__17189 (
            .O(N__87651),
            .I(N__87624));
    LocalMux I__17188 (
            .O(N__87648),
            .I(N__87619));
    LocalMux I__17187 (
            .O(N__87645),
            .I(N__87619));
    Span12Mux_v I__17186 (
            .O(N__87642),
            .I(N__87614));
    Span12Mux_h I__17185 (
            .O(N__87639),
            .I(N__87614));
    InMux I__17184 (
            .O(N__87636),
            .I(N__87605));
    InMux I__17183 (
            .O(N__87635),
            .I(N__87605));
    InMux I__17182 (
            .O(N__87634),
            .I(N__87605));
    InMux I__17181 (
            .O(N__87633),
            .I(N__87605));
    Span4Mux_h I__17180 (
            .O(N__87630),
            .I(N__87602));
    Span4Mux_h I__17179 (
            .O(N__87627),
            .I(N__87595));
    Span4Mux_h I__17178 (
            .O(N__87624),
            .I(N__87595));
    Span4Mux_v I__17177 (
            .O(N__87619),
            .I(N__87595));
    Odrv12 I__17176 (
            .O(N__87614),
            .I(rco_c_162));
    LocalMux I__17175 (
            .O(N__87605),
            .I(rco_c_162));
    Odrv4 I__17174 (
            .O(N__87602),
            .I(rco_c_162));
    Odrv4 I__17173 (
            .O(N__87595),
            .I(rco_c_162));
    IoInMux I__17172 (
            .O(N__87586),
            .I(N__87583));
    LocalMux I__17171 (
            .O(N__87583),
            .I(N__87580));
    Span4Mux_s3_h I__17170 (
            .O(N__87580),
            .I(N__87577));
    Odrv4 I__17169 (
            .O(N__87577),
            .I(rco_c_163));
    InMux I__17168 (
            .O(N__87574),
            .I(N__87571));
    LocalMux I__17167 (
            .O(N__87571),
            .I(shift_srl_168Z0Z_0));
    InMux I__17166 (
            .O(N__87568),
            .I(N__87565));
    LocalMux I__17165 (
            .O(N__87565),
            .I(shift_srl_168Z0Z_1));
    InMux I__17164 (
            .O(N__87562),
            .I(N__87559));
    LocalMux I__17163 (
            .O(N__87559),
            .I(shift_srl_168Z0Z_2));
    InMux I__17162 (
            .O(N__87556),
            .I(N__87553));
    LocalMux I__17161 (
            .O(N__87553),
            .I(shift_srl_168Z0Z_3));
    InMux I__17160 (
            .O(N__87550),
            .I(N__87547));
    LocalMux I__17159 (
            .O(N__87547),
            .I(shift_srl_168Z0Z_4));
    InMux I__17158 (
            .O(N__87544),
            .I(N__87541));
    LocalMux I__17157 (
            .O(N__87541),
            .I(shift_srl_168Z0Z_5));
    InMux I__17156 (
            .O(N__87538),
            .I(N__87535));
    LocalMux I__17155 (
            .O(N__87535),
            .I(shift_srl_164Z0Z_3));
    InMux I__17154 (
            .O(N__87532),
            .I(N__87529));
    LocalMux I__17153 (
            .O(N__87529),
            .I(shift_srl_164Z0Z_4));
    InMux I__17152 (
            .O(N__87526),
            .I(N__87523));
    LocalMux I__17151 (
            .O(N__87523),
            .I(shift_srl_164Z0Z_5));
    InMux I__17150 (
            .O(N__87520),
            .I(N__87517));
    LocalMux I__17149 (
            .O(N__87517),
            .I(shift_srl_164Z0Z_11));
    InMux I__17148 (
            .O(N__87514),
            .I(N__87511));
    LocalMux I__17147 (
            .O(N__87511),
            .I(shift_srl_164Z0Z_12));
    IoInMux I__17146 (
            .O(N__87508),
            .I(N__87505));
    LocalMux I__17145 (
            .O(N__87505),
            .I(N__87502));
    Span12Mux_s4_h I__17144 (
            .O(N__87502),
            .I(N__87499));
    Odrv12 I__17143 (
            .O(N__87499),
            .I(rco_c_171));
    InMux I__17142 (
            .O(N__87496),
            .I(N__87491));
    InMux I__17141 (
            .O(N__87495),
            .I(N__87488));
    InMux I__17140 (
            .O(N__87494),
            .I(N__87485));
    LocalMux I__17139 (
            .O(N__87491),
            .I(N__87480));
    LocalMux I__17138 (
            .O(N__87488),
            .I(N__87480));
    LocalMux I__17137 (
            .O(N__87485),
            .I(shift_srl_171Z0Z_15));
    Odrv12 I__17136 (
            .O(N__87480),
            .I(shift_srl_171Z0Z_15));
    InMux I__17135 (
            .O(N__87475),
            .I(N__87472));
    LocalMux I__17134 (
            .O(N__87472),
            .I(shift_srl_171_RNIVSP62Z0Z_15));
    CascadeMux I__17133 (
            .O(N__87469),
            .I(shift_srl_171_RNIVSP62Z0Z_15_cascade_));
    InMux I__17132 (
            .O(N__87466),
            .I(N__87463));
    LocalMux I__17131 (
            .O(N__87463),
            .I(N__87458));
    InMux I__17130 (
            .O(N__87462),
            .I(N__87453));
    InMux I__17129 (
            .O(N__87461),
            .I(N__87453));
    Span4Mux_h I__17128 (
            .O(N__87458),
            .I(N__87450));
    LocalMux I__17127 (
            .O(N__87453),
            .I(N__87447));
    Odrv4 I__17126 (
            .O(N__87450),
            .I(shift_srl_170_RNIRM2S1Z0Z_15));
    Odrv4 I__17125 (
            .O(N__87447),
            .I(shift_srl_170_RNIRM2S1Z0Z_15));
    IoInMux I__17124 (
            .O(N__87442),
            .I(N__87439));
    LocalMux I__17123 (
            .O(N__87439),
            .I(N__87436));
    Span4Mux_s3_h I__17122 (
            .O(N__87436),
            .I(N__87433));
    Odrv4 I__17121 (
            .O(N__87433),
            .I(rco_c_170));
    CascadeMux I__17120 (
            .O(N__87430),
            .I(N__87426));
    InMux I__17119 (
            .O(N__87429),
            .I(N__87420));
    InMux I__17118 (
            .O(N__87426),
            .I(N__87420));
    CascadeMux I__17117 (
            .O(N__87425),
            .I(N__87416));
    LocalMux I__17116 (
            .O(N__87420),
            .I(N__87411));
    InMux I__17115 (
            .O(N__87419),
            .I(N__87406));
    InMux I__17114 (
            .O(N__87416),
            .I(N__87406));
    InMux I__17113 (
            .O(N__87415),
            .I(N__87401));
    InMux I__17112 (
            .O(N__87414),
            .I(N__87401));
    Span4Mux_v I__17111 (
            .O(N__87411),
            .I(N__87398));
    LocalMux I__17110 (
            .O(N__87406),
            .I(N__87395));
    LocalMux I__17109 (
            .O(N__87401),
            .I(shift_srl_163_RNI3MR51Z0Z_15));
    Odrv4 I__17108 (
            .O(N__87398),
            .I(shift_srl_163_RNI3MR51Z0Z_15));
    Odrv4 I__17107 (
            .O(N__87395),
            .I(shift_srl_163_RNI3MR51Z0Z_15));
    IoInMux I__17106 (
            .O(N__87388),
            .I(N__87385));
    LocalMux I__17105 (
            .O(N__87385),
            .I(N__87382));
    IoSpan4Mux I__17104 (
            .O(N__87382),
            .I(N__87379));
    Span4Mux_s0_h I__17103 (
            .O(N__87379),
            .I(N__87376));
    Odrv4 I__17102 (
            .O(N__87376),
            .I(rco_c_167));
    InMux I__17101 (
            .O(N__87373),
            .I(N__87370));
    LocalMux I__17100 (
            .O(N__87370),
            .I(shift_srl_32Z0Z_8));
    IoInMux I__17099 (
            .O(N__87367),
            .I(N__87364));
    LocalMux I__17098 (
            .O(N__87364),
            .I(N__87360));
    InMux I__17097 (
            .O(N__87363),
            .I(N__87357));
    Span4Mux_s2_v I__17096 (
            .O(N__87360),
            .I(N__87354));
    LocalMux I__17095 (
            .O(N__87357),
            .I(N__87351));
    Span4Mux_v I__17094 (
            .O(N__87354),
            .I(N__87348));
    Span4Mux_h I__17093 (
            .O(N__87351),
            .I(N__87344));
    Span4Mux_v I__17092 (
            .O(N__87348),
            .I(N__87341));
    InMux I__17091 (
            .O(N__87347),
            .I(N__87338));
    Span4Mux_h I__17090 (
            .O(N__87344),
            .I(N__87335));
    Span4Mux_v I__17089 (
            .O(N__87341),
            .I(N__87330));
    LocalMux I__17088 (
            .O(N__87338),
            .I(N__87330));
    Odrv4 I__17087 (
            .O(N__87335),
            .I(rco_c_31));
    Odrv4 I__17086 (
            .O(N__87330),
            .I(rco_c_31));
    InMux I__17085 (
            .O(N__87325),
            .I(N__87320));
    InMux I__17084 (
            .O(N__87324),
            .I(N__87313));
    InMux I__17083 (
            .O(N__87323),
            .I(N__87313));
    LocalMux I__17082 (
            .O(N__87320),
            .I(N__87310));
    InMux I__17081 (
            .O(N__87319),
            .I(N__87305));
    InMux I__17080 (
            .O(N__87318),
            .I(N__87305));
    LocalMux I__17079 (
            .O(N__87313),
            .I(N__87302));
    Span4Mux_h I__17078 (
            .O(N__87310),
            .I(N__87299));
    LocalMux I__17077 (
            .O(N__87305),
            .I(N__87295));
    Span4Mux_v I__17076 (
            .O(N__87302),
            .I(N__87292));
    Span4Mux_h I__17075 (
            .O(N__87299),
            .I(N__87289));
    InMux I__17074 (
            .O(N__87298),
            .I(N__87286));
    Span4Mux_v I__17073 (
            .O(N__87295),
            .I(N__87283));
    Sp12to4 I__17072 (
            .O(N__87292),
            .I(N__87280));
    Span4Mux_h I__17071 (
            .O(N__87289),
            .I(N__87277));
    LocalMux I__17070 (
            .O(N__87286),
            .I(shift_srl_32Z0Z_15));
    Odrv4 I__17069 (
            .O(N__87283),
            .I(shift_srl_32Z0Z_15));
    Odrv12 I__17068 (
            .O(N__87280),
            .I(shift_srl_32Z0Z_15));
    Odrv4 I__17067 (
            .O(N__87277),
            .I(shift_srl_32Z0Z_15));
    InMux I__17066 (
            .O(N__87268),
            .I(N__87265));
    LocalMux I__17065 (
            .O(N__87265),
            .I(shift_srl_32Z0Z_0));
    InMux I__17064 (
            .O(N__87262),
            .I(N__87259));
    LocalMux I__17063 (
            .O(N__87259),
            .I(shift_srl_32Z0Z_1));
    InMux I__17062 (
            .O(N__87256),
            .I(N__87252));
    InMux I__17061 (
            .O(N__87255),
            .I(N__87249));
    LocalMux I__17060 (
            .O(N__87252),
            .I(N__87246));
    LocalMux I__17059 (
            .O(N__87249),
            .I(N__87243));
    Span4Mux_h I__17058 (
            .O(N__87246),
            .I(N__87239));
    Span4Mux_h I__17057 (
            .O(N__87243),
            .I(N__87236));
    InMux I__17056 (
            .O(N__87242),
            .I(N__87233));
    Odrv4 I__17055 (
            .O(N__87239),
            .I(shift_srl_164Z0Z_15));
    Odrv4 I__17054 (
            .O(N__87236),
            .I(shift_srl_164Z0Z_15));
    LocalMux I__17053 (
            .O(N__87233),
            .I(shift_srl_164Z0Z_15));
    InMux I__17052 (
            .O(N__87226),
            .I(N__87223));
    LocalMux I__17051 (
            .O(N__87223),
            .I(shift_srl_164Z0Z_0));
    InMux I__17050 (
            .O(N__87220),
            .I(N__87217));
    LocalMux I__17049 (
            .O(N__87217),
            .I(shift_srl_164Z0Z_1));
    InMux I__17048 (
            .O(N__87214),
            .I(N__87211));
    LocalMux I__17047 (
            .O(N__87211),
            .I(shift_srl_164Z0Z_2));
    InMux I__17046 (
            .O(N__87208),
            .I(N__87205));
    LocalMux I__17045 (
            .O(N__87205),
            .I(shift_srl_54Z0Z_8));
    InMux I__17044 (
            .O(N__87202),
            .I(N__87199));
    LocalMux I__17043 (
            .O(N__87199),
            .I(N__87196));
    Span4Mux_v I__17042 (
            .O(N__87196),
            .I(N__87193));
    Span4Mux_h I__17041 (
            .O(N__87193),
            .I(N__87190));
    Odrv4 I__17040 (
            .O(N__87190),
            .I(shift_srl_54Z0Z_9));
    CEMux I__17039 (
            .O(N__87187),
            .I(N__87183));
    CEMux I__17038 (
            .O(N__87186),
            .I(N__87180));
    LocalMux I__17037 (
            .O(N__87183),
            .I(N__87177));
    LocalMux I__17036 (
            .O(N__87180),
            .I(N__87174));
    Span4Mux_v I__17035 (
            .O(N__87177),
            .I(N__87171));
    Span12Mux_v I__17034 (
            .O(N__87174),
            .I(N__87167));
    Span4Mux_h I__17033 (
            .O(N__87171),
            .I(N__87164));
    CEMux I__17032 (
            .O(N__87170),
            .I(N__87161));
    Odrv12 I__17031 (
            .O(N__87167),
            .I(clk_en_54));
    Odrv4 I__17030 (
            .O(N__87164),
            .I(clk_en_54));
    LocalMux I__17029 (
            .O(N__87161),
            .I(clk_en_54));
    InMux I__17028 (
            .O(N__87154),
            .I(N__87151));
    LocalMux I__17027 (
            .O(N__87151),
            .I(N__87148));
    Odrv4 I__17026 (
            .O(N__87148),
            .I(shift_srl_34Z0Z_7));
    InMux I__17025 (
            .O(N__87145),
            .I(N__87142));
    LocalMux I__17024 (
            .O(N__87142),
            .I(N__87139));
    Odrv12 I__17023 (
            .O(N__87139),
            .I(shift_srl_34Z0Z_8));
    CEMux I__17022 (
            .O(N__87136),
            .I(N__87132));
    CEMux I__17021 (
            .O(N__87135),
            .I(N__87128));
    LocalMux I__17020 (
            .O(N__87132),
            .I(N__87125));
    CEMux I__17019 (
            .O(N__87131),
            .I(N__87122));
    LocalMux I__17018 (
            .O(N__87128),
            .I(N__87117));
    Span4Mux_h I__17017 (
            .O(N__87125),
            .I(N__87112));
    LocalMux I__17016 (
            .O(N__87122),
            .I(N__87112));
    CEMux I__17015 (
            .O(N__87121),
            .I(N__87109));
    CEMux I__17014 (
            .O(N__87120),
            .I(N__87106));
    Span4Mux_v I__17013 (
            .O(N__87117),
            .I(N__87103));
    Span4Mux_h I__17012 (
            .O(N__87112),
            .I(N__87100));
    LocalMux I__17011 (
            .O(N__87109),
            .I(N__87097));
    LocalMux I__17010 (
            .O(N__87106),
            .I(N__87094));
    Odrv4 I__17009 (
            .O(N__87103),
            .I(clk_en_34));
    Odrv4 I__17008 (
            .O(N__87100),
            .I(clk_en_34));
    Odrv12 I__17007 (
            .O(N__87097),
            .I(clk_en_34));
    Odrv4 I__17006 (
            .O(N__87094),
            .I(clk_en_34));
    InMux I__17005 (
            .O(N__87085),
            .I(N__87082));
    LocalMux I__17004 (
            .O(N__87082),
            .I(shift_srl_32Z0Z_10));
    InMux I__17003 (
            .O(N__87079),
            .I(N__87076));
    LocalMux I__17002 (
            .O(N__87076),
            .I(shift_srl_32Z0Z_11));
    InMux I__17001 (
            .O(N__87073),
            .I(N__87070));
    LocalMux I__17000 (
            .O(N__87070),
            .I(shift_srl_32Z0Z_12));
    InMux I__16999 (
            .O(N__87067),
            .I(N__87064));
    LocalMux I__16998 (
            .O(N__87064),
            .I(shift_srl_32Z0Z_13));
    InMux I__16997 (
            .O(N__87061),
            .I(N__87058));
    LocalMux I__16996 (
            .O(N__87058),
            .I(shift_srl_32Z0Z_14));
    InMux I__16995 (
            .O(N__87055),
            .I(N__87052));
    LocalMux I__16994 (
            .O(N__87052),
            .I(shift_srl_32Z0Z_9));
    InMux I__16993 (
            .O(N__87049),
            .I(N__87046));
    LocalMux I__16992 (
            .O(N__87046),
            .I(shift_srl_72Z0Z_12));
    InMux I__16991 (
            .O(N__87043),
            .I(N__87040));
    LocalMux I__16990 (
            .O(N__87040),
            .I(shift_srl_72Z0Z_13));
    InMux I__16989 (
            .O(N__87037),
            .I(N__87034));
    LocalMux I__16988 (
            .O(N__87034),
            .I(shift_srl_72Z0Z_14));
    InMux I__16987 (
            .O(N__87031),
            .I(N__87028));
    LocalMux I__16986 (
            .O(N__87028),
            .I(shift_srl_72Z0Z_9));
    InMux I__16985 (
            .O(N__87025),
            .I(N__87022));
    LocalMux I__16984 (
            .O(N__87022),
            .I(N__87019));
    Odrv4 I__16983 (
            .O(N__87019),
            .I(shift_srl_72Z0Z_7));
    InMux I__16982 (
            .O(N__87016),
            .I(N__87013));
    LocalMux I__16981 (
            .O(N__87013),
            .I(shift_srl_72Z0Z_8));
    CEMux I__16980 (
            .O(N__87010),
            .I(N__87007));
    LocalMux I__16979 (
            .O(N__87007),
            .I(N__87004));
    Span4Mux_v I__16978 (
            .O(N__87004),
            .I(N__86999));
    CEMux I__16977 (
            .O(N__87003),
            .I(N__86996));
    CEMux I__16976 (
            .O(N__87002),
            .I(N__86993));
    Odrv4 I__16975 (
            .O(N__86999),
            .I(clk_en_72));
    LocalMux I__16974 (
            .O(N__86996),
            .I(clk_en_72));
    LocalMux I__16973 (
            .O(N__86993),
            .I(clk_en_72));
    InMux I__16972 (
            .O(N__86986),
            .I(N__86983));
    LocalMux I__16971 (
            .O(N__86983),
            .I(N__86980));
    Odrv4 I__16970 (
            .O(N__86980),
            .I(shift_srl_34Z0Z_6));
    InMux I__16969 (
            .O(N__86977),
            .I(N__86974));
    LocalMux I__16968 (
            .O(N__86974),
            .I(N__86971));
    Span4Mux_h I__16967 (
            .O(N__86971),
            .I(N__86968));
    Span4Mux_h I__16966 (
            .O(N__86968),
            .I(N__86965));
    Odrv4 I__16965 (
            .O(N__86965),
            .I(shift_srl_54Z0Z_4));
    InMux I__16964 (
            .O(N__86962),
            .I(N__86959));
    LocalMux I__16963 (
            .O(N__86959),
            .I(shift_srl_54Z0Z_5));
    InMux I__16962 (
            .O(N__86956),
            .I(N__86953));
    LocalMux I__16961 (
            .O(N__86953),
            .I(shift_srl_54Z0Z_6));
    InMux I__16960 (
            .O(N__86950),
            .I(N__86947));
    LocalMux I__16959 (
            .O(N__86947),
            .I(shift_srl_54Z0Z_7));
    InMux I__16958 (
            .O(N__86944),
            .I(N__86941));
    LocalMux I__16957 (
            .O(N__86941),
            .I(shift_srl_72Z0Z_6));
    CEMux I__16956 (
            .O(N__86938),
            .I(N__86935));
    LocalMux I__16955 (
            .O(N__86935),
            .I(N__86931));
    CEMux I__16954 (
            .O(N__86934),
            .I(N__86928));
    Span4Mux_v I__16953 (
            .O(N__86931),
            .I(N__86920));
    LocalMux I__16952 (
            .O(N__86928),
            .I(N__86920));
    CEMux I__16951 (
            .O(N__86927),
            .I(N__86917));
    InMux I__16950 (
            .O(N__86926),
            .I(N__86914));
    InMux I__16949 (
            .O(N__86925),
            .I(N__86911));
    Span4Mux_h I__16948 (
            .O(N__86920),
            .I(N__86908));
    LocalMux I__16947 (
            .O(N__86917),
            .I(N__86901));
    LocalMux I__16946 (
            .O(N__86914),
            .I(N__86901));
    LocalMux I__16945 (
            .O(N__86911),
            .I(N__86901));
    Odrv4 I__16944 (
            .O(N__86908),
            .I(clk_en_67));
    Odrv12 I__16943 (
            .O(N__86901),
            .I(clk_en_67));
    InMux I__16942 (
            .O(N__86896),
            .I(N__86893));
    LocalMux I__16941 (
            .O(N__86893),
            .I(N__86888));
    InMux I__16940 (
            .O(N__86892),
            .I(N__86885));
    InMux I__16939 (
            .O(N__86891),
            .I(N__86882));
    Span4Mux_v I__16938 (
            .O(N__86888),
            .I(N__86879));
    LocalMux I__16937 (
            .O(N__86885),
            .I(N__86876));
    LocalMux I__16936 (
            .O(N__86882),
            .I(shift_srl_68Z0Z_15));
    Odrv4 I__16935 (
            .O(N__86879),
            .I(shift_srl_68Z0Z_15));
    Odrv4 I__16934 (
            .O(N__86876),
            .I(shift_srl_68Z0Z_15));
    CascadeMux I__16933 (
            .O(N__86869),
            .I(N__86865));
    CascadeMux I__16932 (
            .O(N__86868),
            .I(N__86862));
    InMux I__16931 (
            .O(N__86865),
            .I(N__86857));
    InMux I__16930 (
            .O(N__86862),
            .I(N__86853));
    InMux I__16929 (
            .O(N__86861),
            .I(N__86848));
    InMux I__16928 (
            .O(N__86860),
            .I(N__86848));
    LocalMux I__16927 (
            .O(N__86857),
            .I(N__86845));
    InMux I__16926 (
            .O(N__86856),
            .I(N__86842));
    LocalMux I__16925 (
            .O(N__86853),
            .I(N__86839));
    LocalMux I__16924 (
            .O(N__86848),
            .I(N__86834));
    Span4Mux_h I__16923 (
            .O(N__86845),
            .I(N__86834));
    LocalMux I__16922 (
            .O(N__86842),
            .I(N__86829));
    Span4Mux_v I__16921 (
            .O(N__86839),
            .I(N__86829));
    Odrv4 I__16920 (
            .O(N__86834),
            .I(shift_srl_67Z0Z_15));
    Odrv4 I__16919 (
            .O(N__86829),
            .I(shift_srl_67Z0Z_15));
    CascadeMux I__16918 (
            .O(N__86824),
            .I(shift_srl_74_RNIS4SRZ0Z_15_cascade_));
    InMux I__16917 (
            .O(N__86821),
            .I(N__86818));
    LocalMux I__16916 (
            .O(N__86818),
            .I(N__86812));
    InMux I__16915 (
            .O(N__86817),
            .I(N__86806));
    InMux I__16914 (
            .O(N__86816),
            .I(N__86801));
    InMux I__16913 (
            .O(N__86815),
            .I(N__86797));
    Span4Mux_h I__16912 (
            .O(N__86812),
            .I(N__86794));
    InMux I__16911 (
            .O(N__86811),
            .I(N__86791));
    InMux I__16910 (
            .O(N__86810),
            .I(N__86786));
    InMux I__16909 (
            .O(N__86809),
            .I(N__86786));
    LocalMux I__16908 (
            .O(N__86806),
            .I(N__86783));
    InMux I__16907 (
            .O(N__86805),
            .I(N__86778));
    InMux I__16906 (
            .O(N__86804),
            .I(N__86778));
    LocalMux I__16905 (
            .O(N__86801),
            .I(N__86775));
    InMux I__16904 (
            .O(N__86800),
            .I(N__86772));
    LocalMux I__16903 (
            .O(N__86797),
            .I(N__86769));
    Span4Mux_v I__16902 (
            .O(N__86794),
            .I(N__86766));
    LocalMux I__16901 (
            .O(N__86791),
            .I(N__86763));
    LocalMux I__16900 (
            .O(N__86786),
            .I(N__86760));
    Span4Mux_v I__16899 (
            .O(N__86783),
            .I(N__86755));
    LocalMux I__16898 (
            .O(N__86778),
            .I(N__86755));
    Span12Mux_v I__16897 (
            .O(N__86775),
            .I(N__86751));
    LocalMux I__16896 (
            .O(N__86772),
            .I(N__86742));
    Span4Mux_v I__16895 (
            .O(N__86769),
            .I(N__86742));
    Span4Mux_h I__16894 (
            .O(N__86766),
            .I(N__86742));
    Span4Mux_v I__16893 (
            .O(N__86763),
            .I(N__86742));
    Span4Mux_v I__16892 (
            .O(N__86760),
            .I(N__86737));
    Span4Mux_h I__16891 (
            .O(N__86755),
            .I(N__86737));
    InMux I__16890 (
            .O(N__86754),
            .I(N__86734));
    Span12Mux_h I__16889 (
            .O(N__86751),
            .I(N__86731));
    Span4Mux_h I__16888 (
            .O(N__86742),
            .I(N__86728));
    Odrv4 I__16887 (
            .O(N__86737),
            .I(rco_int_0_a3_0_a2_0_74));
    LocalMux I__16886 (
            .O(N__86734),
            .I(rco_int_0_a3_0_a2_0_74));
    Odrv12 I__16885 (
            .O(N__86731),
            .I(rco_int_0_a3_0_a2_0_74));
    Odrv4 I__16884 (
            .O(N__86728),
            .I(rco_int_0_a3_0_a2_0_74));
    InMux I__16883 (
            .O(N__86719),
            .I(N__86715));
    InMux I__16882 (
            .O(N__86718),
            .I(N__86711));
    LocalMux I__16881 (
            .O(N__86715),
            .I(N__86708));
    InMux I__16880 (
            .O(N__86714),
            .I(N__86705));
    LocalMux I__16879 (
            .O(N__86711),
            .I(shift_srl_71Z0Z_15));
    Odrv4 I__16878 (
            .O(N__86708),
            .I(shift_srl_71Z0Z_15));
    LocalMux I__16877 (
            .O(N__86705),
            .I(shift_srl_71Z0Z_15));
    InMux I__16876 (
            .O(N__86698),
            .I(N__86689));
    InMux I__16875 (
            .O(N__86697),
            .I(N__86689));
    InMux I__16874 (
            .O(N__86696),
            .I(N__86686));
    InMux I__16873 (
            .O(N__86695),
            .I(N__86683));
    InMux I__16872 (
            .O(N__86694),
            .I(N__86680));
    LocalMux I__16871 (
            .O(N__86689),
            .I(N__86677));
    LocalMux I__16870 (
            .O(N__86686),
            .I(N__86672));
    LocalMux I__16869 (
            .O(N__86683),
            .I(N__86672));
    LocalMux I__16868 (
            .O(N__86680),
            .I(shift_srl_70Z0Z_15));
    Odrv12 I__16867 (
            .O(N__86677),
            .I(shift_srl_70Z0Z_15));
    Odrv4 I__16866 (
            .O(N__86672),
            .I(shift_srl_70Z0Z_15));
    InMux I__16865 (
            .O(N__86665),
            .I(N__86661));
    InMux I__16864 (
            .O(N__86664),
            .I(N__86657));
    LocalMux I__16863 (
            .O(N__86661),
            .I(N__86651));
    InMux I__16862 (
            .O(N__86660),
            .I(N__86648));
    LocalMux I__16861 (
            .O(N__86657),
            .I(N__86645));
    InMux I__16860 (
            .O(N__86656),
            .I(N__86640));
    InMux I__16859 (
            .O(N__86655),
            .I(N__86640));
    InMux I__16858 (
            .O(N__86654),
            .I(N__86637));
    Odrv4 I__16857 (
            .O(N__86651),
            .I(shift_srl_69Z0Z_15));
    LocalMux I__16856 (
            .O(N__86648),
            .I(shift_srl_69Z0Z_15));
    Odrv4 I__16855 (
            .O(N__86645),
            .I(shift_srl_69Z0Z_15));
    LocalMux I__16854 (
            .O(N__86640),
            .I(shift_srl_69Z0Z_15));
    LocalMux I__16853 (
            .O(N__86637),
            .I(shift_srl_69Z0Z_15));
    InMux I__16852 (
            .O(N__86626),
            .I(N__86623));
    LocalMux I__16851 (
            .O(N__86623),
            .I(rco_int_0_a3_0_a2_0_1_74));
    InMux I__16850 (
            .O(N__86620),
            .I(N__86617));
    LocalMux I__16849 (
            .O(N__86617),
            .I(shift_srl_72Z0Z_10));
    InMux I__16848 (
            .O(N__86614),
            .I(N__86611));
    LocalMux I__16847 (
            .O(N__86611),
            .I(shift_srl_72Z0Z_11));
    InMux I__16846 (
            .O(N__86608),
            .I(N__86605));
    LocalMux I__16845 (
            .O(N__86605),
            .I(shift_srl_68Z0Z_9));
    InMux I__16844 (
            .O(N__86602),
            .I(N__86599));
    LocalMux I__16843 (
            .O(N__86599),
            .I(shift_srl_68Z0Z_7));
    InMux I__16842 (
            .O(N__86596),
            .I(N__86593));
    LocalMux I__16841 (
            .O(N__86593),
            .I(shift_srl_68Z0Z_8));
    CEMux I__16840 (
            .O(N__86590),
            .I(N__86586));
    CEMux I__16839 (
            .O(N__86589),
            .I(N__86583));
    LocalMux I__16838 (
            .O(N__86586),
            .I(N__86580));
    LocalMux I__16837 (
            .O(N__86583),
            .I(N__86577));
    Odrv4 I__16836 (
            .O(N__86580),
            .I(clk_en_68));
    Odrv4 I__16835 (
            .O(N__86577),
            .I(clk_en_68));
    InMux I__16834 (
            .O(N__86572),
            .I(N__86569));
    LocalMux I__16833 (
            .O(N__86569),
            .I(shift_srl_72Z0Z_0));
    InMux I__16832 (
            .O(N__86566),
            .I(N__86563));
    LocalMux I__16831 (
            .O(N__86563),
            .I(shift_srl_72Z0Z_1));
    InMux I__16830 (
            .O(N__86560),
            .I(N__86557));
    LocalMux I__16829 (
            .O(N__86557),
            .I(shift_srl_72Z0Z_2));
    InMux I__16828 (
            .O(N__86554),
            .I(N__86551));
    LocalMux I__16827 (
            .O(N__86551),
            .I(shift_srl_72Z0Z_3));
    InMux I__16826 (
            .O(N__86548),
            .I(N__86545));
    LocalMux I__16825 (
            .O(N__86545),
            .I(shift_srl_72Z0Z_4));
    InMux I__16824 (
            .O(N__86542),
            .I(N__86539));
    LocalMux I__16823 (
            .O(N__86539),
            .I(shift_srl_72Z0Z_5));
    InMux I__16822 (
            .O(N__86536),
            .I(N__86533));
    LocalMux I__16821 (
            .O(N__86533),
            .I(shift_srl_77Z0Z_14));
    InMux I__16820 (
            .O(N__86530),
            .I(N__86527));
    LocalMux I__16819 (
            .O(N__86527),
            .I(shift_srl_77Z0Z_9));
    InMux I__16818 (
            .O(N__86524),
            .I(N__86521));
    LocalMux I__16817 (
            .O(N__86521),
            .I(shift_srl_77Z0Z_8));
    InMux I__16816 (
            .O(N__86518),
            .I(N__86515));
    LocalMux I__16815 (
            .O(N__86515),
            .I(shift_srl_68Z0Z_10));
    InMux I__16814 (
            .O(N__86512),
            .I(N__86509));
    LocalMux I__16813 (
            .O(N__86509),
            .I(shift_srl_68Z0Z_11));
    InMux I__16812 (
            .O(N__86506),
            .I(N__86503));
    LocalMux I__16811 (
            .O(N__86503),
            .I(shift_srl_68Z0Z_12));
    InMux I__16810 (
            .O(N__86500),
            .I(N__86497));
    LocalMux I__16809 (
            .O(N__86497),
            .I(shift_srl_68Z0Z_13));
    InMux I__16808 (
            .O(N__86494),
            .I(N__86491));
    LocalMux I__16807 (
            .O(N__86491),
            .I(shift_srl_68Z0Z_14));
    InMux I__16806 (
            .O(N__86488),
            .I(N__86485));
    LocalMux I__16805 (
            .O(N__86485),
            .I(shift_srl_79Z0Z_13));
    InMux I__16804 (
            .O(N__86482),
            .I(N__86479));
    LocalMux I__16803 (
            .O(N__86479),
            .I(shift_srl_79Z0Z_14));
    InMux I__16802 (
            .O(N__86476),
            .I(N__86471));
    InMux I__16801 (
            .O(N__86475),
            .I(N__86465));
    InMux I__16800 (
            .O(N__86474),
            .I(N__86465));
    LocalMux I__16799 (
            .O(N__86471),
            .I(N__86462));
    InMux I__16798 (
            .O(N__86470),
            .I(N__86459));
    LocalMux I__16797 (
            .O(N__86465),
            .I(shift_srl_79Z0Z_15));
    Odrv12 I__16796 (
            .O(N__86462),
            .I(shift_srl_79Z0Z_15));
    LocalMux I__16795 (
            .O(N__86459),
            .I(shift_srl_79Z0Z_15));
    InMux I__16794 (
            .O(N__86452),
            .I(N__86449));
    LocalMux I__16793 (
            .O(N__86449),
            .I(shift_srl_79Z0Z_9));
    InMux I__16792 (
            .O(N__86446),
            .I(N__86443));
    LocalMux I__16791 (
            .O(N__86443),
            .I(N__86440));
    Odrv4 I__16790 (
            .O(N__86440),
            .I(shift_srl_79Z0Z_7));
    InMux I__16789 (
            .O(N__86437),
            .I(N__86434));
    LocalMux I__16788 (
            .O(N__86434),
            .I(shift_srl_79Z0Z_8));
    CEMux I__16787 (
            .O(N__86431),
            .I(N__86428));
    LocalMux I__16786 (
            .O(N__86428),
            .I(N__86423));
    CEMux I__16785 (
            .O(N__86427),
            .I(N__86420));
    CEMux I__16784 (
            .O(N__86426),
            .I(N__86417));
    Span4Mux_v I__16783 (
            .O(N__86423),
            .I(N__86414));
    LocalMux I__16782 (
            .O(N__86420),
            .I(N__86411));
    LocalMux I__16781 (
            .O(N__86417),
            .I(N__86408));
    Span4Mux_s3_h I__16780 (
            .O(N__86414),
            .I(N__86403));
    Span4Mux_v I__16779 (
            .O(N__86411),
            .I(N__86403));
    Span4Mux_h I__16778 (
            .O(N__86408),
            .I(N__86400));
    Odrv4 I__16777 (
            .O(N__86403),
            .I(clk_en_79));
    Odrv4 I__16776 (
            .O(N__86400),
            .I(clk_en_79));
    InMux I__16775 (
            .O(N__86395),
            .I(N__86392));
    LocalMux I__16774 (
            .O(N__86392),
            .I(shift_srl_77Z0Z_10));
    InMux I__16773 (
            .O(N__86389),
            .I(N__86386));
    LocalMux I__16772 (
            .O(N__86386),
            .I(shift_srl_77Z0Z_11));
    InMux I__16771 (
            .O(N__86383),
            .I(N__86380));
    LocalMux I__16770 (
            .O(N__86380),
            .I(shift_srl_77Z0Z_12));
    InMux I__16769 (
            .O(N__86377),
            .I(N__86374));
    LocalMux I__16768 (
            .O(N__86374),
            .I(shift_srl_77Z0Z_13));
    InMux I__16767 (
            .O(N__86371),
            .I(N__86368));
    LocalMux I__16766 (
            .O(N__86368),
            .I(shift_srl_81Z0Z_12));
    InMux I__16765 (
            .O(N__86365),
            .I(N__86362));
    LocalMux I__16764 (
            .O(N__86362),
            .I(shift_srl_81Z0Z_13));
    InMux I__16763 (
            .O(N__86359),
            .I(N__86356));
    LocalMux I__16762 (
            .O(N__86356),
            .I(shift_srl_81Z0Z_14));
    CascadeMux I__16761 (
            .O(N__86353),
            .I(N__86350));
    InMux I__16760 (
            .O(N__86350),
            .I(N__86344));
    InMux I__16759 (
            .O(N__86349),
            .I(N__86339));
    InMux I__16758 (
            .O(N__86348),
            .I(N__86339));
    InMux I__16757 (
            .O(N__86347),
            .I(N__86335));
    LocalMux I__16756 (
            .O(N__86344),
            .I(N__86331));
    LocalMux I__16755 (
            .O(N__86339),
            .I(N__86328));
    CascadeMux I__16754 (
            .O(N__86338),
            .I(N__86325));
    LocalMux I__16753 (
            .O(N__86335),
            .I(N__86322));
    InMux I__16752 (
            .O(N__86334),
            .I(N__86319));
    Span4Mux_v I__16751 (
            .O(N__86331),
            .I(N__86314));
    Span4Mux_v I__16750 (
            .O(N__86328),
            .I(N__86314));
    InMux I__16749 (
            .O(N__86325),
            .I(N__86311));
    Odrv4 I__16748 (
            .O(N__86322),
            .I(shift_srl_81Z0Z_15));
    LocalMux I__16747 (
            .O(N__86319),
            .I(shift_srl_81Z0Z_15));
    Odrv4 I__16746 (
            .O(N__86314),
            .I(shift_srl_81Z0Z_15));
    LocalMux I__16745 (
            .O(N__86311),
            .I(shift_srl_81Z0Z_15));
    InMux I__16744 (
            .O(N__86302),
            .I(N__86299));
    LocalMux I__16743 (
            .O(N__86299),
            .I(shift_srl_81Z0Z_9));
    InMux I__16742 (
            .O(N__86296),
            .I(N__86293));
    LocalMux I__16741 (
            .O(N__86293),
            .I(shift_srl_81Z0Z_7));
    InMux I__16740 (
            .O(N__86290),
            .I(N__86287));
    LocalMux I__16739 (
            .O(N__86287),
            .I(shift_srl_81Z0Z_8));
    CEMux I__16738 (
            .O(N__86284),
            .I(N__86280));
    CEMux I__16737 (
            .O(N__86283),
            .I(N__86277));
    LocalMux I__16736 (
            .O(N__86280),
            .I(N_786));
    LocalMux I__16735 (
            .O(N__86277),
            .I(N_786));
    InMux I__16734 (
            .O(N__86272),
            .I(N__86269));
    LocalMux I__16733 (
            .O(N__86269),
            .I(shift_srl_79Z0Z_10));
    InMux I__16732 (
            .O(N__86266),
            .I(N__86263));
    LocalMux I__16731 (
            .O(N__86263),
            .I(shift_srl_79Z0Z_11));
    InMux I__16730 (
            .O(N__86260),
            .I(N__86257));
    LocalMux I__16729 (
            .O(N__86257),
            .I(shift_srl_79Z0Z_12));
    InMux I__16728 (
            .O(N__86254),
            .I(N__86251));
    LocalMux I__16727 (
            .O(N__86251),
            .I(shift_srl_79Z0Z_1));
    InMux I__16726 (
            .O(N__86248),
            .I(N__86245));
    LocalMux I__16725 (
            .O(N__86245),
            .I(shift_srl_79Z0Z_2));
    InMux I__16724 (
            .O(N__86242),
            .I(N__86239));
    LocalMux I__16723 (
            .O(N__86239),
            .I(shift_srl_79Z0Z_3));
    InMux I__16722 (
            .O(N__86236),
            .I(N__86233));
    LocalMux I__16721 (
            .O(N__86233),
            .I(shift_srl_79Z0Z_4));
    InMux I__16720 (
            .O(N__86230),
            .I(N__86227));
    LocalMux I__16719 (
            .O(N__86227),
            .I(shift_srl_79Z0Z_5));
    InMux I__16718 (
            .O(N__86224),
            .I(N__86221));
    LocalMux I__16717 (
            .O(N__86221),
            .I(shift_srl_79Z0Z_6));
    InMux I__16716 (
            .O(N__86218),
            .I(N__86215));
    LocalMux I__16715 (
            .O(N__86215),
            .I(shift_srl_81Z0Z_10));
    InMux I__16714 (
            .O(N__86212),
            .I(N__86209));
    LocalMux I__16713 (
            .O(N__86209),
            .I(shift_srl_81Z0Z_11));
    InMux I__16712 (
            .O(N__86206),
            .I(N__86203));
    LocalMux I__16711 (
            .O(N__86203),
            .I(shift_srl_191Z0Z_2));
    InMux I__16710 (
            .O(N__86200),
            .I(N__86197));
    LocalMux I__16709 (
            .O(N__86197),
            .I(shift_srl_191Z0Z_3));
    InMux I__16708 (
            .O(N__86194),
            .I(N__86191));
    LocalMux I__16707 (
            .O(N__86191),
            .I(shift_srl_191Z0Z_4));
    InMux I__16706 (
            .O(N__86188),
            .I(N__86185));
    LocalMux I__16705 (
            .O(N__86185),
            .I(shift_srl_191Z0Z_5));
    InMux I__16704 (
            .O(N__86182),
            .I(N__86179));
    LocalMux I__16703 (
            .O(N__86179),
            .I(shift_srl_191Z0Z_6));
    InMux I__16702 (
            .O(N__86176),
            .I(N__86173));
    LocalMux I__16701 (
            .O(N__86173),
            .I(shift_srl_191Z0Z_7));
    CascadeMux I__16700 (
            .O(N__86170),
            .I(N__86166));
    CascadeMux I__16699 (
            .O(N__86169),
            .I(N__86163));
    InMux I__16698 (
            .O(N__86166),
            .I(N__86159));
    InMux I__16697 (
            .O(N__86163),
            .I(N__86156));
    InMux I__16696 (
            .O(N__86162),
            .I(N__86153));
    LocalMux I__16695 (
            .O(N__86159),
            .I(N__86150));
    LocalMux I__16694 (
            .O(N__86156),
            .I(N__86147));
    LocalMux I__16693 (
            .O(N__86153),
            .I(shift_srl_187Z0Z_15));
    Odrv12 I__16692 (
            .O(N__86150),
            .I(shift_srl_187Z0Z_15));
    Odrv4 I__16691 (
            .O(N__86147),
            .I(shift_srl_187Z0Z_15));
    InMux I__16690 (
            .O(N__86140),
            .I(N__86137));
    LocalMux I__16689 (
            .O(N__86137),
            .I(N__86132));
    InMux I__16688 (
            .O(N__86136),
            .I(N__86129));
    InMux I__16687 (
            .O(N__86135),
            .I(N__86126));
    Span4Mux_h I__16686 (
            .O(N__86132),
            .I(N__86123));
    LocalMux I__16685 (
            .O(N__86129),
            .I(N__86120));
    LocalMux I__16684 (
            .O(N__86126),
            .I(N__86117));
    Span4Mux_h I__16683 (
            .O(N__86123),
            .I(N__86112));
    Span4Mux_h I__16682 (
            .O(N__86120),
            .I(N__86112));
    Odrv4 I__16681 (
            .O(N__86117),
            .I(shift_srl_189Z0Z_15));
    Odrv4 I__16680 (
            .O(N__86112),
            .I(shift_srl_189Z0Z_15));
    CascadeMux I__16679 (
            .O(N__86107),
            .I(clk_en_0_a3_0_a2_0_sx_190_cascade_));
    InMux I__16678 (
            .O(N__86104),
            .I(N__86100));
    InMux I__16677 (
            .O(N__86103),
            .I(N__86097));
    LocalMux I__16676 (
            .O(N__86100),
            .I(N__86091));
    LocalMux I__16675 (
            .O(N__86097),
            .I(N__86088));
    InMux I__16674 (
            .O(N__86096),
            .I(N__86085));
    InMux I__16673 (
            .O(N__86095),
            .I(N__86080));
    InMux I__16672 (
            .O(N__86094),
            .I(N__86080));
    Span4Mux_h I__16671 (
            .O(N__86091),
            .I(N__86077));
    Span4Mux_h I__16670 (
            .O(N__86088),
            .I(N__86074));
    LocalMux I__16669 (
            .O(N__86085),
            .I(shift_srl_188Z0Z_15));
    LocalMux I__16668 (
            .O(N__86080),
            .I(shift_srl_188Z0Z_15));
    Odrv4 I__16667 (
            .O(N__86077),
            .I(shift_srl_188Z0Z_15));
    Odrv4 I__16666 (
            .O(N__86074),
            .I(shift_srl_188Z0Z_15));
    CascadeMux I__16665 (
            .O(N__86065),
            .I(N_4175_cascade_));
    CEMux I__16664 (
            .O(N__86062),
            .I(N__86058));
    CEMux I__16663 (
            .O(N__86061),
            .I(N__86055));
    LocalMux I__16662 (
            .O(N__86058),
            .I(clk_en_191));
    LocalMux I__16661 (
            .O(N__86055),
            .I(clk_en_191));
    InMux I__16660 (
            .O(N__86050),
            .I(N__86047));
    LocalMux I__16659 (
            .O(N__86047),
            .I(N__86044));
    Span4Mux_v I__16658 (
            .O(N__86044),
            .I(N__86041));
    Span4Mux_h I__16657 (
            .O(N__86041),
            .I(N__86031));
    InMux I__16656 (
            .O(N__86040),
            .I(N__86018));
    InMux I__16655 (
            .O(N__86039),
            .I(N__86018));
    InMux I__16654 (
            .O(N__86038),
            .I(N__86018));
    InMux I__16653 (
            .O(N__86037),
            .I(N__86018));
    InMux I__16652 (
            .O(N__86036),
            .I(N__86018));
    InMux I__16651 (
            .O(N__86035),
            .I(N__86018));
    InMux I__16650 (
            .O(N__86034),
            .I(N__86015));
    Span4Mux_h I__16649 (
            .O(N__86031),
            .I(N__86010));
    LocalMux I__16648 (
            .O(N__86018),
            .I(N__86010));
    LocalMux I__16647 (
            .O(N__86015),
            .I(N__86006));
    Span4Mux_v I__16646 (
            .O(N__86010),
            .I(N__86003));
    InMux I__16645 (
            .O(N__86009),
            .I(N__86000));
    Odrv4 I__16644 (
            .O(N__86006),
            .I(rco_int_0_a3_0_a2_0_183));
    Odrv4 I__16643 (
            .O(N__86003),
            .I(rco_int_0_a3_0_a2_0_183));
    LocalMux I__16642 (
            .O(N__86000),
            .I(rco_int_0_a3_0_a2_0_183));
    IoInMux I__16641 (
            .O(N__85993),
            .I(N__85986));
    InMux I__16640 (
            .O(N__85992),
            .I(N__85975));
    InMux I__16639 (
            .O(N__85991),
            .I(N__85975));
    InMux I__16638 (
            .O(N__85990),
            .I(N__85975));
    InMux I__16637 (
            .O(N__85989),
            .I(N__85975));
    LocalMux I__16636 (
            .O(N__85986),
            .I(N__85972));
    CascadeMux I__16635 (
            .O(N__85985),
            .I(N__85965));
    InMux I__16634 (
            .O(N__85984),
            .I(N__85961));
    LocalMux I__16633 (
            .O(N__85975),
            .I(N__85958));
    Span4Mux_s2_v I__16632 (
            .O(N__85972),
            .I(N__85955));
    InMux I__16631 (
            .O(N__85971),
            .I(N__85952));
    CascadeMux I__16630 (
            .O(N__85970),
            .I(N__85949));
    InMux I__16629 (
            .O(N__85969),
            .I(N__85945));
    CascadeMux I__16628 (
            .O(N__85968),
            .I(N__85942));
    InMux I__16627 (
            .O(N__85965),
            .I(N__85936));
    InMux I__16626 (
            .O(N__85964),
            .I(N__85936));
    LocalMux I__16625 (
            .O(N__85961),
            .I(N__85933));
    Span12Mux_h I__16624 (
            .O(N__85958),
            .I(N__85927));
    Span4Mux_h I__16623 (
            .O(N__85955),
            .I(N__85922));
    LocalMux I__16622 (
            .O(N__85952),
            .I(N__85922));
    InMux I__16621 (
            .O(N__85949),
            .I(N__85917));
    InMux I__16620 (
            .O(N__85948),
            .I(N__85917));
    LocalMux I__16619 (
            .O(N__85945),
            .I(N__85914));
    InMux I__16618 (
            .O(N__85942),
            .I(N__85909));
    InMux I__16617 (
            .O(N__85941),
            .I(N__85909));
    LocalMux I__16616 (
            .O(N__85936),
            .I(N__85904));
    Span4Mux_h I__16615 (
            .O(N__85933),
            .I(N__85904));
    CascadeMux I__16614 (
            .O(N__85932),
            .I(N__85901));
    CascadeMux I__16613 (
            .O(N__85931),
            .I(N__85896));
    CascadeMux I__16612 (
            .O(N__85930),
            .I(N__85892));
    Span12Mux_v I__16611 (
            .O(N__85927),
            .I(N__85889));
    Span4Mux_v I__16610 (
            .O(N__85922),
            .I(N__85886));
    LocalMux I__16609 (
            .O(N__85917),
            .I(N__85883));
    Span4Mux_v I__16608 (
            .O(N__85914),
            .I(N__85878));
    LocalMux I__16607 (
            .O(N__85909),
            .I(N__85878));
    Span4Mux_h I__16606 (
            .O(N__85904),
            .I(N__85875));
    InMux I__16605 (
            .O(N__85901),
            .I(N__85862));
    InMux I__16604 (
            .O(N__85900),
            .I(N__85862));
    InMux I__16603 (
            .O(N__85899),
            .I(N__85862));
    InMux I__16602 (
            .O(N__85896),
            .I(N__85862));
    InMux I__16601 (
            .O(N__85895),
            .I(N__85862));
    InMux I__16600 (
            .O(N__85892),
            .I(N__85862));
    Odrv12 I__16599 (
            .O(N__85889),
            .I(rco_c_172));
    Odrv4 I__16598 (
            .O(N__85886),
            .I(rco_c_172));
    Odrv4 I__16597 (
            .O(N__85883),
            .I(rco_c_172));
    Odrv4 I__16596 (
            .O(N__85878),
            .I(rco_c_172));
    Odrv4 I__16595 (
            .O(N__85875),
            .I(rco_c_172));
    LocalMux I__16594 (
            .O(N__85862),
            .I(rco_c_172));
    InMux I__16593 (
            .O(N__85849),
            .I(N__85846));
    LocalMux I__16592 (
            .O(N__85846),
            .I(shift_srl_163Z0Z_1));
    InMux I__16591 (
            .O(N__85843),
            .I(N__85840));
    LocalMux I__16590 (
            .O(N__85840),
            .I(shift_srl_163Z0Z_2));
    InMux I__16589 (
            .O(N__85837),
            .I(N__85834));
    LocalMux I__16588 (
            .O(N__85834),
            .I(shift_srl_163Z0Z_3));
    InMux I__16587 (
            .O(N__85831),
            .I(N__85828));
    LocalMux I__16586 (
            .O(N__85828),
            .I(shift_srl_163Z0Z_4));
    InMux I__16585 (
            .O(N__85825),
            .I(N__85822));
    LocalMux I__16584 (
            .O(N__85822),
            .I(shift_srl_163Z0Z_5));
    InMux I__16583 (
            .O(N__85819),
            .I(N__85816));
    LocalMux I__16582 (
            .O(N__85816),
            .I(shift_srl_163Z0Z_6));
    InMux I__16581 (
            .O(N__85813),
            .I(N__85810));
    LocalMux I__16580 (
            .O(N__85810),
            .I(shift_srl_163Z0Z_7));
    CEMux I__16579 (
            .O(N__85807),
            .I(N__85804));
    LocalMux I__16578 (
            .O(N__85804),
            .I(N__85800));
    CEMux I__16577 (
            .O(N__85803),
            .I(N__85797));
    Span4Mux_h I__16576 (
            .O(N__85800),
            .I(N__85791));
    LocalMux I__16575 (
            .O(N__85797),
            .I(N__85791));
    InMux I__16574 (
            .O(N__85796),
            .I(N__85788));
    Odrv4 I__16573 (
            .O(N__85791),
            .I(clk_en_163));
    LocalMux I__16572 (
            .O(N__85788),
            .I(clk_en_163));
    CascadeMux I__16571 (
            .O(N__85783),
            .I(N__85780));
    InMux I__16570 (
            .O(N__85780),
            .I(N__85777));
    LocalMux I__16569 (
            .O(N__85777),
            .I(N__85773));
    InMux I__16568 (
            .O(N__85776),
            .I(N__85770));
    Span4Mux_h I__16567 (
            .O(N__85773),
            .I(N__85767));
    LocalMux I__16566 (
            .O(N__85770),
            .I(shift_srl_191Z0Z_15));
    Odrv4 I__16565 (
            .O(N__85767),
            .I(shift_srl_191Z0Z_15));
    InMux I__16564 (
            .O(N__85762),
            .I(N__85759));
    LocalMux I__16563 (
            .O(N__85759),
            .I(shift_srl_191Z0Z_0));
    InMux I__16562 (
            .O(N__85756),
            .I(N__85753));
    LocalMux I__16561 (
            .O(N__85753),
            .I(shift_srl_191Z0Z_1));
    InMux I__16560 (
            .O(N__85750),
            .I(N__85747));
    LocalMux I__16559 (
            .O(N__85747),
            .I(shift_srl_164Z0Z_10));
    InMux I__16558 (
            .O(N__85744),
            .I(N__85741));
    LocalMux I__16557 (
            .O(N__85741),
            .I(shift_srl_164Z0Z_13));
    InMux I__16556 (
            .O(N__85738),
            .I(N__85735));
    LocalMux I__16555 (
            .O(N__85735),
            .I(shift_srl_164Z0Z_14));
    InMux I__16554 (
            .O(N__85732),
            .I(N__85729));
    LocalMux I__16553 (
            .O(N__85729),
            .I(shift_srl_164Z0Z_8));
    InMux I__16552 (
            .O(N__85726),
            .I(N__85723));
    LocalMux I__16551 (
            .O(N__85723),
            .I(shift_srl_164Z0Z_9));
    InMux I__16550 (
            .O(N__85720),
            .I(N__85717));
    LocalMux I__16549 (
            .O(N__85717),
            .I(shift_srl_164Z0Z_6));
    InMux I__16548 (
            .O(N__85714),
            .I(N__85711));
    LocalMux I__16547 (
            .O(N__85711),
            .I(shift_srl_164Z0Z_7));
    InMux I__16546 (
            .O(N__85708),
            .I(N__85705));
    LocalMux I__16545 (
            .O(N__85705),
            .I(shift_srl_163Z0Z_0));
    InMux I__16544 (
            .O(N__85702),
            .I(N__85699));
    LocalMux I__16543 (
            .O(N__85699),
            .I(shift_srl_33Z0Z_10));
    InMux I__16542 (
            .O(N__85696),
            .I(N__85693));
    LocalMux I__16541 (
            .O(N__85693),
            .I(shift_srl_33Z0Z_11));
    InMux I__16540 (
            .O(N__85690),
            .I(N__85687));
    LocalMux I__16539 (
            .O(N__85687),
            .I(shift_srl_33Z0Z_12));
    InMux I__16538 (
            .O(N__85684),
            .I(N__85681));
    LocalMux I__16537 (
            .O(N__85681),
            .I(shift_srl_33Z0Z_4));
    InMux I__16536 (
            .O(N__85678),
            .I(N__85675));
    LocalMux I__16535 (
            .O(N__85675),
            .I(shift_srl_33Z0Z_5));
    InMux I__16534 (
            .O(N__85672),
            .I(N__85669));
    LocalMux I__16533 (
            .O(N__85669),
            .I(shift_srl_33Z0Z_6));
    InMux I__16532 (
            .O(N__85666),
            .I(N__85663));
    LocalMux I__16531 (
            .O(N__85663),
            .I(shift_srl_33Z0Z_9));
    InMux I__16530 (
            .O(N__85660),
            .I(N__85657));
    LocalMux I__16529 (
            .O(N__85657),
            .I(shift_srl_33Z0Z_7));
    InMux I__16528 (
            .O(N__85654),
            .I(N__85651));
    LocalMux I__16527 (
            .O(N__85651),
            .I(shift_srl_33Z0Z_8));
    CEMux I__16526 (
            .O(N__85648),
            .I(N__85645));
    LocalMux I__16525 (
            .O(N__85645),
            .I(N__85641));
    CEMux I__16524 (
            .O(N__85644),
            .I(N__85638));
    Span4Mux_h I__16523 (
            .O(N__85641),
            .I(N__85635));
    LocalMux I__16522 (
            .O(N__85638),
            .I(N__85632));
    Odrv4 I__16521 (
            .O(N__85635),
            .I(clk_en_33));
    Odrv4 I__16520 (
            .O(N__85632),
            .I(clk_en_33));
    InMux I__16519 (
            .O(N__85627),
            .I(N__85624));
    LocalMux I__16518 (
            .O(N__85624),
            .I(shift_srl_37Z0Z_7));
    InMux I__16517 (
            .O(N__85621),
            .I(N__85618));
    LocalMux I__16516 (
            .O(N__85618),
            .I(shift_srl_37Z0Z_8));
    InMux I__16515 (
            .O(N__85615),
            .I(N__85612));
    LocalMux I__16514 (
            .O(N__85612),
            .I(shift_srl_33Z0Z_0));
    InMux I__16513 (
            .O(N__85609),
            .I(N__85606));
    LocalMux I__16512 (
            .O(N__85606),
            .I(shift_srl_33Z0Z_1));
    InMux I__16511 (
            .O(N__85603),
            .I(N__85600));
    LocalMux I__16510 (
            .O(N__85600),
            .I(shift_srl_33Z0Z_2));
    InMux I__16509 (
            .O(N__85597),
            .I(N__85594));
    LocalMux I__16508 (
            .O(N__85594),
            .I(shift_srl_33Z0Z_3));
    InMux I__16507 (
            .O(N__85591),
            .I(N__85588));
    LocalMux I__16506 (
            .O(N__85588),
            .I(shift_srl_33Z0Z_13));
    InMux I__16505 (
            .O(N__85585),
            .I(N__85582));
    LocalMux I__16504 (
            .O(N__85582),
            .I(shift_srl_33Z0Z_14));
    CascadeMux I__16503 (
            .O(N__85579),
            .I(N__85576));
    InMux I__16502 (
            .O(N__85576),
            .I(N__85569));
    InMux I__16501 (
            .O(N__85575),
            .I(N__85569));
    InMux I__16500 (
            .O(N__85574),
            .I(N__85566));
    LocalMux I__16499 (
            .O(N__85569),
            .I(N__85563));
    LocalMux I__16498 (
            .O(N__85566),
            .I(N__85560));
    Span4Mux_h I__16497 (
            .O(N__85563),
            .I(N__85557));
    Span4Mux_h I__16496 (
            .O(N__85560),
            .I(N__85552));
    Span4Mux_v I__16495 (
            .O(N__85557),
            .I(N__85549));
    InMux I__16494 (
            .O(N__85556),
            .I(N__85546));
    InMux I__16493 (
            .O(N__85555),
            .I(N__85543));
    Span4Mux_h I__16492 (
            .O(N__85552),
            .I(N__85540));
    Span4Mux_h I__16491 (
            .O(N__85549),
            .I(N__85537));
    LocalMux I__16490 (
            .O(N__85546),
            .I(shift_srl_33Z0Z_15));
    LocalMux I__16489 (
            .O(N__85543),
            .I(shift_srl_33Z0Z_15));
    Odrv4 I__16488 (
            .O(N__85540),
            .I(shift_srl_33Z0Z_15));
    Odrv4 I__16487 (
            .O(N__85537),
            .I(shift_srl_33Z0Z_15));
    InMux I__16486 (
            .O(N__85528),
            .I(N__85525));
    LocalMux I__16485 (
            .O(N__85525),
            .I(shift_srl_70Z0Z_8));
    InMux I__16484 (
            .O(N__85522),
            .I(N__85519));
    LocalMux I__16483 (
            .O(N__85519),
            .I(shift_srl_70Z0Z_9));
    InMux I__16482 (
            .O(N__85516),
            .I(N__85513));
    LocalMux I__16481 (
            .O(N__85513),
            .I(shift_srl_70Z0Z_0));
    CEMux I__16480 (
            .O(N__85510),
            .I(N__85506));
    CEMux I__16479 (
            .O(N__85509),
            .I(N__85503));
    LocalMux I__16478 (
            .O(N__85506),
            .I(clk_en_70));
    LocalMux I__16477 (
            .O(N__85503),
            .I(clk_en_70));
    InMux I__16476 (
            .O(N__85498),
            .I(N__85495));
    LocalMux I__16475 (
            .O(N__85495),
            .I(shift_srl_34Z0Z_4));
    InMux I__16474 (
            .O(N__85492),
            .I(N__85489));
    LocalMux I__16473 (
            .O(N__85489),
            .I(shift_srl_34Z0Z_5));
    InMux I__16472 (
            .O(N__85486),
            .I(N__85483));
    LocalMux I__16471 (
            .O(N__85483),
            .I(shift_srl_37Z0Z_12));
    InMux I__16470 (
            .O(N__85480),
            .I(N__85477));
    LocalMux I__16469 (
            .O(N__85477),
            .I(shift_srl_37Z0Z_13));
    InMux I__16468 (
            .O(N__85474),
            .I(N__85471));
    LocalMux I__16467 (
            .O(N__85471),
            .I(shift_srl_37Z0Z_5));
    InMux I__16466 (
            .O(N__85468),
            .I(N__85465));
    LocalMux I__16465 (
            .O(N__85465),
            .I(shift_srl_37Z0Z_6));
    InMux I__16464 (
            .O(N__85462),
            .I(N__85459));
    LocalMux I__16463 (
            .O(N__85459),
            .I(shift_srl_37Z0Z_9));
    InMux I__16462 (
            .O(N__85456),
            .I(N__85453));
    LocalMux I__16461 (
            .O(N__85453),
            .I(N__85450));
    Span4Mux_v I__16460 (
            .O(N__85450),
            .I(N__85447));
    Odrv4 I__16459 (
            .O(N__85447),
            .I(shift_srl_69Z0Z_6));
    InMux I__16458 (
            .O(N__85444),
            .I(N__85441));
    LocalMux I__16457 (
            .O(N__85441),
            .I(shift_srl_69Z0Z_7));
    InMux I__16456 (
            .O(N__85438),
            .I(N__85435));
    LocalMux I__16455 (
            .O(N__85435),
            .I(shift_srl_69Z0Z_8));
    InMux I__16454 (
            .O(N__85432),
            .I(N__85429));
    LocalMux I__16453 (
            .O(N__85429),
            .I(N__85426));
    Odrv4 I__16452 (
            .O(N__85426),
            .I(shift_srl_69Z0Z_9));
    CEMux I__16451 (
            .O(N__85423),
            .I(N__85418));
    CEMux I__16450 (
            .O(N__85422),
            .I(N__85415));
    CEMux I__16449 (
            .O(N__85421),
            .I(N__85412));
    LocalMux I__16448 (
            .O(N__85418),
            .I(N__85407));
    LocalMux I__16447 (
            .O(N__85415),
            .I(N__85407));
    LocalMux I__16446 (
            .O(N__85412),
            .I(N__85404));
    Span4Mux_v I__16445 (
            .O(N__85407),
            .I(N__85401));
    Span4Mux_h I__16444 (
            .O(N__85404),
            .I(N__85398));
    Span4Mux_h I__16443 (
            .O(N__85401),
            .I(N__85395));
    Odrv4 I__16442 (
            .O(N__85398),
            .I(clk_en_69));
    Odrv4 I__16441 (
            .O(N__85395),
            .I(clk_en_69));
    InMux I__16440 (
            .O(N__85390),
            .I(N__85387));
    LocalMux I__16439 (
            .O(N__85387),
            .I(shift_srl_70Z0Z_10));
    InMux I__16438 (
            .O(N__85384),
            .I(N__85381));
    LocalMux I__16437 (
            .O(N__85381),
            .I(shift_srl_70Z0Z_11));
    InMux I__16436 (
            .O(N__85378),
            .I(N__85375));
    LocalMux I__16435 (
            .O(N__85375),
            .I(shift_srl_70Z0Z_12));
    InMux I__16434 (
            .O(N__85372),
            .I(N__85369));
    LocalMux I__16433 (
            .O(N__85369),
            .I(shift_srl_70Z0Z_13));
    InMux I__16432 (
            .O(N__85366),
            .I(N__85363));
    LocalMux I__16431 (
            .O(N__85363),
            .I(shift_srl_70Z0Z_14));
    InMux I__16430 (
            .O(N__85360),
            .I(N__85357));
    LocalMux I__16429 (
            .O(N__85357),
            .I(shift_srl_69Z0Z_10));
    InMux I__16428 (
            .O(N__85354),
            .I(N__85351));
    LocalMux I__16427 (
            .O(N__85351),
            .I(shift_srl_71Z0Z_4));
    InMux I__16426 (
            .O(N__85348),
            .I(N__85345));
    LocalMux I__16425 (
            .O(N__85345),
            .I(shift_srl_71Z0Z_5));
    InMux I__16424 (
            .O(N__85342),
            .I(N__85339));
    LocalMux I__16423 (
            .O(N__85339),
            .I(shift_srl_71Z0Z_6));
    InMux I__16422 (
            .O(N__85336),
            .I(N__85333));
    LocalMux I__16421 (
            .O(N__85333),
            .I(shift_srl_71Z0Z_13));
    InMux I__16420 (
            .O(N__85330),
            .I(N__85327));
    LocalMux I__16419 (
            .O(N__85327),
            .I(shift_srl_71Z0Z_14));
    InMux I__16418 (
            .O(N__85324),
            .I(N__85321));
    LocalMux I__16417 (
            .O(N__85321),
            .I(shift_srl_71Z0Z_11));
    InMux I__16416 (
            .O(N__85318),
            .I(N__85315));
    LocalMux I__16415 (
            .O(N__85315),
            .I(shift_srl_71Z0Z_12));
    InMux I__16414 (
            .O(N__85312),
            .I(N__85309));
    LocalMux I__16413 (
            .O(N__85309),
            .I(shift_srl_71Z0Z_7));
    InMux I__16412 (
            .O(N__85306),
            .I(N__85303));
    LocalMux I__16411 (
            .O(N__85303),
            .I(shift_srl_71Z0Z_8));
    CEMux I__16410 (
            .O(N__85300),
            .I(N__85297));
    LocalMux I__16409 (
            .O(N__85297),
            .I(N__85293));
    CEMux I__16408 (
            .O(N__85296),
            .I(N__85290));
    Span4Mux_h I__16407 (
            .O(N__85293),
            .I(N__85285));
    LocalMux I__16406 (
            .O(N__85290),
            .I(N__85285));
    Span4Mux_h I__16405 (
            .O(N__85285),
            .I(N__85282));
    Odrv4 I__16404 (
            .O(N__85282),
            .I(clk_en_71));
    InMux I__16403 (
            .O(N__85279),
            .I(N__85276));
    LocalMux I__16402 (
            .O(N__85276),
            .I(N__85273));
    Span12Mux_h I__16401 (
            .O(N__85273),
            .I(N__85270));
    Odrv12 I__16400 (
            .O(N__85270),
            .I(rco_int_0_a2_1_a2_sx_59));
    CascadeMux I__16399 (
            .O(N__85267),
            .I(N__85262));
    InMux I__16398 (
            .O(N__85266),
            .I(N__85258));
    InMux I__16397 (
            .O(N__85265),
            .I(N__85255));
    InMux I__16396 (
            .O(N__85262),
            .I(N__85250));
    InMux I__16395 (
            .O(N__85261),
            .I(N__85250));
    LocalMux I__16394 (
            .O(N__85258),
            .I(N__85247));
    LocalMux I__16393 (
            .O(N__85255),
            .I(N__85244));
    LocalMux I__16392 (
            .O(N__85250),
            .I(N__85241));
    Span4Mux_h I__16391 (
            .O(N__85247),
            .I(N__85238));
    Odrv4 I__16390 (
            .O(N__85244),
            .I(rco_int_0_a2_1_a2_sx_44));
    Odrv12 I__16389 (
            .O(N__85241),
            .I(rco_int_0_a2_1_a2_sx_44));
    Odrv4 I__16388 (
            .O(N__85238),
            .I(rco_int_0_a2_1_a2_sx_44));
    IoInMux I__16387 (
            .O(N__85231),
            .I(N__85221));
    CascadeMux I__16386 (
            .O(N__85230),
            .I(N__85218));
    InMux I__16385 (
            .O(N__85229),
            .I(N__85204));
    InMux I__16384 (
            .O(N__85228),
            .I(N__85204));
    InMux I__16383 (
            .O(N__85227),
            .I(N__85204));
    InMux I__16382 (
            .O(N__85226),
            .I(N__85204));
    InMux I__16381 (
            .O(N__85225),
            .I(N__85204));
    InMux I__16380 (
            .O(N__85224),
            .I(N__85201));
    LocalMux I__16379 (
            .O(N__85221),
            .I(N__85198));
    InMux I__16378 (
            .O(N__85218),
            .I(N__85191));
    InMux I__16377 (
            .O(N__85217),
            .I(N__85186));
    InMux I__16376 (
            .O(N__85216),
            .I(N__85186));
    InMux I__16375 (
            .O(N__85215),
            .I(N__85183));
    LocalMux I__16374 (
            .O(N__85204),
            .I(N__85180));
    LocalMux I__16373 (
            .O(N__85201),
            .I(N__85173));
    IoSpan4Mux I__16372 (
            .O(N__85198),
            .I(N__85169));
    InMux I__16371 (
            .O(N__85197),
            .I(N__85166));
    InMux I__16370 (
            .O(N__85196),
            .I(N__85161));
    InMux I__16369 (
            .O(N__85195),
            .I(N__85161));
    InMux I__16368 (
            .O(N__85194),
            .I(N__85157));
    LocalMux I__16367 (
            .O(N__85191),
            .I(N__85152));
    LocalMux I__16366 (
            .O(N__85186),
            .I(N__85152));
    LocalMux I__16365 (
            .O(N__85183),
            .I(N__85149));
    Span4Mux_v I__16364 (
            .O(N__85180),
            .I(N__85146));
    InMux I__16363 (
            .O(N__85179),
            .I(N__85143));
    InMux I__16362 (
            .O(N__85178),
            .I(N__85136));
    InMux I__16361 (
            .O(N__85177),
            .I(N__85136));
    InMux I__16360 (
            .O(N__85176),
            .I(N__85136));
    Span4Mux_v I__16359 (
            .O(N__85173),
            .I(N__85133));
    InMux I__16358 (
            .O(N__85172),
            .I(N__85130));
    Span4Mux_s2_h I__16357 (
            .O(N__85169),
            .I(N__85126));
    LocalMux I__16356 (
            .O(N__85166),
            .I(N__85123));
    LocalMux I__16355 (
            .O(N__85161),
            .I(N__85120));
    InMux I__16354 (
            .O(N__85160),
            .I(N__85117));
    LocalMux I__16353 (
            .O(N__85157),
            .I(N__85113));
    Span4Mux_v I__16352 (
            .O(N__85152),
            .I(N__85110));
    Span4Mux_v I__16351 (
            .O(N__85149),
            .I(N__85105));
    Span4Mux_h I__16350 (
            .O(N__85146),
            .I(N__85105));
    LocalMux I__16349 (
            .O(N__85143),
            .I(N__85100));
    LocalMux I__16348 (
            .O(N__85136),
            .I(N__85100));
    Span4Mux_v I__16347 (
            .O(N__85133),
            .I(N__85097));
    LocalMux I__16346 (
            .O(N__85130),
            .I(N__85094));
    InMux I__16345 (
            .O(N__85129),
            .I(N__85091));
    Span4Mux_h I__16344 (
            .O(N__85126),
            .I(N__85087));
    Span4Mux_h I__16343 (
            .O(N__85123),
            .I(N__85084));
    Span12Mux_h I__16342 (
            .O(N__85120),
            .I(N__85081));
    LocalMux I__16341 (
            .O(N__85117),
            .I(N__85078));
    InMux I__16340 (
            .O(N__85116),
            .I(N__85075));
    Span4Mux_v I__16339 (
            .O(N__85113),
            .I(N__85066));
    Span4Mux_v I__16338 (
            .O(N__85110),
            .I(N__85066));
    Span4Mux_h I__16337 (
            .O(N__85105),
            .I(N__85066));
    Span4Mux_v I__16336 (
            .O(N__85100),
            .I(N__85066));
    Sp12to4 I__16335 (
            .O(N__85097),
            .I(N__85063));
    Sp12to4 I__16334 (
            .O(N__85094),
            .I(N__85058));
    LocalMux I__16333 (
            .O(N__85091),
            .I(N__85058));
    InMux I__16332 (
            .O(N__85090),
            .I(N__85055));
    Span4Mux_v I__16331 (
            .O(N__85087),
            .I(N__85052));
    Span4Mux_h I__16330 (
            .O(N__85084),
            .I(N__85049));
    Span12Mux_h I__16329 (
            .O(N__85081),
            .I(N__85044));
    Span12Mux_h I__16328 (
            .O(N__85078),
            .I(N__85044));
    LocalMux I__16327 (
            .O(N__85075),
            .I(N__85033));
    Sp12to4 I__16326 (
            .O(N__85066),
            .I(N__85033));
    Span12Mux_h I__16325 (
            .O(N__85063),
            .I(N__85033));
    Span12Mux_v I__16324 (
            .O(N__85058),
            .I(N__85033));
    LocalMux I__16323 (
            .O(N__85055),
            .I(N__85033));
    Odrv4 I__16322 (
            .O(N__85052),
            .I(N_4016_i));
    Odrv4 I__16321 (
            .O(N__85049),
            .I(N_4016_i));
    Odrv12 I__16320 (
            .O(N__85044),
            .I(N_4016_i));
    Odrv12 I__16319 (
            .O(N__85033),
            .I(N_4016_i));
    CascadeMux I__16318 (
            .O(N__85024),
            .I(rco_c_59_cascade_));
    InMux I__16317 (
            .O(N__85021),
            .I(N__85009));
    InMux I__16316 (
            .O(N__85020),
            .I(N__85009));
    InMux I__16315 (
            .O(N__85019),
            .I(N__85009));
    InMux I__16314 (
            .O(N__85018),
            .I(N__85009));
    LocalMux I__16313 (
            .O(N__85009),
            .I(N__85005));
    InMux I__16312 (
            .O(N__85008),
            .I(N__85000));
    Span4Mux_v I__16311 (
            .O(N__85005),
            .I(N__84994));
    InMux I__16310 (
            .O(N__85004),
            .I(N__84991));
    InMux I__16309 (
            .O(N__85003),
            .I(N__84988));
    LocalMux I__16308 (
            .O(N__85000),
            .I(N__84985));
    InMux I__16307 (
            .O(N__84999),
            .I(N__84982));
    InMux I__16306 (
            .O(N__84998),
            .I(N__84979));
    InMux I__16305 (
            .O(N__84997),
            .I(N__84976));
    Span4Mux_h I__16304 (
            .O(N__84994),
            .I(N__84971));
    LocalMux I__16303 (
            .O(N__84991),
            .I(N__84971));
    LocalMux I__16302 (
            .O(N__84988),
            .I(N__84968));
    Span4Mux_v I__16301 (
            .O(N__84985),
            .I(N__84965));
    LocalMux I__16300 (
            .O(N__84982),
            .I(N__84962));
    LocalMux I__16299 (
            .O(N__84979),
            .I(N__84957));
    LocalMux I__16298 (
            .O(N__84976),
            .I(N__84957));
    Span4Mux_h I__16297 (
            .O(N__84971),
            .I(N__84952));
    Span4Mux_h I__16296 (
            .O(N__84968),
            .I(N__84952));
    Span4Mux_h I__16295 (
            .O(N__84965),
            .I(N__84948));
    Span4Mux_v I__16294 (
            .O(N__84962),
            .I(N__84945));
    Span12Mux_v I__16293 (
            .O(N__84957),
            .I(N__84942));
    Span4Mux_v I__16292 (
            .O(N__84952),
            .I(N__84939));
    InMux I__16291 (
            .O(N__84951),
            .I(N__84936));
    Odrv4 I__16290 (
            .O(N__84948),
            .I(rco_int_0_a3_0_a2_0_66));
    Odrv4 I__16289 (
            .O(N__84945),
            .I(rco_int_0_a3_0_a2_0_66));
    Odrv12 I__16288 (
            .O(N__84942),
            .I(rco_int_0_a3_0_a2_0_66));
    Odrv4 I__16287 (
            .O(N__84939),
            .I(rco_int_0_a3_0_a2_0_66));
    LocalMux I__16286 (
            .O(N__84936),
            .I(rco_int_0_a3_0_a2_0_66));
    InMux I__16285 (
            .O(N__84925),
            .I(N__84912));
    InMux I__16284 (
            .O(N__84924),
            .I(N__84912));
    InMux I__16283 (
            .O(N__84923),
            .I(N__84912));
    InMux I__16282 (
            .O(N__84922),
            .I(N__84912));
    IoInMux I__16281 (
            .O(N__84921),
            .I(N__84909));
    LocalMux I__16280 (
            .O(N__84912),
            .I(N__84906));
    LocalMux I__16279 (
            .O(N__84909),
            .I(N__84899));
    Span4Mux_h I__16278 (
            .O(N__84906),
            .I(N__84896));
    InMux I__16277 (
            .O(N__84905),
            .I(N__84890));
    InMux I__16276 (
            .O(N__84904),
            .I(N__84890));
    InMux I__16275 (
            .O(N__84903),
            .I(N__84887));
    InMux I__16274 (
            .O(N__84902),
            .I(N__84884));
    IoSpan4Mux I__16273 (
            .O(N__84899),
            .I(N__84881));
    Span4Mux_h I__16272 (
            .O(N__84896),
            .I(N__84878));
    InMux I__16271 (
            .O(N__84895),
            .I(N__84875));
    LocalMux I__16270 (
            .O(N__84890),
            .I(N__84870));
    LocalMux I__16269 (
            .O(N__84887),
            .I(N__84870));
    LocalMux I__16268 (
            .O(N__84884),
            .I(N__84867));
    Span4Mux_s1_h I__16267 (
            .O(N__84881),
            .I(N__84861));
    Span4Mux_v I__16266 (
            .O(N__84878),
            .I(N__84856));
    LocalMux I__16265 (
            .O(N__84875),
            .I(N__84856));
    Span4Mux_v I__16264 (
            .O(N__84870),
            .I(N__84851));
    Span4Mux_v I__16263 (
            .O(N__84867),
            .I(N__84851));
    InMux I__16262 (
            .O(N__84866),
            .I(N__84844));
    InMux I__16261 (
            .O(N__84865),
            .I(N__84844));
    InMux I__16260 (
            .O(N__84864),
            .I(N__84844));
    Odrv4 I__16259 (
            .O(N__84861),
            .I(rco_c_59));
    Odrv4 I__16258 (
            .O(N__84856),
            .I(rco_c_59));
    Odrv4 I__16257 (
            .O(N__84851),
            .I(rco_c_59));
    LocalMux I__16256 (
            .O(N__84844),
            .I(rco_c_59));
    CascadeMux I__16255 (
            .O(N__84835),
            .I(N__84829));
    CascadeMux I__16254 (
            .O(N__84834),
            .I(N__84825));
    CascadeMux I__16253 (
            .O(N__84833),
            .I(N__84822));
    InMux I__16252 (
            .O(N__84832),
            .I(N__84819));
    InMux I__16251 (
            .O(N__84829),
            .I(N__84816));
    InMux I__16250 (
            .O(N__84828),
            .I(N__84809));
    InMux I__16249 (
            .O(N__84825),
            .I(N__84809));
    InMux I__16248 (
            .O(N__84822),
            .I(N__84809));
    LocalMux I__16247 (
            .O(N__84819),
            .I(N__84802));
    LocalMux I__16246 (
            .O(N__84816),
            .I(N__84802));
    LocalMux I__16245 (
            .O(N__84809),
            .I(N__84802));
    Odrv4 I__16244 (
            .O(N__84802),
            .I(shift_srl_68_RNIHDC4Z0Z_15));
    InMux I__16243 (
            .O(N__84799),
            .I(N__84796));
    LocalMux I__16242 (
            .O(N__84796),
            .I(shift_srl_69Z0Z_14));
    InMux I__16241 (
            .O(N__84793),
            .I(N__84790));
    LocalMux I__16240 (
            .O(N__84790),
            .I(shift_srl_69Z0Z_13));
    InMux I__16239 (
            .O(N__84787),
            .I(N__84784));
    LocalMux I__16238 (
            .O(N__84784),
            .I(shift_srl_69Z0Z_12));
    InMux I__16237 (
            .O(N__84781),
            .I(N__84778));
    LocalMux I__16236 (
            .O(N__84778),
            .I(shift_srl_69Z0Z_11));
    InMux I__16235 (
            .O(N__84775),
            .I(N__84772));
    LocalMux I__16234 (
            .O(N__84772),
            .I(shift_srl_68Z0Z_2));
    InMux I__16233 (
            .O(N__84769),
            .I(N__84766));
    LocalMux I__16232 (
            .O(N__84766),
            .I(shift_srl_68Z0Z_3));
    InMux I__16231 (
            .O(N__84763),
            .I(N__84760));
    LocalMux I__16230 (
            .O(N__84760),
            .I(shift_srl_68Z0Z_4));
    InMux I__16229 (
            .O(N__84757),
            .I(N__84754));
    LocalMux I__16228 (
            .O(N__84754),
            .I(shift_srl_68Z0Z_5));
    InMux I__16227 (
            .O(N__84751),
            .I(N__84748));
    LocalMux I__16226 (
            .O(N__84748),
            .I(shift_srl_68Z0Z_6));
    IoInMux I__16225 (
            .O(N__84745),
            .I(N__84742));
    LocalMux I__16224 (
            .O(N__84742),
            .I(N__84739));
    Span12Mux_s5_h I__16223 (
            .O(N__84739),
            .I(N__84736));
    Odrv12 I__16222 (
            .O(N__84736),
            .I(rco_c_70));
    CascadeMux I__16221 (
            .O(N__84733),
            .I(shift_srl_71_RNIGP6RZ0Z_15_cascade_));
    CEMux I__16220 (
            .O(N__84730),
            .I(N__84726));
    CEMux I__16219 (
            .O(N__84729),
            .I(N__84723));
    LocalMux I__16218 (
            .O(N__84726),
            .I(clk_en_78));
    LocalMux I__16217 (
            .O(N__84723),
            .I(clk_en_78));
    InMux I__16216 (
            .O(N__84718),
            .I(N__84715));
    LocalMux I__16215 (
            .O(N__84715),
            .I(shift_srl_75Z0Z_14));
    InMux I__16214 (
            .O(N__84712),
            .I(N__84709));
    LocalMux I__16213 (
            .O(N__84709),
            .I(shift_srl_75Z0Z_13));
    InMux I__16212 (
            .O(N__84706),
            .I(N__84703));
    LocalMux I__16211 (
            .O(N__84703),
            .I(shift_srl_75Z0Z_12));
    InMux I__16210 (
            .O(N__84700),
            .I(N__84697));
    LocalMux I__16209 (
            .O(N__84697),
            .I(shift_srl_75Z0Z_11));
    InMux I__16208 (
            .O(N__84694),
            .I(N__84691));
    LocalMux I__16207 (
            .O(N__84691),
            .I(shift_srl_68Z0Z_0));
    InMux I__16206 (
            .O(N__84688),
            .I(N__84685));
    LocalMux I__16205 (
            .O(N__84685),
            .I(shift_srl_68Z0Z_1));
    CascadeMux I__16204 (
            .O(N__84682),
            .I(N__84679));
    InMux I__16203 (
            .O(N__84679),
            .I(N__84675));
    InMux I__16202 (
            .O(N__84678),
            .I(N__84671));
    LocalMux I__16201 (
            .O(N__84675),
            .I(N__84668));
    InMux I__16200 (
            .O(N__84674),
            .I(N__84665));
    LocalMux I__16199 (
            .O(N__84671),
            .I(shift_srl_80Z0Z_15));
    Odrv12 I__16198 (
            .O(N__84668),
            .I(shift_srl_80Z0Z_15));
    LocalMux I__16197 (
            .O(N__84665),
            .I(shift_srl_80Z0Z_15));
    InMux I__16196 (
            .O(N__84658),
            .I(N__84655));
    LocalMux I__16195 (
            .O(N__84655),
            .I(shift_srl_80Z0Z_14));
    InMux I__16194 (
            .O(N__84652),
            .I(N__84649));
    LocalMux I__16193 (
            .O(N__84649),
            .I(shift_srl_80Z0Z_13));
    InMux I__16192 (
            .O(N__84646),
            .I(N__84643));
    LocalMux I__16191 (
            .O(N__84643),
            .I(shift_srl_80Z0Z_12));
    InMux I__16190 (
            .O(N__84640),
            .I(N__84637));
    LocalMux I__16189 (
            .O(N__84637),
            .I(shift_srl_80Z0Z_11));
    InMux I__16188 (
            .O(N__84634),
            .I(N__84631));
    LocalMux I__16187 (
            .O(N__84631),
            .I(shift_srl_80Z0Z_10));
    InMux I__16186 (
            .O(N__84628),
            .I(N__84625));
    LocalMux I__16185 (
            .O(N__84625),
            .I(N__84622));
    Odrv4 I__16184 (
            .O(N__84622),
            .I(shift_srl_80Z0Z_8));
    InMux I__16183 (
            .O(N__84619),
            .I(N__84616));
    LocalMux I__16182 (
            .O(N__84616),
            .I(shift_srl_80Z0Z_9));
    CEMux I__16181 (
            .O(N__84613),
            .I(N__84609));
    CEMux I__16180 (
            .O(N__84612),
            .I(N__84606));
    LocalMux I__16179 (
            .O(N__84609),
            .I(N__84602));
    LocalMux I__16178 (
            .O(N__84606),
            .I(N__84599));
    CEMux I__16177 (
            .O(N__84605),
            .I(N__84596));
    Span4Mux_v I__16176 (
            .O(N__84602),
            .I(N__84593));
    Span4Mux_h I__16175 (
            .O(N__84599),
            .I(N__84590));
    LocalMux I__16174 (
            .O(N__84596),
            .I(N__84587));
    Odrv4 I__16173 (
            .O(N__84593),
            .I(clk_en_80));
    Odrv4 I__16172 (
            .O(N__84590),
            .I(clk_en_80));
    Odrv4 I__16171 (
            .O(N__84587),
            .I(clk_en_80));
    InMux I__16170 (
            .O(N__84580),
            .I(N__84577));
    LocalMux I__16169 (
            .O(N__84577),
            .I(N__84573));
    InMux I__16168 (
            .O(N__84576),
            .I(N__84569));
    Span4Mux_h I__16167 (
            .O(N__84573),
            .I(N__84566));
    InMux I__16166 (
            .O(N__84572),
            .I(N__84563));
    LocalMux I__16165 (
            .O(N__84569),
            .I(shift_srl_76Z0Z_15));
    Odrv4 I__16164 (
            .O(N__84566),
            .I(shift_srl_76Z0Z_15));
    LocalMux I__16163 (
            .O(N__84563),
            .I(shift_srl_76Z0Z_15));
    CascadeMux I__16162 (
            .O(N__84556),
            .I(shift_srl_76_RNIF788Z0Z_15_cascade_));
    InMux I__16161 (
            .O(N__84553),
            .I(N__84550));
    LocalMux I__16160 (
            .O(N__84550),
            .I(shift_srl_81Z0Z_5));
    InMux I__16159 (
            .O(N__84547),
            .I(N__84544));
    LocalMux I__16158 (
            .O(N__84544),
            .I(shift_srl_81Z0Z_6));
    InMux I__16157 (
            .O(N__84541),
            .I(N__84538));
    LocalMux I__16156 (
            .O(N__84538),
            .I(N__84535));
    Odrv12 I__16155 (
            .O(N__84535),
            .I(shift_srl_79_RNITG241Z0Z_15));
    CascadeMux I__16154 (
            .O(N__84532),
            .I(shift_srl_79_RNITG241Z0Z_15_cascade_));
    IoInMux I__16153 (
            .O(N__84529),
            .I(N__84526));
    LocalMux I__16152 (
            .O(N__84526),
            .I(N__84523));
    Span4Mux_s1_v I__16151 (
            .O(N__84523),
            .I(N__84520));
    Span4Mux_v I__16150 (
            .O(N__84520),
            .I(N__84517));
    Odrv4 I__16149 (
            .O(N__84517),
            .I(rco_c_78));
    InMux I__16148 (
            .O(N__84514),
            .I(N__84511));
    LocalMux I__16147 (
            .O(N__84511),
            .I(shift_srl_79Z0Z_0));
    InMux I__16146 (
            .O(N__84508),
            .I(N__84501));
    InMux I__16145 (
            .O(N__84507),
            .I(N__84497));
    InMux I__16144 (
            .O(N__84506),
            .I(N__84490));
    InMux I__16143 (
            .O(N__84505),
            .I(N__84490));
    InMux I__16142 (
            .O(N__84504),
            .I(N__84490));
    LocalMux I__16141 (
            .O(N__84501),
            .I(N__84487));
    InMux I__16140 (
            .O(N__84500),
            .I(N__84484));
    LocalMux I__16139 (
            .O(N__84497),
            .I(shift_srl_78Z0Z_15));
    LocalMux I__16138 (
            .O(N__84490),
            .I(shift_srl_78Z0Z_15));
    Odrv4 I__16137 (
            .O(N__84487),
            .I(shift_srl_78Z0Z_15));
    LocalMux I__16136 (
            .O(N__84484),
            .I(shift_srl_78Z0Z_15));
    InMux I__16135 (
            .O(N__84475),
            .I(N__84472));
    LocalMux I__16134 (
            .O(N__84472),
            .I(N__84469));
    Odrv12 I__16133 (
            .O(N__84469),
            .I(rco_int_0_a2_0_a2_0_1_83));
    InMux I__16132 (
            .O(N__84466),
            .I(N__84463));
    LocalMux I__16131 (
            .O(N__84463),
            .I(N__84460));
    Span4Mux_v I__16130 (
            .O(N__84460),
            .I(N__84457));
    Odrv4 I__16129 (
            .O(N__84457),
            .I(shift_srl_36Z0Z_5));
    InMux I__16128 (
            .O(N__84454),
            .I(N__84451));
    LocalMux I__16127 (
            .O(N__84451),
            .I(N__84448));
    Odrv4 I__16126 (
            .O(N__84448),
            .I(shift_srl_36Z0Z_6));
    IoInMux I__16125 (
            .O(N__84445),
            .I(N__84442));
    LocalMux I__16124 (
            .O(N__84442),
            .I(N__84439));
    Span4Mux_s0_v I__16123 (
            .O(N__84439),
            .I(N__84436));
    Odrv4 I__16122 (
            .O(N__84436),
            .I(rco_c_79));
    IoInMux I__16121 (
            .O(N__84433),
            .I(N__84430));
    LocalMux I__16120 (
            .O(N__84430),
            .I(N__84427));
    Odrv4 I__16119 (
            .O(N__84427),
            .I(N_785));
    InMux I__16118 (
            .O(N__84424),
            .I(N__84421));
    LocalMux I__16117 (
            .O(N__84421),
            .I(shift_srl_81Z0Z_0));
    InMux I__16116 (
            .O(N__84418),
            .I(N__84415));
    LocalMux I__16115 (
            .O(N__84415),
            .I(shift_srl_81Z0Z_1));
    InMux I__16114 (
            .O(N__84412),
            .I(N__84409));
    LocalMux I__16113 (
            .O(N__84409),
            .I(shift_srl_81Z0Z_2));
    InMux I__16112 (
            .O(N__84406),
            .I(N__84403));
    LocalMux I__16111 (
            .O(N__84403),
            .I(shift_srl_81Z0Z_3));
    InMux I__16110 (
            .O(N__84400),
            .I(N__84397));
    LocalMux I__16109 (
            .O(N__84397),
            .I(shift_srl_81Z0Z_4));
    InMux I__16108 (
            .O(N__84394),
            .I(N__84391));
    LocalMux I__16107 (
            .O(N__84391),
            .I(shift_srl_36Z0Z_7));
    InMux I__16106 (
            .O(N__84388),
            .I(N__84385));
    LocalMux I__16105 (
            .O(N__84385),
            .I(shift_srl_191Z0Z_10));
    InMux I__16104 (
            .O(N__84382),
            .I(N__84379));
    LocalMux I__16103 (
            .O(N__84379),
            .I(shift_srl_191Z0Z_11));
    InMux I__16102 (
            .O(N__84376),
            .I(N__84373));
    LocalMux I__16101 (
            .O(N__84373),
            .I(shift_srl_191Z0Z_12));
    InMux I__16100 (
            .O(N__84370),
            .I(N__84367));
    LocalMux I__16099 (
            .O(N__84367),
            .I(shift_srl_191Z0Z_13));
    InMux I__16098 (
            .O(N__84364),
            .I(N__84361));
    LocalMux I__16097 (
            .O(N__84361),
            .I(shift_srl_191Z0Z_14));
    InMux I__16096 (
            .O(N__84358),
            .I(N__84355));
    LocalMux I__16095 (
            .O(N__84355),
            .I(shift_srl_191Z0Z_9));
    InMux I__16094 (
            .O(N__84352),
            .I(N__84349));
    LocalMux I__16093 (
            .O(N__84349),
            .I(shift_srl_191Z0Z_8));
    InMux I__16092 (
            .O(N__84346),
            .I(N__84343));
    LocalMux I__16091 (
            .O(N__84343),
            .I(shift_srl_163Z0Z_14));
    InMux I__16090 (
            .O(N__84340),
            .I(N__84337));
    LocalMux I__16089 (
            .O(N__84337),
            .I(shift_srl_163Z0Z_9));
    InMux I__16088 (
            .O(N__84334),
            .I(N__84331));
    LocalMux I__16087 (
            .O(N__84331),
            .I(shift_srl_163Z0Z_8));
    InMux I__16086 (
            .O(N__84328),
            .I(N__84325));
    LocalMux I__16085 (
            .O(N__84325),
            .I(shift_srl_36Z0Z_10));
    InMux I__16084 (
            .O(N__84322),
            .I(N__84319));
    LocalMux I__16083 (
            .O(N__84319),
            .I(shift_srl_36Z0Z_11));
    InMux I__16082 (
            .O(N__84316),
            .I(N__84313));
    LocalMux I__16081 (
            .O(N__84313),
            .I(shift_srl_36Z0Z_12));
    InMux I__16080 (
            .O(N__84310),
            .I(N__84307));
    LocalMux I__16079 (
            .O(N__84307),
            .I(shift_srl_36Z0Z_9));
    InMux I__16078 (
            .O(N__84304),
            .I(N__84301));
    LocalMux I__16077 (
            .O(N__84301),
            .I(shift_srl_36Z0Z_8));
    CascadeMux I__16076 (
            .O(N__84298),
            .I(shift_srl_167_RNIUC2TZ0Z_15_cascade_));
    InMux I__16075 (
            .O(N__84295),
            .I(N__84292));
    LocalMux I__16074 (
            .O(N__84292),
            .I(N__84289));
    Span4Mux_h I__16073 (
            .O(N__84289),
            .I(N__84285));
    InMux I__16072 (
            .O(N__84288),
            .I(N__84282));
    Span4Mux_h I__16071 (
            .O(N__84285),
            .I(N__84279));
    LocalMux I__16070 (
            .O(N__84282),
            .I(shift_srl_170Z0Z_15));
    Odrv4 I__16069 (
            .O(N__84279),
            .I(shift_srl_170Z0Z_15));
    InMux I__16068 (
            .O(N__84274),
            .I(N__84268));
    InMux I__16067 (
            .O(N__84273),
            .I(N__84265));
    InMux I__16066 (
            .O(N__84272),
            .I(N__84260));
    InMux I__16065 (
            .O(N__84271),
            .I(N__84260));
    LocalMux I__16064 (
            .O(N__84268),
            .I(N__84255));
    LocalMux I__16063 (
            .O(N__84265),
            .I(N__84255));
    LocalMux I__16062 (
            .O(N__84260),
            .I(shift_srl_169Z0Z_15));
    Odrv4 I__16061 (
            .O(N__84255),
            .I(shift_srl_169Z0Z_15));
    CascadeMux I__16060 (
            .O(N__84250),
            .I(shift_srl_163_RNI3MR51Z0Z_15_cascade_));
    CascadeMux I__16059 (
            .O(N__84247),
            .I(shift_srl_170_RNIRM2S1Z0Z_15_cascade_));
    InMux I__16058 (
            .O(N__84244),
            .I(N__84241));
    LocalMux I__16057 (
            .O(N__84241),
            .I(N__84237));
    CascadeMux I__16056 (
            .O(N__84240),
            .I(N__84231));
    Span4Mux_v I__16055 (
            .O(N__84237),
            .I(N__84227));
    InMux I__16054 (
            .O(N__84236),
            .I(N__84224));
    CascadeMux I__16053 (
            .O(N__84235),
            .I(N__84221));
    InMux I__16052 (
            .O(N__84234),
            .I(N__84213));
    InMux I__16051 (
            .O(N__84231),
            .I(N__84213));
    InMux I__16050 (
            .O(N__84230),
            .I(N__84213));
    Span4Mux_h I__16049 (
            .O(N__84227),
            .I(N__84206));
    LocalMux I__16048 (
            .O(N__84224),
            .I(N__84206));
    InMux I__16047 (
            .O(N__84221),
            .I(N__84203));
    InMux I__16046 (
            .O(N__84220),
            .I(N__84200));
    LocalMux I__16045 (
            .O(N__84213),
            .I(N__84197));
    InMux I__16044 (
            .O(N__84212),
            .I(N__84192));
    InMux I__16043 (
            .O(N__84211),
            .I(N__84192));
    Span4Mux_v I__16042 (
            .O(N__84206),
            .I(N__84187));
    LocalMux I__16041 (
            .O(N__84203),
            .I(N__84187));
    LocalMux I__16040 (
            .O(N__84200),
            .I(N__84184));
    Span4Mux_h I__16039 (
            .O(N__84197),
            .I(N__84181));
    LocalMux I__16038 (
            .O(N__84192),
            .I(N__84176));
    Span4Mux_h I__16037 (
            .O(N__84187),
            .I(N__84176));
    Span12Mux_h I__16036 (
            .O(N__84184),
            .I(N__84173));
    Span4Mux_h I__16035 (
            .O(N__84181),
            .I(N__84168));
    Span4Mux_h I__16034 (
            .O(N__84176),
            .I(N__84168));
    Odrv12 I__16033 (
            .O(N__84173),
            .I(rco_int_0_a3_0_a2_0_172));
    Odrv4 I__16032 (
            .O(N__84168),
            .I(rco_int_0_a3_0_a2_0_172));
    CascadeMux I__16031 (
            .O(N__84163),
            .I(rco_int_0_a3_0_a2_0_172_cascade_));
    CascadeMux I__16030 (
            .O(N__84160),
            .I(N__84156));
    InMux I__16029 (
            .O(N__84159),
            .I(N__84151));
    InMux I__16028 (
            .O(N__84156),
            .I(N__84146));
    InMux I__16027 (
            .O(N__84155),
            .I(N__84146));
    InMux I__16026 (
            .O(N__84154),
            .I(N__84143));
    LocalMux I__16025 (
            .O(N__84151),
            .I(N__84140));
    LocalMux I__16024 (
            .O(N__84146),
            .I(N__84137));
    LocalMux I__16023 (
            .O(N__84143),
            .I(N__84134));
    Span4Mux_v I__16022 (
            .O(N__84140),
            .I(N__84131));
    Span4Mux_h I__16021 (
            .O(N__84137),
            .I(N__84128));
    Span4Mux_v I__16020 (
            .O(N__84134),
            .I(N__84125));
    Span4Mux_h I__16019 (
            .O(N__84131),
            .I(N__84120));
    Span4Mux_h I__16018 (
            .O(N__84128),
            .I(N__84120));
    Span4Mux_h I__16017 (
            .O(N__84125),
            .I(N__84117));
    Odrv4 I__16016 (
            .O(N__84120),
            .I(clk_en_0_a3_0_a2cf1_1_176));
    Odrv4 I__16015 (
            .O(N__84117),
            .I(clk_en_0_a3_0_a2cf1_1_176));
    InMux I__16014 (
            .O(N__84112),
            .I(N__84109));
    LocalMux I__16013 (
            .O(N__84109),
            .I(shift_srl_163Z0Z_10));
    InMux I__16012 (
            .O(N__84106),
            .I(N__84103));
    LocalMux I__16011 (
            .O(N__84103),
            .I(shift_srl_163Z0Z_11));
    InMux I__16010 (
            .O(N__84100),
            .I(N__84097));
    LocalMux I__16009 (
            .O(N__84097),
            .I(shift_srl_163Z0Z_12));
    InMux I__16008 (
            .O(N__84094),
            .I(N__84091));
    LocalMux I__16007 (
            .O(N__84091),
            .I(shift_srl_163Z0Z_13));
    InMux I__16006 (
            .O(N__84088),
            .I(N__84085));
    LocalMux I__16005 (
            .O(N__84085),
            .I(shift_srl_36Z0Z_0));
    InMux I__16004 (
            .O(N__84082),
            .I(N__84079));
    LocalMux I__16003 (
            .O(N__84079),
            .I(shift_srl_36Z0Z_1));
    InMux I__16002 (
            .O(N__84076),
            .I(N__84073));
    LocalMux I__16001 (
            .O(N__84073),
            .I(shift_srl_36Z0Z_2));
    InMux I__16000 (
            .O(N__84070),
            .I(N__84067));
    LocalMux I__15999 (
            .O(N__84067),
            .I(shift_srl_36Z0Z_3));
    InMux I__15998 (
            .O(N__84064),
            .I(N__84061));
    LocalMux I__15997 (
            .O(N__84061),
            .I(shift_srl_36Z0Z_4));
    IoInMux I__15996 (
            .O(N__84058),
            .I(N__84055));
    LocalMux I__15995 (
            .O(N__84055),
            .I(N__84052));
    IoSpan4Mux I__15994 (
            .O(N__84052),
            .I(N__84049));
    Span4Mux_s0_v I__15993 (
            .O(N__84049),
            .I(N__84046));
    Sp12to4 I__15992 (
            .O(N__84046),
            .I(N__84043));
    Span12Mux_v I__15991 (
            .O(N__84043),
            .I(N__84040));
    Odrv12 I__15990 (
            .O(N__84040),
            .I(rco_c_169));
    IoInMux I__15989 (
            .O(N__84037),
            .I(N__84034));
    LocalMux I__15988 (
            .O(N__84034),
            .I(N__84031));
    IoSpan4Mux I__15987 (
            .O(N__84031),
            .I(N__84028));
    Span4Mux_s2_v I__15986 (
            .O(N__84028),
            .I(N__84025));
    Span4Mux_h I__15985 (
            .O(N__84025),
            .I(N__84022));
    Sp12to4 I__15984 (
            .O(N__84022),
            .I(N__84019));
    Odrv12 I__15983 (
            .O(N__84019),
            .I(rco_c_168));
    InMux I__15982 (
            .O(N__84016),
            .I(N__84013));
    LocalMux I__15981 (
            .O(N__84013),
            .I(N__84007));
    InMux I__15980 (
            .O(N__84012),
            .I(N__84004));
    InMux I__15979 (
            .O(N__84011),
            .I(N__84001));
    InMux I__15978 (
            .O(N__84010),
            .I(N__83998));
    Span4Mux_v I__15977 (
            .O(N__84007),
            .I(N__83995));
    LocalMux I__15976 (
            .O(N__84004),
            .I(N__83992));
    LocalMux I__15975 (
            .O(N__84001),
            .I(shift_srl_166Z0Z_15));
    LocalMux I__15974 (
            .O(N__83998),
            .I(shift_srl_166Z0Z_15));
    Odrv4 I__15973 (
            .O(N__83995),
            .I(shift_srl_166Z0Z_15));
    Odrv12 I__15972 (
            .O(N__83992),
            .I(shift_srl_166Z0Z_15));
    InMux I__15971 (
            .O(N__83983),
            .I(N__83980));
    LocalMux I__15970 (
            .O(N__83980),
            .I(N__83977));
    Span4Mux_v I__15969 (
            .O(N__83977),
            .I(N__83974));
    Span4Mux_v I__15968 (
            .O(N__83974),
            .I(N__83971));
    Span4Mux_v I__15967 (
            .O(N__83971),
            .I(N__83966));
    InMux I__15966 (
            .O(N__83970),
            .I(N__83959));
    InMux I__15965 (
            .O(N__83969),
            .I(N__83959));
    Span4Mux_v I__15964 (
            .O(N__83966),
            .I(N__83956));
    InMux I__15963 (
            .O(N__83965),
            .I(N__83953));
    InMux I__15962 (
            .O(N__83964),
            .I(N__83950));
    LocalMux I__15961 (
            .O(N__83959),
            .I(N__83946));
    Span4Mux_h I__15960 (
            .O(N__83956),
            .I(N__83943));
    LocalMux I__15959 (
            .O(N__83953),
            .I(N__83940));
    LocalMux I__15958 (
            .O(N__83950),
            .I(N__83937));
    InMux I__15957 (
            .O(N__83949),
            .I(N__83934));
    Span4Mux_v I__15956 (
            .O(N__83946),
            .I(N__83931));
    Span4Mux_h I__15955 (
            .O(N__83943),
            .I(N__83926));
    Span4Mux_v I__15954 (
            .O(N__83940),
            .I(N__83926));
    Span4Mux_h I__15953 (
            .O(N__83937),
            .I(N__83923));
    LocalMux I__15952 (
            .O(N__83934),
            .I(shift_srl_165Z0Z_15));
    Odrv4 I__15951 (
            .O(N__83931),
            .I(shift_srl_165Z0Z_15));
    Odrv4 I__15950 (
            .O(N__83926),
            .I(shift_srl_165Z0Z_15));
    Odrv4 I__15949 (
            .O(N__83923),
            .I(shift_srl_165Z0Z_15));
    CascadeMux I__15948 (
            .O(N__83914),
            .I(N__83911));
    InMux I__15947 (
            .O(N__83911),
            .I(N__83907));
    InMux I__15946 (
            .O(N__83910),
            .I(N__83904));
    LocalMux I__15945 (
            .O(N__83907),
            .I(N__83901));
    LocalMux I__15944 (
            .O(N__83904),
            .I(shift_srl_167Z0Z_15));
    Odrv4 I__15943 (
            .O(N__83901),
            .I(shift_srl_167Z0Z_15));
    CascadeMux I__15942 (
            .O(N__83896),
            .I(rco_c_32_cascade_));
    InMux I__15941 (
            .O(N__83893),
            .I(N__83889));
    CascadeMux I__15940 (
            .O(N__83892),
            .I(N__83885));
    LocalMux I__15939 (
            .O(N__83889),
            .I(N__83880));
    InMux I__15938 (
            .O(N__83888),
            .I(N__83877));
    InMux I__15937 (
            .O(N__83885),
            .I(N__83872));
    InMux I__15936 (
            .O(N__83884),
            .I(N__83872));
    InMux I__15935 (
            .O(N__83883),
            .I(N__83869));
    Span4Mux_v I__15934 (
            .O(N__83880),
            .I(N__83866));
    LocalMux I__15933 (
            .O(N__83877),
            .I(N__83861));
    LocalMux I__15932 (
            .O(N__83872),
            .I(N__83861));
    LocalMux I__15931 (
            .O(N__83869),
            .I(N__83856));
    Sp12to4 I__15930 (
            .O(N__83866),
            .I(N__83856));
    Span4Mux_h I__15929 (
            .O(N__83861),
            .I(N__83853));
    Odrv12 I__15928 (
            .O(N__83856),
            .I(shift_srl_29Z0Z_15));
    Odrv4 I__15927 (
            .O(N__83853),
            .I(shift_srl_29Z0Z_15));
    InMux I__15926 (
            .O(N__83848),
            .I(N__83845));
    LocalMux I__15925 (
            .O(N__83845),
            .I(N__83842));
    Span4Mux_v I__15924 (
            .O(N__83842),
            .I(N__83834));
    InMux I__15923 (
            .O(N__83841),
            .I(N__83829));
    InMux I__15922 (
            .O(N__83840),
            .I(N__83829));
    InMux I__15921 (
            .O(N__83839),
            .I(N__83826));
    InMux I__15920 (
            .O(N__83838),
            .I(N__83823));
    InMux I__15919 (
            .O(N__83837),
            .I(N__83820));
    Sp12to4 I__15918 (
            .O(N__83834),
            .I(N__83817));
    LocalMux I__15917 (
            .O(N__83829),
            .I(N__83814));
    LocalMux I__15916 (
            .O(N__83826),
            .I(shift_srl_28Z0Z_15));
    LocalMux I__15915 (
            .O(N__83823),
            .I(shift_srl_28Z0Z_15));
    LocalMux I__15914 (
            .O(N__83820),
            .I(shift_srl_28Z0Z_15));
    Odrv12 I__15913 (
            .O(N__83817),
            .I(shift_srl_28Z0Z_15));
    Odrv4 I__15912 (
            .O(N__83814),
            .I(shift_srl_28Z0Z_15));
    InMux I__15911 (
            .O(N__83803),
            .I(N__83797));
    InMux I__15910 (
            .O(N__83802),
            .I(N__83797));
    LocalMux I__15909 (
            .O(N__83797),
            .I(N__83787));
    InMux I__15908 (
            .O(N__83796),
            .I(N__83784));
    InMux I__15907 (
            .O(N__83795),
            .I(N__83779));
    InMux I__15906 (
            .O(N__83794),
            .I(N__83779));
    InMux I__15905 (
            .O(N__83793),
            .I(N__83776));
    InMux I__15904 (
            .O(N__83792),
            .I(N__83773));
    InMux I__15903 (
            .O(N__83791),
            .I(N__83770));
    InMux I__15902 (
            .O(N__83790),
            .I(N__83767));
    Span4Mux_h I__15901 (
            .O(N__83787),
            .I(N__83764));
    LocalMux I__15900 (
            .O(N__83784),
            .I(N__83761));
    LocalMux I__15899 (
            .O(N__83779),
            .I(N__83758));
    LocalMux I__15898 (
            .O(N__83776),
            .I(N__83755));
    LocalMux I__15897 (
            .O(N__83773),
            .I(N__83750));
    LocalMux I__15896 (
            .O(N__83770),
            .I(N__83750));
    LocalMux I__15895 (
            .O(N__83767),
            .I(N__83747));
    Span4Mux_h I__15894 (
            .O(N__83764),
            .I(N__83742));
    Span4Mux_h I__15893 (
            .O(N__83761),
            .I(N__83742));
    Span4Mux_h I__15892 (
            .O(N__83758),
            .I(N__83739));
    Span12Mux_v I__15891 (
            .O(N__83755),
            .I(N__83736));
    Span4Mux_v I__15890 (
            .O(N__83750),
            .I(N__83733));
    Odrv4 I__15889 (
            .O(N__83747),
            .I(shift_srl_24Z0Z_15));
    Odrv4 I__15888 (
            .O(N__83742),
            .I(shift_srl_24Z0Z_15));
    Odrv4 I__15887 (
            .O(N__83739),
            .I(shift_srl_24Z0Z_15));
    Odrv12 I__15886 (
            .O(N__83736),
            .I(shift_srl_24Z0Z_15));
    Odrv4 I__15885 (
            .O(N__83733),
            .I(shift_srl_24Z0Z_15));
    InMux I__15884 (
            .O(N__83722),
            .I(N__83713));
    InMux I__15883 (
            .O(N__83721),
            .I(N__83713));
    InMux I__15882 (
            .O(N__83720),
            .I(N__83708));
    InMux I__15881 (
            .O(N__83719),
            .I(N__83708));
    InMux I__15880 (
            .O(N__83718),
            .I(N__83705));
    LocalMux I__15879 (
            .O(N__83713),
            .I(N__83700));
    LocalMux I__15878 (
            .O(N__83708),
            .I(N__83700));
    LocalMux I__15877 (
            .O(N__83705),
            .I(N__83696));
    Span4Mux_v I__15876 (
            .O(N__83700),
            .I(N__83693));
    InMux I__15875 (
            .O(N__83699),
            .I(N__83690));
    Span4Mux_v I__15874 (
            .O(N__83696),
            .I(N__83685));
    Span4Mux_h I__15873 (
            .O(N__83693),
            .I(N__83685));
    LocalMux I__15872 (
            .O(N__83690),
            .I(shift_srl_30Z0Z_15));
    Odrv4 I__15871 (
            .O(N__83685),
            .I(shift_srl_30Z0Z_15));
    InMux I__15870 (
            .O(N__83680),
            .I(N__83677));
    LocalMux I__15869 (
            .O(N__83677),
            .I(N__83674));
    Span4Mux_v I__15868 (
            .O(N__83674),
            .I(N__83671));
    Sp12to4 I__15867 (
            .O(N__83671),
            .I(N__83668));
    Odrv12 I__15866 (
            .O(N__83668),
            .I(shift_srl_27_RNIP5TNZ0Z_15));
    CascadeMux I__15865 (
            .O(N__83665),
            .I(shift_srl_29_RNISHF41Z0Z_15_cascade_));
    CascadeMux I__15864 (
            .O(N__83662),
            .I(N__83658));
    InMux I__15863 (
            .O(N__83661),
            .I(N__83652));
    InMux I__15862 (
            .O(N__83658),
            .I(N__83652));
    InMux I__15861 (
            .O(N__83657),
            .I(N__83648));
    LocalMux I__15860 (
            .O(N__83652),
            .I(N__83645));
    InMux I__15859 (
            .O(N__83651),
            .I(N__83642));
    LocalMux I__15858 (
            .O(N__83648),
            .I(N__83639));
    Span4Mux_h I__15857 (
            .O(N__83645),
            .I(N__83636));
    LocalMux I__15856 (
            .O(N__83642),
            .I(shift_srl_31Z0Z_15));
    Odrv12 I__15855 (
            .O(N__83639),
            .I(shift_srl_31Z0Z_15));
    Odrv4 I__15854 (
            .O(N__83636),
            .I(shift_srl_31Z0Z_15));
    CascadeMux I__15853 (
            .O(N__83629),
            .I(rco_int_0_a2_0_a2_out_4_cascade_));
    IoInMux I__15852 (
            .O(N__83626),
            .I(N__83623));
    LocalMux I__15851 (
            .O(N__83623),
            .I(N__83620));
    Span4Mux_s2_v I__15850 (
            .O(N__83620),
            .I(N__83617));
    Sp12to4 I__15849 (
            .O(N__83617),
            .I(N__83613));
    InMux I__15848 (
            .O(N__83616),
            .I(N__83610));
    Span12Mux_s6_h I__15847 (
            .O(N__83613),
            .I(N__83606));
    LocalMux I__15846 (
            .O(N__83610),
            .I(N__83603));
    InMux I__15845 (
            .O(N__83609),
            .I(N__83600));
    Span12Mux_v I__15844 (
            .O(N__83606),
            .I(N__83597));
    Span4Mux_v I__15843 (
            .O(N__83603),
            .I(N__83594));
    LocalMux I__15842 (
            .O(N__83600),
            .I(N__83591));
    Odrv12 I__15841 (
            .O(N__83597),
            .I(rco_c_33));
    Odrv4 I__15840 (
            .O(N__83594),
            .I(rco_c_33));
    Odrv4 I__15839 (
            .O(N__83591),
            .I(rco_c_33));
    CascadeMux I__15838 (
            .O(N__83584),
            .I(N__83579));
    InMux I__15837 (
            .O(N__83583),
            .I(N__83573));
    InMux I__15836 (
            .O(N__83582),
            .I(N__83573));
    InMux I__15835 (
            .O(N__83579),
            .I(N__83568));
    InMux I__15834 (
            .O(N__83578),
            .I(N__83568));
    LocalMux I__15833 (
            .O(N__83573),
            .I(rco_int_0_a2_0_a2_out_4));
    LocalMux I__15832 (
            .O(N__83568),
            .I(rco_int_0_a2_0_a2_out_4));
    CascadeMux I__15831 (
            .O(N__83563),
            .I(N__83560));
    InMux I__15830 (
            .O(N__83560),
            .I(N__83554));
    InMux I__15829 (
            .O(N__83559),
            .I(N__83554));
    LocalMux I__15828 (
            .O(N__83554),
            .I(N__83551));
    Span4Mux_h I__15827 (
            .O(N__83551),
            .I(N__83548));
    Span4Mux_h I__15826 (
            .O(N__83548),
            .I(N__83545));
    Odrv4 I__15825 (
            .O(N__83545),
            .I(rco_int_0_a2_0_a2_s_0_0_35));
    IoInMux I__15824 (
            .O(N__83542),
            .I(N__83539));
    LocalMux I__15823 (
            .O(N__83539),
            .I(N__83536));
    IoSpan4Mux I__15822 (
            .O(N__83536),
            .I(N__83533));
    Sp12to4 I__15821 (
            .O(N__83533),
            .I(N__83530));
    Span12Mux_s9_h I__15820 (
            .O(N__83530),
            .I(N__83527));
    Span12Mux_v I__15819 (
            .O(N__83527),
            .I(N__83523));
    InMux I__15818 (
            .O(N__83526),
            .I(N__83520));
    Odrv12 I__15817 (
            .O(N__83523),
            .I(rco_c_36));
    LocalMux I__15816 (
            .O(N__83520),
            .I(rco_c_36));
    IoInMux I__15815 (
            .O(N__83515),
            .I(N__83512));
    LocalMux I__15814 (
            .O(N__83512),
            .I(N__83509));
    Span4Mux_s2_v I__15813 (
            .O(N__83509),
            .I(N__83506));
    Sp12to4 I__15812 (
            .O(N__83506),
            .I(N__83503));
    Span12Mux_s8_h I__15811 (
            .O(N__83503),
            .I(N__83500));
    Span12Mux_v I__15810 (
            .O(N__83500),
            .I(N__83496));
    InMux I__15809 (
            .O(N__83499),
            .I(N__83493));
    Odrv12 I__15808 (
            .O(N__83496),
            .I(rco_c_35));
    LocalMux I__15807 (
            .O(N__83493),
            .I(rco_c_35));
    InMux I__15806 (
            .O(N__83488),
            .I(N__83485));
    LocalMux I__15805 (
            .O(N__83485),
            .I(N__83481));
    InMux I__15804 (
            .O(N__83484),
            .I(N__83478));
    Span4Mux_v I__15803 (
            .O(N__83481),
            .I(N__83473));
    LocalMux I__15802 (
            .O(N__83478),
            .I(N__83473));
    Span4Mux_h I__15801 (
            .O(N__83473),
            .I(N__83470));
    Span4Mux_h I__15800 (
            .O(N__83470),
            .I(N__83465));
    InMux I__15799 (
            .O(N__83469),
            .I(N__83462));
    InMux I__15798 (
            .O(N__83468),
            .I(N__83459));
    Odrv4 I__15797 (
            .O(N__83465),
            .I(shift_srl_36Z0Z_15));
    LocalMux I__15796 (
            .O(N__83462),
            .I(shift_srl_36Z0Z_15));
    LocalMux I__15795 (
            .O(N__83459),
            .I(shift_srl_36Z0Z_15));
    InMux I__15794 (
            .O(N__83452),
            .I(N__83449));
    LocalMux I__15793 (
            .O(N__83449),
            .I(shift_srl_37Z0Z_14));
    CascadeMux I__15792 (
            .O(N__83446),
            .I(N__83442));
    InMux I__15791 (
            .O(N__83445),
            .I(N__83437));
    InMux I__15790 (
            .O(N__83442),
            .I(N__83437));
    LocalMux I__15789 (
            .O(N__83437),
            .I(N__83434));
    Span4Mux_h I__15788 (
            .O(N__83434),
            .I(N__83430));
    InMux I__15787 (
            .O(N__83433),
            .I(N__83427));
    Span4Mux_h I__15786 (
            .O(N__83430),
            .I(N__83424));
    LocalMux I__15785 (
            .O(N__83427),
            .I(shift_srl_37Z0Z_15));
    Odrv4 I__15784 (
            .O(N__83424),
            .I(shift_srl_37Z0Z_15));
    InMux I__15783 (
            .O(N__83419),
            .I(N__83416));
    LocalMux I__15782 (
            .O(N__83416),
            .I(shift_srl_37Z0Z_0));
    InMux I__15781 (
            .O(N__83413),
            .I(N__83410));
    LocalMux I__15780 (
            .O(N__83410),
            .I(shift_srl_37Z0Z_1));
    InMux I__15779 (
            .O(N__83407),
            .I(N__83404));
    LocalMux I__15778 (
            .O(N__83404),
            .I(shift_srl_37Z0Z_2));
    InMux I__15777 (
            .O(N__83401),
            .I(N__83398));
    LocalMux I__15776 (
            .O(N__83398),
            .I(shift_srl_37Z0Z_3));
    InMux I__15775 (
            .O(N__83395),
            .I(N__83392));
    LocalMux I__15774 (
            .O(N__83392),
            .I(shift_srl_37Z0Z_4));
    IoInMux I__15773 (
            .O(N__83389),
            .I(N__83386));
    LocalMux I__15772 (
            .O(N__83386),
            .I(N__83383));
    Span4Mux_s2_v I__15771 (
            .O(N__83383),
            .I(N__83380));
    Span4Mux_v I__15770 (
            .O(N__83380),
            .I(N__83377));
    Span4Mux_v I__15769 (
            .O(N__83377),
            .I(N__83374));
    Span4Mux_v I__15768 (
            .O(N__83374),
            .I(N__83371));
    Odrv4 I__15767 (
            .O(N__83371),
            .I(rco_c_32));
    InMux I__15766 (
            .O(N__83368),
            .I(N__83365));
    LocalMux I__15765 (
            .O(N__83365),
            .I(shift_srl_70Z0Z_5));
    InMux I__15764 (
            .O(N__83362),
            .I(N__83359));
    LocalMux I__15763 (
            .O(N__83359),
            .I(shift_srl_70Z0Z_6));
    InMux I__15762 (
            .O(N__83356),
            .I(N__83353));
    LocalMux I__15761 (
            .O(N__83353),
            .I(shift_srl_70Z0Z_7));
    InMux I__15760 (
            .O(N__83350),
            .I(N__83343));
    InMux I__15759 (
            .O(N__83349),
            .I(N__83343));
    InMux I__15758 (
            .O(N__83348),
            .I(N__83340));
    LocalMux I__15757 (
            .O(N__83343),
            .I(N__83335));
    LocalMux I__15756 (
            .O(N__83340),
            .I(N__83332));
    InMux I__15755 (
            .O(N__83339),
            .I(N__83329));
    InMux I__15754 (
            .O(N__83338),
            .I(N__83326));
    Span4Mux_v I__15753 (
            .O(N__83335),
            .I(N__83323));
    Span4Mux_h I__15752 (
            .O(N__83332),
            .I(N__83320));
    LocalMux I__15751 (
            .O(N__83329),
            .I(N__83313));
    LocalMux I__15750 (
            .O(N__83326),
            .I(N__83313));
    Span4Mux_h I__15749 (
            .O(N__83323),
            .I(N__83313));
    Span4Mux_h I__15748 (
            .O(N__83320),
            .I(N__83310));
    Odrv4 I__15747 (
            .O(N__83313),
            .I(shift_srl_34Z0Z_15));
    Odrv4 I__15746 (
            .O(N__83310),
            .I(shift_srl_34Z0Z_15));
    InMux I__15745 (
            .O(N__83305),
            .I(N__83302));
    LocalMux I__15744 (
            .O(N__83302),
            .I(shift_srl_34Z0Z_0));
    InMux I__15743 (
            .O(N__83299),
            .I(N__83296));
    LocalMux I__15742 (
            .O(N__83296),
            .I(shift_srl_34Z0Z_1));
    InMux I__15741 (
            .O(N__83293),
            .I(N__83290));
    LocalMux I__15740 (
            .O(N__83290),
            .I(shift_srl_34Z0Z_2));
    InMux I__15739 (
            .O(N__83287),
            .I(N__83284));
    LocalMux I__15738 (
            .O(N__83284),
            .I(shift_srl_34Z0Z_3));
    InMux I__15737 (
            .O(N__83281),
            .I(N__83278));
    LocalMux I__15736 (
            .O(N__83278),
            .I(shift_srl_67Z0Z_14));
    InMux I__15735 (
            .O(N__83275),
            .I(N__83272));
    LocalMux I__15734 (
            .O(N__83272),
            .I(shift_srl_67Z0Z_13));
    InMux I__15733 (
            .O(N__83269),
            .I(N__83266));
    LocalMux I__15732 (
            .O(N__83266),
            .I(shift_srl_67Z0Z_12));
    InMux I__15731 (
            .O(N__83263),
            .I(N__83260));
    LocalMux I__15730 (
            .O(N__83260),
            .I(N__83257));
    Odrv12 I__15729 (
            .O(N__83257),
            .I(shift_srl_67Z0Z_10));
    InMux I__15728 (
            .O(N__83254),
            .I(N__83251));
    LocalMux I__15727 (
            .O(N__83251),
            .I(shift_srl_67Z0Z_11));
    InMux I__15726 (
            .O(N__83248),
            .I(N__83245));
    LocalMux I__15725 (
            .O(N__83245),
            .I(shift_srl_70Z0Z_1));
    InMux I__15724 (
            .O(N__83242),
            .I(N__83239));
    LocalMux I__15723 (
            .O(N__83239),
            .I(shift_srl_70Z0Z_2));
    InMux I__15722 (
            .O(N__83236),
            .I(N__83233));
    LocalMux I__15721 (
            .O(N__83233),
            .I(shift_srl_70Z0Z_3));
    InMux I__15720 (
            .O(N__83230),
            .I(N__83227));
    LocalMux I__15719 (
            .O(N__83227),
            .I(shift_srl_70Z0Z_4));
    InMux I__15718 (
            .O(N__83224),
            .I(N__83221));
    LocalMux I__15717 (
            .O(N__83221),
            .I(shift_srl_71Z0Z_3));
    InMux I__15716 (
            .O(N__83218),
            .I(N__83215));
    LocalMux I__15715 (
            .O(N__83215),
            .I(shift_srl_71Z0Z_9));
    InMux I__15714 (
            .O(N__83212),
            .I(N__83209));
    LocalMux I__15713 (
            .O(N__83209),
            .I(shift_srl_71Z0Z_0));
    InMux I__15712 (
            .O(N__83206),
            .I(N__83203));
    LocalMux I__15711 (
            .O(N__83203),
            .I(shift_srl_71Z0Z_1));
    InMux I__15710 (
            .O(N__83200),
            .I(N__83197));
    LocalMux I__15709 (
            .O(N__83197),
            .I(shift_srl_71Z0Z_2));
    CascadeMux I__15708 (
            .O(N__83194),
            .I(shift_srl_68_RNIHDC4Z0Z_15_cascade_));
    InMux I__15707 (
            .O(N__83191),
            .I(N__83188));
    LocalMux I__15706 (
            .O(N__83188),
            .I(N__83185));
    Odrv12 I__15705 (
            .O(N__83185),
            .I(shift_srl_69_RNIBQRCZ0Z_15));
    CascadeMux I__15704 (
            .O(N__83182),
            .I(shift_srl_69_RNIBQRCZ0Z_15_cascade_));
    IoInMux I__15703 (
            .O(N__83179),
            .I(N__83176));
    LocalMux I__15702 (
            .O(N__83176),
            .I(N__83173));
    Span12Mux_s9_v I__15701 (
            .O(N__83173),
            .I(N__83170));
    Span12Mux_v I__15700 (
            .O(N__83170),
            .I(N__83167));
    Span12Mux_h I__15699 (
            .O(N__83167),
            .I(N__83164));
    Odrv12 I__15698 (
            .O(N__83164),
            .I(rco_c_69));
    InMux I__15697 (
            .O(N__83161),
            .I(N__83158));
    LocalMux I__15696 (
            .O(N__83158),
            .I(shift_srl_67Z0Z_0));
    InMux I__15695 (
            .O(N__83155),
            .I(N__83152));
    LocalMux I__15694 (
            .O(N__83152),
            .I(shift_srl_67Z0Z_1));
    InMux I__15693 (
            .O(N__83149),
            .I(N__83146));
    LocalMux I__15692 (
            .O(N__83146),
            .I(shift_srl_67Z0Z_2));
    InMux I__15691 (
            .O(N__83143),
            .I(N__83140));
    LocalMux I__15690 (
            .O(N__83140),
            .I(shift_srl_67Z0Z_3));
    InMux I__15689 (
            .O(N__83137),
            .I(N__83134));
    LocalMux I__15688 (
            .O(N__83134),
            .I(shift_srl_67Z0Z_4));
    InMux I__15687 (
            .O(N__83131),
            .I(N__83128));
    LocalMux I__15686 (
            .O(N__83128),
            .I(shift_srl_71Z0Z_10));
    InMux I__15685 (
            .O(N__83125),
            .I(N__83122));
    LocalMux I__15684 (
            .O(N__83122),
            .I(shift_srl_69Z0Z_4));
    InMux I__15683 (
            .O(N__83119),
            .I(N__83116));
    LocalMux I__15682 (
            .O(N__83116),
            .I(shift_srl_69Z0Z_5));
    InMux I__15681 (
            .O(N__83113),
            .I(N__83110));
    LocalMux I__15680 (
            .O(N__83110),
            .I(shift_srl_67Z0Z_9));
    InMux I__15679 (
            .O(N__83107),
            .I(N__83104));
    LocalMux I__15678 (
            .O(N__83104),
            .I(shift_srl_67Z0Z_8));
    InMux I__15677 (
            .O(N__83101),
            .I(N__83098));
    LocalMux I__15676 (
            .O(N__83098),
            .I(shift_srl_67Z0Z_7));
    InMux I__15675 (
            .O(N__83095),
            .I(N__83092));
    LocalMux I__15674 (
            .O(N__83092),
            .I(shift_srl_67Z0Z_6));
    InMux I__15673 (
            .O(N__83089),
            .I(N__83086));
    LocalMux I__15672 (
            .O(N__83086),
            .I(shift_srl_67Z0Z_5));
    IoInMux I__15671 (
            .O(N__83083),
            .I(N__83080));
    LocalMux I__15670 (
            .O(N__83080),
            .I(N__83077));
    Span4Mux_s1_v I__15669 (
            .O(N__83077),
            .I(N__83074));
    Sp12to4 I__15668 (
            .O(N__83074),
            .I(N__83071));
    Span12Mux_h I__15667 (
            .O(N__83071),
            .I(N__83068));
    Span12Mux_h I__15666 (
            .O(N__83068),
            .I(N__83065));
    Span12Mux_v I__15665 (
            .O(N__83065),
            .I(N__83062));
    Odrv12 I__15664 (
            .O(N__83062),
            .I(rco_c_67));
    IoInMux I__15663 (
            .O(N__83059),
            .I(N__83056));
    LocalMux I__15662 (
            .O(N__83056),
            .I(N__83053));
    IoSpan4Mux I__15661 (
            .O(N__83053),
            .I(N__83050));
    IoSpan4Mux I__15660 (
            .O(N__83050),
            .I(N__83047));
    Sp12to4 I__15659 (
            .O(N__83047),
            .I(N__83044));
    Span12Mux_v I__15658 (
            .O(N__83044),
            .I(N__83041));
    Span12Mux_h I__15657 (
            .O(N__83041),
            .I(N__83038));
    Odrv12 I__15656 (
            .O(N__83038),
            .I(rco_c_68));
    InMux I__15655 (
            .O(N__83035),
            .I(N__83032));
    LocalMux I__15654 (
            .O(N__83032),
            .I(shift_srl_78Z0Z_3));
    InMux I__15653 (
            .O(N__83029),
            .I(N__83026));
    LocalMux I__15652 (
            .O(N__83026),
            .I(shift_srl_78Z0Z_4));
    InMux I__15651 (
            .O(N__83023),
            .I(N__83020));
    LocalMux I__15650 (
            .O(N__83020),
            .I(shift_srl_78Z0Z_5));
    InMux I__15649 (
            .O(N__83017),
            .I(N__83014));
    LocalMux I__15648 (
            .O(N__83014),
            .I(shift_srl_78Z0Z_6));
    InMux I__15647 (
            .O(N__83011),
            .I(N__83008));
    LocalMux I__15646 (
            .O(N__83008),
            .I(shift_srl_78Z0Z_7));
    InMux I__15645 (
            .O(N__83005),
            .I(N__83002));
    LocalMux I__15644 (
            .O(N__83002),
            .I(shift_srl_69Z0Z_0));
    InMux I__15643 (
            .O(N__82999),
            .I(N__82996));
    LocalMux I__15642 (
            .O(N__82996),
            .I(shift_srl_69Z0Z_1));
    InMux I__15641 (
            .O(N__82993),
            .I(N__82990));
    LocalMux I__15640 (
            .O(N__82990),
            .I(shift_srl_69Z0Z_2));
    InMux I__15639 (
            .O(N__82987),
            .I(N__82984));
    LocalMux I__15638 (
            .O(N__82984),
            .I(shift_srl_69Z0Z_3));
    InMux I__15637 (
            .O(N__82981),
            .I(N__82978));
    LocalMux I__15636 (
            .O(N__82978),
            .I(shift_srl_78Z0Z_12));
    InMux I__15635 (
            .O(N__82975),
            .I(N__82972));
    LocalMux I__15634 (
            .O(N__82972),
            .I(shift_srl_78Z0Z_13));
    InMux I__15633 (
            .O(N__82969),
            .I(N__82966));
    LocalMux I__15632 (
            .O(N__82966),
            .I(shift_srl_78Z0Z_14));
    InMux I__15631 (
            .O(N__82963),
            .I(N__82960));
    LocalMux I__15630 (
            .O(N__82960),
            .I(shift_srl_78Z0Z_9));
    InMux I__15629 (
            .O(N__82957),
            .I(N__82954));
    LocalMux I__15628 (
            .O(N__82954),
            .I(shift_srl_78Z0Z_8));
    InMux I__15627 (
            .O(N__82951),
            .I(N__82948));
    LocalMux I__15626 (
            .O(N__82948),
            .I(shift_srl_78Z0Z_0));
    InMux I__15625 (
            .O(N__82945),
            .I(N__82942));
    LocalMux I__15624 (
            .O(N__82942),
            .I(shift_srl_78Z0Z_1));
    InMux I__15623 (
            .O(N__82939),
            .I(N__82936));
    LocalMux I__15622 (
            .O(N__82936),
            .I(shift_srl_78Z0Z_2));
    InMux I__15621 (
            .O(N__82933),
            .I(N__82930));
    LocalMux I__15620 (
            .O(N__82930),
            .I(shift_srl_80Z0Z_1));
    InMux I__15619 (
            .O(N__82927),
            .I(N__82924));
    LocalMux I__15618 (
            .O(N__82924),
            .I(shift_srl_80Z0Z_2));
    InMux I__15617 (
            .O(N__82921),
            .I(N__82918));
    LocalMux I__15616 (
            .O(N__82918),
            .I(shift_srl_80Z0Z_3));
    InMux I__15615 (
            .O(N__82915),
            .I(N__82912));
    LocalMux I__15614 (
            .O(N__82912),
            .I(shift_srl_80Z0Z_4));
    InMux I__15613 (
            .O(N__82909),
            .I(N__82906));
    LocalMux I__15612 (
            .O(N__82906),
            .I(shift_srl_80Z0Z_5));
    InMux I__15611 (
            .O(N__82903),
            .I(N__82900));
    LocalMux I__15610 (
            .O(N__82900),
            .I(shift_srl_80Z0Z_6));
    InMux I__15609 (
            .O(N__82897),
            .I(N__82894));
    LocalMux I__15608 (
            .O(N__82894),
            .I(shift_srl_80Z0Z_7));
    InMux I__15607 (
            .O(N__82891),
            .I(N__82888));
    LocalMux I__15606 (
            .O(N__82888),
            .I(shift_srl_78Z0Z_10));
    InMux I__15605 (
            .O(N__82885),
            .I(N__82882));
    LocalMux I__15604 (
            .O(N__82882),
            .I(shift_srl_78Z0Z_11));
    InMux I__15603 (
            .O(N__82879),
            .I(N__82876));
    LocalMux I__15602 (
            .O(N__82876),
            .I(shift_srl_189Z0Z_3));
    InMux I__15601 (
            .O(N__82873),
            .I(N__82870));
    LocalMux I__15600 (
            .O(N__82870),
            .I(shift_srl_189Z0Z_4));
    InMux I__15599 (
            .O(N__82867),
            .I(N__82864));
    LocalMux I__15598 (
            .O(N__82864),
            .I(shift_srl_189Z0Z_5));
    InMux I__15597 (
            .O(N__82861),
            .I(N__82858));
    LocalMux I__15596 (
            .O(N__82858),
            .I(shift_srl_189Z0Z_6));
    InMux I__15595 (
            .O(N__82855),
            .I(N__82852));
    LocalMux I__15594 (
            .O(N__82852),
            .I(N__82849));
    Odrv4 I__15593 (
            .O(N__82849),
            .I(shift_srl_189Z0Z_7));
    CEMux I__15592 (
            .O(N__82846),
            .I(N__82842));
    CEMux I__15591 (
            .O(N__82845),
            .I(N__82839));
    LocalMux I__15590 (
            .O(N__82842),
            .I(N__82836));
    LocalMux I__15589 (
            .O(N__82839),
            .I(N__82833));
    Span4Mux_v I__15588 (
            .O(N__82836),
            .I(N__82830));
    Odrv12 I__15587 (
            .O(N__82833),
            .I(clk_en_189));
    Odrv4 I__15586 (
            .O(N__82830),
            .I(clk_en_189));
    InMux I__15585 (
            .O(N__82825),
            .I(N__82822));
    LocalMux I__15584 (
            .O(N__82822),
            .I(N__82819));
    Odrv4 I__15583 (
            .O(N__82819),
            .I(shift_srl_188Z0Z_7));
    InMux I__15582 (
            .O(N__82816),
            .I(N__82813));
    LocalMux I__15581 (
            .O(N__82813),
            .I(shift_srl_188Z0Z_8));
    InMux I__15580 (
            .O(N__82810),
            .I(N__82807));
    LocalMux I__15579 (
            .O(N__82807),
            .I(shift_srl_188Z0Z_9));
    CEMux I__15578 (
            .O(N__82804),
            .I(N__82801));
    LocalMux I__15577 (
            .O(N__82801),
            .I(N__82798));
    Span4Mux_v I__15576 (
            .O(N__82798),
            .I(N__82793));
    CEMux I__15575 (
            .O(N__82797),
            .I(N__82790));
    CEMux I__15574 (
            .O(N__82796),
            .I(N__82787));
    Span4Mux_v I__15573 (
            .O(N__82793),
            .I(N__82782));
    LocalMux I__15572 (
            .O(N__82790),
            .I(N__82782));
    LocalMux I__15571 (
            .O(N__82787),
            .I(N__82779));
    Span4Mux_h I__15570 (
            .O(N__82782),
            .I(N__82776));
    Odrv12 I__15569 (
            .O(N__82779),
            .I(clk_en_188));
    Odrv4 I__15568 (
            .O(N__82776),
            .I(clk_en_188));
    InMux I__15567 (
            .O(N__82771),
            .I(N__82768));
    LocalMux I__15566 (
            .O(N__82768),
            .I(shift_srl_80Z0Z_0));
    InMux I__15565 (
            .O(N__82765),
            .I(N__82762));
    LocalMux I__15564 (
            .O(N__82762),
            .I(shift_srl_180Z0Z_13));
    InMux I__15563 (
            .O(N__82759),
            .I(N__82756));
    LocalMux I__15562 (
            .O(N__82756),
            .I(shift_srl_180Z0Z_14));
    InMux I__15561 (
            .O(N__82753),
            .I(N__82743));
    InMux I__15560 (
            .O(N__82752),
            .I(N__82743));
    InMux I__15559 (
            .O(N__82751),
            .I(N__82743));
    CascadeMux I__15558 (
            .O(N__82750),
            .I(N__82739));
    LocalMux I__15557 (
            .O(N__82743),
            .I(N__82736));
    InMux I__15556 (
            .O(N__82742),
            .I(N__82731));
    InMux I__15555 (
            .O(N__82739),
            .I(N__82731));
    Span4Mux_h I__15554 (
            .O(N__82736),
            .I(N__82725));
    LocalMux I__15553 (
            .O(N__82731),
            .I(N__82725));
    InMux I__15552 (
            .O(N__82730),
            .I(N__82722));
    Span4Mux_h I__15551 (
            .O(N__82725),
            .I(N__82719));
    LocalMux I__15550 (
            .O(N__82722),
            .I(shift_srl_180Z0Z_15));
    Odrv4 I__15549 (
            .O(N__82719),
            .I(shift_srl_180Z0Z_15));
    InMux I__15548 (
            .O(N__82714),
            .I(N__82711));
    LocalMux I__15547 (
            .O(N__82711),
            .I(shift_srl_180Z0Z_11));
    InMux I__15546 (
            .O(N__82708),
            .I(N__82705));
    LocalMux I__15545 (
            .O(N__82705),
            .I(shift_srl_180Z0Z_12));
    InMux I__15544 (
            .O(N__82702),
            .I(N__82699));
    LocalMux I__15543 (
            .O(N__82699),
            .I(shift_srl_180Z0Z_8));
    InMux I__15542 (
            .O(N__82696),
            .I(N__82693));
    LocalMux I__15541 (
            .O(N__82693),
            .I(shift_srl_180Z0Z_9));
    CEMux I__15540 (
            .O(N__82690),
            .I(N__82686));
    CEMux I__15539 (
            .O(N__82689),
            .I(N__82683));
    LocalMux I__15538 (
            .O(N__82686),
            .I(N__82680));
    LocalMux I__15537 (
            .O(N__82683),
            .I(N__82677));
    Span4Mux_h I__15536 (
            .O(N__82680),
            .I(N__82674));
    Span4Mux_h I__15535 (
            .O(N__82677),
            .I(N__82671));
    Odrv4 I__15534 (
            .O(N__82674),
            .I(clk_en_180));
    Odrv4 I__15533 (
            .O(N__82671),
            .I(clk_en_180));
    InMux I__15532 (
            .O(N__82666),
            .I(N__82663));
    LocalMux I__15531 (
            .O(N__82663),
            .I(shift_srl_189Z0Z_0));
    InMux I__15530 (
            .O(N__82660),
            .I(N__82657));
    LocalMux I__15529 (
            .O(N__82657),
            .I(shift_srl_189Z0Z_1));
    InMux I__15528 (
            .O(N__82654),
            .I(N__82651));
    LocalMux I__15527 (
            .O(N__82651),
            .I(shift_srl_189Z0Z_2));
    InMux I__15526 (
            .O(N__82648),
            .I(N__82645));
    LocalMux I__15525 (
            .O(N__82645),
            .I(shift_srl_177Z0Z_10));
    InMux I__15524 (
            .O(N__82642),
            .I(N__82639));
    LocalMux I__15523 (
            .O(N__82639),
            .I(shift_srl_177Z0Z_11));
    InMux I__15522 (
            .O(N__82636),
            .I(N__82633));
    LocalMux I__15521 (
            .O(N__82633),
            .I(shift_srl_177Z0Z_12));
    InMux I__15520 (
            .O(N__82630),
            .I(N__82627));
    LocalMux I__15519 (
            .O(N__82627),
            .I(shift_srl_177Z0Z_6));
    InMux I__15518 (
            .O(N__82624),
            .I(N__82621));
    LocalMux I__15517 (
            .O(N__82621),
            .I(shift_srl_177Z0Z_9));
    InMux I__15516 (
            .O(N__82618),
            .I(N__82615));
    LocalMux I__15515 (
            .O(N__82615),
            .I(shift_srl_177Z0Z_7));
    InMux I__15514 (
            .O(N__82612),
            .I(N__82609));
    LocalMux I__15513 (
            .O(N__82609),
            .I(shift_srl_177Z0Z_8));
    CEMux I__15512 (
            .O(N__82606),
            .I(N__82603));
    LocalMux I__15511 (
            .O(N__82603),
            .I(N__82600));
    Span4Mux_h I__15510 (
            .O(N__82600),
            .I(N__82595));
    CEMux I__15509 (
            .O(N__82599),
            .I(N__82592));
    CEMux I__15508 (
            .O(N__82598),
            .I(N__82589));
    Odrv4 I__15507 (
            .O(N__82595),
            .I(clk_en_177));
    LocalMux I__15506 (
            .O(N__82592),
            .I(clk_en_177));
    LocalMux I__15505 (
            .O(N__82589),
            .I(clk_en_177));
    InMux I__15504 (
            .O(N__82582),
            .I(N__82579));
    LocalMux I__15503 (
            .O(N__82579),
            .I(shift_srl_180Z0Z_10));
    InMux I__15502 (
            .O(N__82576),
            .I(N__82573));
    LocalMux I__15501 (
            .O(N__82573),
            .I(shift_srl_180Z0Z_4));
    InMux I__15500 (
            .O(N__82570),
            .I(N__82567));
    LocalMux I__15499 (
            .O(N__82567),
            .I(shift_srl_180Z0Z_5));
    InMux I__15498 (
            .O(N__82564),
            .I(N__82561));
    LocalMux I__15497 (
            .O(N__82561),
            .I(shift_srl_169Z0Z_0));
    InMux I__15496 (
            .O(N__82558),
            .I(N__82555));
    LocalMux I__15495 (
            .O(N__82555),
            .I(N__82552));
    Odrv4 I__15494 (
            .O(N__82552),
            .I(shift_srl_169Z0Z_1));
    CEMux I__15493 (
            .O(N__82549),
            .I(N__82546));
    LocalMux I__15492 (
            .O(N__82546),
            .I(N__82541));
    CEMux I__15491 (
            .O(N__82545),
            .I(N__82538));
    CEMux I__15490 (
            .O(N__82544),
            .I(N__82535));
    Odrv4 I__15489 (
            .O(N__82541),
            .I(clk_en_169));
    LocalMux I__15488 (
            .O(N__82538),
            .I(clk_en_169));
    LocalMux I__15487 (
            .O(N__82535),
            .I(clk_en_169));
    InMux I__15486 (
            .O(N__82528),
            .I(N__82525));
    LocalMux I__15485 (
            .O(N__82525),
            .I(shift_srl_170Z0Z_10));
    InMux I__15484 (
            .O(N__82522),
            .I(N__82519));
    LocalMux I__15483 (
            .O(N__82519),
            .I(shift_srl_170Z0Z_11));
    InMux I__15482 (
            .O(N__82516),
            .I(N__82513));
    LocalMux I__15481 (
            .O(N__82513),
            .I(shift_srl_170Z0Z_12));
    InMux I__15480 (
            .O(N__82510),
            .I(N__82507));
    LocalMux I__15479 (
            .O(N__82507),
            .I(shift_srl_170Z0Z_13));
    InMux I__15478 (
            .O(N__82504),
            .I(N__82501));
    LocalMux I__15477 (
            .O(N__82501),
            .I(shift_srl_170Z0Z_14));
    InMux I__15476 (
            .O(N__82498),
            .I(N__82495));
    LocalMux I__15475 (
            .O(N__82495),
            .I(shift_srl_170Z0Z_9));
    InMux I__15474 (
            .O(N__82492),
            .I(N__82489));
    LocalMux I__15473 (
            .O(N__82489),
            .I(shift_srl_170Z0Z_7));
    InMux I__15472 (
            .O(N__82486),
            .I(N__82483));
    LocalMux I__15471 (
            .O(N__82483),
            .I(shift_srl_170Z0Z_8));
    CEMux I__15470 (
            .O(N__82480),
            .I(N__82476));
    CEMux I__15469 (
            .O(N__82479),
            .I(N__82473));
    LocalMux I__15468 (
            .O(N__82476),
            .I(clk_en_170));
    LocalMux I__15467 (
            .O(N__82473),
            .I(clk_en_170));
    InMux I__15466 (
            .O(N__82468),
            .I(N__82465));
    LocalMux I__15465 (
            .O(N__82465),
            .I(shift_srl_169Z0Z_13));
    InMux I__15464 (
            .O(N__82462),
            .I(N__82459));
    LocalMux I__15463 (
            .O(N__82459),
            .I(shift_srl_169Z0Z_14));
    InMux I__15462 (
            .O(N__82456),
            .I(N__82453));
    LocalMux I__15461 (
            .O(N__82453),
            .I(shift_srl_169Z0Z_9));
    InMux I__15460 (
            .O(N__82450),
            .I(N__82447));
    LocalMux I__15459 (
            .O(N__82447),
            .I(N__82444));
    Odrv4 I__15458 (
            .O(N__82444),
            .I(shift_srl_169Z0Z_7));
    InMux I__15457 (
            .O(N__82441),
            .I(N__82438));
    LocalMux I__15456 (
            .O(N__82438),
            .I(shift_srl_169Z0Z_8));
    InMux I__15455 (
            .O(N__82435),
            .I(N__82432));
    LocalMux I__15454 (
            .O(N__82432),
            .I(N__82429));
    Span4Mux_s3_v I__15453 (
            .O(N__82429),
            .I(N__82422));
    InMux I__15452 (
            .O(N__82428),
            .I(N__82419));
    CascadeMux I__15451 (
            .O(N__82427),
            .I(N__82416));
    CascadeMux I__15450 (
            .O(N__82426),
            .I(N__82412));
    CascadeMux I__15449 (
            .O(N__82425),
            .I(N__82409));
    Sp12to4 I__15448 (
            .O(N__82422),
            .I(N__82404));
    LocalMux I__15447 (
            .O(N__82419),
            .I(N__82404));
    InMux I__15446 (
            .O(N__82416),
            .I(N__82401));
    InMux I__15445 (
            .O(N__82415),
            .I(N__82396));
    InMux I__15444 (
            .O(N__82412),
            .I(N__82396));
    InMux I__15443 (
            .O(N__82409),
            .I(N__82393));
    Span12Mux_h I__15442 (
            .O(N__82404),
            .I(N__82390));
    LocalMux I__15441 (
            .O(N__82401),
            .I(N__82387));
    LocalMux I__15440 (
            .O(N__82396),
            .I(N__82382));
    LocalMux I__15439 (
            .O(N__82393),
            .I(N__82382));
    Span12Mux_v I__15438 (
            .O(N__82390),
            .I(N__82379));
    Span4Mux_v I__15437 (
            .O(N__82387),
            .I(N__82376));
    Span4Mux_h I__15436 (
            .O(N__82382),
            .I(N__82373));
    Odrv12 I__15435 (
            .O(N__82379),
            .I(shift_srl_164_RNIBMOLZ0Z_15));
    Odrv4 I__15434 (
            .O(N__82376),
            .I(shift_srl_164_RNIBMOLZ0Z_15));
    Odrv4 I__15433 (
            .O(N__82373),
            .I(shift_srl_164_RNIBMOLZ0Z_15));
    CEMux I__15432 (
            .O(N__82366),
            .I(N__82363));
    LocalMux I__15431 (
            .O(N__82363),
            .I(N__82359));
    CEMux I__15430 (
            .O(N__82362),
            .I(N__82356));
    Span4Mux_v I__15429 (
            .O(N__82359),
            .I(N__82353));
    LocalMux I__15428 (
            .O(N__82356),
            .I(N__82350));
    Span4Mux_v I__15427 (
            .O(N__82353),
            .I(N__82345));
    Span4Mux_v I__15426 (
            .O(N__82350),
            .I(N__82345));
    Odrv4 I__15425 (
            .O(N__82345),
            .I(clk_en_167));
    InMux I__15424 (
            .O(N__82342),
            .I(N__82336));
    CascadeMux I__15423 (
            .O(N__82341),
            .I(N__82331));
    InMux I__15422 (
            .O(N__82340),
            .I(N__82328));
    InMux I__15421 (
            .O(N__82339),
            .I(N__82324));
    LocalMux I__15420 (
            .O(N__82336),
            .I(N__82321));
    InMux I__15419 (
            .O(N__82335),
            .I(N__82316));
    InMux I__15418 (
            .O(N__82334),
            .I(N__82316));
    InMux I__15417 (
            .O(N__82331),
            .I(N__82313));
    LocalMux I__15416 (
            .O(N__82328),
            .I(N__82309));
    InMux I__15415 (
            .O(N__82327),
            .I(N__82306));
    LocalMux I__15414 (
            .O(N__82324),
            .I(N__82303));
    Span4Mux_v I__15413 (
            .O(N__82321),
            .I(N__82296));
    LocalMux I__15412 (
            .O(N__82316),
            .I(N__82296));
    LocalMux I__15411 (
            .O(N__82313),
            .I(N__82296));
    InMux I__15410 (
            .O(N__82312),
            .I(N__82289));
    Span4Mux_v I__15409 (
            .O(N__82309),
            .I(N__82285));
    LocalMux I__15408 (
            .O(N__82306),
            .I(N__82282));
    Span4Mux_h I__15407 (
            .O(N__82303),
            .I(N__82279));
    Span4Mux_v I__15406 (
            .O(N__82296),
            .I(N__82276));
    InMux I__15405 (
            .O(N__82295),
            .I(N__82267));
    InMux I__15404 (
            .O(N__82294),
            .I(N__82267));
    InMux I__15403 (
            .O(N__82293),
            .I(N__82267));
    InMux I__15402 (
            .O(N__82292),
            .I(N__82267));
    LocalMux I__15401 (
            .O(N__82289),
            .I(N__82264));
    InMux I__15400 (
            .O(N__82288),
            .I(N__82261));
    Span4Mux_h I__15399 (
            .O(N__82285),
            .I(N__82256));
    Span4Mux_v I__15398 (
            .O(N__82282),
            .I(N__82256));
    Span4Mux_v I__15397 (
            .O(N__82279),
            .I(N__82253));
    Span4Mux_h I__15396 (
            .O(N__82276),
            .I(N__82250));
    LocalMux I__15395 (
            .O(N__82267),
            .I(N__82245));
    Span4Mux_v I__15394 (
            .O(N__82264),
            .I(N__82245));
    LocalMux I__15393 (
            .O(N__82261),
            .I(N__82242));
    Sp12to4 I__15392 (
            .O(N__82256),
            .I(N__82237));
    Sp12to4 I__15391 (
            .O(N__82253),
            .I(N__82237));
    Span4Mux_h I__15390 (
            .O(N__82250),
            .I(N__82234));
    Span4Mux_h I__15389 (
            .O(N__82245),
            .I(N__82231));
    Odrv12 I__15388 (
            .O(N__82242),
            .I(rco_int_0_a2_0_a2_0_153));
    Odrv12 I__15387 (
            .O(N__82237),
            .I(rco_int_0_a2_0_a2_0_153));
    Odrv4 I__15386 (
            .O(N__82234),
            .I(rco_int_0_a2_0_a2_0_153));
    Odrv4 I__15385 (
            .O(N__82231),
            .I(rco_int_0_a2_0_a2_0_153));
    InMux I__15384 (
            .O(N__82222),
            .I(N__82217));
    IoInMux I__15383 (
            .O(N__82221),
            .I(N__82213));
    InMux I__15382 (
            .O(N__82220),
            .I(N__82209));
    LocalMux I__15381 (
            .O(N__82217),
            .I(N__82206));
    InMux I__15380 (
            .O(N__82216),
            .I(N__82203));
    LocalMux I__15379 (
            .O(N__82213),
            .I(N__82199));
    CascadeMux I__15378 (
            .O(N__82212),
            .I(N__82195));
    LocalMux I__15377 (
            .O(N__82209),
            .I(N__82191));
    Span4Mux_h I__15376 (
            .O(N__82206),
            .I(N__82186));
    LocalMux I__15375 (
            .O(N__82203),
            .I(N__82186));
    InMux I__15374 (
            .O(N__82202),
            .I(N__82182));
    Span4Mux_s2_v I__15373 (
            .O(N__82199),
            .I(N__82179));
    InMux I__15372 (
            .O(N__82198),
            .I(N__82176));
    InMux I__15371 (
            .O(N__82195),
            .I(N__82170));
    InMux I__15370 (
            .O(N__82194),
            .I(N__82170));
    Span4Mux_v I__15369 (
            .O(N__82191),
            .I(N__82167));
    Span4Mux_v I__15368 (
            .O(N__82186),
            .I(N__82164));
    InMux I__15367 (
            .O(N__82185),
            .I(N__82161));
    LocalMux I__15366 (
            .O(N__82182),
            .I(N__82157));
    Span4Mux_h I__15365 (
            .O(N__82179),
            .I(N__82152));
    LocalMux I__15364 (
            .O(N__82176),
            .I(N__82152));
    InMux I__15363 (
            .O(N__82175),
            .I(N__82149));
    LocalMux I__15362 (
            .O(N__82170),
            .I(N__82142));
    Span4Mux_v I__15361 (
            .O(N__82167),
            .I(N__82139));
    Span4Mux_v I__15360 (
            .O(N__82164),
            .I(N__82134));
    LocalMux I__15359 (
            .O(N__82161),
            .I(N__82134));
    InMux I__15358 (
            .O(N__82160),
            .I(N__82131));
    Span4Mux_v I__15357 (
            .O(N__82157),
            .I(N__82128));
    Sp12to4 I__15356 (
            .O(N__82152),
            .I(N__82125));
    LocalMux I__15355 (
            .O(N__82149),
            .I(N__82122));
    InMux I__15354 (
            .O(N__82148),
            .I(N__82113));
    InMux I__15353 (
            .O(N__82147),
            .I(N__82113));
    InMux I__15352 (
            .O(N__82146),
            .I(N__82113));
    InMux I__15351 (
            .O(N__82145),
            .I(N__82113));
    Span4Mux_h I__15350 (
            .O(N__82142),
            .I(N__82110));
    Span4Mux_h I__15349 (
            .O(N__82139),
            .I(N__82105));
    Span4Mux_h I__15348 (
            .O(N__82134),
            .I(N__82105));
    LocalMux I__15347 (
            .O(N__82131),
            .I(N__82102));
    Span4Mux_h I__15346 (
            .O(N__82128),
            .I(N__82099));
    Span12Mux_v I__15345 (
            .O(N__82125),
            .I(N__82096));
    Span12Mux_v I__15344 (
            .O(N__82122),
            .I(N__82091));
    LocalMux I__15343 (
            .O(N__82113),
            .I(N__82091));
    Span4Mux_h I__15342 (
            .O(N__82110),
            .I(N__82086));
    Span4Mux_v I__15341 (
            .O(N__82105),
            .I(N__82086));
    Span12Mux_h I__15340 (
            .O(N__82102),
            .I(N__82083));
    Span4Mux_v I__15339 (
            .O(N__82099),
            .I(N__82080));
    Odrv12 I__15338 (
            .O(N__82096),
            .I(rco_c_145));
    Odrv12 I__15337 (
            .O(N__82091),
            .I(rco_c_145));
    Odrv4 I__15336 (
            .O(N__82086),
            .I(rco_c_145));
    Odrv12 I__15335 (
            .O(N__82083),
            .I(rco_c_145));
    Odrv4 I__15334 (
            .O(N__82080),
            .I(rco_c_145));
    CascadeMux I__15333 (
            .O(N__82069),
            .I(clk_en_163_cascade_));
    InMux I__15332 (
            .O(N__82066),
            .I(N__82063));
    LocalMux I__15331 (
            .O(N__82063),
            .I(shift_srl_169Z0Z_5));
    InMux I__15330 (
            .O(N__82060),
            .I(N__82057));
    LocalMux I__15329 (
            .O(N__82057),
            .I(shift_srl_169Z0Z_6));
    InMux I__15328 (
            .O(N__82054),
            .I(N__82051));
    LocalMux I__15327 (
            .O(N__82051),
            .I(N__82048));
    Odrv4 I__15326 (
            .O(N__82048),
            .I(shift_srl_39Z0Z_7));
    InMux I__15325 (
            .O(N__82045),
            .I(N__82042));
    LocalMux I__15324 (
            .O(N__82042),
            .I(N__82039));
    Span4Mux_v I__15323 (
            .O(N__82039),
            .I(N__82036));
    Span4Mux_h I__15322 (
            .O(N__82036),
            .I(N__82033));
    Odrv4 I__15321 (
            .O(N__82033),
            .I(shift_srl_39Z0Z_8));
    CEMux I__15320 (
            .O(N__82030),
            .I(N__82027));
    LocalMux I__15319 (
            .O(N__82027),
            .I(N__82024));
    Span4Mux_v I__15318 (
            .O(N__82024),
            .I(N__82020));
    CEMux I__15317 (
            .O(N__82023),
            .I(N__82017));
    Span4Mux_h I__15316 (
            .O(N__82020),
            .I(N__82013));
    LocalMux I__15315 (
            .O(N__82017),
            .I(N__82010));
    CEMux I__15314 (
            .O(N__82016),
            .I(N__82007));
    Odrv4 I__15313 (
            .O(N__82013),
            .I(clk_en_39));
    Odrv4 I__15312 (
            .O(N__82010),
            .I(clk_en_39));
    LocalMux I__15311 (
            .O(N__82007),
            .I(clk_en_39));
    InMux I__15310 (
            .O(N__82000),
            .I(N__81997));
    LocalMux I__15309 (
            .O(N__81997),
            .I(shift_srl_169Z0Z_10));
    InMux I__15308 (
            .O(N__81994),
            .I(N__81991));
    LocalMux I__15307 (
            .O(N__81991),
            .I(N__81988));
    Odrv4 I__15306 (
            .O(N__81988),
            .I(shift_srl_169Z0Z_11));
    InMux I__15305 (
            .O(N__81985),
            .I(N__81982));
    LocalMux I__15304 (
            .O(N__81982),
            .I(N__81979));
    Odrv4 I__15303 (
            .O(N__81979),
            .I(shift_srl_169Z0Z_2));
    InMux I__15302 (
            .O(N__81976),
            .I(N__81973));
    LocalMux I__15301 (
            .O(N__81973),
            .I(N__81970));
    Odrv4 I__15300 (
            .O(N__81970),
            .I(shift_srl_169Z0Z_3));
    InMux I__15299 (
            .O(N__81967),
            .I(N__81964));
    LocalMux I__15298 (
            .O(N__81964),
            .I(N__81961));
    Odrv4 I__15297 (
            .O(N__81961),
            .I(shift_srl_169Z0Z_12));
    InMux I__15296 (
            .O(N__81958),
            .I(N__81955));
    LocalMux I__15295 (
            .O(N__81955),
            .I(shift_srl_39Z0Z_0));
    InMux I__15294 (
            .O(N__81952),
            .I(N__81949));
    LocalMux I__15293 (
            .O(N__81949),
            .I(shift_srl_39Z0Z_1));
    InMux I__15292 (
            .O(N__81946),
            .I(N__81943));
    LocalMux I__15291 (
            .O(N__81943),
            .I(shift_srl_39Z0Z_2));
    InMux I__15290 (
            .O(N__81940),
            .I(N__81937));
    LocalMux I__15289 (
            .O(N__81937),
            .I(shift_srl_39Z0Z_3));
    InMux I__15288 (
            .O(N__81934),
            .I(N__81931));
    LocalMux I__15287 (
            .O(N__81931),
            .I(shift_srl_39Z0Z_4));
    InMux I__15286 (
            .O(N__81928),
            .I(N__81925));
    LocalMux I__15285 (
            .O(N__81925),
            .I(shift_srl_39Z0Z_5));
    InMux I__15284 (
            .O(N__81922),
            .I(N__81919));
    LocalMux I__15283 (
            .O(N__81919),
            .I(shift_srl_39Z0Z_6));
    InMux I__15282 (
            .O(N__81916),
            .I(N__81913));
    LocalMux I__15281 (
            .O(N__81913),
            .I(shift_srl_169Z0Z_4));
    CascadeMux I__15280 (
            .O(N__81910),
            .I(N__81907));
    InMux I__15279 (
            .O(N__81907),
            .I(N__81904));
    LocalMux I__15278 (
            .O(N__81904),
            .I(N__81899));
    InMux I__15277 (
            .O(N__81903),
            .I(N__81896));
    InMux I__15276 (
            .O(N__81902),
            .I(N__81893));
    Span4Mux_h I__15275 (
            .O(N__81899),
            .I(N__81890));
    LocalMux I__15274 (
            .O(N__81896),
            .I(N__81887));
    LocalMux I__15273 (
            .O(N__81893),
            .I(N__81882));
    Span4Mux_h I__15272 (
            .O(N__81890),
            .I(N__81882));
    Odrv12 I__15271 (
            .O(N__81887),
            .I(shift_srl_35Z0Z_15));
    Odrv4 I__15270 (
            .O(N__81882),
            .I(shift_srl_35Z0Z_15));
    InMux I__15269 (
            .O(N__81877),
            .I(N__81874));
    LocalMux I__15268 (
            .O(N__81874),
            .I(shift_srl_35Z0Z_0));
    InMux I__15267 (
            .O(N__81871),
            .I(N__81868));
    LocalMux I__15266 (
            .O(N__81868),
            .I(shift_srl_35Z0Z_1));
    InMux I__15265 (
            .O(N__81865),
            .I(N__81862));
    LocalMux I__15264 (
            .O(N__81862),
            .I(shift_srl_35Z0Z_2));
    InMux I__15263 (
            .O(N__81859),
            .I(N__81856));
    LocalMux I__15262 (
            .O(N__81856),
            .I(shift_srl_35Z0Z_3));
    InMux I__15261 (
            .O(N__81853),
            .I(N__81850));
    LocalMux I__15260 (
            .O(N__81850),
            .I(shift_srl_35Z0Z_4));
    InMux I__15259 (
            .O(N__81847),
            .I(N__81844));
    LocalMux I__15258 (
            .O(N__81844),
            .I(shift_srl_35Z0Z_5));
    InMux I__15257 (
            .O(N__81841),
            .I(N__81838));
    LocalMux I__15256 (
            .O(N__81838),
            .I(shift_srl_35Z0Z_6));
    InMux I__15255 (
            .O(N__81835),
            .I(N__81832));
    LocalMux I__15254 (
            .O(N__81832),
            .I(N__81829));
    Odrv4 I__15253 (
            .O(N__81829),
            .I(shift_srl_35Z0Z_7));
    CEMux I__15252 (
            .O(N__81826),
            .I(N__81823));
    LocalMux I__15251 (
            .O(N__81823),
            .I(N__81819));
    CEMux I__15250 (
            .O(N__81822),
            .I(N__81816));
    Sp12to4 I__15249 (
            .O(N__81819),
            .I(N__81811));
    LocalMux I__15248 (
            .O(N__81816),
            .I(N__81811));
    Odrv12 I__15247 (
            .O(N__81811),
            .I(clk_en_35));
    InMux I__15246 (
            .O(N__81808),
            .I(N__81805));
    LocalMux I__15245 (
            .O(N__81805),
            .I(N__81801));
    InMux I__15244 (
            .O(N__81804),
            .I(N__81798));
    Span4Mux_v I__15243 (
            .O(N__81801),
            .I(N__81794));
    LocalMux I__15242 (
            .O(N__81798),
            .I(N__81791));
    CascadeMux I__15241 (
            .O(N__81797),
            .I(N__81788));
    Span4Mux_h I__15240 (
            .O(N__81794),
            .I(N__81783));
    Span4Mux_v I__15239 (
            .O(N__81791),
            .I(N__81783));
    InMux I__15238 (
            .O(N__81788),
            .I(N__81780));
    Odrv4 I__15237 (
            .O(N__81783),
            .I(shift_srl_39Z0Z_15));
    LocalMux I__15236 (
            .O(N__81780),
            .I(shift_srl_39Z0Z_15));
    InMux I__15235 (
            .O(N__81775),
            .I(N__81772));
    LocalMux I__15234 (
            .O(N__81772),
            .I(shift_srl_35Z0Z_9));
    InMux I__15233 (
            .O(N__81769),
            .I(N__81766));
    LocalMux I__15232 (
            .O(N__81766),
            .I(shift_srl_35Z0Z_8));
    InMux I__15231 (
            .O(N__81763),
            .I(N__81760));
    LocalMux I__15230 (
            .O(N__81760),
            .I(shift_srl_34Z0Z_14));
    InMux I__15229 (
            .O(N__81757),
            .I(N__81754));
    LocalMux I__15228 (
            .O(N__81754),
            .I(shift_srl_34Z0Z_13));
    InMux I__15227 (
            .O(N__81751),
            .I(N__81748));
    LocalMux I__15226 (
            .O(N__81748),
            .I(shift_srl_34Z0Z_12));
    InMux I__15225 (
            .O(N__81745),
            .I(N__81742));
    LocalMux I__15224 (
            .O(N__81742),
            .I(shift_srl_34Z0Z_11));
    InMux I__15223 (
            .O(N__81739),
            .I(N__81736));
    LocalMux I__15222 (
            .O(N__81736),
            .I(shift_srl_34Z0Z_10));
    InMux I__15221 (
            .O(N__81733),
            .I(N__81730));
    LocalMux I__15220 (
            .O(N__81730),
            .I(shift_srl_34Z0Z_9));
    InMux I__15219 (
            .O(N__81727),
            .I(N__81724));
    LocalMux I__15218 (
            .O(N__81724),
            .I(shift_srl_66Z0Z_14));
    InMux I__15217 (
            .O(N__81721),
            .I(N__81718));
    LocalMux I__15216 (
            .O(N__81718),
            .I(N__81714));
    InMux I__15215 (
            .O(N__81717),
            .I(N__81711));
    Span4Mux_h I__15214 (
            .O(N__81714),
            .I(N__81708));
    LocalMux I__15213 (
            .O(N__81711),
            .I(shift_srl_66Z0Z_15));
    Odrv4 I__15212 (
            .O(N__81708),
            .I(shift_srl_66Z0Z_15));
    InMux I__15211 (
            .O(N__81703),
            .I(N__81700));
    LocalMux I__15210 (
            .O(N__81700),
            .I(shift_srl_66Z0Z_9));
    InMux I__15209 (
            .O(N__81697),
            .I(N__81694));
    LocalMux I__15208 (
            .O(N__81694),
            .I(shift_srl_66Z0Z_7));
    InMux I__15207 (
            .O(N__81691),
            .I(N__81688));
    LocalMux I__15206 (
            .O(N__81688),
            .I(shift_srl_66Z0Z_8));
    CEMux I__15205 (
            .O(N__81685),
            .I(N__81682));
    LocalMux I__15204 (
            .O(N__81682),
            .I(N__81678));
    CEMux I__15203 (
            .O(N__81681),
            .I(N__81675));
    Odrv12 I__15202 (
            .O(N__81678),
            .I(clk_en_66));
    LocalMux I__15201 (
            .O(N__81675),
            .I(clk_en_66));
    InMux I__15200 (
            .O(N__81670),
            .I(N__81667));
    LocalMux I__15199 (
            .O(N__81667),
            .I(shift_srl_35Z0Z_10));
    InMux I__15198 (
            .O(N__81664),
            .I(N__81661));
    LocalMux I__15197 (
            .O(N__81661),
            .I(shift_srl_35Z0Z_11));
    InMux I__15196 (
            .O(N__81658),
            .I(N__81655));
    LocalMux I__15195 (
            .O(N__81655),
            .I(shift_srl_35Z0Z_12));
    InMux I__15194 (
            .O(N__81652),
            .I(N__81649));
    LocalMux I__15193 (
            .O(N__81649),
            .I(shift_srl_35Z0Z_13));
    InMux I__15192 (
            .O(N__81646),
            .I(N__81643));
    LocalMux I__15191 (
            .O(N__81643),
            .I(shift_srl_35Z0Z_14));
    InMux I__15190 (
            .O(N__81640),
            .I(N__81637));
    LocalMux I__15189 (
            .O(N__81637),
            .I(shift_srl_66Z0Z_3));
    InMux I__15188 (
            .O(N__81634),
            .I(N__81631));
    LocalMux I__15187 (
            .O(N__81631),
            .I(shift_srl_66Z0Z_4));
    InMux I__15186 (
            .O(N__81628),
            .I(N__81625));
    LocalMux I__15185 (
            .O(N__81625),
            .I(shift_srl_66Z0Z_5));
    InMux I__15184 (
            .O(N__81622),
            .I(N__81619));
    LocalMux I__15183 (
            .O(N__81619),
            .I(shift_srl_66Z0Z_6));
    InMux I__15182 (
            .O(N__81616),
            .I(N__81613));
    LocalMux I__15181 (
            .O(N__81613),
            .I(shift_srl_66Z0Z_10));
    InMux I__15180 (
            .O(N__81610),
            .I(N__81607));
    LocalMux I__15179 (
            .O(N__81607),
            .I(shift_srl_66Z0Z_11));
    InMux I__15178 (
            .O(N__81604),
            .I(N__81601));
    LocalMux I__15177 (
            .O(N__81601),
            .I(shift_srl_66Z0Z_12));
    InMux I__15176 (
            .O(N__81598),
            .I(N__81595));
    LocalMux I__15175 (
            .O(N__81595),
            .I(shift_srl_66Z0Z_13));
    CascadeMux I__15174 (
            .O(N__81592),
            .I(shift_srl_65_RNILFDF1Z0Z_15_cascade_));
    InMux I__15173 (
            .O(N__81589),
            .I(N__81583));
    InMux I__15172 (
            .O(N__81588),
            .I(N__81580));
    CascadeMux I__15171 (
            .O(N__81587),
            .I(N__81577));
    InMux I__15170 (
            .O(N__81586),
            .I(N__81574));
    LocalMux I__15169 (
            .O(N__81583),
            .I(N__81571));
    LocalMux I__15168 (
            .O(N__81580),
            .I(N__81568));
    InMux I__15167 (
            .O(N__81577),
            .I(N__81565));
    LocalMux I__15166 (
            .O(N__81574),
            .I(N__81558));
    Span4Mux_h I__15165 (
            .O(N__81571),
            .I(N__81558));
    Span4Mux_v I__15164 (
            .O(N__81568),
            .I(N__81558));
    LocalMux I__15163 (
            .O(N__81565),
            .I(shift_srl_59Z0Z_15));
    Odrv4 I__15162 (
            .O(N__81558),
            .I(shift_srl_59Z0Z_15));
    InMux I__15161 (
            .O(N__81553),
            .I(N__81544));
    InMux I__15160 (
            .O(N__81552),
            .I(N__81544));
    InMux I__15159 (
            .O(N__81551),
            .I(N__81541));
    InMux I__15158 (
            .O(N__81550),
            .I(N__81536));
    InMux I__15157 (
            .O(N__81549),
            .I(N__81533));
    LocalMux I__15156 (
            .O(N__81544),
            .I(N__81527));
    LocalMux I__15155 (
            .O(N__81541),
            .I(N__81527));
    InMux I__15154 (
            .O(N__81540),
            .I(N__81523));
    InMux I__15153 (
            .O(N__81539),
            .I(N__81520));
    LocalMux I__15152 (
            .O(N__81536),
            .I(N__81515));
    LocalMux I__15151 (
            .O(N__81533),
            .I(N__81515));
    InMux I__15150 (
            .O(N__81532),
            .I(N__81512));
    Span4Mux_h I__15149 (
            .O(N__81527),
            .I(N__81509));
    InMux I__15148 (
            .O(N__81526),
            .I(N__81506));
    LocalMux I__15147 (
            .O(N__81523),
            .I(N__81499));
    LocalMux I__15146 (
            .O(N__81520),
            .I(N__81499));
    Span4Mux_v I__15145 (
            .O(N__81515),
            .I(N__81499));
    LocalMux I__15144 (
            .O(N__81512),
            .I(rco_int_0_a2_1_a2_0_53));
    Odrv4 I__15143 (
            .O(N__81509),
            .I(rco_int_0_a2_1_a2_0_53));
    LocalMux I__15142 (
            .O(N__81506),
            .I(rco_int_0_a2_1_a2_0_53));
    Odrv4 I__15141 (
            .O(N__81499),
            .I(rco_int_0_a2_1_a2_0_53));
    InMux I__15140 (
            .O(N__81490),
            .I(N__81486));
    CascadeMux I__15139 (
            .O(N__81489),
            .I(N__81483));
    LocalMux I__15138 (
            .O(N__81486),
            .I(N__81480));
    InMux I__15137 (
            .O(N__81483),
            .I(N__81475));
    Span12Mux_h I__15136 (
            .O(N__81480),
            .I(N__81472));
    InMux I__15135 (
            .O(N__81479),
            .I(N__81469));
    InMux I__15134 (
            .O(N__81478),
            .I(N__81466));
    LocalMux I__15133 (
            .O(N__81475),
            .I(N__81463));
    Span12Mux_v I__15132 (
            .O(N__81472),
            .I(N__81460));
    LocalMux I__15131 (
            .O(N__81469),
            .I(N__81455));
    LocalMux I__15130 (
            .O(N__81466),
            .I(N__81455));
    Span4Mux_v I__15129 (
            .O(N__81463),
            .I(N__81452));
    Odrv12 I__15128 (
            .O(N__81460),
            .I(shift_srl_54_RNIEAU71Z0Z_15));
    Odrv12 I__15127 (
            .O(N__81455),
            .I(shift_srl_54_RNIEAU71Z0Z_15));
    Odrv4 I__15126 (
            .O(N__81452),
            .I(shift_srl_54_RNIEAU71Z0Z_15));
    InMux I__15125 (
            .O(N__81445),
            .I(N__81437));
    InMux I__15124 (
            .O(N__81444),
            .I(N__81432));
    InMux I__15123 (
            .O(N__81443),
            .I(N__81432));
    CascadeMux I__15122 (
            .O(N__81442),
            .I(N__81429));
    InMux I__15121 (
            .O(N__81441),
            .I(N__81424));
    InMux I__15120 (
            .O(N__81440),
            .I(N__81424));
    LocalMux I__15119 (
            .O(N__81437),
            .I(N__81418));
    LocalMux I__15118 (
            .O(N__81432),
            .I(N__81418));
    InMux I__15117 (
            .O(N__81429),
            .I(N__81415));
    LocalMux I__15116 (
            .O(N__81424),
            .I(N__81411));
    InMux I__15115 (
            .O(N__81423),
            .I(N__81408));
    Span4Mux_v I__15114 (
            .O(N__81418),
            .I(N__81403));
    LocalMux I__15113 (
            .O(N__81415),
            .I(N__81403));
    InMux I__15112 (
            .O(N__81414),
            .I(N__81400));
    Span4Mux_h I__15111 (
            .O(N__81411),
            .I(N__81397));
    LocalMux I__15110 (
            .O(N__81408),
            .I(N__81394));
    Span4Mux_h I__15109 (
            .O(N__81403),
            .I(N__81391));
    LocalMux I__15108 (
            .O(N__81400),
            .I(rco_int_0_a2_1_a2_0_0_59));
    Odrv4 I__15107 (
            .O(N__81397),
            .I(rco_int_0_a2_1_a2_0_0_59));
    Odrv4 I__15106 (
            .O(N__81394),
            .I(rco_int_0_a2_1_a2_0_0_59));
    Odrv4 I__15105 (
            .O(N__81391),
            .I(rco_int_0_a2_1_a2_0_0_59));
    InMux I__15104 (
            .O(N__81382),
            .I(N__81379));
    LocalMux I__15103 (
            .O(N__81379),
            .I(N__81376));
    Span4Mux_v I__15102 (
            .O(N__81376),
            .I(N__81373));
    Span4Mux_h I__15101 (
            .O(N__81373),
            .I(N__81370));
    Odrv4 I__15100 (
            .O(N__81370),
            .I(rco_int_0_a3_0_a2cf1_1_66));
    InMux I__15099 (
            .O(N__81367),
            .I(N__81364));
    LocalMux I__15098 (
            .O(N__81364),
            .I(N__81360));
    CascadeMux I__15097 (
            .O(N__81363),
            .I(N__81357));
    Span4Mux_v I__15096 (
            .O(N__81360),
            .I(N__81354));
    InMux I__15095 (
            .O(N__81357),
            .I(N__81351));
    Odrv4 I__15094 (
            .O(N__81354),
            .I(rco_int_0_a2_1_a2_1_48));
    LocalMux I__15093 (
            .O(N__81351),
            .I(rco_int_0_a2_1_a2_1_48));
    CascadeMux I__15092 (
            .O(N__81346),
            .I(rco_int_0_a2_1_a2_0_0_59_cascade_));
    CascadeMux I__15091 (
            .O(N__81343),
            .I(rco_int_0_a3_0_a2cf1_66_cascade_));
    IoInMux I__15090 (
            .O(N__81340),
            .I(N__81337));
    LocalMux I__15089 (
            .O(N__81337),
            .I(N__81334));
    IoSpan4Mux I__15088 (
            .O(N__81334),
            .I(N__81328));
    InMux I__15087 (
            .O(N__81333),
            .I(N__81324));
    InMux I__15086 (
            .O(N__81332),
            .I(N__81319));
    InMux I__15085 (
            .O(N__81331),
            .I(N__81316));
    Span4Mux_s3_h I__15084 (
            .O(N__81328),
            .I(N__81313));
    InMux I__15083 (
            .O(N__81327),
            .I(N__81310));
    LocalMux I__15082 (
            .O(N__81324),
            .I(N__81307));
    InMux I__15081 (
            .O(N__81323),
            .I(N__81304));
    InMux I__15080 (
            .O(N__81322),
            .I(N__81301));
    LocalMux I__15079 (
            .O(N__81319),
            .I(N__81298));
    LocalMux I__15078 (
            .O(N__81316),
            .I(N__81295));
    Span4Mux_h I__15077 (
            .O(N__81313),
            .I(N__81290));
    LocalMux I__15076 (
            .O(N__81310),
            .I(N__81290));
    Span4Mux_v I__15075 (
            .O(N__81307),
            .I(N__81285));
    LocalMux I__15074 (
            .O(N__81304),
            .I(N__81282));
    LocalMux I__15073 (
            .O(N__81301),
            .I(N__81279));
    Span4Mux_v I__15072 (
            .O(N__81298),
            .I(N__81272));
    Span4Mux_v I__15071 (
            .O(N__81295),
            .I(N__81272));
    Span4Mux_h I__15070 (
            .O(N__81290),
            .I(N__81272));
    InMux I__15069 (
            .O(N__81289),
            .I(N__81269));
    InMux I__15068 (
            .O(N__81288),
            .I(N__81266));
    Span4Mux_h I__15067 (
            .O(N__81285),
            .I(N__81261));
    Span4Mux_h I__15066 (
            .O(N__81282),
            .I(N__81261));
    Odrv12 I__15065 (
            .O(N__81279),
            .I(rco_c_37));
    Odrv4 I__15064 (
            .O(N__81272),
            .I(rco_c_37));
    LocalMux I__15063 (
            .O(N__81269),
            .I(rco_c_37));
    LocalMux I__15062 (
            .O(N__81266),
            .I(rco_c_37));
    Odrv4 I__15061 (
            .O(N__81261),
            .I(rco_c_37));
    CascadeMux I__15060 (
            .O(N__81250),
            .I(rco_c_66_cascade_));
    CEMux I__15059 (
            .O(N__81247),
            .I(N__81243));
    CEMux I__15058 (
            .O(N__81246),
            .I(N__81240));
    LocalMux I__15057 (
            .O(N__81243),
            .I(N__81237));
    LocalMux I__15056 (
            .O(N__81240),
            .I(N__81234));
    Odrv12 I__15055 (
            .O(N__81237),
            .I(clk_en_76));
    Odrv4 I__15054 (
            .O(N__81234),
            .I(clk_en_76));
    InMux I__15053 (
            .O(N__81229),
            .I(N__81226));
    LocalMux I__15052 (
            .O(N__81226),
            .I(shift_srl_66Z0Z_0));
    InMux I__15051 (
            .O(N__81223),
            .I(N__81220));
    LocalMux I__15050 (
            .O(N__81220),
            .I(shift_srl_66Z0Z_1));
    InMux I__15049 (
            .O(N__81217),
            .I(N__81214));
    LocalMux I__15048 (
            .O(N__81214),
            .I(shift_srl_66Z0Z_2));
    InMux I__15047 (
            .O(N__81211),
            .I(N__81208));
    LocalMux I__15046 (
            .O(N__81208),
            .I(shift_srl_76Z0Z_2));
    InMux I__15045 (
            .O(N__81205),
            .I(N__81202));
    LocalMux I__15044 (
            .O(N__81202),
            .I(shift_srl_76Z0Z_3));
    InMux I__15043 (
            .O(N__81199),
            .I(N__81196));
    LocalMux I__15042 (
            .O(N__81196),
            .I(shift_srl_76Z0Z_4));
    InMux I__15041 (
            .O(N__81193),
            .I(N__81190));
    LocalMux I__15040 (
            .O(N__81190),
            .I(shift_srl_76Z0Z_5));
    InMux I__15039 (
            .O(N__81187),
            .I(N__81184));
    LocalMux I__15038 (
            .O(N__81184),
            .I(shift_srl_76Z0Z_6));
    InMux I__15037 (
            .O(N__81181),
            .I(N__81178));
    LocalMux I__15036 (
            .O(N__81178),
            .I(shift_srl_76Z0Z_7));
    IoInMux I__15035 (
            .O(N__81175),
            .I(N__81172));
    LocalMux I__15034 (
            .O(N__81172),
            .I(N__81169));
    Span4Mux_s3_h I__15033 (
            .O(N__81169),
            .I(N__81166));
    Span4Mux_v I__15032 (
            .O(N__81166),
            .I(N__81163));
    Span4Mux_h I__15031 (
            .O(N__81163),
            .I(N__81160));
    Odrv4 I__15030 (
            .O(N__81160),
            .I(rco_c_64));
    IoInMux I__15029 (
            .O(N__81157),
            .I(N__81154));
    LocalMux I__15028 (
            .O(N__81154),
            .I(N__81151));
    IoSpan4Mux I__15027 (
            .O(N__81151),
            .I(N__81148));
    Span4Mux_s3_h I__15026 (
            .O(N__81148),
            .I(N__81145));
    Span4Mux_h I__15025 (
            .O(N__81145),
            .I(N__81142));
    Odrv4 I__15024 (
            .O(N__81142),
            .I(rco_c_63));
    CascadeMux I__15023 (
            .O(N__81139),
            .I(N__81134));
    InMux I__15022 (
            .O(N__81138),
            .I(N__81129));
    InMux I__15021 (
            .O(N__81137),
            .I(N__81126));
    InMux I__15020 (
            .O(N__81134),
            .I(N__81117));
    InMux I__15019 (
            .O(N__81133),
            .I(N__81117));
    InMux I__15018 (
            .O(N__81132),
            .I(N__81117));
    LocalMux I__15017 (
            .O(N__81129),
            .I(N__81112));
    LocalMux I__15016 (
            .O(N__81126),
            .I(N__81112));
    InMux I__15015 (
            .O(N__81125),
            .I(N__81107));
    InMux I__15014 (
            .O(N__81124),
            .I(N__81107));
    LocalMux I__15013 (
            .O(N__81117),
            .I(N__81104));
    Span4Mux_h I__15012 (
            .O(N__81112),
            .I(N__81101));
    LocalMux I__15011 (
            .O(N__81107),
            .I(shift_srl_63Z0Z_15));
    Odrv4 I__15010 (
            .O(N__81104),
            .I(shift_srl_63Z0Z_15));
    Odrv4 I__15009 (
            .O(N__81101),
            .I(shift_srl_63Z0Z_15));
    InMux I__15008 (
            .O(N__81094),
            .I(N__81087));
    InMux I__15007 (
            .O(N__81093),
            .I(N__81087));
    InMux I__15006 (
            .O(N__81092),
            .I(N__81084));
    LocalMux I__15005 (
            .O(N__81087),
            .I(N__81079));
    LocalMux I__15004 (
            .O(N__81084),
            .I(N__81076));
    InMux I__15003 (
            .O(N__81083),
            .I(N__81073));
    InMux I__15002 (
            .O(N__81082),
            .I(N__81070));
    Span4Mux_v I__15001 (
            .O(N__81079),
            .I(N__81065));
    Span4Mux_v I__15000 (
            .O(N__81076),
            .I(N__81065));
    LocalMux I__14999 (
            .O(N__81073),
            .I(shift_srl_64Z0Z_15));
    LocalMux I__14998 (
            .O(N__81070),
            .I(shift_srl_64Z0Z_15));
    Odrv4 I__14997 (
            .O(N__81065),
            .I(shift_srl_64Z0Z_15));
    CascadeMux I__14996 (
            .O(N__81058),
            .I(N__81051));
    CascadeMux I__14995 (
            .O(N__81057),
            .I(N__81048));
    CascadeMux I__14994 (
            .O(N__81056),
            .I(N__81045));
    InMux I__14993 (
            .O(N__81055),
            .I(N__81038));
    InMux I__14992 (
            .O(N__81054),
            .I(N__81038));
    InMux I__14991 (
            .O(N__81051),
            .I(N__81038));
    InMux I__14990 (
            .O(N__81048),
            .I(N__81033));
    InMux I__14989 (
            .O(N__81045),
            .I(N__81033));
    LocalMux I__14988 (
            .O(N__81038),
            .I(N__81029));
    LocalMux I__14987 (
            .O(N__81033),
            .I(N__81025));
    CascadeMux I__14986 (
            .O(N__81032),
            .I(N__81022));
    Span4Mux_h I__14985 (
            .O(N__81029),
            .I(N__81019));
    InMux I__14984 (
            .O(N__81028),
            .I(N__81016));
    Span4Mux_v I__14983 (
            .O(N__81025),
            .I(N__81013));
    InMux I__14982 (
            .O(N__81022),
            .I(N__81010));
    Span4Mux_v I__14981 (
            .O(N__81019),
            .I(N__81007));
    LocalMux I__14980 (
            .O(N__81016),
            .I(shift_srl_62_RNIM5RKZ0Z_15));
    Odrv4 I__14979 (
            .O(N__81013),
            .I(shift_srl_62_RNIM5RKZ0Z_15));
    LocalMux I__14978 (
            .O(N__81010),
            .I(shift_srl_62_RNIM5RKZ0Z_15));
    Odrv4 I__14977 (
            .O(N__81007),
            .I(shift_srl_62_RNIM5RKZ0Z_15));
    InMux I__14976 (
            .O(N__80998),
            .I(N__80995));
    LocalMux I__14975 (
            .O(N__80995),
            .I(N__80991));
    InMux I__14974 (
            .O(N__80994),
            .I(N__80987));
    Span4Mux_h I__14973 (
            .O(N__80991),
            .I(N__80984));
    InMux I__14972 (
            .O(N__80990),
            .I(N__80981));
    LocalMux I__14971 (
            .O(N__80987),
            .I(shift_srl_65Z0Z_15));
    Odrv4 I__14970 (
            .O(N__80984),
            .I(shift_srl_65Z0Z_15));
    LocalMux I__14969 (
            .O(N__80981),
            .I(shift_srl_65Z0Z_15));
    InMux I__14968 (
            .O(N__80974),
            .I(N__80971));
    LocalMux I__14967 (
            .O(N__80971),
            .I(N__80968));
    Span4Mux_h I__14966 (
            .O(N__80968),
            .I(N__80965));
    Sp12to4 I__14965 (
            .O(N__80965),
            .I(N__80962));
    Odrv12 I__14964 (
            .O(N__80962),
            .I(shift_srl_65_RNILFDF1Z0Z_15));
    InMux I__14963 (
            .O(N__80959),
            .I(N__80956));
    LocalMux I__14962 (
            .O(N__80956),
            .I(shift_srl_76Z0Z_10));
    InMux I__14961 (
            .O(N__80953),
            .I(N__80950));
    LocalMux I__14960 (
            .O(N__80950),
            .I(shift_srl_76Z0Z_11));
    InMux I__14959 (
            .O(N__80947),
            .I(N__80944));
    LocalMux I__14958 (
            .O(N__80944),
            .I(shift_srl_76Z0Z_12));
    InMux I__14957 (
            .O(N__80941),
            .I(N__80938));
    LocalMux I__14956 (
            .O(N__80938),
            .I(shift_srl_76Z0Z_13));
    InMux I__14955 (
            .O(N__80935),
            .I(N__80932));
    LocalMux I__14954 (
            .O(N__80932),
            .I(shift_srl_76Z0Z_14));
    InMux I__14953 (
            .O(N__80929),
            .I(N__80926));
    LocalMux I__14952 (
            .O(N__80926),
            .I(shift_srl_76Z0Z_9));
    InMux I__14951 (
            .O(N__80923),
            .I(N__80920));
    LocalMux I__14950 (
            .O(N__80920),
            .I(shift_srl_76Z0Z_8));
    InMux I__14949 (
            .O(N__80917),
            .I(N__80914));
    LocalMux I__14948 (
            .O(N__80914),
            .I(shift_srl_76Z0Z_0));
    InMux I__14947 (
            .O(N__80911),
            .I(N__80908));
    LocalMux I__14946 (
            .O(N__80908),
            .I(shift_srl_76Z0Z_1));
    InMux I__14945 (
            .O(N__80905),
            .I(N__80902));
    LocalMux I__14944 (
            .O(N__80902),
            .I(shift_srl_82Z0Z_7));
    InMux I__14943 (
            .O(N__80899),
            .I(N__80896));
    LocalMux I__14942 (
            .O(N__80896),
            .I(shift_srl_82Z0Z_8));
    IoInMux I__14941 (
            .O(N__80893),
            .I(N__80890));
    LocalMux I__14940 (
            .O(N__80890),
            .I(N__80887));
    Span4Mux_s2_v I__14939 (
            .O(N__80887),
            .I(N__80884));
    Span4Mux_v I__14938 (
            .O(N__80884),
            .I(N__80881));
    Odrv4 I__14937 (
            .O(N__80881),
            .I(N_3998_i));
    CascadeMux I__14936 (
            .O(N__80878),
            .I(shift_srl_80_RNIG3FB1Z0Z_15_cascade_));
    CascadeMux I__14935 (
            .O(N__80875),
            .I(clk_en_0_a3_0_a2_0_83_cascade_));
    CEMux I__14934 (
            .O(N__80872),
            .I(N__80869));
    LocalMux I__14933 (
            .O(N__80869),
            .I(N__80865));
    CEMux I__14932 (
            .O(N__80868),
            .I(N__80861));
    Span4Mux_v I__14931 (
            .O(N__80865),
            .I(N__80858));
    CEMux I__14930 (
            .O(N__80864),
            .I(N__80855));
    LocalMux I__14929 (
            .O(N__80861),
            .I(N__80852));
    Odrv4 I__14928 (
            .O(N__80858),
            .I(clk_en_83));
    LocalMux I__14927 (
            .O(N__80855),
            .I(clk_en_83));
    Odrv12 I__14926 (
            .O(N__80852),
            .I(clk_en_83));
    CEMux I__14925 (
            .O(N__80845),
            .I(N__80842));
    LocalMux I__14924 (
            .O(N__80842),
            .I(N__80838));
    CEMux I__14923 (
            .O(N__80841),
            .I(N__80835));
    Span4Mux_h I__14922 (
            .O(N__80838),
            .I(N__80832));
    LocalMux I__14921 (
            .O(N__80835),
            .I(N__80829));
    Odrv4 I__14920 (
            .O(N__80832),
            .I(N_787));
    Odrv4 I__14919 (
            .O(N__80829),
            .I(N_787));
    InMux I__14918 (
            .O(N__80824),
            .I(N__80814));
    InMux I__14917 (
            .O(N__80823),
            .I(N__80814));
    InMux I__14916 (
            .O(N__80822),
            .I(N__80814));
    InMux I__14915 (
            .O(N__80821),
            .I(N__80811));
    LocalMux I__14914 (
            .O(N__80814),
            .I(N__80808));
    LocalMux I__14913 (
            .O(N__80811),
            .I(shift_srl_82Z0Z_15));
    Odrv4 I__14912 (
            .O(N__80808),
            .I(shift_srl_82Z0Z_15));
    CascadeMux I__14911 (
            .O(N__80803),
            .I(N__80800));
    InMux I__14910 (
            .O(N__80800),
            .I(N__80796));
    InMux I__14909 (
            .O(N__80799),
            .I(N__80793));
    LocalMux I__14908 (
            .O(N__80796),
            .I(N__80790));
    LocalMux I__14907 (
            .O(N__80793),
            .I(shift_srl_83Z0Z_15));
    Odrv4 I__14906 (
            .O(N__80790),
            .I(shift_srl_83Z0Z_15));
    InMux I__14905 (
            .O(N__80785),
            .I(N__80782));
    LocalMux I__14904 (
            .O(N__80782),
            .I(N__80779));
    Span4Mux_h I__14903 (
            .O(N__80779),
            .I(N__80776));
    Span4Mux_h I__14902 (
            .O(N__80776),
            .I(N__80771));
    InMux I__14901 (
            .O(N__80775),
            .I(N__80768));
    InMux I__14900 (
            .O(N__80774),
            .I(N__80765));
    Sp12to4 I__14899 (
            .O(N__80771),
            .I(N__80760));
    LocalMux I__14898 (
            .O(N__80768),
            .I(N__80760));
    LocalMux I__14897 (
            .O(N__80765),
            .I(N__80757));
    Span12Mux_v I__14896 (
            .O(N__80760),
            .I(N__80754));
    Odrv12 I__14895 (
            .O(N__80757),
            .I(rco_int_0_a2_0_a2_0_83));
    Odrv12 I__14894 (
            .O(N__80754),
            .I(rco_int_0_a2_0_a2_0_83));
    InMux I__14893 (
            .O(N__80749),
            .I(N__80746));
    LocalMux I__14892 (
            .O(N__80746),
            .I(shift_srl_83Z0Z_10));
    InMux I__14891 (
            .O(N__80743),
            .I(N__80740));
    LocalMux I__14890 (
            .O(N__80740),
            .I(shift_srl_83Z0Z_8));
    InMux I__14889 (
            .O(N__80737),
            .I(N__80734));
    LocalMux I__14888 (
            .O(N__80734),
            .I(shift_srl_83Z0Z_9));
    InMux I__14887 (
            .O(N__80731),
            .I(N__80728));
    LocalMux I__14886 (
            .O(N__80728),
            .I(shift_srl_82Z0Z_10));
    InMux I__14885 (
            .O(N__80725),
            .I(N__80722));
    LocalMux I__14884 (
            .O(N__80722),
            .I(shift_srl_82Z0Z_11));
    InMux I__14883 (
            .O(N__80719),
            .I(N__80716));
    LocalMux I__14882 (
            .O(N__80716),
            .I(shift_srl_82Z0Z_12));
    InMux I__14881 (
            .O(N__80713),
            .I(N__80710));
    LocalMux I__14880 (
            .O(N__80710),
            .I(shift_srl_82Z0Z_13));
    InMux I__14879 (
            .O(N__80707),
            .I(N__80704));
    LocalMux I__14878 (
            .O(N__80704),
            .I(shift_srl_82Z0Z_14));
    InMux I__14877 (
            .O(N__80701),
            .I(N__80698));
    LocalMux I__14876 (
            .O(N__80698),
            .I(shift_srl_82Z0Z_9));
    InMux I__14875 (
            .O(N__80695),
            .I(N__80692));
    LocalMux I__14874 (
            .O(N__80692),
            .I(shift_srl_192Z0Z_8));
    InMux I__14873 (
            .O(N__80689),
            .I(N__80686));
    LocalMux I__14872 (
            .O(N__80686),
            .I(N__80683));
    Span4Mux_h I__14871 (
            .O(N__80683),
            .I(N__80680));
    Odrv4 I__14870 (
            .O(N__80680),
            .I(shift_srl_192Z0Z_9));
    CEMux I__14869 (
            .O(N__80677),
            .I(N__80674));
    LocalMux I__14868 (
            .O(N__80674),
            .I(N__80669));
    CEMux I__14867 (
            .O(N__80673),
            .I(N__80666));
    CEMux I__14866 (
            .O(N__80672),
            .I(N__80663));
    Span4Mux_h I__14865 (
            .O(N__80669),
            .I(N__80658));
    LocalMux I__14864 (
            .O(N__80666),
            .I(N__80658));
    LocalMux I__14863 (
            .O(N__80663),
            .I(N__80655));
    Span4Mux_v I__14862 (
            .O(N__80658),
            .I(N__80652));
    Odrv4 I__14861 (
            .O(N__80655),
            .I(clk_en_192));
    Odrv4 I__14860 (
            .O(N__80652),
            .I(clk_en_192));
    InMux I__14859 (
            .O(N__80647),
            .I(N__80644));
    LocalMux I__14858 (
            .O(N__80644),
            .I(shift_srl_173Z0Z_10));
    InMux I__14857 (
            .O(N__80641),
            .I(N__80638));
    LocalMux I__14856 (
            .O(N__80638),
            .I(shift_srl_173Z0Z_11));
    InMux I__14855 (
            .O(N__80635),
            .I(N__80632));
    LocalMux I__14854 (
            .O(N__80632),
            .I(shift_srl_173Z0Z_12));
    InMux I__14853 (
            .O(N__80629),
            .I(N__80626));
    LocalMux I__14852 (
            .O(N__80626),
            .I(shift_srl_173Z0Z_13));
    InMux I__14851 (
            .O(N__80623),
            .I(N__80620));
    LocalMux I__14850 (
            .O(N__80620),
            .I(N__80617));
    Span4Mux_h I__14849 (
            .O(N__80617),
            .I(N__80614));
    Odrv4 I__14848 (
            .O(N__80614),
            .I(shift_srl_173Z0Z_14));
    InMux I__14847 (
            .O(N__80611),
            .I(N__80608));
    LocalMux I__14846 (
            .O(N__80608),
            .I(shift_srl_173Z0Z_9));
    InMux I__14845 (
            .O(N__80605),
            .I(N__80602));
    LocalMux I__14844 (
            .O(N__80602),
            .I(N__80599));
    Span4Mux_h I__14843 (
            .O(N__80599),
            .I(N__80596));
    Span4Mux_h I__14842 (
            .O(N__80596),
            .I(N__80593));
    Odrv4 I__14841 (
            .O(N__80593),
            .I(shift_srl_173Z0Z_7));
    InMux I__14840 (
            .O(N__80590),
            .I(N__80587));
    LocalMux I__14839 (
            .O(N__80587),
            .I(shift_srl_173Z0Z_8));
    CEMux I__14838 (
            .O(N__80584),
            .I(N__80580));
    CEMux I__14837 (
            .O(N__80583),
            .I(N__80576));
    LocalMux I__14836 (
            .O(N__80580),
            .I(N__80573));
    CEMux I__14835 (
            .O(N__80579),
            .I(N__80570));
    LocalMux I__14834 (
            .O(N__80576),
            .I(N__80567));
    Span4Mux_v I__14833 (
            .O(N__80573),
            .I(N__80564));
    LocalMux I__14832 (
            .O(N__80570),
            .I(N__80561));
    Span4Mux_h I__14831 (
            .O(N__80567),
            .I(N__80558));
    Span4Mux_h I__14830 (
            .O(N__80564),
            .I(N__80553));
    Span4Mux_h I__14829 (
            .O(N__80561),
            .I(N__80553));
    Odrv4 I__14828 (
            .O(N__80558),
            .I(clk_en_173));
    Odrv4 I__14827 (
            .O(N__80553),
            .I(clk_en_173));
    InMux I__14826 (
            .O(N__80548),
            .I(N__80545));
    LocalMux I__14825 (
            .O(N__80545),
            .I(N__80540));
    CascadeMux I__14824 (
            .O(N__80544),
            .I(N__80535));
    CascadeMux I__14823 (
            .O(N__80543),
            .I(N__80532));
    Span4Mux_v I__14822 (
            .O(N__80540),
            .I(N__80529));
    CascadeMux I__14821 (
            .O(N__80539),
            .I(N__80526));
    InMux I__14820 (
            .O(N__80538),
            .I(N__80523));
    InMux I__14819 (
            .O(N__80535),
            .I(N__80517));
    InMux I__14818 (
            .O(N__80532),
            .I(N__80517));
    Sp12to4 I__14817 (
            .O(N__80529),
            .I(N__80514));
    InMux I__14816 (
            .O(N__80526),
            .I(N__80511));
    LocalMux I__14815 (
            .O(N__80523),
            .I(N__80508));
    InMux I__14814 (
            .O(N__80522),
            .I(N__80505));
    LocalMux I__14813 (
            .O(N__80517),
            .I(N__80502));
    Span12Mux_h I__14812 (
            .O(N__80514),
            .I(N__80497));
    LocalMux I__14811 (
            .O(N__80511),
            .I(N__80497));
    Span4Mux_v I__14810 (
            .O(N__80508),
            .I(N__80494));
    LocalMux I__14809 (
            .O(N__80505),
            .I(N__80491));
    Span4Mux_h I__14808 (
            .O(N__80502),
            .I(N__80488));
    Span12Mux_v I__14807 (
            .O(N__80497),
            .I(N__80485));
    Odrv4 I__14806 (
            .O(N__80494),
            .I(shift_srl_176_RNIUGI51Z0Z_15));
    Odrv4 I__14805 (
            .O(N__80491),
            .I(shift_srl_176_RNIUGI51Z0Z_15));
    Odrv4 I__14804 (
            .O(N__80488),
            .I(shift_srl_176_RNIUGI51Z0Z_15));
    Odrv12 I__14803 (
            .O(N__80485),
            .I(shift_srl_176_RNIUGI51Z0Z_15));
    InMux I__14802 (
            .O(N__80476),
            .I(N__80471));
    InMux I__14801 (
            .O(N__80475),
            .I(N__80468));
    InMux I__14800 (
            .O(N__80474),
            .I(N__80465));
    LocalMux I__14799 (
            .O(N__80471),
            .I(N__80462));
    LocalMux I__14798 (
            .O(N__80468),
            .I(N__80459));
    LocalMux I__14797 (
            .O(N__80465),
            .I(N__80456));
    Span4Mux_h I__14796 (
            .O(N__80462),
            .I(N__80452));
    Span4Mux_v I__14795 (
            .O(N__80459),
            .I(N__80446));
    Span4Mux_v I__14794 (
            .O(N__80456),
            .I(N__80443));
    InMux I__14793 (
            .O(N__80455),
            .I(N__80440));
    Span4Mux_v I__14792 (
            .O(N__80452),
            .I(N__80437));
    InMux I__14791 (
            .O(N__80451),
            .I(N__80430));
    InMux I__14790 (
            .O(N__80450),
            .I(N__80430));
    InMux I__14789 (
            .O(N__80449),
            .I(N__80430));
    Odrv4 I__14788 (
            .O(N__80446),
            .I(shift_srl_177Z0Z_15));
    Odrv4 I__14787 (
            .O(N__80443),
            .I(shift_srl_177Z0Z_15));
    LocalMux I__14786 (
            .O(N__80440),
            .I(shift_srl_177Z0Z_15));
    Odrv4 I__14785 (
            .O(N__80437),
            .I(shift_srl_177Z0Z_15));
    LocalMux I__14784 (
            .O(N__80430),
            .I(shift_srl_177Z0Z_15));
    CascadeMux I__14783 (
            .O(N__80419),
            .I(N__80416));
    InMux I__14782 (
            .O(N__80416),
            .I(N__80412));
    InMux I__14781 (
            .O(N__80415),
            .I(N__80409));
    LocalMux I__14780 (
            .O(N__80412),
            .I(N__80406));
    LocalMux I__14779 (
            .O(N__80409),
            .I(N__80402));
    Span4Mux_v I__14778 (
            .O(N__80406),
            .I(N__80397));
    InMux I__14777 (
            .O(N__80405),
            .I(N__80394));
    Span4Mux_v I__14776 (
            .O(N__80402),
            .I(N__80391));
    InMux I__14775 (
            .O(N__80401),
            .I(N__80386));
    InMux I__14774 (
            .O(N__80400),
            .I(N__80386));
    Odrv4 I__14773 (
            .O(N__80397),
            .I(shift_srl_178Z0Z_15));
    LocalMux I__14772 (
            .O(N__80394),
            .I(shift_srl_178Z0Z_15));
    Odrv4 I__14771 (
            .O(N__80391),
            .I(shift_srl_178Z0Z_15));
    LocalMux I__14770 (
            .O(N__80386),
            .I(shift_srl_178Z0Z_15));
    IoInMux I__14769 (
            .O(N__80377),
            .I(N__80374));
    LocalMux I__14768 (
            .O(N__80374),
            .I(N__80371));
    IoSpan4Mux I__14767 (
            .O(N__80371),
            .I(N__80368));
    Span4Mux_s0_v I__14766 (
            .O(N__80368),
            .I(N__80365));
    Span4Mux_v I__14765 (
            .O(N__80365),
            .I(N__80362));
    Odrv4 I__14764 (
            .O(N__80362),
            .I(rco_c_178));
    InMux I__14763 (
            .O(N__80359),
            .I(N__80356));
    LocalMux I__14762 (
            .O(N__80356),
            .I(N__80351));
    InMux I__14761 (
            .O(N__80355),
            .I(N__80346));
    InMux I__14760 (
            .O(N__80354),
            .I(N__80346));
    Span4Mux_v I__14759 (
            .O(N__80351),
            .I(N__80342));
    LocalMux I__14758 (
            .O(N__80346),
            .I(N__80339));
    InMux I__14757 (
            .O(N__80345),
            .I(N__80336));
    Span4Mux_h I__14756 (
            .O(N__80342),
            .I(N__80329));
    Span4Mux_v I__14755 (
            .O(N__80339),
            .I(N__80329));
    LocalMux I__14754 (
            .O(N__80336),
            .I(N__80326));
    InMux I__14753 (
            .O(N__80335),
            .I(N__80321));
    InMux I__14752 (
            .O(N__80334),
            .I(N__80321));
    Odrv4 I__14751 (
            .O(N__80329),
            .I(N_4173));
    Odrv4 I__14750 (
            .O(N__80326),
            .I(N_4173));
    LocalMux I__14749 (
            .O(N__80321),
            .I(N_4173));
    IoInMux I__14748 (
            .O(N__80314),
            .I(N__80311));
    LocalMux I__14747 (
            .O(N__80311),
            .I(N__80308));
    Span4Mux_s3_v I__14746 (
            .O(N__80308),
            .I(N__80305));
    Span4Mux_v I__14745 (
            .O(N__80305),
            .I(N__80302));
    Odrv4 I__14744 (
            .O(N__80302),
            .I(rco_c_188));
    InMux I__14743 (
            .O(N__80299),
            .I(N__80296));
    LocalMux I__14742 (
            .O(N__80296),
            .I(shift_srl_188Z0Z_14));
    InMux I__14741 (
            .O(N__80293),
            .I(N__80290));
    LocalMux I__14740 (
            .O(N__80290),
            .I(shift_srl_188Z0Z_13));
    InMux I__14739 (
            .O(N__80287),
            .I(N__80284));
    LocalMux I__14738 (
            .O(N__80284),
            .I(shift_srl_188Z0Z_12));
    InMux I__14737 (
            .O(N__80281),
            .I(N__80278));
    LocalMux I__14736 (
            .O(N__80278),
            .I(shift_srl_188Z0Z_11));
    InMux I__14735 (
            .O(N__80275),
            .I(N__80272));
    LocalMux I__14734 (
            .O(N__80272),
            .I(shift_srl_188Z0Z_10));
    InMux I__14733 (
            .O(N__80269),
            .I(N__80266));
    LocalMux I__14732 (
            .O(N__80266),
            .I(N__80263));
    Span4Mux_h I__14731 (
            .O(N__80263),
            .I(N__80260));
    Odrv4 I__14730 (
            .O(N__80260),
            .I(shift_srl_192Z0Z_7));
    InMux I__14729 (
            .O(N__80257),
            .I(N__80254));
    LocalMux I__14728 (
            .O(N__80254),
            .I(shift_srl_177Z0Z_13));
    InMux I__14727 (
            .O(N__80251),
            .I(N__80248));
    LocalMux I__14726 (
            .O(N__80248),
            .I(shift_srl_180Z0Z_0));
    InMux I__14725 (
            .O(N__80245),
            .I(N__80242));
    LocalMux I__14724 (
            .O(N__80242),
            .I(shift_srl_180Z0Z_1));
    InMux I__14723 (
            .O(N__80239),
            .I(N__80236));
    LocalMux I__14722 (
            .O(N__80236),
            .I(shift_srl_180Z0Z_2));
    InMux I__14721 (
            .O(N__80233),
            .I(N__80230));
    LocalMux I__14720 (
            .O(N__80230),
            .I(shift_srl_180Z0Z_3));
    InMux I__14719 (
            .O(N__80227),
            .I(N__80224));
    LocalMux I__14718 (
            .O(N__80224),
            .I(shift_srl_180Z0Z_7));
    InMux I__14717 (
            .O(N__80221),
            .I(N__80218));
    LocalMux I__14716 (
            .O(N__80218),
            .I(shift_srl_180Z0Z_6));
    InMux I__14715 (
            .O(N__80215),
            .I(N__80212));
    LocalMux I__14714 (
            .O(N__80212),
            .I(shift_srl_170Z0Z_5));
    InMux I__14713 (
            .O(N__80209),
            .I(N__80206));
    LocalMux I__14712 (
            .O(N__80206),
            .I(shift_srl_170Z0Z_6));
    InMux I__14711 (
            .O(N__80203),
            .I(N__80200));
    LocalMux I__14710 (
            .O(N__80200),
            .I(shift_srl_177Z0Z_0));
    InMux I__14709 (
            .O(N__80197),
            .I(N__80194));
    LocalMux I__14708 (
            .O(N__80194),
            .I(shift_srl_177Z0Z_1));
    InMux I__14707 (
            .O(N__80191),
            .I(N__80188));
    LocalMux I__14706 (
            .O(N__80188),
            .I(shift_srl_177Z0Z_2));
    InMux I__14705 (
            .O(N__80185),
            .I(N__80182));
    LocalMux I__14704 (
            .O(N__80182),
            .I(shift_srl_177Z0Z_3));
    InMux I__14703 (
            .O(N__80179),
            .I(N__80176));
    LocalMux I__14702 (
            .O(N__80176),
            .I(shift_srl_177Z0Z_4));
    InMux I__14701 (
            .O(N__80173),
            .I(N__80170));
    LocalMux I__14700 (
            .O(N__80170),
            .I(shift_srl_177Z0Z_5));
    InMux I__14699 (
            .O(N__80167),
            .I(N__80164));
    LocalMux I__14698 (
            .O(N__80164),
            .I(shift_srl_167Z0Z_3));
    InMux I__14697 (
            .O(N__80161),
            .I(N__80158));
    LocalMux I__14696 (
            .O(N__80158),
            .I(shift_srl_167Z0Z_4));
    InMux I__14695 (
            .O(N__80155),
            .I(N__80152));
    LocalMux I__14694 (
            .O(N__80152),
            .I(shift_srl_167Z0Z_5));
    InMux I__14693 (
            .O(N__80149),
            .I(N__80146));
    LocalMux I__14692 (
            .O(N__80146),
            .I(shift_srl_167Z0Z_6));
    InMux I__14691 (
            .O(N__80143),
            .I(N__80140));
    LocalMux I__14690 (
            .O(N__80140),
            .I(shift_srl_167Z0Z_7));
    InMux I__14689 (
            .O(N__80137),
            .I(N__80134));
    LocalMux I__14688 (
            .O(N__80134),
            .I(shift_srl_170Z0Z_0));
    InMux I__14687 (
            .O(N__80131),
            .I(N__80128));
    LocalMux I__14686 (
            .O(N__80128),
            .I(shift_srl_170Z0Z_1));
    InMux I__14685 (
            .O(N__80125),
            .I(N__80122));
    LocalMux I__14684 (
            .O(N__80122),
            .I(shift_srl_170Z0Z_2));
    InMux I__14683 (
            .O(N__80119),
            .I(N__80116));
    LocalMux I__14682 (
            .O(N__80116),
            .I(shift_srl_170Z0Z_3));
    InMux I__14681 (
            .O(N__80113),
            .I(N__80110));
    LocalMux I__14680 (
            .O(N__80110),
            .I(shift_srl_170Z0Z_4));
    InMux I__14679 (
            .O(N__80107),
            .I(N__80104));
    LocalMux I__14678 (
            .O(N__80104),
            .I(shift_srl_167Z0Z_12));
    InMux I__14677 (
            .O(N__80101),
            .I(N__80098));
    LocalMux I__14676 (
            .O(N__80098),
            .I(shift_srl_167Z0Z_13));
    InMux I__14675 (
            .O(N__80095),
            .I(N__80092));
    LocalMux I__14674 (
            .O(N__80092),
            .I(shift_srl_167Z0Z_14));
    InMux I__14673 (
            .O(N__80089),
            .I(N__80086));
    LocalMux I__14672 (
            .O(N__80086),
            .I(shift_srl_167Z0Z_9));
    InMux I__14671 (
            .O(N__80083),
            .I(N__80080));
    LocalMux I__14670 (
            .O(N__80080),
            .I(shift_srl_167Z0Z_8));
    InMux I__14669 (
            .O(N__80077),
            .I(N__80074));
    LocalMux I__14668 (
            .O(N__80074),
            .I(shift_srl_167Z0Z_0));
    InMux I__14667 (
            .O(N__80071),
            .I(N__80068));
    LocalMux I__14666 (
            .O(N__80068),
            .I(shift_srl_167Z0Z_1));
    InMux I__14665 (
            .O(N__80065),
            .I(N__80062));
    LocalMux I__14664 (
            .O(N__80062),
            .I(shift_srl_167Z0Z_2));
    InMux I__14663 (
            .O(N__80059),
            .I(N__80056));
    LocalMux I__14662 (
            .O(N__80056),
            .I(shift_srl_165Z0Z_1));
    InMux I__14661 (
            .O(N__80053),
            .I(N__80050));
    LocalMux I__14660 (
            .O(N__80050),
            .I(shift_srl_165Z0Z_2));
    InMux I__14659 (
            .O(N__80047),
            .I(N__80044));
    LocalMux I__14658 (
            .O(N__80044),
            .I(shift_srl_165Z0Z_3));
    InMux I__14657 (
            .O(N__80041),
            .I(N__80038));
    LocalMux I__14656 (
            .O(N__80038),
            .I(shift_srl_165Z0Z_4));
    InMux I__14655 (
            .O(N__80035),
            .I(N__80032));
    LocalMux I__14654 (
            .O(N__80032),
            .I(shift_srl_165Z0Z_5));
    InMux I__14653 (
            .O(N__80029),
            .I(N__80026));
    LocalMux I__14652 (
            .O(N__80026),
            .I(shift_srl_165Z0Z_6));
    InMux I__14651 (
            .O(N__80023),
            .I(N__80020));
    LocalMux I__14650 (
            .O(N__80020),
            .I(shift_srl_165Z0Z_7));
    CEMux I__14649 (
            .O(N__80017),
            .I(N__80014));
    LocalMux I__14648 (
            .O(N__80014),
            .I(N__80011));
    Span4Mux_v I__14647 (
            .O(N__80011),
            .I(N__80007));
    CEMux I__14646 (
            .O(N__80010),
            .I(N__80004));
    Sp12to4 I__14645 (
            .O(N__80007),
            .I(N__79999));
    LocalMux I__14644 (
            .O(N__80004),
            .I(N__79999));
    Odrv12 I__14643 (
            .O(N__79999),
            .I(clk_en_165));
    InMux I__14642 (
            .O(N__79996),
            .I(N__79993));
    LocalMux I__14641 (
            .O(N__79993),
            .I(shift_srl_167Z0Z_10));
    InMux I__14640 (
            .O(N__79990),
            .I(N__79987));
    LocalMux I__14639 (
            .O(N__79987),
            .I(shift_srl_167Z0Z_11));
    InMux I__14638 (
            .O(N__79984),
            .I(N__79981));
    LocalMux I__14637 (
            .O(N__79981),
            .I(shift_srl_165Z0Z_10));
    InMux I__14636 (
            .O(N__79978),
            .I(N__79975));
    LocalMux I__14635 (
            .O(N__79975),
            .I(shift_srl_165Z0Z_11));
    InMux I__14634 (
            .O(N__79972),
            .I(N__79969));
    LocalMux I__14633 (
            .O(N__79969),
            .I(shift_srl_165Z0Z_12));
    InMux I__14632 (
            .O(N__79966),
            .I(N__79963));
    LocalMux I__14631 (
            .O(N__79963),
            .I(shift_srl_165Z0Z_13));
    InMux I__14630 (
            .O(N__79960),
            .I(N__79957));
    LocalMux I__14629 (
            .O(N__79957),
            .I(shift_srl_165Z0Z_14));
    InMux I__14628 (
            .O(N__79954),
            .I(N__79951));
    LocalMux I__14627 (
            .O(N__79951),
            .I(shift_srl_165Z0Z_9));
    InMux I__14626 (
            .O(N__79948),
            .I(N__79945));
    LocalMux I__14625 (
            .O(N__79945),
            .I(shift_srl_165Z0Z_8));
    InMux I__14624 (
            .O(N__79942),
            .I(N__79939));
    LocalMux I__14623 (
            .O(N__79939),
            .I(shift_srl_165Z0Z_0));
    IoInMux I__14622 (
            .O(N__79936),
            .I(N__79933));
    LocalMux I__14621 (
            .O(N__79933),
            .I(N__79930));
    Span4Mux_s1_h I__14620 (
            .O(N__79930),
            .I(N__79926));
    InMux I__14619 (
            .O(N__79929),
            .I(N__79923));
    Sp12to4 I__14618 (
            .O(N__79926),
            .I(N__79920));
    LocalMux I__14617 (
            .O(N__79923),
            .I(N__79917));
    Span12Mux_v I__14616 (
            .O(N__79920),
            .I(N__79913));
    Span4Mux_v I__14615 (
            .O(N__79917),
            .I(N__79910));
    InMux I__14614 (
            .O(N__79916),
            .I(N__79907));
    Span12Mux_h I__14613 (
            .O(N__79913),
            .I(N__79900));
    Sp12to4 I__14612 (
            .O(N__79910),
            .I(N__79900));
    LocalMux I__14611 (
            .O(N__79907),
            .I(N__79900));
    Odrv12 I__14610 (
            .O(N__79900),
            .I(rco_c_29));
    CEMux I__14609 (
            .O(N__79897),
            .I(N__79894));
    LocalMux I__14608 (
            .O(N__79894),
            .I(N__79890));
    CEMux I__14607 (
            .O(N__79893),
            .I(N__79887));
    Span4Mux_v I__14606 (
            .O(N__79890),
            .I(N__79882));
    LocalMux I__14605 (
            .O(N__79887),
            .I(N__79882));
    Span4Mux_v I__14604 (
            .O(N__79882),
            .I(N__79879));
    Odrv4 I__14603 (
            .O(N__79879),
            .I(clk_en_31));
    InMux I__14602 (
            .O(N__79876),
            .I(N__79873));
    LocalMux I__14601 (
            .O(N__79873),
            .I(shift_srl_30Z0Z_14));
    InMux I__14600 (
            .O(N__79870),
            .I(N__79867));
    LocalMux I__14599 (
            .O(N__79867),
            .I(shift_srl_30Z0Z_13));
    InMux I__14598 (
            .O(N__79864),
            .I(N__79861));
    LocalMux I__14597 (
            .O(N__79861),
            .I(shift_srl_30Z0Z_12));
    InMux I__14596 (
            .O(N__79858),
            .I(N__79855));
    LocalMux I__14595 (
            .O(N__79855),
            .I(shift_srl_30Z0Z_11));
    InMux I__14594 (
            .O(N__79852),
            .I(N__79849));
    LocalMux I__14593 (
            .O(N__79849),
            .I(shift_srl_30Z0Z_10));
    InMux I__14592 (
            .O(N__79846),
            .I(N__79843));
    LocalMux I__14591 (
            .O(N__79843),
            .I(shift_srl_30Z0Z_8));
    InMux I__14590 (
            .O(N__79840),
            .I(N__79837));
    LocalMux I__14589 (
            .O(N__79837),
            .I(shift_srl_30Z0Z_9));
    CEMux I__14588 (
            .O(N__79834),
            .I(N__79831));
    LocalMux I__14587 (
            .O(N__79831),
            .I(N__79827));
    CEMux I__14586 (
            .O(N__79830),
            .I(N__79824));
    Span4Mux_h I__14585 (
            .O(N__79827),
            .I(N__79820));
    LocalMux I__14584 (
            .O(N__79824),
            .I(N__79817));
    CEMux I__14583 (
            .O(N__79823),
            .I(N__79814));
    Span4Mux_v I__14582 (
            .O(N__79820),
            .I(N__79811));
    Span4Mux_h I__14581 (
            .O(N__79817),
            .I(N__79808));
    LocalMux I__14580 (
            .O(N__79814),
            .I(N__79805));
    Odrv4 I__14579 (
            .O(N__79811),
            .I(clk_en_30));
    Odrv4 I__14578 (
            .O(N__79808),
            .I(clk_en_30));
    Odrv4 I__14577 (
            .O(N__79805),
            .I(clk_en_30));
    InMux I__14576 (
            .O(N__79798),
            .I(N__79795));
    LocalMux I__14575 (
            .O(N__79795),
            .I(shift_srl_65Z0Z_6));
    InMux I__14574 (
            .O(N__79792),
            .I(N__79789));
    LocalMux I__14573 (
            .O(N__79789),
            .I(shift_srl_65Z0Z_7));
    CEMux I__14572 (
            .O(N__79786),
            .I(N__79782));
    CEMux I__14571 (
            .O(N__79785),
            .I(N__79779));
    LocalMux I__14570 (
            .O(N__79782),
            .I(clk_en_65));
    LocalMux I__14569 (
            .O(N__79779),
            .I(clk_en_65));
    InMux I__14568 (
            .O(N__79774),
            .I(N__79771));
    LocalMux I__14567 (
            .O(N__79771),
            .I(N__79768));
    Span4Mux_h I__14566 (
            .O(N__79768),
            .I(N__79765));
    Odrv4 I__14565 (
            .O(N__79765),
            .I(shift_srl_30Z0Z_6));
    InMux I__14564 (
            .O(N__79762),
            .I(N__79758));
    InMux I__14563 (
            .O(N__79761),
            .I(N__79755));
    LocalMux I__14562 (
            .O(N__79758),
            .I(N__79751));
    LocalMux I__14561 (
            .O(N__79755),
            .I(N__79748));
    InMux I__14560 (
            .O(N__79754),
            .I(N__79745));
    Span4Mux_h I__14559 (
            .O(N__79751),
            .I(N__79741));
    Sp12to4 I__14558 (
            .O(N__79748),
            .I(N__79738));
    LocalMux I__14557 (
            .O(N__79745),
            .I(N__79735));
    InMux I__14556 (
            .O(N__79744),
            .I(N__79732));
    Span4Mux_h I__14555 (
            .O(N__79741),
            .I(N__79729));
    Span12Mux_v I__14554 (
            .O(N__79738),
            .I(N__79726));
    Span4Mux_h I__14553 (
            .O(N__79735),
            .I(N__79723));
    LocalMux I__14552 (
            .O(N__79732),
            .I(shift_srl_38Z0Z_15));
    Odrv4 I__14551 (
            .O(N__79729),
            .I(shift_srl_38Z0Z_15));
    Odrv12 I__14550 (
            .O(N__79726),
            .I(shift_srl_38Z0Z_15));
    Odrv4 I__14549 (
            .O(N__79723),
            .I(shift_srl_38Z0Z_15));
    IoInMux I__14548 (
            .O(N__79714),
            .I(N__79711));
    LocalMux I__14547 (
            .O(N__79711),
            .I(N__79708));
    Span12Mux_s9_h I__14546 (
            .O(N__79708),
            .I(N__79705));
    Odrv12 I__14545 (
            .O(N__79705),
            .I(rco_c_38));
    CascadeMux I__14544 (
            .O(N__79702),
            .I(rco_c_38_cascade_));
    InMux I__14543 (
            .O(N__79699),
            .I(N__79696));
    LocalMux I__14542 (
            .O(N__79696),
            .I(shift_srl_30Z0Z_7));
    InMux I__14541 (
            .O(N__79693),
            .I(N__79690));
    LocalMux I__14540 (
            .O(N__79690),
            .I(N__79685));
    InMux I__14539 (
            .O(N__79689),
            .I(N__79682));
    CascadeMux I__14538 (
            .O(N__79688),
            .I(N__79679));
    Span12Mux_h I__14537 (
            .O(N__79685),
            .I(N__79670));
    LocalMux I__14536 (
            .O(N__79682),
            .I(N__79667));
    InMux I__14535 (
            .O(N__79679),
            .I(N__79658));
    InMux I__14534 (
            .O(N__79678),
            .I(N__79658));
    InMux I__14533 (
            .O(N__79677),
            .I(N__79658));
    InMux I__14532 (
            .O(N__79676),
            .I(N__79658));
    InMux I__14531 (
            .O(N__79675),
            .I(N__79651));
    InMux I__14530 (
            .O(N__79674),
            .I(N__79651));
    InMux I__14529 (
            .O(N__79673),
            .I(N__79651));
    Odrv12 I__14528 (
            .O(N__79670),
            .I(shift_srl_100Z0Z_15));
    Odrv4 I__14527 (
            .O(N__79667),
            .I(shift_srl_100Z0Z_15));
    LocalMux I__14526 (
            .O(N__79658),
            .I(shift_srl_100Z0Z_15));
    LocalMux I__14525 (
            .O(N__79651),
            .I(shift_srl_100Z0Z_15));
    InMux I__14524 (
            .O(N__79642),
            .I(N__79639));
    LocalMux I__14523 (
            .O(N__79639),
            .I(N__79635));
    IoInMux I__14522 (
            .O(N__79638),
            .I(N__79632));
    Span4Mux_v I__14521 (
            .O(N__79635),
            .I(N__79629));
    LocalMux I__14520 (
            .O(N__79632),
            .I(N__79626));
    Sp12to4 I__14519 (
            .O(N__79629),
            .I(N__79623));
    IoSpan4Mux I__14518 (
            .O(N__79626),
            .I(N__79620));
    Span12Mux_h I__14517 (
            .O(N__79623),
            .I(N__79617));
    Span4Mux_s2_h I__14516 (
            .O(N__79620),
            .I(N__79614));
    Span12Mux_v I__14515 (
            .O(N__79617),
            .I(N__79609));
    Sp12to4 I__14514 (
            .O(N__79614),
            .I(N__79609));
    Odrv12 I__14513 (
            .O(N__79609),
            .I(rco_c_100));
    InMux I__14512 (
            .O(N__79606),
            .I(N__79603));
    LocalMux I__14511 (
            .O(N__79603),
            .I(N__79600));
    Span4Mux_v I__14510 (
            .O(N__79600),
            .I(N__79597));
    Sp12to4 I__14509 (
            .O(N__79597),
            .I(N__79592));
    InMux I__14508 (
            .O(N__79596),
            .I(N__79587));
    InMux I__14507 (
            .O(N__79595),
            .I(N__79587));
    Span12Mux_h I__14506 (
            .O(N__79592),
            .I(N__79579));
    LocalMux I__14505 (
            .O(N__79587),
            .I(N__79579));
    InMux I__14504 (
            .O(N__79586),
            .I(N__79572));
    InMux I__14503 (
            .O(N__79585),
            .I(N__79572));
    InMux I__14502 (
            .O(N__79584),
            .I(N__79572));
    Odrv12 I__14501 (
            .O(N__79579),
            .I(rco_int_0_a3_0_a2_out_0));
    LocalMux I__14500 (
            .O(N__79572),
            .I(rco_int_0_a3_0_a2_out_0));
    IoInMux I__14499 (
            .O(N__79567),
            .I(N__79564));
    LocalMux I__14498 (
            .O(N__79564),
            .I(N__79560));
    InMux I__14497 (
            .O(N__79563),
            .I(N__79557));
    Span4Mux_s2_v I__14496 (
            .O(N__79560),
            .I(N__79552));
    LocalMux I__14495 (
            .O(N__79557),
            .I(N__79538));
    InMux I__14494 (
            .O(N__79556),
            .I(N__79533));
    InMux I__14493 (
            .O(N__79555),
            .I(N__79533));
    Span4Mux_h I__14492 (
            .O(N__79552),
            .I(N__79522));
    InMux I__14491 (
            .O(N__79551),
            .I(N__79519));
    InMux I__14490 (
            .O(N__79550),
            .I(N__79512));
    InMux I__14489 (
            .O(N__79549),
            .I(N__79512));
    InMux I__14488 (
            .O(N__79548),
            .I(N__79512));
    InMux I__14487 (
            .O(N__79547),
            .I(N__79499));
    InMux I__14486 (
            .O(N__79546),
            .I(N__79499));
    InMux I__14485 (
            .O(N__79545),
            .I(N__79499));
    InMux I__14484 (
            .O(N__79544),
            .I(N__79499));
    InMux I__14483 (
            .O(N__79543),
            .I(N__79499));
    InMux I__14482 (
            .O(N__79542),
            .I(N__79493));
    InMux I__14481 (
            .O(N__79541),
            .I(N__79490));
    Span4Mux_h I__14480 (
            .O(N__79538),
            .I(N__79487));
    LocalMux I__14479 (
            .O(N__79533),
            .I(N__79484));
    InMux I__14478 (
            .O(N__79532),
            .I(N__79479));
    InMux I__14477 (
            .O(N__79531),
            .I(N__79476));
    InMux I__14476 (
            .O(N__79530),
            .I(N__79467));
    InMux I__14475 (
            .O(N__79529),
            .I(N__79467));
    InMux I__14474 (
            .O(N__79528),
            .I(N__79467));
    InMux I__14473 (
            .O(N__79527),
            .I(N__79467));
    InMux I__14472 (
            .O(N__79526),
            .I(N__79459));
    InMux I__14471 (
            .O(N__79525),
            .I(N__79459));
    Span4Mux_h I__14470 (
            .O(N__79522),
            .I(N__79456));
    LocalMux I__14469 (
            .O(N__79519),
            .I(N__79452));
    LocalMux I__14468 (
            .O(N__79512),
            .I(N__79449));
    InMux I__14467 (
            .O(N__79511),
            .I(N__79446));
    InMux I__14466 (
            .O(N__79510),
            .I(N__79443));
    LocalMux I__14465 (
            .O(N__79499),
            .I(N__79440));
    InMux I__14464 (
            .O(N__79498),
            .I(N__79437));
    InMux I__14463 (
            .O(N__79497),
            .I(N__79432));
    InMux I__14462 (
            .O(N__79496),
            .I(N__79432));
    LocalMux I__14461 (
            .O(N__79493),
            .I(N__79427));
    LocalMux I__14460 (
            .O(N__79490),
            .I(N__79427));
    Span4Mux_v I__14459 (
            .O(N__79487),
            .I(N__79422));
    Span4Mux_h I__14458 (
            .O(N__79484),
            .I(N__79422));
    InMux I__14457 (
            .O(N__79483),
            .I(N__79417));
    InMux I__14456 (
            .O(N__79482),
            .I(N__79417));
    LocalMux I__14455 (
            .O(N__79479),
            .I(N__79412));
    LocalMux I__14454 (
            .O(N__79476),
            .I(N__79409));
    LocalMux I__14453 (
            .O(N__79467),
            .I(N__79406));
    InMux I__14452 (
            .O(N__79466),
            .I(N__79399));
    InMux I__14451 (
            .O(N__79465),
            .I(N__79399));
    InMux I__14450 (
            .O(N__79464),
            .I(N__79399));
    LocalMux I__14449 (
            .O(N__79459),
            .I(N__79393));
    Sp12to4 I__14448 (
            .O(N__79456),
            .I(N__79386));
    InMux I__14447 (
            .O(N__79455),
            .I(N__79383));
    Span4Mux_h I__14446 (
            .O(N__79452),
            .I(N__79380));
    Span4Mux_v I__14445 (
            .O(N__79449),
            .I(N__79375));
    LocalMux I__14444 (
            .O(N__79446),
            .I(N__79375));
    LocalMux I__14443 (
            .O(N__79443),
            .I(N__79366));
    Span4Mux_v I__14442 (
            .O(N__79440),
            .I(N__79366));
    LocalMux I__14441 (
            .O(N__79437),
            .I(N__79366));
    LocalMux I__14440 (
            .O(N__79432),
            .I(N__79366));
    Span4Mux_v I__14439 (
            .O(N__79427),
            .I(N__79359));
    Span4Mux_v I__14438 (
            .O(N__79422),
            .I(N__79359));
    LocalMux I__14437 (
            .O(N__79417),
            .I(N__79359));
    InMux I__14436 (
            .O(N__79416),
            .I(N__79356));
    InMux I__14435 (
            .O(N__79415),
            .I(N__79353));
    Span4Mux_h I__14434 (
            .O(N__79412),
            .I(N__79348));
    Span4Mux_v I__14433 (
            .O(N__79409),
            .I(N__79348));
    Span4Mux_v I__14432 (
            .O(N__79406),
            .I(N__79343));
    LocalMux I__14431 (
            .O(N__79399),
            .I(N__79343));
    InMux I__14430 (
            .O(N__79398),
            .I(N__79336));
    InMux I__14429 (
            .O(N__79397),
            .I(N__79336));
    InMux I__14428 (
            .O(N__79396),
            .I(N__79336));
    Span4Mux_v I__14427 (
            .O(N__79393),
            .I(N__79331));
    InMux I__14426 (
            .O(N__79392),
            .I(N__79328));
    InMux I__14425 (
            .O(N__79391),
            .I(N__79325));
    InMux I__14424 (
            .O(N__79390),
            .I(N__79322));
    InMux I__14423 (
            .O(N__79389),
            .I(N__79317));
    Span12Mux_v I__14422 (
            .O(N__79386),
            .I(N__79314));
    LocalMux I__14421 (
            .O(N__79383),
            .I(N__79311));
    Span4Mux_h I__14420 (
            .O(N__79380),
            .I(N__79300));
    Span4Mux_v I__14419 (
            .O(N__79375),
            .I(N__79300));
    Span4Mux_v I__14418 (
            .O(N__79366),
            .I(N__79300));
    Span4Mux_v I__14417 (
            .O(N__79359),
            .I(N__79300));
    LocalMux I__14416 (
            .O(N__79356),
            .I(N__79300));
    LocalMux I__14415 (
            .O(N__79353),
            .I(N__79291));
    Span4Mux_h I__14414 (
            .O(N__79348),
            .I(N__79291));
    Span4Mux_v I__14413 (
            .O(N__79343),
            .I(N__79291));
    LocalMux I__14412 (
            .O(N__79336),
            .I(N__79291));
    InMux I__14411 (
            .O(N__79335),
            .I(N__79286));
    InMux I__14410 (
            .O(N__79334),
            .I(N__79286));
    Sp12to4 I__14409 (
            .O(N__79331),
            .I(N__79277));
    LocalMux I__14408 (
            .O(N__79328),
            .I(N__79277));
    LocalMux I__14407 (
            .O(N__79325),
            .I(N__79277));
    LocalMux I__14406 (
            .O(N__79322),
            .I(N__79277));
    InMux I__14405 (
            .O(N__79321),
            .I(N__79272));
    InMux I__14404 (
            .O(N__79320),
            .I(N__79272));
    LocalMux I__14403 (
            .O(N__79317),
            .I(N__79269));
    Odrv12 I__14402 (
            .O(N__79314),
            .I(rco_c_99));
    Odrv4 I__14401 (
            .O(N__79311),
            .I(rco_c_99));
    Odrv4 I__14400 (
            .O(N__79300),
            .I(rco_c_99));
    Odrv4 I__14399 (
            .O(N__79291),
            .I(rco_c_99));
    LocalMux I__14398 (
            .O(N__79286),
            .I(rco_c_99));
    Odrv12 I__14397 (
            .O(N__79277),
            .I(rco_c_99));
    LocalMux I__14396 (
            .O(N__79272),
            .I(rco_c_99));
    Odrv12 I__14395 (
            .O(N__79269),
            .I(rco_c_99));
    InMux I__14394 (
            .O(N__79252),
            .I(N__79249));
    LocalMux I__14393 (
            .O(N__79249),
            .I(N__79245));
    IoInMux I__14392 (
            .O(N__79248),
            .I(N__79242));
    Span4Mux_v I__14391 (
            .O(N__79245),
            .I(N__79239));
    LocalMux I__14390 (
            .O(N__79242),
            .I(N__79236));
    Sp12to4 I__14389 (
            .O(N__79239),
            .I(N__79233));
    Span4Mux_s1_h I__14388 (
            .O(N__79236),
            .I(N__79230));
    Span12Mux_h I__14387 (
            .O(N__79233),
            .I(N__79227));
    Span4Mux_h I__14386 (
            .O(N__79230),
            .I(N__79224));
    Span12Mux_v I__14385 (
            .O(N__79227),
            .I(N__79221));
    Span4Mux_h I__14384 (
            .O(N__79224),
            .I(N__79218));
    Odrv12 I__14383 (
            .O(N__79221),
            .I(rco_c_104));
    Odrv4 I__14382 (
            .O(N__79218),
            .I(rco_c_104));
    InMux I__14381 (
            .O(N__79213),
            .I(N__79210));
    LocalMux I__14380 (
            .O(N__79210),
            .I(shift_srl_63Z0Z_11));
    InMux I__14379 (
            .O(N__79207),
            .I(N__79204));
    LocalMux I__14378 (
            .O(N__79204),
            .I(N__79201));
    Odrv4 I__14377 (
            .O(N__79201),
            .I(shift_srl_63Z0Z_9));
    InMux I__14376 (
            .O(N__79198),
            .I(N__79195));
    LocalMux I__14375 (
            .O(N__79195),
            .I(shift_srl_63Z0Z_10));
    CEMux I__14374 (
            .O(N__79192),
            .I(N__79188));
    CEMux I__14373 (
            .O(N__79191),
            .I(N__79185));
    LocalMux I__14372 (
            .O(N__79188),
            .I(N__79181));
    LocalMux I__14371 (
            .O(N__79185),
            .I(N__79178));
    CEMux I__14370 (
            .O(N__79184),
            .I(N__79175));
    Span4Mux_h I__14369 (
            .O(N__79181),
            .I(N__79172));
    Span4Mux_h I__14368 (
            .O(N__79178),
            .I(N__79167));
    LocalMux I__14367 (
            .O(N__79175),
            .I(N__79167));
    Odrv4 I__14366 (
            .O(N__79172),
            .I(clk_en_63));
    Odrv4 I__14365 (
            .O(N__79167),
            .I(clk_en_63));
    InMux I__14364 (
            .O(N__79162),
            .I(N__79159));
    LocalMux I__14363 (
            .O(N__79159),
            .I(shift_srl_65Z0Z_0));
    InMux I__14362 (
            .O(N__79156),
            .I(N__79153));
    LocalMux I__14361 (
            .O(N__79153),
            .I(shift_srl_65Z0Z_1));
    InMux I__14360 (
            .O(N__79150),
            .I(N__79147));
    LocalMux I__14359 (
            .O(N__79147),
            .I(shift_srl_65Z0Z_2));
    InMux I__14358 (
            .O(N__79144),
            .I(N__79141));
    LocalMux I__14357 (
            .O(N__79141),
            .I(shift_srl_65Z0Z_3));
    InMux I__14356 (
            .O(N__79138),
            .I(N__79135));
    LocalMux I__14355 (
            .O(N__79135),
            .I(shift_srl_65Z0Z_4));
    InMux I__14354 (
            .O(N__79132),
            .I(N__79129));
    LocalMux I__14353 (
            .O(N__79129),
            .I(shift_srl_65Z0Z_5));
    InMux I__14352 (
            .O(N__79126),
            .I(N__79123));
    LocalMux I__14351 (
            .O(N__79123),
            .I(shift_srl_64Z0Z_4));
    InMux I__14350 (
            .O(N__79120),
            .I(N__79117));
    LocalMux I__14349 (
            .O(N__79117),
            .I(shift_srl_64Z0Z_5));
    InMux I__14348 (
            .O(N__79114),
            .I(N__79111));
    LocalMux I__14347 (
            .O(N__79111),
            .I(shift_srl_64Z0Z_6));
    InMux I__14346 (
            .O(N__79108),
            .I(N__79105));
    LocalMux I__14345 (
            .O(N__79105),
            .I(shift_srl_64Z0Z_7));
    CEMux I__14344 (
            .O(N__79102),
            .I(N__79098));
    CEMux I__14343 (
            .O(N__79101),
            .I(N__79095));
    LocalMux I__14342 (
            .O(N__79098),
            .I(N__79092));
    LocalMux I__14341 (
            .O(N__79095),
            .I(N__79089));
    Span4Mux_v I__14340 (
            .O(N__79092),
            .I(N__79086));
    Odrv12 I__14339 (
            .O(N__79089),
            .I(clk_en_64));
    Odrv4 I__14338 (
            .O(N__79086),
            .I(clk_en_64));
    CEMux I__14337 (
            .O(N__79081),
            .I(N__79076));
    CEMux I__14336 (
            .O(N__79080),
            .I(N__79072));
    InMux I__14335 (
            .O(N__79079),
            .I(N__79069));
    LocalMux I__14334 (
            .O(N__79076),
            .I(N__79066));
    CEMux I__14333 (
            .O(N__79075),
            .I(N__79063));
    LocalMux I__14332 (
            .O(N__79072),
            .I(N__79060));
    LocalMux I__14331 (
            .O(N__79069),
            .I(N__79057));
    Span4Mux_v I__14330 (
            .O(N__79066),
            .I(N__79054));
    LocalMux I__14329 (
            .O(N__79063),
            .I(N__79051));
    Span4Mux_h I__14328 (
            .O(N__79060),
            .I(N__79048));
    Span4Mux_v I__14327 (
            .O(N__79057),
            .I(N__79045));
    Odrv4 I__14326 (
            .O(N__79054),
            .I(clk_en_60));
    Odrv12 I__14325 (
            .O(N__79051),
            .I(clk_en_60));
    Odrv4 I__14324 (
            .O(N__79048),
            .I(clk_en_60));
    Odrv4 I__14323 (
            .O(N__79045),
            .I(clk_en_60));
    InMux I__14322 (
            .O(N__79036),
            .I(N__79033));
    LocalMux I__14321 (
            .O(N__79033),
            .I(shift_srl_63Z0Z_14));
    InMux I__14320 (
            .O(N__79030),
            .I(N__79027));
    LocalMux I__14319 (
            .O(N__79027),
            .I(shift_srl_63Z0Z_13));
    InMux I__14318 (
            .O(N__79024),
            .I(N__79021));
    LocalMux I__14317 (
            .O(N__79021),
            .I(shift_srl_63Z0Z_12));
    InMux I__14316 (
            .O(N__79018),
            .I(N__79015));
    LocalMux I__14315 (
            .O(N__79015),
            .I(shift_srl_58Z0Z_13));
    InMux I__14314 (
            .O(N__79012),
            .I(N__79009));
    LocalMux I__14313 (
            .O(N__79009),
            .I(shift_srl_58Z0Z_14));
    InMux I__14312 (
            .O(N__79006),
            .I(N__79003));
    LocalMux I__14311 (
            .O(N__79003),
            .I(N__78999));
    InMux I__14310 (
            .O(N__79002),
            .I(N__78996));
    Span4Mux_h I__14309 (
            .O(N__78999),
            .I(N__78993));
    LocalMux I__14308 (
            .O(N__78996),
            .I(shift_srl_58Z0Z_15));
    Odrv4 I__14307 (
            .O(N__78993),
            .I(shift_srl_58Z0Z_15));
    InMux I__14306 (
            .O(N__78988),
            .I(N__78985));
    LocalMux I__14305 (
            .O(N__78985),
            .I(shift_srl_58Z0Z_9));
    InMux I__14304 (
            .O(N__78982),
            .I(N__78979));
    LocalMux I__14303 (
            .O(N__78979),
            .I(shift_srl_58Z0Z_7));
    InMux I__14302 (
            .O(N__78976),
            .I(N__78973));
    LocalMux I__14301 (
            .O(N__78973),
            .I(shift_srl_58Z0Z_8));
    CEMux I__14300 (
            .O(N__78970),
            .I(N__78966));
    CEMux I__14299 (
            .O(N__78969),
            .I(N__78963));
    LocalMux I__14298 (
            .O(N__78966),
            .I(clk_en_58));
    LocalMux I__14297 (
            .O(N__78963),
            .I(clk_en_58));
    InMux I__14296 (
            .O(N__78958),
            .I(N__78955));
    LocalMux I__14295 (
            .O(N__78955),
            .I(shift_srl_64Z0Z_0));
    InMux I__14294 (
            .O(N__78952),
            .I(N__78949));
    LocalMux I__14293 (
            .O(N__78949),
            .I(shift_srl_64Z0Z_1));
    InMux I__14292 (
            .O(N__78946),
            .I(N__78943));
    LocalMux I__14291 (
            .O(N__78943),
            .I(shift_srl_64Z0Z_2));
    InMux I__14290 (
            .O(N__78940),
            .I(N__78937));
    LocalMux I__14289 (
            .O(N__78937),
            .I(shift_srl_64Z0Z_3));
    InMux I__14288 (
            .O(N__78934),
            .I(N__78931));
    LocalMux I__14287 (
            .O(N__78931),
            .I(shift_srl_58Z0Z_1));
    InMux I__14286 (
            .O(N__78928),
            .I(N__78925));
    LocalMux I__14285 (
            .O(N__78925),
            .I(shift_srl_58Z0Z_2));
    InMux I__14284 (
            .O(N__78922),
            .I(N__78919));
    LocalMux I__14283 (
            .O(N__78919),
            .I(shift_srl_58Z0Z_3));
    InMux I__14282 (
            .O(N__78916),
            .I(N__78913));
    LocalMux I__14281 (
            .O(N__78913),
            .I(shift_srl_58Z0Z_4));
    InMux I__14280 (
            .O(N__78910),
            .I(N__78907));
    LocalMux I__14279 (
            .O(N__78907),
            .I(shift_srl_58Z0Z_5));
    InMux I__14278 (
            .O(N__78904),
            .I(N__78901));
    LocalMux I__14277 (
            .O(N__78901),
            .I(shift_srl_58Z0Z_6));
    InMux I__14276 (
            .O(N__78898),
            .I(N__78895));
    LocalMux I__14275 (
            .O(N__78895),
            .I(shift_srl_58Z0Z_10));
    InMux I__14274 (
            .O(N__78892),
            .I(N__78889));
    LocalMux I__14273 (
            .O(N__78889),
            .I(shift_srl_58Z0Z_11));
    InMux I__14272 (
            .O(N__78886),
            .I(N__78883));
    LocalMux I__14271 (
            .O(N__78883),
            .I(shift_srl_58Z0Z_12));
    InMux I__14270 (
            .O(N__78880),
            .I(N__78877));
    LocalMux I__14269 (
            .O(N__78877),
            .I(shift_srl_56Z0Z_1));
    InMux I__14268 (
            .O(N__78874),
            .I(N__78871));
    LocalMux I__14267 (
            .O(N__78871),
            .I(shift_srl_56Z0Z_6));
    InMux I__14266 (
            .O(N__78868),
            .I(N__78865));
    LocalMux I__14265 (
            .O(N__78865),
            .I(shift_srl_56Z0Z_2));
    InMux I__14264 (
            .O(N__78862),
            .I(N__78859));
    LocalMux I__14263 (
            .O(N__78859),
            .I(shift_srl_56Z0Z_5));
    InMux I__14262 (
            .O(N__78856),
            .I(N__78853));
    LocalMux I__14261 (
            .O(N__78853),
            .I(shift_srl_56Z0Z_3));
    InMux I__14260 (
            .O(N__78850),
            .I(N__78847));
    LocalMux I__14259 (
            .O(N__78847),
            .I(shift_srl_56Z0Z_4));
    InMux I__14258 (
            .O(N__78844),
            .I(N__78841));
    LocalMux I__14257 (
            .O(N__78841),
            .I(shift_srl_56Z0Z_7));
    InMux I__14256 (
            .O(N__78838),
            .I(N__78835));
    LocalMux I__14255 (
            .O(N__78835),
            .I(N__78832));
    Odrv4 I__14254 (
            .O(N__78832),
            .I(shift_srl_56Z0Z_8));
    CEMux I__14253 (
            .O(N__78829),
            .I(N__78825));
    CEMux I__14252 (
            .O(N__78828),
            .I(N__78822));
    LocalMux I__14251 (
            .O(N__78825),
            .I(N__78819));
    LocalMux I__14250 (
            .O(N__78822),
            .I(N__78816));
    Span4Mux_h I__14249 (
            .O(N__78819),
            .I(N__78813));
    Sp12to4 I__14248 (
            .O(N__78816),
            .I(N__78810));
    Odrv4 I__14247 (
            .O(N__78813),
            .I(clk_en_56));
    Odrv12 I__14246 (
            .O(N__78810),
            .I(clk_en_56));
    InMux I__14245 (
            .O(N__78805),
            .I(N__78802));
    LocalMux I__14244 (
            .O(N__78802),
            .I(shift_srl_58Z0Z_0));
    InMux I__14243 (
            .O(N__78799),
            .I(N__78794));
    InMux I__14242 (
            .O(N__78798),
            .I(N__78790));
    InMux I__14241 (
            .O(N__78797),
            .I(N__78787));
    LocalMux I__14240 (
            .O(N__78794),
            .I(N__78783));
    InMux I__14239 (
            .O(N__78793),
            .I(N__78780));
    LocalMux I__14238 (
            .O(N__78790),
            .I(N__78775));
    LocalMux I__14237 (
            .O(N__78787),
            .I(N__78772));
    InMux I__14236 (
            .O(N__78786),
            .I(N__78769));
    Span4Mux_v I__14235 (
            .O(N__78783),
            .I(N__78764));
    LocalMux I__14234 (
            .O(N__78780),
            .I(N__78764));
    InMux I__14233 (
            .O(N__78779),
            .I(N__78759));
    InMux I__14232 (
            .O(N__78778),
            .I(N__78759));
    Span4Mux_h I__14231 (
            .O(N__78775),
            .I(N__78754));
    Span4Mux_v I__14230 (
            .O(N__78772),
            .I(N__78754));
    LocalMux I__14229 (
            .O(N__78769),
            .I(shift_srl_41Z0Z_15));
    Odrv4 I__14228 (
            .O(N__78764),
            .I(shift_srl_41Z0Z_15));
    LocalMux I__14227 (
            .O(N__78759),
            .I(shift_srl_41Z0Z_15));
    Odrv4 I__14226 (
            .O(N__78754),
            .I(shift_srl_41Z0Z_15));
    InMux I__14225 (
            .O(N__78745),
            .I(N__78742));
    LocalMux I__14224 (
            .O(N__78742),
            .I(shift_srl_41Z0Z_0));
    InMux I__14223 (
            .O(N__78739),
            .I(N__78736));
    LocalMux I__14222 (
            .O(N__78736),
            .I(shift_srl_41Z0Z_1));
    InMux I__14221 (
            .O(N__78733),
            .I(N__78730));
    LocalMux I__14220 (
            .O(N__78730),
            .I(shift_srl_41Z0Z_2));
    InMux I__14219 (
            .O(N__78727),
            .I(N__78724));
    LocalMux I__14218 (
            .O(N__78724),
            .I(shift_srl_41Z0Z_3));
    InMux I__14217 (
            .O(N__78721),
            .I(N__78718));
    LocalMux I__14216 (
            .O(N__78718),
            .I(shift_srl_41Z0Z_4));
    InMux I__14215 (
            .O(N__78715),
            .I(N__78712));
    LocalMux I__14214 (
            .O(N__78712),
            .I(shift_srl_41Z0Z_5));
    InMux I__14213 (
            .O(N__78709),
            .I(N__78706));
    LocalMux I__14212 (
            .O(N__78706),
            .I(shift_srl_41Z0Z_6));
    InMux I__14211 (
            .O(N__78703),
            .I(N__78700));
    LocalMux I__14210 (
            .O(N__78700),
            .I(N__78697));
    Span4Mux_h I__14209 (
            .O(N__78697),
            .I(N__78694));
    Odrv4 I__14208 (
            .O(N__78694),
            .I(shift_srl_41Z0Z_7));
    CEMux I__14207 (
            .O(N__78691),
            .I(N__78688));
    LocalMux I__14206 (
            .O(N__78688),
            .I(N__78684));
    CEMux I__14205 (
            .O(N__78687),
            .I(N__78681));
    Span4Mux_h I__14204 (
            .O(N__78684),
            .I(N__78676));
    LocalMux I__14203 (
            .O(N__78681),
            .I(N__78676));
    Span4Mux_v I__14202 (
            .O(N__78676),
            .I(N__78673));
    Odrv4 I__14201 (
            .O(N__78673),
            .I(clk_en_41));
    InMux I__14200 (
            .O(N__78670),
            .I(N__78667));
    LocalMux I__14199 (
            .O(N__78667),
            .I(N__78664));
    Odrv12 I__14198 (
            .O(N__78664),
            .I(shift_srl_56Z0Z_0));
    InMux I__14197 (
            .O(N__78661),
            .I(N__78658));
    LocalMux I__14196 (
            .O(N__78658),
            .I(shift_srl_83Z0Z_5));
    InMux I__14195 (
            .O(N__78655),
            .I(N__78652));
    LocalMux I__14194 (
            .O(N__78652),
            .I(shift_srl_83Z0Z_6));
    InMux I__14193 (
            .O(N__78649),
            .I(N__78646));
    LocalMux I__14192 (
            .O(N__78646),
            .I(shift_srl_82Z0Z_0));
    InMux I__14191 (
            .O(N__78643),
            .I(N__78640));
    LocalMux I__14190 (
            .O(N__78640),
            .I(shift_srl_82Z0Z_1));
    InMux I__14189 (
            .O(N__78637),
            .I(N__78634));
    LocalMux I__14188 (
            .O(N__78634),
            .I(shift_srl_82Z0Z_2));
    InMux I__14187 (
            .O(N__78631),
            .I(N__78628));
    LocalMux I__14186 (
            .O(N__78628),
            .I(shift_srl_82Z0Z_3));
    InMux I__14185 (
            .O(N__78625),
            .I(N__78622));
    LocalMux I__14184 (
            .O(N__78622),
            .I(shift_srl_82Z0Z_4));
    InMux I__14183 (
            .O(N__78619),
            .I(N__78616));
    LocalMux I__14182 (
            .O(N__78616),
            .I(shift_srl_82Z0Z_5));
    InMux I__14181 (
            .O(N__78613),
            .I(N__78610));
    LocalMux I__14180 (
            .O(N__78610),
            .I(shift_srl_82Z0Z_6));
    InMux I__14179 (
            .O(N__78607),
            .I(N__78604));
    LocalMux I__14178 (
            .O(N__78604),
            .I(shift_srl_83Z0Z_14));
    InMux I__14177 (
            .O(N__78601),
            .I(N__78598));
    LocalMux I__14176 (
            .O(N__78598),
            .I(shift_srl_83Z0Z_11));
    InMux I__14175 (
            .O(N__78595),
            .I(N__78592));
    LocalMux I__14174 (
            .O(N__78592),
            .I(shift_srl_83Z0Z_0));
    InMux I__14173 (
            .O(N__78589),
            .I(N__78586));
    LocalMux I__14172 (
            .O(N__78586),
            .I(shift_srl_83Z0Z_1));
    InMux I__14171 (
            .O(N__78583),
            .I(N__78580));
    LocalMux I__14170 (
            .O(N__78580),
            .I(shift_srl_83Z0Z_2));
    InMux I__14169 (
            .O(N__78577),
            .I(N__78574));
    LocalMux I__14168 (
            .O(N__78574),
            .I(shift_srl_83Z0Z_3));
    InMux I__14167 (
            .O(N__78571),
            .I(N__78568));
    LocalMux I__14166 (
            .O(N__78568),
            .I(shift_srl_83Z0Z_7));
    InMux I__14165 (
            .O(N__78565),
            .I(N__78562));
    LocalMux I__14164 (
            .O(N__78562),
            .I(shift_srl_83Z0Z_4));
    InMux I__14163 (
            .O(N__78559),
            .I(N__78556));
    LocalMux I__14162 (
            .O(N__78556),
            .I(shift_srl_176Z0Z_4));
    InMux I__14161 (
            .O(N__78553),
            .I(N__78550));
    LocalMux I__14160 (
            .O(N__78550),
            .I(shift_srl_176Z0Z_5));
    InMux I__14159 (
            .O(N__78547),
            .I(N__78544));
    LocalMux I__14158 (
            .O(N__78544),
            .I(shift_srl_176Z0Z_6));
    InMux I__14157 (
            .O(N__78541),
            .I(N__78538));
    LocalMux I__14156 (
            .O(N__78538),
            .I(N__78535));
    Odrv4 I__14155 (
            .O(N__78535),
            .I(shift_srl_176Z0Z_7));
    CEMux I__14154 (
            .O(N__78532),
            .I(N__78528));
    CEMux I__14153 (
            .O(N__78531),
            .I(N__78525));
    LocalMux I__14152 (
            .O(N__78528),
            .I(clk_en_176));
    LocalMux I__14151 (
            .O(N__78525),
            .I(clk_en_176));
    InMux I__14150 (
            .O(N__78520),
            .I(N__78516));
    IoInMux I__14149 (
            .O(N__78519),
            .I(N__78513));
    LocalMux I__14148 (
            .O(N__78516),
            .I(N__78510));
    LocalMux I__14147 (
            .O(N__78513),
            .I(N__78505));
    Span4Mux_v I__14146 (
            .O(N__78510),
            .I(N__78502));
    InMux I__14145 (
            .O(N__78509),
            .I(N__78497));
    InMux I__14144 (
            .O(N__78508),
            .I(N__78497));
    Span12Mux_s3_v I__14143 (
            .O(N__78505),
            .I(N__78492));
    Sp12to4 I__14142 (
            .O(N__78502),
            .I(N__78492));
    LocalMux I__14141 (
            .O(N__78497),
            .I(N__78489));
    Span12Mux_h I__14140 (
            .O(N__78492),
            .I(N__78486));
    Span4Mux_v I__14139 (
            .O(N__78489),
            .I(N__78483));
    Odrv12 I__14138 (
            .O(N__78486),
            .I(rco_c_120));
    Odrv4 I__14137 (
            .O(N__78483),
            .I(rco_c_120));
    InMux I__14136 (
            .O(N__78478),
            .I(N__78475));
    LocalMux I__14135 (
            .O(N__78475),
            .I(N__78469));
    InMux I__14134 (
            .O(N__78474),
            .I(N__78466));
    InMux I__14133 (
            .O(N__78473),
            .I(N__78463));
    CascadeMux I__14132 (
            .O(N__78472),
            .I(N__78460));
    Span12Mux_s7_v I__14131 (
            .O(N__78469),
            .I(N__78457));
    LocalMux I__14130 (
            .O(N__78466),
            .I(N__78454));
    LocalMux I__14129 (
            .O(N__78463),
            .I(N__78451));
    InMux I__14128 (
            .O(N__78460),
            .I(N__78448));
    Span12Mux_h I__14127 (
            .O(N__78457),
            .I(N__78443));
    Span12Mux_v I__14126 (
            .O(N__78454),
            .I(N__78440));
    Span4Mux_h I__14125 (
            .O(N__78451),
            .I(N__78437));
    LocalMux I__14124 (
            .O(N__78448),
            .I(N__78434));
    InMux I__14123 (
            .O(N__78447),
            .I(N__78431));
    InMux I__14122 (
            .O(N__78446),
            .I(N__78428));
    Odrv12 I__14121 (
            .O(N__78443),
            .I(shift_srl_121Z0Z_15));
    Odrv12 I__14120 (
            .O(N__78440),
            .I(shift_srl_121Z0Z_15));
    Odrv4 I__14119 (
            .O(N__78437),
            .I(shift_srl_121Z0Z_15));
    Odrv4 I__14118 (
            .O(N__78434),
            .I(shift_srl_121Z0Z_15));
    LocalMux I__14117 (
            .O(N__78431),
            .I(shift_srl_121Z0Z_15));
    LocalMux I__14116 (
            .O(N__78428),
            .I(shift_srl_121Z0Z_15));
    IoInMux I__14115 (
            .O(N__78415),
            .I(N__78412));
    LocalMux I__14114 (
            .O(N__78412),
            .I(N__78409));
    Span4Mux_s1_v I__14113 (
            .O(N__78409),
            .I(N__78406));
    Odrv4 I__14112 (
            .O(N__78406),
            .I(rco_c_121));
    IoInMux I__14111 (
            .O(N__78403),
            .I(N__78400));
    LocalMux I__14110 (
            .O(N__78400),
            .I(N__78397));
    Span4Mux_s3_v I__14109 (
            .O(N__78397),
            .I(N__78394));
    Span4Mux_h I__14108 (
            .O(N__78394),
            .I(N__78391));
    Odrv4 I__14107 (
            .O(N__78391),
            .I(rco_c_177));
    InMux I__14106 (
            .O(N__78388),
            .I(N__78385));
    LocalMux I__14105 (
            .O(N__78385),
            .I(shift_srl_83Z0Z_12));
    InMux I__14104 (
            .O(N__78382),
            .I(N__78379));
    LocalMux I__14103 (
            .O(N__78379),
            .I(shift_srl_83Z0Z_13));
    InMux I__14102 (
            .O(N__78376),
            .I(N__78373));
    LocalMux I__14101 (
            .O(N__78373),
            .I(shift_srl_188Z0Z_3));
    InMux I__14100 (
            .O(N__78370),
            .I(N__78367));
    LocalMux I__14099 (
            .O(N__78367),
            .I(shift_srl_188Z0Z_4));
    InMux I__14098 (
            .O(N__78364),
            .I(N__78361));
    LocalMux I__14097 (
            .O(N__78361),
            .I(shift_srl_188Z0Z_5));
    InMux I__14096 (
            .O(N__78358),
            .I(N__78355));
    LocalMux I__14095 (
            .O(N__78355),
            .I(shift_srl_188Z0Z_6));
    CascadeMux I__14094 (
            .O(N__78352),
            .I(N__78347));
    InMux I__14093 (
            .O(N__78351),
            .I(N__78344));
    InMux I__14092 (
            .O(N__78350),
            .I(N__78339));
    InMux I__14091 (
            .O(N__78347),
            .I(N__78339));
    LocalMux I__14090 (
            .O(N__78344),
            .I(N__78334));
    LocalMux I__14089 (
            .O(N__78339),
            .I(N__78334));
    Odrv4 I__14088 (
            .O(N__78334),
            .I(shift_srl_176Z0Z_15));
    InMux I__14087 (
            .O(N__78331),
            .I(N__78328));
    LocalMux I__14086 (
            .O(N__78328),
            .I(shift_srl_176Z0Z_0));
    InMux I__14085 (
            .O(N__78325),
            .I(N__78322));
    LocalMux I__14084 (
            .O(N__78322),
            .I(shift_srl_176Z0Z_1));
    InMux I__14083 (
            .O(N__78319),
            .I(N__78316));
    LocalMux I__14082 (
            .O(N__78316),
            .I(shift_srl_176Z0Z_2));
    InMux I__14081 (
            .O(N__78313),
            .I(N__78310));
    LocalMux I__14080 (
            .O(N__78310),
            .I(shift_srl_176Z0Z_3));
    InMux I__14079 (
            .O(N__78307),
            .I(N__78304));
    LocalMux I__14078 (
            .O(N__78304),
            .I(shift_srl_189Z0Z_12));
    InMux I__14077 (
            .O(N__78301),
            .I(N__78298));
    LocalMux I__14076 (
            .O(N__78298),
            .I(shift_srl_189Z0Z_13));
    InMux I__14075 (
            .O(N__78295),
            .I(N__78292));
    LocalMux I__14074 (
            .O(N__78292),
            .I(shift_srl_189Z0Z_14));
    InMux I__14073 (
            .O(N__78289),
            .I(N__78286));
    LocalMux I__14072 (
            .O(N__78286),
            .I(shift_srl_189Z0Z_9));
    InMux I__14071 (
            .O(N__78283),
            .I(N__78280));
    LocalMux I__14070 (
            .O(N__78280),
            .I(shift_srl_189Z0Z_8));
    InMux I__14069 (
            .O(N__78277),
            .I(N__78274));
    LocalMux I__14068 (
            .O(N__78274),
            .I(shift_srl_188Z0Z_0));
    InMux I__14067 (
            .O(N__78271),
            .I(N__78268));
    LocalMux I__14066 (
            .O(N__78268),
            .I(shift_srl_188Z0Z_1));
    InMux I__14065 (
            .O(N__78265),
            .I(N__78262));
    LocalMux I__14064 (
            .O(N__78262),
            .I(shift_srl_188Z0Z_2));
    InMux I__14063 (
            .O(N__78259),
            .I(N__78256));
    LocalMux I__14062 (
            .O(N__78256),
            .I(shift_srl_181Z0Z_11));
    InMux I__14061 (
            .O(N__78253),
            .I(N__78250));
    LocalMux I__14060 (
            .O(N__78250),
            .I(shift_srl_181Z0Z_12));
    InMux I__14059 (
            .O(N__78247),
            .I(N__78244));
    LocalMux I__14058 (
            .O(N__78244),
            .I(shift_srl_181Z0Z_6));
    InMux I__14057 (
            .O(N__78241),
            .I(N__78238));
    LocalMux I__14056 (
            .O(N__78238),
            .I(shift_srl_181Z0Z_13));
    InMux I__14055 (
            .O(N__78235),
            .I(N__78232));
    LocalMux I__14054 (
            .O(N__78232),
            .I(shift_srl_181Z0Z_14));
    InMux I__14053 (
            .O(N__78229),
            .I(N__78226));
    LocalMux I__14052 (
            .O(N__78226),
            .I(shift_srl_181Z0Z_9));
    InMux I__14051 (
            .O(N__78223),
            .I(N__78220));
    LocalMux I__14050 (
            .O(N__78220),
            .I(shift_srl_181Z0Z_7));
    InMux I__14049 (
            .O(N__78217),
            .I(N__78214));
    LocalMux I__14048 (
            .O(N__78214),
            .I(shift_srl_181Z0Z_8));
    CEMux I__14047 (
            .O(N__78211),
            .I(N__78207));
    CEMux I__14046 (
            .O(N__78210),
            .I(N__78204));
    LocalMux I__14045 (
            .O(N__78207),
            .I(clk_en_181));
    LocalMux I__14044 (
            .O(N__78204),
            .I(clk_en_181));
    InMux I__14043 (
            .O(N__78199),
            .I(N__78196));
    LocalMux I__14042 (
            .O(N__78196),
            .I(shift_srl_189Z0Z_10));
    InMux I__14041 (
            .O(N__78193),
            .I(N__78190));
    LocalMux I__14040 (
            .O(N__78190),
            .I(shift_srl_189Z0Z_11));
    CascadeMux I__14039 (
            .O(N__78187),
            .I(N__78184));
    InMux I__14038 (
            .O(N__78184),
            .I(N__78181));
    LocalMux I__14037 (
            .O(N__78181),
            .I(N__78178));
    Odrv4 I__14036 (
            .O(N__78178),
            .I(rco_int_0_a2_1_a2_0_sx_179));
    CascadeMux I__14035 (
            .O(N__78175),
            .I(shift_srl_179_RNIVNOT1Z0Z_15_cascade_));
    InMux I__14034 (
            .O(N__78172),
            .I(N__78169));
    LocalMux I__14033 (
            .O(N__78169),
            .I(N__78166));
    Sp12to4 I__14032 (
            .O(N__78166),
            .I(N__78163));
    Span12Mux_s10_v I__14031 (
            .O(N__78163),
            .I(N__78156));
    InMux I__14030 (
            .O(N__78162),
            .I(N__78153));
    InMux I__14029 (
            .O(N__78161),
            .I(N__78148));
    InMux I__14028 (
            .O(N__78160),
            .I(N__78148));
    InMux I__14027 (
            .O(N__78159),
            .I(N__78145));
    Span12Mux_v I__14026 (
            .O(N__78156),
            .I(N__78138));
    LocalMux I__14025 (
            .O(N__78153),
            .I(N__78138));
    LocalMux I__14024 (
            .O(N__78148),
            .I(N__78138));
    LocalMux I__14023 (
            .O(N__78145),
            .I(shift_srl_179_RNIVNOT1Z0Z_15));
    Odrv12 I__14022 (
            .O(N__78138),
            .I(shift_srl_179_RNIVNOT1Z0Z_15));
    InMux I__14021 (
            .O(N__78133),
            .I(N__78126));
    InMux I__14020 (
            .O(N__78132),
            .I(N__78126));
    InMux I__14019 (
            .O(N__78131),
            .I(N__78123));
    LocalMux I__14018 (
            .O(N__78126),
            .I(N__78120));
    LocalMux I__14017 (
            .O(N__78123),
            .I(shift_srl_179Z0Z_15));
    Odrv4 I__14016 (
            .O(N__78120),
            .I(shift_srl_179Z0Z_15));
    InMux I__14015 (
            .O(N__78115),
            .I(N__78112));
    LocalMux I__14014 (
            .O(N__78112),
            .I(N__78109));
    Odrv4 I__14013 (
            .O(N__78109),
            .I(rco_int_0_a2_1_a2_0_sx_182));
    CEMux I__14012 (
            .O(N__78106),
            .I(N__78103));
    LocalMux I__14011 (
            .O(N__78103),
            .I(N__78099));
    CEMux I__14010 (
            .O(N__78102),
            .I(N__78096));
    Span4Mux_h I__14009 (
            .O(N__78099),
            .I(N__78093));
    LocalMux I__14008 (
            .O(N__78096),
            .I(N__78090));
    Odrv4 I__14007 (
            .O(N__78093),
            .I(clk_en_178));
    Odrv12 I__14006 (
            .O(N__78090),
            .I(clk_en_178));
    InMux I__14005 (
            .O(N__78085),
            .I(N__78082));
    LocalMux I__14004 (
            .O(N__78082),
            .I(shift_srl_177Z0Z_14));
    InMux I__14003 (
            .O(N__78079),
            .I(N__78076));
    LocalMux I__14002 (
            .O(N__78076),
            .I(shift_srl_181Z0Z_10));
    InMux I__14001 (
            .O(N__78073),
            .I(N__78070));
    LocalMux I__14000 (
            .O(N__78070),
            .I(shift_srl_179Z0Z_7));
    InMux I__13999 (
            .O(N__78067),
            .I(N__78064));
    LocalMux I__13998 (
            .O(N__78064),
            .I(shift_srl_179Z0Z_8));
    CEMux I__13997 (
            .O(N__78061),
            .I(N__78057));
    CEMux I__13996 (
            .O(N__78060),
            .I(N__78054));
    LocalMux I__13995 (
            .O(N__78057),
            .I(N__78051));
    LocalMux I__13994 (
            .O(N__78054),
            .I(N__78048));
    Span4Mux_v I__13993 (
            .O(N__78051),
            .I(N__78045));
    Span4Mux_v I__13992 (
            .O(N__78048),
            .I(N__78042));
    Span4Mux_h I__13991 (
            .O(N__78045),
            .I(N__78039));
    Odrv4 I__13990 (
            .O(N__78042),
            .I(clk_en_179));
    Odrv4 I__13989 (
            .O(N__78039),
            .I(clk_en_179));
    InMux I__13988 (
            .O(N__78034),
            .I(N__78031));
    LocalMux I__13987 (
            .O(N__78031),
            .I(shift_srl_178Z0Z_5));
    InMux I__13986 (
            .O(N__78028),
            .I(N__78025));
    LocalMux I__13985 (
            .O(N__78025),
            .I(shift_srl_178Z0Z_10));
    InMux I__13984 (
            .O(N__78022),
            .I(N__78019));
    LocalMux I__13983 (
            .O(N__78019),
            .I(shift_srl_178Z0Z_11));
    InMux I__13982 (
            .O(N__78016),
            .I(N__78013));
    LocalMux I__13981 (
            .O(N__78013),
            .I(shift_srl_178Z0Z_12));
    InMux I__13980 (
            .O(N__78010),
            .I(N__78007));
    LocalMux I__13979 (
            .O(N__78007),
            .I(shift_srl_178Z0Z_6));
    InMux I__13978 (
            .O(N__78004),
            .I(N__78001));
    LocalMux I__13977 (
            .O(N__78001),
            .I(shift_srl_178Z0Z_13));
    InMux I__13976 (
            .O(N__77998),
            .I(N__77995));
    LocalMux I__13975 (
            .O(N__77995),
            .I(shift_srl_178Z0Z_14));
    InMux I__13974 (
            .O(N__77992),
            .I(N__77989));
    LocalMux I__13973 (
            .O(N__77989),
            .I(shift_srl_178Z0Z_7));
    InMux I__13972 (
            .O(N__77986),
            .I(N__77983));
    LocalMux I__13971 (
            .O(N__77983),
            .I(shift_srl_178Z0Z_8));
    InMux I__13970 (
            .O(N__77980),
            .I(N__77977));
    LocalMux I__13969 (
            .O(N__77977),
            .I(shift_srl_171Z0Z_8));
    InMux I__13968 (
            .O(N__77974),
            .I(N__77971));
    LocalMux I__13967 (
            .O(N__77971),
            .I(shift_srl_171Z0Z_9));
    InMux I__13966 (
            .O(N__77968),
            .I(N__77965));
    LocalMux I__13965 (
            .O(N__77965),
            .I(shift_srl_171Z0Z_0));
    InMux I__13964 (
            .O(N__77962),
            .I(N__77959));
    LocalMux I__13963 (
            .O(N__77959),
            .I(shift_srl_171Z0Z_1));
    CEMux I__13962 (
            .O(N__77956),
            .I(N__77952));
    CEMux I__13961 (
            .O(N__77955),
            .I(N__77949));
    LocalMux I__13960 (
            .O(N__77952),
            .I(clk_en_171));
    LocalMux I__13959 (
            .O(N__77949),
            .I(clk_en_171));
    InMux I__13958 (
            .O(N__77944),
            .I(N__77941));
    LocalMux I__13957 (
            .O(N__77941),
            .I(shift_srl_179Z0Z_10));
    InMux I__13956 (
            .O(N__77938),
            .I(N__77935));
    LocalMux I__13955 (
            .O(N__77935),
            .I(shift_srl_179Z0Z_11));
    InMux I__13954 (
            .O(N__77932),
            .I(N__77929));
    LocalMux I__13953 (
            .O(N__77929),
            .I(shift_srl_179Z0Z_12));
    InMux I__13952 (
            .O(N__77926),
            .I(N__77923));
    LocalMux I__13951 (
            .O(N__77923),
            .I(shift_srl_179Z0Z_13));
    InMux I__13950 (
            .O(N__77920),
            .I(N__77917));
    LocalMux I__13949 (
            .O(N__77917),
            .I(shift_srl_179Z0Z_14));
    InMux I__13948 (
            .O(N__77914),
            .I(N__77911));
    LocalMux I__13947 (
            .O(N__77911),
            .I(shift_srl_179Z0Z_9));
    CascadeMux I__13946 (
            .O(N__77908),
            .I(N__77904));
    CascadeMux I__13945 (
            .O(N__77907),
            .I(N__77899));
    InMux I__13944 (
            .O(N__77904),
            .I(N__77895));
    InMux I__13943 (
            .O(N__77903),
            .I(N__77892));
    InMux I__13942 (
            .O(N__77902),
            .I(N__77887));
    InMux I__13941 (
            .O(N__77899),
            .I(N__77887));
    InMux I__13940 (
            .O(N__77898),
            .I(N__77884));
    LocalMux I__13939 (
            .O(N__77895),
            .I(N__77881));
    LocalMux I__13938 (
            .O(N__77892),
            .I(N__77876));
    LocalMux I__13937 (
            .O(N__77887),
            .I(N__77876));
    LocalMux I__13936 (
            .O(N__77884),
            .I(N__77873));
    Span4Mux_v I__13935 (
            .O(N__77881),
            .I(N__77868));
    Span4Mux_v I__13934 (
            .O(N__77876),
            .I(N__77865));
    Span4Mux_v I__13933 (
            .O(N__77873),
            .I(N__77862));
    InMux I__13932 (
            .O(N__77872),
            .I(N__77859));
    InMux I__13931 (
            .O(N__77871),
            .I(N__77856));
    Span4Mux_v I__13930 (
            .O(N__77868),
            .I(N__77853));
    Span4Mux_v I__13929 (
            .O(N__77865),
            .I(N__77850));
    Span4Mux_v I__13928 (
            .O(N__77862),
            .I(N__77847));
    LocalMux I__13927 (
            .O(N__77859),
            .I(N__77844));
    LocalMux I__13926 (
            .O(N__77856),
            .I(N__77833));
    Sp12to4 I__13925 (
            .O(N__77853),
            .I(N__77833));
    Sp12to4 I__13924 (
            .O(N__77850),
            .I(N__77833));
    Sp12to4 I__13923 (
            .O(N__77847),
            .I(N__77833));
    Span12Mux_v I__13922 (
            .O(N__77844),
            .I(N__77833));
    Odrv12 I__13921 (
            .O(N__77833),
            .I(shift_srl_157Z0Z_15));
    InMux I__13920 (
            .O(N__77830),
            .I(N__77827));
    LocalMux I__13919 (
            .O(N__77827),
            .I(N__77817));
    InMux I__13918 (
            .O(N__77826),
            .I(N__77812));
    CascadeMux I__13917 (
            .O(N__77825),
            .I(N__77809));
    CascadeMux I__13916 (
            .O(N__77824),
            .I(N__77806));
    InMux I__13915 (
            .O(N__77823),
            .I(N__77801));
    InMux I__13914 (
            .O(N__77822),
            .I(N__77796));
    InMux I__13913 (
            .O(N__77821),
            .I(N__77796));
    InMux I__13912 (
            .O(N__77820),
            .I(N__77793));
    Span4Mux_h I__13911 (
            .O(N__77817),
            .I(N__77790));
    InMux I__13910 (
            .O(N__77816),
            .I(N__77785));
    InMux I__13909 (
            .O(N__77815),
            .I(N__77785));
    LocalMux I__13908 (
            .O(N__77812),
            .I(N__77782));
    InMux I__13907 (
            .O(N__77809),
            .I(N__77775));
    InMux I__13906 (
            .O(N__77806),
            .I(N__77775));
    InMux I__13905 (
            .O(N__77805),
            .I(N__77775));
    InMux I__13904 (
            .O(N__77804),
            .I(N__77771));
    LocalMux I__13903 (
            .O(N__77801),
            .I(N__77768));
    LocalMux I__13902 (
            .O(N__77796),
            .I(N__77765));
    LocalMux I__13901 (
            .O(N__77793),
            .I(N__77757));
    Span4Mux_h I__13900 (
            .O(N__77790),
            .I(N__77757));
    LocalMux I__13899 (
            .O(N__77785),
            .I(N__77757));
    Span4Mux_v I__13898 (
            .O(N__77782),
            .I(N__77752));
    LocalMux I__13897 (
            .O(N__77775),
            .I(N__77752));
    InMux I__13896 (
            .O(N__77774),
            .I(N__77749));
    LocalMux I__13895 (
            .O(N__77771),
            .I(N__77746));
    Span4Mux_v I__13894 (
            .O(N__77768),
            .I(N__77743));
    Span4Mux_v I__13893 (
            .O(N__77765),
            .I(N__77740));
    InMux I__13892 (
            .O(N__77764),
            .I(N__77737));
    Span4Mux_h I__13891 (
            .O(N__77757),
            .I(N__77734));
    Span4Mux_v I__13890 (
            .O(N__77752),
            .I(N__77729));
    LocalMux I__13889 (
            .O(N__77749),
            .I(N__77729));
    Span12Mux_h I__13888 (
            .O(N__77746),
            .I(N__77720));
    Sp12to4 I__13887 (
            .O(N__77743),
            .I(N__77720));
    Sp12to4 I__13886 (
            .O(N__77740),
            .I(N__77720));
    LocalMux I__13885 (
            .O(N__77737),
            .I(N__77720));
    Span4Mux_v I__13884 (
            .O(N__77734),
            .I(N__77717));
    Odrv4 I__13883 (
            .O(N__77729),
            .I(rco_int_0_a2_0_a2_1_145));
    Odrv12 I__13882 (
            .O(N__77720),
            .I(rco_int_0_a2_0_a2_1_145));
    Odrv4 I__13881 (
            .O(N__77717),
            .I(rco_int_0_a2_0_a2_1_145));
    CascadeMux I__13880 (
            .O(N__77710),
            .I(clk_en_0_a3_0_a2_sx_159_cascade_));
    CEMux I__13879 (
            .O(N__77707),
            .I(N__77703));
    CEMux I__13878 (
            .O(N__77706),
            .I(N__77699));
    LocalMux I__13877 (
            .O(N__77703),
            .I(N__77696));
    CEMux I__13876 (
            .O(N__77702),
            .I(N__77693));
    LocalMux I__13875 (
            .O(N__77699),
            .I(N__77690));
    Span4Mux_h I__13874 (
            .O(N__77696),
            .I(N__77687));
    LocalMux I__13873 (
            .O(N__77693),
            .I(N__77684));
    Span4Mux_v I__13872 (
            .O(N__77690),
            .I(N__77681));
    Odrv4 I__13871 (
            .O(N__77687),
            .I(clk_en_159));
    Odrv12 I__13870 (
            .O(N__77684),
            .I(clk_en_159));
    Odrv4 I__13869 (
            .O(N__77681),
            .I(clk_en_159));
    InMux I__13868 (
            .O(N__77674),
            .I(N__77671));
    LocalMux I__13867 (
            .O(N__77671),
            .I(N__77667));
    InMux I__13866 (
            .O(N__77670),
            .I(N__77664));
    Span4Mux_h I__13865 (
            .O(N__77667),
            .I(N__77661));
    LocalMux I__13864 (
            .O(N__77664),
            .I(shift_srl_156Z0Z_15));
    Odrv4 I__13863 (
            .O(N__77661),
            .I(shift_srl_156Z0Z_15));
    InMux I__13862 (
            .O(N__77656),
            .I(N__77653));
    LocalMux I__13861 (
            .O(N__77653),
            .I(N__77648));
    InMux I__13860 (
            .O(N__77652),
            .I(N__77645));
    InMux I__13859 (
            .O(N__77651),
            .I(N__77642));
    Span4Mux_v I__13858 (
            .O(N__77648),
            .I(N__77639));
    LocalMux I__13857 (
            .O(N__77645),
            .I(N__77636));
    LocalMux I__13856 (
            .O(N__77642),
            .I(N__77633));
    Span4Mux_h I__13855 (
            .O(N__77639),
            .I(N__77629));
    Span4Mux_v I__13854 (
            .O(N__77636),
            .I(N__77624));
    Span4Mux_v I__13853 (
            .O(N__77633),
            .I(N__77624));
    InMux I__13852 (
            .O(N__77632),
            .I(N__77621));
    Sp12to4 I__13851 (
            .O(N__77629),
            .I(N__77616));
    Sp12to4 I__13850 (
            .O(N__77624),
            .I(N__77616));
    LocalMux I__13849 (
            .O(N__77621),
            .I(shift_srl_155Z0Z_15));
    Odrv12 I__13848 (
            .O(N__77616),
            .I(shift_srl_155Z0Z_15));
    InMux I__13847 (
            .O(N__77611),
            .I(N__77608));
    LocalMux I__13846 (
            .O(N__77608),
            .I(N__77601));
    InMux I__13845 (
            .O(N__77607),
            .I(N__77598));
    InMux I__13844 (
            .O(N__77606),
            .I(N__77591));
    InMux I__13843 (
            .O(N__77605),
            .I(N__77591));
    InMux I__13842 (
            .O(N__77604),
            .I(N__77591));
    Span4Mux_v I__13841 (
            .O(N__77601),
            .I(N__77588));
    LocalMux I__13840 (
            .O(N__77598),
            .I(N__77585));
    LocalMux I__13839 (
            .O(N__77591),
            .I(N__77582));
    Span4Mux_v I__13838 (
            .O(N__77588),
            .I(N__77578));
    Sp12to4 I__13837 (
            .O(N__77585),
            .I(N__77575));
    Span4Mux_h I__13836 (
            .O(N__77582),
            .I(N__77572));
    InMux I__13835 (
            .O(N__77581),
            .I(N__77569));
    Sp12to4 I__13834 (
            .O(N__77578),
            .I(N__77564));
    Span12Mux_v I__13833 (
            .O(N__77575),
            .I(N__77564));
    Odrv4 I__13832 (
            .O(N__77572),
            .I(shift_srl_154Z0Z_15));
    LocalMux I__13831 (
            .O(N__77569),
            .I(shift_srl_154Z0Z_15));
    Odrv12 I__13830 (
            .O(N__77564),
            .I(shift_srl_154Z0Z_15));
    InMux I__13829 (
            .O(N__77557),
            .I(N__77553));
    CascadeMux I__13828 (
            .O(N__77556),
            .I(N__77548));
    LocalMux I__13827 (
            .O(N__77553),
            .I(N__77544));
    InMux I__13826 (
            .O(N__77552),
            .I(N__77541));
    InMux I__13825 (
            .O(N__77551),
            .I(N__77534));
    InMux I__13824 (
            .O(N__77548),
            .I(N__77534));
    InMux I__13823 (
            .O(N__77547),
            .I(N__77534));
    Span12Mux_v I__13822 (
            .O(N__77544),
            .I(N__77530));
    LocalMux I__13821 (
            .O(N__77541),
            .I(N__77526));
    LocalMux I__13820 (
            .O(N__77534),
            .I(N__77523));
    InMux I__13819 (
            .O(N__77533),
            .I(N__77520));
    Span12Mux_h I__13818 (
            .O(N__77530),
            .I(N__77516));
    InMux I__13817 (
            .O(N__77529),
            .I(N__77513));
    Span12Mux_v I__13816 (
            .O(N__77526),
            .I(N__77510));
    Span4Mux_v I__13815 (
            .O(N__77523),
            .I(N__77505));
    LocalMux I__13814 (
            .O(N__77520),
            .I(N__77505));
    InMux I__13813 (
            .O(N__77519),
            .I(N__77502));
    Odrv12 I__13812 (
            .O(N__77516),
            .I(shift_srl_156_RNII4IKZ0Z_15));
    LocalMux I__13811 (
            .O(N__77513),
            .I(shift_srl_156_RNII4IKZ0Z_15));
    Odrv12 I__13810 (
            .O(N__77510),
            .I(shift_srl_156_RNII4IKZ0Z_15));
    Odrv4 I__13809 (
            .O(N__77505),
            .I(shift_srl_156_RNII4IKZ0Z_15));
    LocalMux I__13808 (
            .O(N__77502),
            .I(shift_srl_156_RNII4IKZ0Z_15));
    InMux I__13807 (
            .O(N__77491),
            .I(N__77488));
    LocalMux I__13806 (
            .O(N__77488),
            .I(shift_srl_171Z0Z_10));
    InMux I__13805 (
            .O(N__77485),
            .I(N__77482));
    LocalMux I__13804 (
            .O(N__77482),
            .I(shift_srl_171Z0Z_11));
    InMux I__13803 (
            .O(N__77479),
            .I(N__77476));
    LocalMux I__13802 (
            .O(N__77476),
            .I(shift_srl_171Z0Z_12));
    InMux I__13801 (
            .O(N__77473),
            .I(N__77470));
    LocalMux I__13800 (
            .O(N__77470),
            .I(shift_srl_171Z0Z_13));
    InMux I__13799 (
            .O(N__77467),
            .I(N__77464));
    LocalMux I__13798 (
            .O(N__77464),
            .I(shift_srl_171Z0Z_14));
    InMux I__13797 (
            .O(N__77461),
            .I(N__77458));
    LocalMux I__13796 (
            .O(N__77458),
            .I(shift_srl_31Z0Z_14));
    InMux I__13795 (
            .O(N__77455),
            .I(N__77452));
    LocalMux I__13794 (
            .O(N__77452),
            .I(shift_srl_31Z0Z_9));
    InMux I__13793 (
            .O(N__77449),
            .I(N__77446));
    LocalMux I__13792 (
            .O(N__77446),
            .I(shift_srl_31Z0Z_7));
    InMux I__13791 (
            .O(N__77443),
            .I(N__77440));
    LocalMux I__13790 (
            .O(N__77440),
            .I(shift_srl_31Z0Z_8));
    CascadeMux I__13789 (
            .O(N__77437),
            .I(N__77434));
    InMux I__13788 (
            .O(N__77434),
            .I(N__77431));
    LocalMux I__13787 (
            .O(N__77431),
            .I(N__77427));
    InMux I__13786 (
            .O(N__77430),
            .I(N__77424));
    Span4Mux_v I__13785 (
            .O(N__77427),
            .I(N__77421));
    LocalMux I__13784 (
            .O(N__77424),
            .I(N__77417));
    Span4Mux_h I__13783 (
            .O(N__77421),
            .I(N__77414));
    InMux I__13782 (
            .O(N__77420),
            .I(N__77411));
    Span12Mux_v I__13781 (
            .O(N__77417),
            .I(N__77408));
    Span4Mux_h I__13780 (
            .O(N__77414),
            .I(N__77405));
    LocalMux I__13779 (
            .O(N__77411),
            .I(shift_srl_160Z0Z_15));
    Odrv12 I__13778 (
            .O(N__77408),
            .I(shift_srl_160Z0Z_15));
    Odrv4 I__13777 (
            .O(N__77405),
            .I(shift_srl_160Z0Z_15));
    InMux I__13776 (
            .O(N__77398),
            .I(N__77395));
    LocalMux I__13775 (
            .O(N__77395),
            .I(N__77392));
    Span4Mux_h I__13774 (
            .O(N__77392),
            .I(N__77388));
    InMux I__13773 (
            .O(N__77391),
            .I(N__77385));
    Span4Mux_h I__13772 (
            .O(N__77388),
            .I(N__77382));
    LocalMux I__13771 (
            .O(N__77385),
            .I(shift_srl_162Z0Z_15));
    Odrv4 I__13770 (
            .O(N__77382),
            .I(shift_srl_162Z0Z_15));
    InMux I__13769 (
            .O(N__77377),
            .I(N__77373));
    InMux I__13768 (
            .O(N__77376),
            .I(N__77370));
    LocalMux I__13767 (
            .O(N__77373),
            .I(N__77366));
    LocalMux I__13766 (
            .O(N__77370),
            .I(N__77363));
    InMux I__13765 (
            .O(N__77369),
            .I(N__77360));
    Span4Mux_h I__13764 (
            .O(N__77366),
            .I(N__77357));
    Span4Mux_h I__13763 (
            .O(N__77363),
            .I(N__77354));
    LocalMux I__13762 (
            .O(N__77360),
            .I(N__77351));
    Span4Mux_h I__13761 (
            .O(N__77357),
            .I(N__77347));
    Span4Mux_h I__13760 (
            .O(N__77354),
            .I(N__77344));
    Span4Mux_v I__13759 (
            .O(N__77351),
            .I(N__77341));
    InMux I__13758 (
            .O(N__77350),
            .I(N__77338));
    Span4Mux_v I__13757 (
            .O(N__77347),
            .I(N__77335));
    Span4Mux_h I__13756 (
            .O(N__77344),
            .I(N__77332));
    Odrv4 I__13755 (
            .O(N__77341),
            .I(shift_srl_161Z0Z_15));
    LocalMux I__13754 (
            .O(N__77338),
            .I(shift_srl_161Z0Z_15));
    Odrv4 I__13753 (
            .O(N__77335),
            .I(shift_srl_161Z0Z_15));
    Odrv4 I__13752 (
            .O(N__77332),
            .I(shift_srl_161Z0Z_15));
    CascadeMux I__13751 (
            .O(N__77323),
            .I(rco_int_0_a3_0_a2_0_sx_162_cascade_));
    CascadeMux I__13750 (
            .O(N__77320),
            .I(rco_int_0_a3_0_a2_0_162_cascade_));
    InMux I__13749 (
            .O(N__77317),
            .I(N__77314));
    LocalMux I__13748 (
            .O(N__77314),
            .I(N__77311));
    Odrv4 I__13747 (
            .O(N__77311),
            .I(shift_srl_159Z0Z_14));
    CascadeMux I__13746 (
            .O(N__77308),
            .I(N__77305));
    InMux I__13745 (
            .O(N__77305),
            .I(N__77301));
    InMux I__13744 (
            .O(N__77304),
            .I(N__77297));
    LocalMux I__13743 (
            .O(N__77301),
            .I(N__77294));
    InMux I__13742 (
            .O(N__77300),
            .I(N__77291));
    LocalMux I__13741 (
            .O(N__77297),
            .I(shift_srl_159Z0Z_15));
    Odrv4 I__13740 (
            .O(N__77294),
            .I(shift_srl_159Z0Z_15));
    LocalMux I__13739 (
            .O(N__77291),
            .I(shift_srl_159Z0Z_15));
    InMux I__13738 (
            .O(N__77284),
            .I(N__77281));
    LocalMux I__13737 (
            .O(N__77281),
            .I(N__77274));
    InMux I__13736 (
            .O(N__77280),
            .I(N__77271));
    InMux I__13735 (
            .O(N__77279),
            .I(N__77268));
    InMux I__13734 (
            .O(N__77278),
            .I(N__77265));
    InMux I__13733 (
            .O(N__77277),
            .I(N__77262));
    Sp12to4 I__13732 (
            .O(N__77274),
            .I(N__77255));
    LocalMux I__13731 (
            .O(N__77271),
            .I(N__77255));
    LocalMux I__13730 (
            .O(N__77268),
            .I(N__77255));
    LocalMux I__13729 (
            .O(N__77265),
            .I(shift_srl_158Z0Z_15));
    LocalMux I__13728 (
            .O(N__77262),
            .I(shift_srl_158Z0Z_15));
    Odrv12 I__13727 (
            .O(N__77255),
            .I(shift_srl_158Z0Z_15));
    InMux I__13726 (
            .O(N__77248),
            .I(N__77245));
    LocalMux I__13725 (
            .O(N__77245),
            .I(shift_srl_31Z0Z_2));
    InMux I__13724 (
            .O(N__77242),
            .I(N__77239));
    LocalMux I__13723 (
            .O(N__77239),
            .I(shift_srl_31Z0Z_3));
    InMux I__13722 (
            .O(N__77236),
            .I(N__77233));
    LocalMux I__13721 (
            .O(N__77233),
            .I(shift_srl_31Z0Z_4));
    InMux I__13720 (
            .O(N__77230),
            .I(N__77227));
    LocalMux I__13719 (
            .O(N__77227),
            .I(shift_srl_31Z0Z_5));
    InMux I__13718 (
            .O(N__77224),
            .I(N__77221));
    LocalMux I__13717 (
            .O(N__77221),
            .I(shift_srl_31Z0Z_6));
    InMux I__13716 (
            .O(N__77218),
            .I(N__77215));
    LocalMux I__13715 (
            .O(N__77215),
            .I(shift_srl_31Z0Z_10));
    InMux I__13714 (
            .O(N__77212),
            .I(N__77209));
    LocalMux I__13713 (
            .O(N__77209),
            .I(shift_srl_31Z0Z_11));
    InMux I__13712 (
            .O(N__77206),
            .I(N__77203));
    LocalMux I__13711 (
            .O(N__77203),
            .I(shift_srl_31Z0Z_12));
    InMux I__13710 (
            .O(N__77200),
            .I(N__77197));
    LocalMux I__13709 (
            .O(N__77197),
            .I(shift_srl_31Z0Z_13));
    InMux I__13708 (
            .O(N__77194),
            .I(N__77191));
    LocalMux I__13707 (
            .O(N__77191),
            .I(shift_srl_65Z0Z_13));
    InMux I__13706 (
            .O(N__77188),
            .I(N__77185));
    LocalMux I__13705 (
            .O(N__77185),
            .I(shift_srl_65Z0Z_14));
    InMux I__13704 (
            .O(N__77182),
            .I(N__77179));
    LocalMux I__13703 (
            .O(N__77179),
            .I(shift_srl_65Z0Z_9));
    InMux I__13702 (
            .O(N__77176),
            .I(N__77173));
    LocalMux I__13701 (
            .O(N__77173),
            .I(shift_srl_65Z0Z_8));
    InMux I__13700 (
            .O(N__77170),
            .I(N__77167));
    LocalMux I__13699 (
            .O(N__77167),
            .I(shift_srl_63Z0Z_7));
    InMux I__13698 (
            .O(N__77164),
            .I(N__77161));
    LocalMux I__13697 (
            .O(N__77161),
            .I(shift_srl_63Z0Z_8));
    InMux I__13696 (
            .O(N__77158),
            .I(N__77155));
    LocalMux I__13695 (
            .O(N__77155),
            .I(shift_srl_31Z0Z_0));
    InMux I__13694 (
            .O(N__77152),
            .I(N__77149));
    LocalMux I__13693 (
            .O(N__77149),
            .I(shift_srl_31Z0Z_1));
    InMux I__13692 (
            .O(N__77146),
            .I(N__77143));
    LocalMux I__13691 (
            .O(N__77143),
            .I(shift_srl_64Z0Z_12));
    InMux I__13690 (
            .O(N__77140),
            .I(N__77137));
    LocalMux I__13689 (
            .O(N__77137),
            .I(shift_srl_64Z0Z_13));
    InMux I__13688 (
            .O(N__77134),
            .I(N__77131));
    LocalMux I__13687 (
            .O(N__77131),
            .I(shift_srl_64Z0Z_14));
    InMux I__13686 (
            .O(N__77128),
            .I(N__77125));
    LocalMux I__13685 (
            .O(N__77125),
            .I(shift_srl_64Z0Z_9));
    InMux I__13684 (
            .O(N__77122),
            .I(N__77119));
    LocalMux I__13683 (
            .O(N__77119),
            .I(shift_srl_64Z0Z_8));
    InMux I__13682 (
            .O(N__77116),
            .I(N__77113));
    LocalMux I__13681 (
            .O(N__77113),
            .I(shift_srl_65Z0Z_10));
    InMux I__13680 (
            .O(N__77110),
            .I(N__77107));
    LocalMux I__13679 (
            .O(N__77107),
            .I(shift_srl_65Z0Z_11));
    InMux I__13678 (
            .O(N__77104),
            .I(N__77101));
    LocalMux I__13677 (
            .O(N__77101),
            .I(shift_srl_65Z0Z_12));
    InMux I__13676 (
            .O(N__77098),
            .I(N__77095));
    LocalMux I__13675 (
            .O(N__77095),
            .I(N__77092));
    Odrv4 I__13674 (
            .O(N__77092),
            .I(rco_int_0_a2_1_a2_sx_53));
    IoInMux I__13673 (
            .O(N__77089),
            .I(N__77086));
    LocalMux I__13672 (
            .O(N__77086),
            .I(N__77083));
    IoSpan4Mux I__13671 (
            .O(N__77083),
            .I(N__77079));
    InMux I__13670 (
            .O(N__77082),
            .I(N__77076));
    IoSpan4Mux I__13669 (
            .O(N__77079),
            .I(N__77073));
    LocalMux I__13668 (
            .O(N__77076),
            .I(N__77070));
    Span4Mux_s3_v I__13667 (
            .O(N__77073),
            .I(N__77064));
    Span4Mux_s3_v I__13666 (
            .O(N__77070),
            .I(N__77064));
    InMux I__13665 (
            .O(N__77069),
            .I(N__77061));
    Span4Mux_v I__13664 (
            .O(N__77064),
            .I(N__77058));
    LocalMux I__13663 (
            .O(N__77061),
            .I(N__77055));
    Sp12to4 I__13662 (
            .O(N__77058),
            .I(N__77052));
    Span4Mux_v I__13661 (
            .O(N__77055),
            .I(N__77049));
    Span12Mux_h I__13660 (
            .O(N__77052),
            .I(N__77041));
    Sp12to4 I__13659 (
            .O(N__77049),
            .I(N__77041));
    InMux I__13658 (
            .O(N__77048),
            .I(N__77034));
    InMux I__13657 (
            .O(N__77047),
            .I(N__77034));
    InMux I__13656 (
            .O(N__77046),
            .I(N__77034));
    Span12Mux_v I__13655 (
            .O(N__77041),
            .I(N__77031));
    LocalMux I__13654 (
            .O(N__77034),
            .I(N__77028));
    Odrv12 I__13653 (
            .O(N__77031),
            .I(rco_c_53));
    Odrv4 I__13652 (
            .O(N__77028),
            .I(rco_c_53));
    InMux I__13651 (
            .O(N__77023),
            .I(N__77020));
    LocalMux I__13650 (
            .O(N__77020),
            .I(N__77017));
    Span4Mux_h I__13649 (
            .O(N__77017),
            .I(N__77014));
    Sp12to4 I__13648 (
            .O(N__77014),
            .I(N__77010));
    InMux I__13647 (
            .O(N__77013),
            .I(N__77007));
    Span12Mux_v I__13646 (
            .O(N__77010),
            .I(N__77001));
    LocalMux I__13645 (
            .O(N__77007),
            .I(N__76998));
    InMux I__13644 (
            .O(N__77006),
            .I(N__76993));
    InMux I__13643 (
            .O(N__77005),
            .I(N__76993));
    InMux I__13642 (
            .O(N__77004),
            .I(N__76990));
    Odrv12 I__13641 (
            .O(N__77001),
            .I(shift_srl_54Z0Z_15));
    Odrv4 I__13640 (
            .O(N__76998),
            .I(shift_srl_54Z0Z_15));
    LocalMux I__13639 (
            .O(N__76993),
            .I(shift_srl_54Z0Z_15));
    LocalMux I__13638 (
            .O(N__76990),
            .I(shift_srl_54Z0Z_15));
    InMux I__13637 (
            .O(N__76981),
            .I(N__76978));
    LocalMux I__13636 (
            .O(N__76978),
            .I(shift_srl_54Z0Z_0));
    InMux I__13635 (
            .O(N__76975),
            .I(N__76972));
    LocalMux I__13634 (
            .O(N__76972),
            .I(shift_srl_54Z0Z_1));
    InMux I__13633 (
            .O(N__76969),
            .I(N__76966));
    LocalMux I__13632 (
            .O(N__76966),
            .I(shift_srl_54Z0Z_2));
    InMux I__13631 (
            .O(N__76963),
            .I(N__76960));
    LocalMux I__13630 (
            .O(N__76960),
            .I(shift_srl_54Z0Z_3));
    InMux I__13629 (
            .O(N__76957),
            .I(N__76954));
    LocalMux I__13628 (
            .O(N__76954),
            .I(shift_srl_64Z0Z_10));
    InMux I__13627 (
            .O(N__76951),
            .I(N__76948));
    LocalMux I__13626 (
            .O(N__76948),
            .I(shift_srl_64Z0Z_11));
    CascadeMux I__13625 (
            .O(N__76945),
            .I(N__76942));
    InMux I__13624 (
            .O(N__76942),
            .I(N__76930));
    InMux I__13623 (
            .O(N__76941),
            .I(N__76930));
    InMux I__13622 (
            .O(N__76940),
            .I(N__76930));
    InMux I__13621 (
            .O(N__76939),
            .I(N__76930));
    LocalMux I__13620 (
            .O(N__76930),
            .I(N__76925));
    InMux I__13619 (
            .O(N__76929),
            .I(N__76922));
    InMux I__13618 (
            .O(N__76928),
            .I(N__76919));
    Odrv4 I__13617 (
            .O(N__76925),
            .I(shift_srl_55_RNI9BJMZ0Z_15));
    LocalMux I__13616 (
            .O(N__76922),
            .I(shift_srl_55_RNI9BJMZ0Z_15));
    LocalMux I__13615 (
            .O(N__76919),
            .I(shift_srl_55_RNI9BJMZ0Z_15));
    IoInMux I__13614 (
            .O(N__76912),
            .I(N__76908));
    InMux I__13613 (
            .O(N__76911),
            .I(N__76903));
    LocalMux I__13612 (
            .O(N__76908),
            .I(N__76900));
    InMux I__13611 (
            .O(N__76907),
            .I(N__76897));
    InMux I__13610 (
            .O(N__76906),
            .I(N__76894));
    LocalMux I__13609 (
            .O(N__76903),
            .I(N__76890));
    Span12Mux_s11_h I__13608 (
            .O(N__76900),
            .I(N__76887));
    LocalMux I__13607 (
            .O(N__76897),
            .I(N__76884));
    LocalMux I__13606 (
            .O(N__76894),
            .I(N__76881));
    InMux I__13605 (
            .O(N__76893),
            .I(N__76878));
    Span4Mux_v I__13604 (
            .O(N__76890),
            .I(N__76875));
    Odrv12 I__13603 (
            .O(N__76887),
            .I(rco_c_44));
    Odrv4 I__13602 (
            .O(N__76884),
            .I(rco_c_44));
    Odrv4 I__13601 (
            .O(N__76881),
            .I(rco_c_44));
    LocalMux I__13600 (
            .O(N__76878),
            .I(rco_c_44));
    Odrv4 I__13599 (
            .O(N__76875),
            .I(rco_c_44));
    CascadeMux I__13598 (
            .O(N__76864),
            .I(clk_en_0_a3_0_a2_sx_57_cascade_));
    InMux I__13597 (
            .O(N__76861),
            .I(N__76858));
    LocalMux I__13596 (
            .O(N__76858),
            .I(N__76851));
    InMux I__13595 (
            .O(N__76857),
            .I(N__76848));
    InMux I__13594 (
            .O(N__76856),
            .I(N__76843));
    InMux I__13593 (
            .O(N__76855),
            .I(N__76843));
    InMux I__13592 (
            .O(N__76854),
            .I(N__76838));
    Span4Mux_h I__13591 (
            .O(N__76851),
            .I(N__76833));
    LocalMux I__13590 (
            .O(N__76848),
            .I(N__76833));
    LocalMux I__13589 (
            .O(N__76843),
            .I(N__76829));
    InMux I__13588 (
            .O(N__76842),
            .I(N__76824));
    InMux I__13587 (
            .O(N__76841),
            .I(N__76824));
    LocalMux I__13586 (
            .O(N__76838),
            .I(N__76821));
    Span4Mux_v I__13585 (
            .O(N__76833),
            .I(N__76818));
    InMux I__13584 (
            .O(N__76832),
            .I(N__76815));
    Span4Mux_v I__13583 (
            .O(N__76829),
            .I(N__76810));
    LocalMux I__13582 (
            .O(N__76824),
            .I(N__76810));
    Span12Mux_v I__13581 (
            .O(N__76821),
            .I(N__76807));
    Odrv4 I__13580 (
            .O(N__76818),
            .I(shift_srl_47_RNIV3QLZ0Z_15));
    LocalMux I__13579 (
            .O(N__76815),
            .I(shift_srl_47_RNIV3QLZ0Z_15));
    Odrv4 I__13578 (
            .O(N__76810),
            .I(shift_srl_47_RNIV3QLZ0Z_15));
    Odrv12 I__13577 (
            .O(N__76807),
            .I(shift_srl_47_RNIV3QLZ0Z_15));
    InMux I__13576 (
            .O(N__76798),
            .I(N__76792));
    InMux I__13575 (
            .O(N__76797),
            .I(N__76789));
    InMux I__13574 (
            .O(N__76796),
            .I(N__76784));
    InMux I__13573 (
            .O(N__76795),
            .I(N__76784));
    LocalMux I__13572 (
            .O(N__76792),
            .I(N__76781));
    LocalMux I__13571 (
            .O(N__76789),
            .I(shift_srl_57Z0Z_15));
    LocalMux I__13570 (
            .O(N__76784),
            .I(shift_srl_57Z0Z_15));
    Odrv4 I__13569 (
            .O(N__76781),
            .I(shift_srl_57Z0Z_15));
    InMux I__13568 (
            .O(N__76774),
            .I(N__76771));
    LocalMux I__13567 (
            .O(N__76771),
            .I(shift_srl_57Z0Z_0));
    InMux I__13566 (
            .O(N__76768),
            .I(N__76765));
    LocalMux I__13565 (
            .O(N__76765),
            .I(shift_srl_57Z0Z_1));
    InMux I__13564 (
            .O(N__76762),
            .I(N__76759));
    LocalMux I__13563 (
            .O(N__76759),
            .I(shift_srl_57Z0Z_2));
    InMux I__13562 (
            .O(N__76756),
            .I(N__76753));
    LocalMux I__13561 (
            .O(N__76753),
            .I(shift_srl_57Z0Z_3));
    InMux I__13560 (
            .O(N__76750),
            .I(N__76747));
    LocalMux I__13559 (
            .O(N__76747),
            .I(shift_srl_57Z0Z_4));
    InMux I__13558 (
            .O(N__76744),
            .I(N__76741));
    LocalMux I__13557 (
            .O(N__76741),
            .I(shift_srl_57Z0Z_5));
    InMux I__13556 (
            .O(N__76738),
            .I(N__76735));
    LocalMux I__13555 (
            .O(N__76735),
            .I(shift_srl_57Z0Z_6));
    InMux I__13554 (
            .O(N__76732),
            .I(N__76729));
    LocalMux I__13553 (
            .O(N__76729),
            .I(shift_srl_57Z0Z_7));
    CEMux I__13552 (
            .O(N__76726),
            .I(N__76722));
    CEMux I__13551 (
            .O(N__76725),
            .I(N__76719));
    LocalMux I__13550 (
            .O(N__76722),
            .I(N__76716));
    LocalMux I__13549 (
            .O(N__76719),
            .I(N__76713));
    Odrv4 I__13548 (
            .O(N__76716),
            .I(clk_en_57));
    Odrv4 I__13547 (
            .O(N__76713),
            .I(clk_en_57));
    InMux I__13546 (
            .O(N__76708),
            .I(N__76705));
    LocalMux I__13545 (
            .O(N__76705),
            .I(shift_srl_52Z0Z_5));
    InMux I__13544 (
            .O(N__76702),
            .I(N__76699));
    LocalMux I__13543 (
            .O(N__76699),
            .I(shift_srl_52Z0Z_6));
    InMux I__13542 (
            .O(N__76696),
            .I(N__76693));
    LocalMux I__13541 (
            .O(N__76693),
            .I(shift_srl_52Z0Z_7));
    CEMux I__13540 (
            .O(N__76690),
            .I(N__76686));
    CEMux I__13539 (
            .O(N__76689),
            .I(N__76683));
    LocalMux I__13538 (
            .O(N__76686),
            .I(clk_en_52));
    LocalMux I__13537 (
            .O(N__76683),
            .I(clk_en_52));
    IoInMux I__13536 (
            .O(N__76678),
            .I(N__76675));
    LocalMux I__13535 (
            .O(N__76675),
            .I(N__76672));
    Span4Mux_s2_h I__13534 (
            .O(N__76672),
            .I(N__76669));
    Sp12to4 I__13533 (
            .O(N__76669),
            .I(N__76666));
    Span12Mux_s10_v I__13532 (
            .O(N__76666),
            .I(N__76663));
    Odrv12 I__13531 (
            .O(N__76663),
            .I(rco_c_57));
    IoInMux I__13530 (
            .O(N__76660),
            .I(N__76657));
    LocalMux I__13529 (
            .O(N__76657),
            .I(N__76654));
    Span4Mux_s3_h I__13528 (
            .O(N__76654),
            .I(N__76651));
    Sp12to4 I__13527 (
            .O(N__76651),
            .I(N__76648));
    Span12Mux_s10_v I__13526 (
            .O(N__76648),
            .I(N__76645));
    Odrv12 I__13525 (
            .O(N__76645),
            .I(rco_c_56));
    CascadeMux I__13524 (
            .O(N__76642),
            .I(clk_en_54_cascade_));
    IoInMux I__13523 (
            .O(N__76639),
            .I(N__76636));
    LocalMux I__13522 (
            .O(N__76636),
            .I(N__76633));
    IoSpan4Mux I__13521 (
            .O(N__76633),
            .I(N__76630));
    Span4Mux_s2_v I__13520 (
            .O(N__76630),
            .I(N__76627));
    Sp12to4 I__13519 (
            .O(N__76627),
            .I(N__76624));
    Span12Mux_s10_h I__13518 (
            .O(N__76624),
            .I(N__76621));
    Odrv12 I__13517 (
            .O(N__76621),
            .I(rco_c_55));
    InMux I__13516 (
            .O(N__76618),
            .I(N__76614));
    InMux I__13515 (
            .O(N__76617),
            .I(N__76609));
    LocalMux I__13514 (
            .O(N__76614),
            .I(N__76605));
    InMux I__13513 (
            .O(N__76613),
            .I(N__76602));
    InMux I__13512 (
            .O(N__76612),
            .I(N__76598));
    LocalMux I__13511 (
            .O(N__76609),
            .I(N__76595));
    InMux I__13510 (
            .O(N__76608),
            .I(N__76589));
    Span4Mux_v I__13509 (
            .O(N__76605),
            .I(N__76584));
    LocalMux I__13508 (
            .O(N__76602),
            .I(N__76584));
    InMux I__13507 (
            .O(N__76601),
            .I(N__76581));
    LocalMux I__13506 (
            .O(N__76598),
            .I(N__76578));
    Span4Mux_h I__13505 (
            .O(N__76595),
            .I(N__76575));
    InMux I__13504 (
            .O(N__76594),
            .I(N__76568));
    InMux I__13503 (
            .O(N__76593),
            .I(N__76568));
    InMux I__13502 (
            .O(N__76592),
            .I(N__76568));
    LocalMux I__13501 (
            .O(N__76589),
            .I(N__76565));
    Span4Mux_v I__13500 (
            .O(N__76584),
            .I(N__76560));
    LocalMux I__13499 (
            .O(N__76581),
            .I(N__76560));
    Odrv4 I__13498 (
            .O(N__76578),
            .I(shift_srl_48Z0Z_15));
    Odrv4 I__13497 (
            .O(N__76575),
            .I(shift_srl_48Z0Z_15));
    LocalMux I__13496 (
            .O(N__76568),
            .I(shift_srl_48Z0Z_15));
    Odrv12 I__13495 (
            .O(N__76565),
            .I(shift_srl_48Z0Z_15));
    Odrv4 I__13494 (
            .O(N__76560),
            .I(shift_srl_48Z0Z_15));
    CascadeMux I__13493 (
            .O(N__76549),
            .I(N__76543));
    InMux I__13492 (
            .O(N__76548),
            .I(N__76538));
    InMux I__13491 (
            .O(N__76547),
            .I(N__76538));
    InMux I__13490 (
            .O(N__76546),
            .I(N__76533));
    InMux I__13489 (
            .O(N__76543),
            .I(N__76533));
    LocalMux I__13488 (
            .O(N__76538),
            .I(N__76527));
    LocalMux I__13487 (
            .O(N__76533),
            .I(N__76527));
    InMux I__13486 (
            .O(N__76532),
            .I(N__76523));
    Span4Mux_v I__13485 (
            .O(N__76527),
            .I(N__76520));
    InMux I__13484 (
            .O(N__76526),
            .I(N__76517));
    LocalMux I__13483 (
            .O(N__76523),
            .I(shift_srl_56Z0Z_15));
    Odrv4 I__13482 (
            .O(N__76520),
            .I(shift_srl_56Z0Z_15));
    LocalMux I__13481 (
            .O(N__76517),
            .I(shift_srl_56Z0Z_15));
    InMux I__13480 (
            .O(N__76510),
            .I(N__76507));
    LocalMux I__13479 (
            .O(N__76507),
            .I(shift_srl_50Z0Z_1));
    InMux I__13478 (
            .O(N__76504),
            .I(N__76501));
    LocalMux I__13477 (
            .O(N__76501),
            .I(shift_srl_50Z0Z_2));
    InMux I__13476 (
            .O(N__76498),
            .I(N__76495));
    LocalMux I__13475 (
            .O(N__76495),
            .I(shift_srl_50Z0Z_3));
    InMux I__13474 (
            .O(N__76492),
            .I(N__76489));
    LocalMux I__13473 (
            .O(N__76489),
            .I(shift_srl_50Z0Z_4));
    CEMux I__13472 (
            .O(N__76486),
            .I(N__76483));
    LocalMux I__13471 (
            .O(N__76483),
            .I(N__76479));
    CEMux I__13470 (
            .O(N__76482),
            .I(N__76476));
    Span4Mux_v I__13469 (
            .O(N__76479),
            .I(N__76469));
    LocalMux I__13468 (
            .O(N__76476),
            .I(N__76469));
    CEMux I__13467 (
            .O(N__76475),
            .I(N__76466));
    CEMux I__13466 (
            .O(N__76474),
            .I(N__76463));
    Sp12to4 I__13465 (
            .O(N__76469),
            .I(N__76458));
    LocalMux I__13464 (
            .O(N__76466),
            .I(N__76458));
    LocalMux I__13463 (
            .O(N__76463),
            .I(N__76455));
    Odrv12 I__13462 (
            .O(N__76458),
            .I(clk_en_50));
    Odrv4 I__13461 (
            .O(N__76455),
            .I(clk_en_50));
    CascadeMux I__13460 (
            .O(N__76450),
            .I(N__76446));
    InMux I__13459 (
            .O(N__76449),
            .I(N__76443));
    InMux I__13458 (
            .O(N__76446),
            .I(N__76438));
    LocalMux I__13457 (
            .O(N__76443),
            .I(N__76435));
    InMux I__13456 (
            .O(N__76442),
            .I(N__76432));
    InMux I__13455 (
            .O(N__76441),
            .I(N__76429));
    LocalMux I__13454 (
            .O(N__76438),
            .I(N__76426));
    Odrv4 I__13453 (
            .O(N__76435),
            .I(shift_srl_52Z0Z_15));
    LocalMux I__13452 (
            .O(N__76432),
            .I(shift_srl_52Z0Z_15));
    LocalMux I__13451 (
            .O(N__76429),
            .I(shift_srl_52Z0Z_15));
    Odrv4 I__13450 (
            .O(N__76426),
            .I(shift_srl_52Z0Z_15));
    InMux I__13449 (
            .O(N__76417),
            .I(N__76414));
    LocalMux I__13448 (
            .O(N__76414),
            .I(shift_srl_52Z0Z_0));
    InMux I__13447 (
            .O(N__76411),
            .I(N__76408));
    LocalMux I__13446 (
            .O(N__76408),
            .I(shift_srl_52Z0Z_1));
    InMux I__13445 (
            .O(N__76405),
            .I(N__76402));
    LocalMux I__13444 (
            .O(N__76402),
            .I(shift_srl_52Z0Z_2));
    InMux I__13443 (
            .O(N__76399),
            .I(N__76396));
    LocalMux I__13442 (
            .O(N__76396),
            .I(shift_srl_52Z0Z_3));
    InMux I__13441 (
            .O(N__76393),
            .I(N__76390));
    LocalMux I__13440 (
            .O(N__76390),
            .I(shift_srl_52Z0Z_4));
    InMux I__13439 (
            .O(N__76387),
            .I(N__76384));
    LocalMux I__13438 (
            .O(N__76384),
            .I(shift_srl_50Z0Z_10));
    InMux I__13437 (
            .O(N__76381),
            .I(N__76378));
    LocalMux I__13436 (
            .O(N__76378),
            .I(shift_srl_50Z0Z_5));
    InMux I__13435 (
            .O(N__76375),
            .I(N__76372));
    LocalMux I__13434 (
            .O(N__76372),
            .I(shift_srl_50Z0Z_6));
    InMux I__13433 (
            .O(N__76369),
            .I(N__76366));
    LocalMux I__13432 (
            .O(N__76366),
            .I(shift_srl_50Z0Z_9));
    InMux I__13431 (
            .O(N__76363),
            .I(N__76360));
    LocalMux I__13430 (
            .O(N__76360),
            .I(shift_srl_50Z0Z_7));
    InMux I__13429 (
            .O(N__76357),
            .I(N__76354));
    LocalMux I__13428 (
            .O(N__76354),
            .I(shift_srl_50Z0Z_8));
    InMux I__13427 (
            .O(N__76351),
            .I(N__76348));
    LocalMux I__13426 (
            .O(N__76348),
            .I(N__76343));
    InMux I__13425 (
            .O(N__76347),
            .I(N__76340));
    InMux I__13424 (
            .O(N__76346),
            .I(N__76337));
    Span4Mux_h I__13423 (
            .O(N__76343),
            .I(N__76334));
    LocalMux I__13422 (
            .O(N__76340),
            .I(shift_srl_50Z0Z_15));
    LocalMux I__13421 (
            .O(N__76337),
            .I(shift_srl_50Z0Z_15));
    Odrv4 I__13420 (
            .O(N__76334),
            .I(shift_srl_50Z0Z_15));
    InMux I__13419 (
            .O(N__76327),
            .I(N__76324));
    LocalMux I__13418 (
            .O(N__76324),
            .I(shift_srl_50Z0Z_0));
    InMux I__13417 (
            .O(N__76321),
            .I(N__76317));
    InMux I__13416 (
            .O(N__76320),
            .I(N__76314));
    LocalMux I__13415 (
            .O(N__76317),
            .I(shift_srl_47Z0Z_15));
    LocalMux I__13414 (
            .O(N__76314),
            .I(shift_srl_47Z0Z_15));
    InMux I__13413 (
            .O(N__76309),
            .I(N__76306));
    LocalMux I__13412 (
            .O(N__76306),
            .I(shift_srl_47Z0Z_10));
    InMux I__13411 (
            .O(N__76303),
            .I(N__76300));
    LocalMux I__13410 (
            .O(N__76300),
            .I(shift_srl_47Z0Z_11));
    InMux I__13409 (
            .O(N__76297),
            .I(N__76294));
    LocalMux I__13408 (
            .O(N__76294),
            .I(shift_srl_47Z0Z_12));
    InMux I__13407 (
            .O(N__76291),
            .I(N__76288));
    LocalMux I__13406 (
            .O(N__76288),
            .I(shift_srl_47Z0Z_13));
    InMux I__13405 (
            .O(N__76285),
            .I(N__76282));
    LocalMux I__13404 (
            .O(N__76282),
            .I(shift_srl_47Z0Z_14));
    InMux I__13403 (
            .O(N__76279),
            .I(N__76276));
    LocalMux I__13402 (
            .O(N__76276),
            .I(shift_srl_47Z0Z_6));
    InMux I__13401 (
            .O(N__76273),
            .I(N__76270));
    LocalMux I__13400 (
            .O(N__76270),
            .I(shift_srl_47Z0Z_9));
    InMux I__13399 (
            .O(N__76267),
            .I(N__76264));
    LocalMux I__13398 (
            .O(N__76264),
            .I(shift_srl_47Z0Z_7));
    InMux I__13397 (
            .O(N__76261),
            .I(N__76258));
    LocalMux I__13396 (
            .O(N__76258),
            .I(shift_srl_47Z0Z_8));
    CEMux I__13395 (
            .O(N__76255),
            .I(N__76251));
    CEMux I__13394 (
            .O(N__76254),
            .I(N__76248));
    LocalMux I__13393 (
            .O(N__76251),
            .I(clk_en_47));
    LocalMux I__13392 (
            .O(N__76248),
            .I(clk_en_47));
    InMux I__13391 (
            .O(N__76243),
            .I(N__76240));
    LocalMux I__13390 (
            .O(N__76240),
            .I(shift_srl_193Z0Z_6));
    InMux I__13389 (
            .O(N__76237),
            .I(N__76234));
    LocalMux I__13388 (
            .O(N__76234),
            .I(shift_srl_193Z0Z_7));
    CEMux I__13387 (
            .O(N__76231),
            .I(N__76228));
    LocalMux I__13386 (
            .O(N__76228),
            .I(N__76225));
    Span4Mux_v I__13385 (
            .O(N__76225),
            .I(N__76221));
    CEMux I__13384 (
            .O(N__76224),
            .I(N__76218));
    Sp12to4 I__13383 (
            .O(N__76221),
            .I(N__76213));
    LocalMux I__13382 (
            .O(N__76218),
            .I(N__76213));
    Odrv12 I__13381 (
            .O(N__76213),
            .I(clk_en_193));
    InMux I__13380 (
            .O(N__76210),
            .I(N__76206));
    InMux I__13379 (
            .O(N__76209),
            .I(N__76203));
    LocalMux I__13378 (
            .O(N__76206),
            .I(N__76196));
    LocalMux I__13377 (
            .O(N__76203),
            .I(N__76196));
    InMux I__13376 (
            .O(N__76202),
            .I(N__76191));
    InMux I__13375 (
            .O(N__76201),
            .I(N__76191));
    Span4Mux_v I__13374 (
            .O(N__76196),
            .I(N__76184));
    LocalMux I__13373 (
            .O(N__76191),
            .I(N__76184));
    InMux I__13372 (
            .O(N__76190),
            .I(N__76181));
    InMux I__13371 (
            .O(N__76189),
            .I(N__76178));
    Span4Mux_v I__13370 (
            .O(N__76184),
            .I(N__76175));
    LocalMux I__13369 (
            .O(N__76181),
            .I(shift_srl_45Z0Z_15));
    LocalMux I__13368 (
            .O(N__76178),
            .I(shift_srl_45Z0Z_15));
    Odrv4 I__13367 (
            .O(N__76175),
            .I(shift_srl_45Z0Z_15));
    IoInMux I__13366 (
            .O(N__76168),
            .I(N__76165));
    LocalMux I__13365 (
            .O(N__76165),
            .I(N__76162));
    Odrv12 I__13364 (
            .O(N__76162),
            .I(rco_c_45));
    InMux I__13363 (
            .O(N__76159),
            .I(N__76156));
    LocalMux I__13362 (
            .O(N__76156),
            .I(shift_srl_47Z0Z_0));
    InMux I__13361 (
            .O(N__76153),
            .I(N__76150));
    LocalMux I__13360 (
            .O(N__76150),
            .I(shift_srl_47Z0Z_1));
    InMux I__13359 (
            .O(N__76147),
            .I(N__76144));
    LocalMux I__13358 (
            .O(N__76144),
            .I(shift_srl_47Z0Z_2));
    InMux I__13357 (
            .O(N__76141),
            .I(N__76138));
    LocalMux I__13356 (
            .O(N__76138),
            .I(shift_srl_47Z0Z_3));
    InMux I__13355 (
            .O(N__76135),
            .I(N__76132));
    LocalMux I__13354 (
            .O(N__76132),
            .I(shift_srl_47Z0Z_4));
    InMux I__13353 (
            .O(N__76129),
            .I(N__76126));
    LocalMux I__13352 (
            .O(N__76126),
            .I(shift_srl_47Z0Z_5));
    InMux I__13351 (
            .O(N__76123),
            .I(N__76120));
    LocalMux I__13350 (
            .O(N__76120),
            .I(shift_srl_193Z0Z_14));
    InMux I__13349 (
            .O(N__76117),
            .I(N__76114));
    LocalMux I__13348 (
            .O(N__76114),
            .I(shift_srl_193Z0Z_9));
    InMux I__13347 (
            .O(N__76111),
            .I(N__76108));
    LocalMux I__13346 (
            .O(N__76108),
            .I(shift_srl_193Z0Z_8));
    InMux I__13345 (
            .O(N__76105),
            .I(N__76102));
    LocalMux I__13344 (
            .O(N__76102),
            .I(N__76098));
    InMux I__13343 (
            .O(N__76101),
            .I(N__76095));
    Span4Mux_h I__13342 (
            .O(N__76098),
            .I(N__76092));
    LocalMux I__13341 (
            .O(N__76095),
            .I(shift_srl_193Z0Z_15));
    Odrv4 I__13340 (
            .O(N__76092),
            .I(shift_srl_193Z0Z_15));
    InMux I__13339 (
            .O(N__76087),
            .I(N__76084));
    LocalMux I__13338 (
            .O(N__76084),
            .I(shift_srl_193Z0Z_0));
    InMux I__13337 (
            .O(N__76081),
            .I(N__76078));
    LocalMux I__13336 (
            .O(N__76078),
            .I(shift_srl_193Z0Z_1));
    InMux I__13335 (
            .O(N__76075),
            .I(N__76072));
    LocalMux I__13334 (
            .O(N__76072),
            .I(shift_srl_193Z0Z_2));
    InMux I__13333 (
            .O(N__76069),
            .I(N__76066));
    LocalMux I__13332 (
            .O(N__76066),
            .I(shift_srl_193Z0Z_3));
    InMux I__13331 (
            .O(N__76063),
            .I(N__76060));
    LocalMux I__13330 (
            .O(N__76060),
            .I(shift_srl_193Z0Z_4));
    InMux I__13329 (
            .O(N__76057),
            .I(N__76054));
    LocalMux I__13328 (
            .O(N__76054),
            .I(shift_srl_193Z0Z_5));
    InMux I__13327 (
            .O(N__76051),
            .I(N__76044));
    InMux I__13326 (
            .O(N__76050),
            .I(N__76035));
    InMux I__13325 (
            .O(N__76049),
            .I(N__76035));
    InMux I__13324 (
            .O(N__76048),
            .I(N__76035));
    InMux I__13323 (
            .O(N__76047),
            .I(N__76035));
    LocalMux I__13322 (
            .O(N__76044),
            .I(N__76032));
    LocalMux I__13321 (
            .O(N__76035),
            .I(N__76029));
    Odrv4 I__13320 (
            .O(N__76032),
            .I(shift_srl_175Z0Z_15));
    Odrv4 I__13319 (
            .O(N__76029),
            .I(shift_srl_175Z0Z_15));
    InMux I__13318 (
            .O(N__76024),
            .I(N__76019));
    InMux I__13317 (
            .O(N__76023),
            .I(N__76016));
    CascadeMux I__13316 (
            .O(N__76022),
            .I(N__76011));
    LocalMux I__13315 (
            .O(N__76019),
            .I(N__76005));
    LocalMux I__13314 (
            .O(N__76016),
            .I(N__76005));
    InMux I__13313 (
            .O(N__76015),
            .I(N__75996));
    InMux I__13312 (
            .O(N__76014),
            .I(N__75996));
    InMux I__13311 (
            .O(N__76011),
            .I(N__75996));
    InMux I__13310 (
            .O(N__76010),
            .I(N__75996));
    Span4Mux_h I__13309 (
            .O(N__76005),
            .I(N__75991));
    LocalMux I__13308 (
            .O(N__75996),
            .I(N__75991));
    Span4Mux_v I__13307 (
            .O(N__75991),
            .I(N__75987));
    InMux I__13306 (
            .O(N__75990),
            .I(N__75984));
    Span4Mux_v I__13305 (
            .O(N__75987),
            .I(N__75981));
    LocalMux I__13304 (
            .O(N__75984),
            .I(shift_srl_174Z0Z_15));
    Odrv4 I__13303 (
            .O(N__75981),
            .I(shift_srl_174Z0Z_15));
    InMux I__13302 (
            .O(N__75976),
            .I(N__75973));
    LocalMux I__13301 (
            .O(N__75973),
            .I(N__75970));
    Span4Mux_v I__13300 (
            .O(N__75970),
            .I(N__75966));
    InMux I__13299 (
            .O(N__75969),
            .I(N__75962));
    Span4Mux_h I__13298 (
            .O(N__75966),
            .I(N__75959));
    InMux I__13297 (
            .O(N__75965),
            .I(N__75956));
    LocalMux I__13296 (
            .O(N__75962),
            .I(N__75953));
    Sp12to4 I__13295 (
            .O(N__75959),
            .I(N__75949));
    LocalMux I__13294 (
            .O(N__75956),
            .I(N__75946));
    Span4Mux_v I__13293 (
            .O(N__75953),
            .I(N__75943));
    InMux I__13292 (
            .O(N__75952),
            .I(N__75940));
    Span12Mux_v I__13291 (
            .O(N__75949),
            .I(N__75932));
    Span4Mux_v I__13290 (
            .O(N__75946),
            .I(N__75929));
    Span4Mux_v I__13289 (
            .O(N__75943),
            .I(N__75924));
    LocalMux I__13288 (
            .O(N__75940),
            .I(N__75924));
    InMux I__13287 (
            .O(N__75939),
            .I(N__75913));
    InMux I__13286 (
            .O(N__75938),
            .I(N__75913));
    InMux I__13285 (
            .O(N__75937),
            .I(N__75913));
    InMux I__13284 (
            .O(N__75936),
            .I(N__75913));
    InMux I__13283 (
            .O(N__75935),
            .I(N__75913));
    Odrv12 I__13282 (
            .O(N__75932),
            .I(shift_srl_173Z0Z_15));
    Odrv4 I__13281 (
            .O(N__75929),
            .I(shift_srl_173Z0Z_15));
    Odrv4 I__13280 (
            .O(N__75924),
            .I(shift_srl_173Z0Z_15));
    LocalMux I__13279 (
            .O(N__75913),
            .I(shift_srl_173Z0Z_15));
    InMux I__13278 (
            .O(N__75904),
            .I(N__75901));
    LocalMux I__13277 (
            .O(N__75901),
            .I(N__75897));
    InMux I__13276 (
            .O(N__75900),
            .I(N__75894));
    Span4Mux_h I__13275 (
            .O(N__75897),
            .I(N__75891));
    LocalMux I__13274 (
            .O(N__75894),
            .I(shift_srl_182Z0Z_15));
    Odrv4 I__13273 (
            .O(N__75891),
            .I(shift_srl_182Z0Z_15));
    CascadeMux I__13272 (
            .O(N__75886),
            .I(N__75882));
    InMux I__13271 (
            .O(N__75885),
            .I(N__75877));
    InMux I__13270 (
            .O(N__75882),
            .I(N__75877));
    LocalMux I__13269 (
            .O(N__75877),
            .I(N__75872));
    InMux I__13268 (
            .O(N__75876),
            .I(N__75869));
    InMux I__13267 (
            .O(N__75875),
            .I(N__75866));
    Span4Mux_v I__13266 (
            .O(N__75872),
            .I(N__75863));
    LocalMux I__13265 (
            .O(N__75869),
            .I(N__75860));
    LocalMux I__13264 (
            .O(N__75866),
            .I(shift_srl_181Z0Z_15));
    Odrv4 I__13263 (
            .O(N__75863),
            .I(shift_srl_181Z0Z_15));
    Odrv4 I__13262 (
            .O(N__75860),
            .I(shift_srl_181Z0Z_15));
    CascadeMux I__13261 (
            .O(N__75853),
            .I(shift_srl_176_RNIUGI51Z0Z_15_cascade_));
    InMux I__13260 (
            .O(N__75850),
            .I(N__75847));
    LocalMux I__13259 (
            .O(N__75847),
            .I(N__75844));
    Span4Mux_v I__13258 (
            .O(N__75844),
            .I(N__75841));
    Span4Mux_v I__13257 (
            .O(N__75841),
            .I(N__75838));
    Span4Mux_v I__13256 (
            .O(N__75838),
            .I(N__75834));
    InMux I__13255 (
            .O(N__75837),
            .I(N__75831));
    Span4Mux_v I__13254 (
            .O(N__75834),
            .I(N__75824));
    LocalMux I__13253 (
            .O(N__75831),
            .I(N__75824));
    InMux I__13252 (
            .O(N__75830),
            .I(N__75819));
    InMux I__13251 (
            .O(N__75829),
            .I(N__75819));
    Span4Mux_h I__13250 (
            .O(N__75824),
            .I(N__75816));
    LocalMux I__13249 (
            .O(N__75819),
            .I(N__75813));
    Span4Mux_v I__13248 (
            .O(N__75816),
            .I(N__75810));
    Span12Mux_v I__13247 (
            .O(N__75813),
            .I(N__75807));
    Odrv4 I__13246 (
            .O(N__75810),
            .I(shift_srl_182_RNIEPSC2Z0Z_15));
    Odrv12 I__13245 (
            .O(N__75807),
            .I(shift_srl_182_RNIEPSC2Z0Z_15));
    InMux I__13244 (
            .O(N__75802),
            .I(N__75799));
    LocalMux I__13243 (
            .O(N__75799),
            .I(shift_srl_193Z0Z_10));
    InMux I__13242 (
            .O(N__75796),
            .I(N__75793));
    LocalMux I__13241 (
            .O(N__75793),
            .I(shift_srl_193Z0Z_11));
    InMux I__13240 (
            .O(N__75790),
            .I(N__75787));
    LocalMux I__13239 (
            .O(N__75787),
            .I(shift_srl_193Z0Z_12));
    InMux I__13238 (
            .O(N__75784),
            .I(N__75781));
    LocalMux I__13237 (
            .O(N__75781),
            .I(shift_srl_193Z0Z_13));
    InMux I__13236 (
            .O(N__75778),
            .I(N__75775));
    LocalMux I__13235 (
            .O(N__75775),
            .I(shift_srl_176Z0Z_12));
    InMux I__13234 (
            .O(N__75772),
            .I(N__75769));
    LocalMux I__13233 (
            .O(N__75769),
            .I(shift_srl_176Z0Z_13));
    InMux I__13232 (
            .O(N__75766),
            .I(N__75763));
    LocalMux I__13231 (
            .O(N__75763),
            .I(shift_srl_176Z0Z_14));
    InMux I__13230 (
            .O(N__75760),
            .I(N__75757));
    LocalMux I__13229 (
            .O(N__75757),
            .I(shift_srl_176Z0Z_9));
    InMux I__13228 (
            .O(N__75754),
            .I(N__75751));
    LocalMux I__13227 (
            .O(N__75751),
            .I(shift_srl_176Z0Z_8));
    IoInMux I__13226 (
            .O(N__75748),
            .I(N__75745));
    LocalMux I__13225 (
            .O(N__75745),
            .I(N__75742));
    Span4Mux_s2_v I__13224 (
            .O(N__75742),
            .I(N__75739));
    Span4Mux_v I__13223 (
            .O(N__75739),
            .I(N__75736));
    Odrv4 I__13222 (
            .O(N__75736),
            .I(rco_c_175));
    IoInMux I__13221 (
            .O(N__75733),
            .I(N__75730));
    LocalMux I__13220 (
            .O(N__75730),
            .I(N__75727));
    IoSpan4Mux I__13219 (
            .O(N__75727),
            .I(N__75724));
    Span4Mux_s0_v I__13218 (
            .O(N__75724),
            .I(N__75721));
    Span4Mux_v I__13217 (
            .O(N__75721),
            .I(N__75718));
    Odrv4 I__13216 (
            .O(N__75718),
            .I(rco_c_174));
    CascadeMux I__13215 (
            .O(N__75715),
            .I(clk_en_0_a3_0_a2cf1_176_cascade_));
    InMux I__13214 (
            .O(N__75712),
            .I(N__75709));
    LocalMux I__13213 (
            .O(N__75709),
            .I(shift_srl_181Z0Z_1));
    InMux I__13212 (
            .O(N__75706),
            .I(N__75703));
    LocalMux I__13211 (
            .O(N__75703),
            .I(shift_srl_181Z0Z_2));
    InMux I__13210 (
            .O(N__75700),
            .I(N__75697));
    LocalMux I__13209 (
            .O(N__75697),
            .I(shift_srl_181Z0Z_3));
    InMux I__13208 (
            .O(N__75694),
            .I(N__75691));
    LocalMux I__13207 (
            .O(N__75691),
            .I(shift_srl_181Z0Z_4));
    InMux I__13206 (
            .O(N__75688),
            .I(N__75685));
    LocalMux I__13205 (
            .O(N__75685),
            .I(shift_srl_181Z0Z_5));
    InMux I__13204 (
            .O(N__75682),
            .I(N__75679));
    LocalMux I__13203 (
            .O(N__75679),
            .I(shift_srl_181Z0Z_0));
    InMux I__13202 (
            .O(N__75676),
            .I(N__75673));
    LocalMux I__13201 (
            .O(N__75673),
            .I(shift_srl_176Z0Z_10));
    InMux I__13200 (
            .O(N__75670),
            .I(N__75667));
    LocalMux I__13199 (
            .O(N__75667),
            .I(shift_srl_176Z0Z_11));
    InMux I__13198 (
            .O(N__75664),
            .I(N__75661));
    LocalMux I__13197 (
            .O(N__75661),
            .I(shift_srl_178Z0Z_0));
    InMux I__13196 (
            .O(N__75658),
            .I(N__75655));
    LocalMux I__13195 (
            .O(N__75655),
            .I(shift_srl_178Z0Z_1));
    InMux I__13194 (
            .O(N__75652),
            .I(N__75649));
    LocalMux I__13193 (
            .O(N__75649),
            .I(shift_srl_178Z0Z_2));
    InMux I__13192 (
            .O(N__75646),
            .I(N__75643));
    LocalMux I__13191 (
            .O(N__75643),
            .I(shift_srl_178Z0Z_3));
    InMux I__13190 (
            .O(N__75640),
            .I(N__75637));
    LocalMux I__13189 (
            .O(N__75637),
            .I(shift_srl_178Z0Z_4));
    InMux I__13188 (
            .O(N__75634),
            .I(N__75631));
    LocalMux I__13187 (
            .O(N__75631),
            .I(shift_srl_178Z0Z_9));
    InMux I__13186 (
            .O(N__75628),
            .I(N__75625));
    LocalMux I__13185 (
            .O(N__75625),
            .I(shift_srl_179Z0Z_6));
    InMux I__13184 (
            .O(N__75622),
            .I(N__75619));
    LocalMux I__13183 (
            .O(N__75619),
            .I(shift_srl_186Z0Z_10));
    InMux I__13182 (
            .O(N__75616),
            .I(N__75613));
    LocalMux I__13181 (
            .O(N__75613),
            .I(shift_srl_186Z0Z_11));
    InMux I__13180 (
            .O(N__75610),
            .I(N__75607));
    LocalMux I__13179 (
            .O(N__75607),
            .I(shift_srl_186Z0Z_12));
    InMux I__13178 (
            .O(N__75604),
            .I(N__75601));
    LocalMux I__13177 (
            .O(N__75601),
            .I(shift_srl_186Z0Z_13));
    InMux I__13176 (
            .O(N__75598),
            .I(N__75595));
    LocalMux I__13175 (
            .O(N__75595),
            .I(shift_srl_186Z0Z_14));
    InMux I__13174 (
            .O(N__75592),
            .I(N__75589));
    LocalMux I__13173 (
            .O(N__75589),
            .I(shift_srl_186Z0Z_9));
    InMux I__13172 (
            .O(N__75586),
            .I(N__75583));
    LocalMux I__13171 (
            .O(N__75583),
            .I(shift_srl_186Z0Z_7));
    InMux I__13170 (
            .O(N__75580),
            .I(N__75577));
    LocalMux I__13169 (
            .O(N__75577),
            .I(shift_srl_186Z0Z_8));
    CEMux I__13168 (
            .O(N__75574),
            .I(N__75571));
    LocalMux I__13167 (
            .O(N__75571),
            .I(N__75568));
    Span4Mux_v I__13166 (
            .O(N__75568),
            .I(N__75564));
    CEMux I__13165 (
            .O(N__75567),
            .I(N__75561));
    Span4Mux_h I__13164 (
            .O(N__75564),
            .I(N__75558));
    LocalMux I__13163 (
            .O(N__75561),
            .I(N__75555));
    Odrv4 I__13162 (
            .O(N__75558),
            .I(clk_en_186));
    Odrv12 I__13161 (
            .O(N__75555),
            .I(clk_en_186));
    InMux I__13160 (
            .O(N__75550),
            .I(N__75547));
    LocalMux I__13159 (
            .O(N__75547),
            .I(shift_srl_171Z0Z_6));
    InMux I__13158 (
            .O(N__75544),
            .I(N__75541));
    LocalMux I__13157 (
            .O(N__75541),
            .I(shift_srl_171Z0Z_7));
    InMux I__13156 (
            .O(N__75538),
            .I(N__75535));
    LocalMux I__13155 (
            .O(N__75535),
            .I(shift_srl_179Z0Z_0));
    InMux I__13154 (
            .O(N__75532),
            .I(N__75529));
    LocalMux I__13153 (
            .O(N__75529),
            .I(shift_srl_179Z0Z_1));
    InMux I__13152 (
            .O(N__75526),
            .I(N__75523));
    LocalMux I__13151 (
            .O(N__75523),
            .I(shift_srl_179Z0Z_2));
    InMux I__13150 (
            .O(N__75520),
            .I(N__75517));
    LocalMux I__13149 (
            .O(N__75517),
            .I(shift_srl_179Z0Z_3));
    InMux I__13148 (
            .O(N__75514),
            .I(N__75511));
    LocalMux I__13147 (
            .O(N__75511),
            .I(shift_srl_179Z0Z_4));
    InMux I__13146 (
            .O(N__75508),
            .I(N__75505));
    LocalMux I__13145 (
            .O(N__75505),
            .I(shift_srl_179Z0Z_5));
    InMux I__13144 (
            .O(N__75502),
            .I(N__75499));
    LocalMux I__13143 (
            .O(N__75499),
            .I(shift_srl_159Z0Z_3));
    InMux I__13142 (
            .O(N__75496),
            .I(N__75493));
    LocalMux I__13141 (
            .O(N__75493),
            .I(shift_srl_159Z0Z_4));
    InMux I__13140 (
            .O(N__75490),
            .I(N__75487));
    LocalMux I__13139 (
            .O(N__75487),
            .I(shift_srl_159Z0Z_7));
    InMux I__13138 (
            .O(N__75484),
            .I(N__75481));
    LocalMux I__13137 (
            .O(N__75481),
            .I(shift_srl_159Z0Z_8));
    InMux I__13136 (
            .O(N__75478),
            .I(N__75475));
    LocalMux I__13135 (
            .O(N__75475),
            .I(shift_srl_159Z0Z_1));
    InMux I__13134 (
            .O(N__75472),
            .I(N__75469));
    LocalMux I__13133 (
            .O(N__75469),
            .I(shift_srl_159Z0Z_2));
    InMux I__13132 (
            .O(N__75466),
            .I(N__75463));
    LocalMux I__13131 (
            .O(N__75463),
            .I(shift_srl_171Z0Z_2));
    InMux I__13130 (
            .O(N__75460),
            .I(N__75457));
    LocalMux I__13129 (
            .O(N__75457),
            .I(shift_srl_171Z0Z_3));
    InMux I__13128 (
            .O(N__75454),
            .I(N__75451));
    LocalMux I__13127 (
            .O(N__75451),
            .I(shift_srl_171Z0Z_4));
    InMux I__13126 (
            .O(N__75448),
            .I(N__75445));
    LocalMux I__13125 (
            .O(N__75445),
            .I(shift_srl_171Z0Z_5));
    InMux I__13124 (
            .O(N__75442),
            .I(N__75439));
    LocalMux I__13123 (
            .O(N__75439),
            .I(shift_srl_159Z0Z_10));
    InMux I__13122 (
            .O(N__75436),
            .I(N__75433));
    LocalMux I__13121 (
            .O(N__75433),
            .I(shift_srl_159Z0Z_9));
    InMux I__13120 (
            .O(N__75430),
            .I(N__75427));
    LocalMux I__13119 (
            .O(N__75427),
            .I(shift_srl_159Z0Z_11));
    InMux I__13118 (
            .O(N__75424),
            .I(N__75421));
    LocalMux I__13117 (
            .O(N__75421),
            .I(shift_srl_159Z0Z_12));
    InMux I__13116 (
            .O(N__75418),
            .I(N__75415));
    LocalMux I__13115 (
            .O(N__75415),
            .I(shift_srl_159Z0Z_5));
    InMux I__13114 (
            .O(N__75412),
            .I(N__75409));
    LocalMux I__13113 (
            .O(N__75409),
            .I(shift_srl_159Z0Z_13));
    InMux I__13112 (
            .O(N__75406),
            .I(N__75403));
    LocalMux I__13111 (
            .O(N__75403),
            .I(shift_srl_159Z0Z_0));
    InMux I__13110 (
            .O(N__75400),
            .I(N__75397));
    LocalMux I__13109 (
            .O(N__75397),
            .I(shift_srl_159Z0Z_6));
    IoInMux I__13108 (
            .O(N__75394),
            .I(N__75391));
    LocalMux I__13107 (
            .O(N__75391),
            .I(N__75388));
    Span12Mux_s6_v I__13106 (
            .O(N__75388),
            .I(N__75385));
    Span12Mux_h I__13105 (
            .O(N__75385),
            .I(N__75382));
    Odrv12 I__13104 (
            .O(N__75382),
            .I(rco_c_61));
    IoInMux I__13103 (
            .O(N__75379),
            .I(N__75376));
    LocalMux I__13102 (
            .O(N__75376),
            .I(N__75373));
    Span4Mux_s1_v I__13101 (
            .O(N__75373),
            .I(N__75370));
    Sp12to4 I__13100 (
            .O(N__75370),
            .I(N__75367));
    Span12Mux_h I__13099 (
            .O(N__75367),
            .I(N__75364));
    Span12Mux_v I__13098 (
            .O(N__75364),
            .I(N__75361));
    Odrv12 I__13097 (
            .O(N__75361),
            .I(rco_c_62));
    IoInMux I__13096 (
            .O(N__75358),
            .I(N__75355));
    LocalMux I__13095 (
            .O(N__75355),
            .I(N__75352));
    IoSpan4Mux I__13094 (
            .O(N__75352),
            .I(N__75349));
    IoSpan4Mux I__13093 (
            .O(N__75349),
            .I(N__75346));
    Span4Mux_s3_v I__13092 (
            .O(N__75346),
            .I(N__75343));
    Span4Mux_h I__13091 (
            .O(N__75343),
            .I(N__75340));
    Sp12to4 I__13090 (
            .O(N__75340),
            .I(N__75337));
    Odrv12 I__13089 (
            .O(N__75337),
            .I(rco_c_65));
    InMux I__13088 (
            .O(N__75334),
            .I(N__75325));
    InMux I__13087 (
            .O(N__75333),
            .I(N__75325));
    InMux I__13086 (
            .O(N__75332),
            .I(N__75318));
    InMux I__13085 (
            .O(N__75331),
            .I(N__75318));
    InMux I__13084 (
            .O(N__75330),
            .I(N__75318));
    LocalMux I__13083 (
            .O(N__75325),
            .I(N__75315));
    LocalMux I__13082 (
            .O(N__75318),
            .I(N__75312));
    Span4Mux_v I__13081 (
            .O(N__75315),
            .I(N__75307));
    Span4Mux_h I__13080 (
            .O(N__75312),
            .I(N__75307));
    Odrv4 I__13079 (
            .O(N__75307),
            .I(shift_srl_60Z0Z_15));
    InMux I__13078 (
            .O(N__75304),
            .I(N__75301));
    LocalMux I__13077 (
            .O(N__75301),
            .I(shift_srl_60Z0Z_0));
    InMux I__13076 (
            .O(N__75298),
            .I(N__75295));
    LocalMux I__13075 (
            .O(N__75295),
            .I(shift_srl_60Z0Z_1));
    InMux I__13074 (
            .O(N__75292),
            .I(N__75289));
    LocalMux I__13073 (
            .O(N__75289),
            .I(shift_srl_60Z0Z_2));
    InMux I__13072 (
            .O(N__75286),
            .I(N__75283));
    LocalMux I__13071 (
            .O(N__75283),
            .I(N__75280));
    Odrv12 I__13070 (
            .O(N__75280),
            .I(shift_srl_60Z0Z_3));
    InMux I__13069 (
            .O(N__75277),
            .I(N__75274));
    LocalMux I__13068 (
            .O(N__75274),
            .I(shift_srl_63Z0Z_0));
    InMux I__13067 (
            .O(N__75271),
            .I(N__75268));
    LocalMux I__13066 (
            .O(N__75268),
            .I(shift_srl_63Z0Z_1));
    InMux I__13065 (
            .O(N__75265),
            .I(N__75262));
    LocalMux I__13064 (
            .O(N__75262),
            .I(shift_srl_63Z0Z_2));
    InMux I__13063 (
            .O(N__75259),
            .I(N__75256));
    LocalMux I__13062 (
            .O(N__75256),
            .I(shift_srl_63Z0Z_3));
    InMux I__13061 (
            .O(N__75253),
            .I(N__75250));
    LocalMux I__13060 (
            .O(N__75250),
            .I(shift_srl_63Z0Z_4));
    InMux I__13059 (
            .O(N__75247),
            .I(N__75244));
    LocalMux I__13058 (
            .O(N__75244),
            .I(shift_srl_63Z0Z_5));
    InMux I__13057 (
            .O(N__75241),
            .I(N__75238));
    LocalMux I__13056 (
            .O(N__75238),
            .I(shift_srl_63Z0Z_6));
    IoInMux I__13055 (
            .O(N__75235),
            .I(N__75232));
    LocalMux I__13054 (
            .O(N__75232),
            .I(N__75229));
    Span12Mux_s3_v I__13053 (
            .O(N__75229),
            .I(N__75226));
    Span12Mux_v I__13052 (
            .O(N__75226),
            .I(N__75223));
    Span12Mux_h I__13051 (
            .O(N__75223),
            .I(N__75220));
    Odrv12 I__13050 (
            .O(N__75220),
            .I(rco_c_60));
    InMux I__13049 (
            .O(N__75217),
            .I(N__75214));
    LocalMux I__13048 (
            .O(N__75214),
            .I(shift_srl_61_RNI3LM9Z0Z_15));
    InMux I__13047 (
            .O(N__75211),
            .I(N__75208));
    LocalMux I__13046 (
            .O(N__75208),
            .I(shift_srl_60Z0Z_4));
    InMux I__13045 (
            .O(N__75205),
            .I(N__75202));
    LocalMux I__13044 (
            .O(N__75202),
            .I(shift_srl_60Z0Z_5));
    InMux I__13043 (
            .O(N__75199),
            .I(N__75196));
    LocalMux I__13042 (
            .O(N__75196),
            .I(shift_srl_60Z0Z_6));
    InMux I__13041 (
            .O(N__75193),
            .I(N__75190));
    LocalMux I__13040 (
            .O(N__75190),
            .I(shift_srl_60Z0Z_7));
    InMux I__13039 (
            .O(N__75187),
            .I(N__75184));
    LocalMux I__13038 (
            .O(N__75184),
            .I(N__75181));
    Span4Mux_h I__13037 (
            .O(N__75181),
            .I(N__75178));
    Span4Mux_v I__13036 (
            .O(N__75178),
            .I(N__75172));
    InMux I__13035 (
            .O(N__75177),
            .I(N__75165));
    InMux I__13034 (
            .O(N__75176),
            .I(N__75165));
    InMux I__13033 (
            .O(N__75175),
            .I(N__75165));
    Odrv4 I__13032 (
            .O(N__75172),
            .I(rco_int_0_a2_0_a2_sx_153));
    LocalMux I__13031 (
            .O(N__75165),
            .I(rco_int_0_a2_0_a2_sx_153));
    CascadeMux I__13030 (
            .O(N__75160),
            .I(clk_en_0_a3_0_a2_sx_179_cascade_));
    InMux I__13029 (
            .O(N__75157),
            .I(N__75154));
    LocalMux I__13028 (
            .O(N__75154),
            .I(N__75151));
    Odrv4 I__13027 (
            .O(N__75151),
            .I(rco_int_0_a2_0_a2_93_m6_0_a2_4_7_0));
    InMux I__13026 (
            .O(N__75148),
            .I(N__75138));
    InMux I__13025 (
            .O(N__75147),
            .I(N__75138));
    InMux I__13024 (
            .O(N__75146),
            .I(N__75138));
    InMux I__13023 (
            .O(N__75145),
            .I(N__75132));
    LocalMux I__13022 (
            .O(N__75138),
            .I(N__75129));
    InMux I__13021 (
            .O(N__75137),
            .I(N__75124));
    InMux I__13020 (
            .O(N__75136),
            .I(N__75124));
    InMux I__13019 (
            .O(N__75135),
            .I(N__75121));
    LocalMux I__13018 (
            .O(N__75132),
            .I(N__75118));
    Span4Mux_v I__13017 (
            .O(N__75129),
            .I(N__75115));
    LocalMux I__13016 (
            .O(N__75124),
            .I(N__75112));
    LocalMux I__13015 (
            .O(N__75121),
            .I(N__75109));
    Span4Mux_v I__13014 (
            .O(N__75118),
            .I(N__75106));
    Odrv4 I__13013 (
            .O(N__75115),
            .I(rco_int_0_a2_1_a2_0_44));
    Odrv4 I__13012 (
            .O(N__75112),
            .I(rco_int_0_a2_1_a2_0_44));
    Odrv12 I__13011 (
            .O(N__75109),
            .I(rco_int_0_a2_1_a2_0_44));
    Odrv4 I__13010 (
            .O(N__75106),
            .I(rco_int_0_a2_1_a2_0_44));
    CascadeMux I__13009 (
            .O(N__75097),
            .I(rco_int_0_a2_0_a2_93_m6_0_a2_4_7_4_sx_cascade_));
    CascadeMux I__13008 (
            .O(N__75094),
            .I(rco_int_0_a2_0_a2_93_m6_0_a2_4_7_4_cascade_));
    InMux I__13007 (
            .O(N__75091),
            .I(N__75082));
    InMux I__13006 (
            .O(N__75090),
            .I(N__75082));
    InMux I__13005 (
            .O(N__75089),
            .I(N__75082));
    LocalMux I__13004 (
            .O(N__75082),
            .I(N__75074));
    InMux I__13003 (
            .O(N__75081),
            .I(N__75071));
    InMux I__13002 (
            .O(N__75080),
            .I(N__75066));
    InMux I__13001 (
            .O(N__75079),
            .I(N__75066));
    InMux I__13000 (
            .O(N__75078),
            .I(N__75063));
    InMux I__12999 (
            .O(N__75077),
            .I(N__75060));
    Span4Mux_v I__12998 (
            .O(N__75074),
            .I(N__75057));
    LocalMux I__12997 (
            .O(N__75071),
            .I(N__75054));
    LocalMux I__12996 (
            .O(N__75066),
            .I(N__75050));
    LocalMux I__12995 (
            .O(N__75063),
            .I(N__75047));
    LocalMux I__12994 (
            .O(N__75060),
            .I(N__75044));
    Span4Mux_h I__12993 (
            .O(N__75057),
            .I(N__75039));
    Span4Mux_h I__12992 (
            .O(N__75054),
            .I(N__75039));
    InMux I__12991 (
            .O(N__75053),
            .I(N__75036));
    Span4Mux_v I__12990 (
            .O(N__75050),
            .I(N__75032));
    Span4Mux_h I__12989 (
            .O(N__75047),
            .I(N__75029));
    Span4Mux_h I__12988 (
            .O(N__75044),
            .I(N__75026));
    Span4Mux_v I__12987 (
            .O(N__75039),
            .I(N__75021));
    LocalMux I__12986 (
            .O(N__75036),
            .I(N__75021));
    InMux I__12985 (
            .O(N__75035),
            .I(N__75018));
    Span4Mux_h I__12984 (
            .O(N__75032),
            .I(N__75011));
    Span4Mux_v I__12983 (
            .O(N__75029),
            .I(N__75011));
    Span4Mux_v I__12982 (
            .O(N__75026),
            .I(N__75011));
    Span4Mux_h I__12981 (
            .O(N__75021),
            .I(N__75008));
    LocalMux I__12980 (
            .O(N__75018),
            .I(rco_int_0_a2_0_a2_93_m6_0_a2_4_7));
    Odrv4 I__12979 (
            .O(N__75011),
            .I(rco_int_0_a2_0_a2_93_m6_0_a2_4_7));
    Odrv4 I__12978 (
            .O(N__75008),
            .I(rco_int_0_a2_0_a2_93_m6_0_a2_4_7));
    InMux I__12977 (
            .O(N__75001),
            .I(N__74998));
    LocalMux I__12976 (
            .O(N__74998),
            .I(rco_int_0_a3_0_a2_0_0_66));
    InMux I__12975 (
            .O(N__74995),
            .I(N__74992));
    LocalMux I__12974 (
            .O(N__74992),
            .I(shift_srl_60Z0Z_10));
    InMux I__12973 (
            .O(N__74989),
            .I(N__74986));
    LocalMux I__12972 (
            .O(N__74986),
            .I(shift_srl_60Z0Z_11));
    InMux I__12971 (
            .O(N__74983),
            .I(N__74980));
    LocalMux I__12970 (
            .O(N__74980),
            .I(shift_srl_60Z0Z_12));
    InMux I__12969 (
            .O(N__74977),
            .I(N__74974));
    LocalMux I__12968 (
            .O(N__74974),
            .I(shift_srl_60Z0Z_13));
    InMux I__12967 (
            .O(N__74971),
            .I(N__74968));
    LocalMux I__12966 (
            .O(N__74968),
            .I(shift_srl_60Z0Z_9));
    InMux I__12965 (
            .O(N__74965),
            .I(N__74962));
    LocalMux I__12964 (
            .O(N__74962),
            .I(shift_srl_60Z0Z_8));
    InMux I__12963 (
            .O(N__74959),
            .I(N__74956));
    LocalMux I__12962 (
            .O(N__74956),
            .I(shift_srl_60Z0Z_14));
    InMux I__12961 (
            .O(N__74953),
            .I(N__74950));
    LocalMux I__12960 (
            .O(N__74950),
            .I(shift_srl_54Z0Z_10));
    InMux I__12959 (
            .O(N__74947),
            .I(N__74944));
    LocalMux I__12958 (
            .O(N__74944),
            .I(shift_srl_57Z0Z_10));
    InMux I__12957 (
            .O(N__74941),
            .I(N__74938));
    LocalMux I__12956 (
            .O(N__74938),
            .I(shift_srl_57Z0Z_11));
    InMux I__12955 (
            .O(N__74935),
            .I(N__74932));
    LocalMux I__12954 (
            .O(N__74932),
            .I(shift_srl_57Z0Z_12));
    InMux I__12953 (
            .O(N__74929),
            .I(N__74926));
    LocalMux I__12952 (
            .O(N__74926),
            .I(shift_srl_57Z0Z_13));
    InMux I__12951 (
            .O(N__74923),
            .I(N__74920));
    LocalMux I__12950 (
            .O(N__74920),
            .I(shift_srl_57Z0Z_14));
    InMux I__12949 (
            .O(N__74917),
            .I(N__74914));
    LocalMux I__12948 (
            .O(N__74914),
            .I(shift_srl_57Z0Z_9));
    InMux I__12947 (
            .O(N__74911),
            .I(N__74908));
    LocalMux I__12946 (
            .O(N__74908),
            .I(shift_srl_57Z0Z_8));
    CascadeMux I__12945 (
            .O(N__74905),
            .I(rco_c_48_cascade_));
    CEMux I__12944 (
            .O(N__74902),
            .I(N__74898));
    CEMux I__12943 (
            .O(N__74901),
            .I(N__74895));
    LocalMux I__12942 (
            .O(N__74898),
            .I(N__74889));
    LocalMux I__12941 (
            .O(N__74895),
            .I(N__74889));
    CEMux I__12940 (
            .O(N__74894),
            .I(N__74886));
    Span4Mux_v I__12939 (
            .O(N__74889),
            .I(N__74881));
    LocalMux I__12938 (
            .O(N__74886),
            .I(N__74881));
    Span4Mux_v I__12937 (
            .O(N__74881),
            .I(N__74878));
    Odrv4 I__12936 (
            .O(N__74878),
            .I(clk_en_55));
    CascadeMux I__12935 (
            .O(N__74875),
            .I(N__74870));
    InMux I__12934 (
            .O(N__74874),
            .I(N__74867));
    InMux I__12933 (
            .O(N__74873),
            .I(N__74864));
    InMux I__12932 (
            .O(N__74870),
            .I(N__74861));
    LocalMux I__12931 (
            .O(N__74867),
            .I(shift_srl_55Z0Z_15));
    LocalMux I__12930 (
            .O(N__74864),
            .I(shift_srl_55Z0Z_15));
    LocalMux I__12929 (
            .O(N__74861),
            .I(shift_srl_55Z0Z_15));
    InMux I__12928 (
            .O(N__74854),
            .I(N__74851));
    LocalMux I__12927 (
            .O(N__74851),
            .I(shift_srl_54Z0Z_14));
    InMux I__12926 (
            .O(N__74848),
            .I(N__74845));
    LocalMux I__12925 (
            .O(N__74845),
            .I(shift_srl_54Z0Z_13));
    InMux I__12924 (
            .O(N__74842),
            .I(N__74839));
    LocalMux I__12923 (
            .O(N__74839),
            .I(shift_srl_54Z0Z_12));
    InMux I__12922 (
            .O(N__74836),
            .I(N__74833));
    LocalMux I__12921 (
            .O(N__74833),
            .I(shift_srl_54Z0Z_11));
    InMux I__12920 (
            .O(N__74830),
            .I(N__74827));
    LocalMux I__12919 (
            .O(N__74827),
            .I(shift_srl_52Z0Z_13));
    InMux I__12918 (
            .O(N__74824),
            .I(N__74821));
    LocalMux I__12917 (
            .O(N__74821),
            .I(shift_srl_52Z0Z_14));
    InMux I__12916 (
            .O(N__74818),
            .I(N__74815));
    LocalMux I__12915 (
            .O(N__74815),
            .I(shift_srl_52Z0Z_9));
    InMux I__12914 (
            .O(N__74812),
            .I(N__74809));
    LocalMux I__12913 (
            .O(N__74809),
            .I(shift_srl_52Z0Z_8));
    IoInMux I__12912 (
            .O(N__74806),
            .I(N__74803));
    LocalMux I__12911 (
            .O(N__74803),
            .I(N__74800));
    IoSpan4Mux I__12910 (
            .O(N__74800),
            .I(N__74797));
    Sp12to4 I__12909 (
            .O(N__74797),
            .I(N__74794));
    Span12Mux_s9_v I__12908 (
            .O(N__74794),
            .I(N__74791));
    Odrv12 I__12907 (
            .O(N__74791),
            .I(rco_c_52));
    IoInMux I__12906 (
            .O(N__74788),
            .I(N__74785));
    LocalMux I__12905 (
            .O(N__74785),
            .I(N__74782));
    IoSpan4Mux I__12904 (
            .O(N__74782),
            .I(N__74779));
    Span4Mux_s2_v I__12903 (
            .O(N__74779),
            .I(N__74776));
    Sp12to4 I__12902 (
            .O(N__74776),
            .I(N__74773));
    Span12Mux_s9_v I__12901 (
            .O(N__74773),
            .I(N__74770));
    Odrv12 I__12900 (
            .O(N__74770),
            .I(rco_c_51));
    InMux I__12899 (
            .O(N__74767),
            .I(N__74764));
    LocalMux I__12898 (
            .O(N__74764),
            .I(N__74760));
    InMux I__12897 (
            .O(N__74763),
            .I(N__74757));
    Span4Mux_v I__12896 (
            .O(N__74760),
            .I(N__74749));
    LocalMux I__12895 (
            .O(N__74757),
            .I(N__74749));
    InMux I__12894 (
            .O(N__74756),
            .I(N__74742));
    InMux I__12893 (
            .O(N__74755),
            .I(N__74742));
    InMux I__12892 (
            .O(N__74754),
            .I(N__74742));
    Span4Mux_v I__12891 (
            .O(N__74749),
            .I(N__74736));
    LocalMux I__12890 (
            .O(N__74742),
            .I(N__74733));
    InMux I__12889 (
            .O(N__74741),
            .I(N__74730));
    InMux I__12888 (
            .O(N__74740),
            .I(N__74725));
    InMux I__12887 (
            .O(N__74739),
            .I(N__74725));
    Odrv4 I__12886 (
            .O(N__74736),
            .I(rco_int_0_a2_0_a2_0_39));
    Odrv12 I__12885 (
            .O(N__74733),
            .I(rco_int_0_a2_0_a2_0_39));
    LocalMux I__12884 (
            .O(N__74730),
            .I(rco_int_0_a2_0_a2_0_39));
    LocalMux I__12883 (
            .O(N__74725),
            .I(rco_int_0_a2_0_a2_0_39));
    CascadeMux I__12882 (
            .O(N__74716),
            .I(N__74711));
    CascadeMux I__12881 (
            .O(N__74715),
            .I(N__74706));
    InMux I__12880 (
            .O(N__74714),
            .I(N__74701));
    InMux I__12879 (
            .O(N__74711),
            .I(N__74697));
    InMux I__12878 (
            .O(N__74710),
            .I(N__74692));
    InMux I__12877 (
            .O(N__74709),
            .I(N__74692));
    InMux I__12876 (
            .O(N__74706),
            .I(N__74689));
    InMux I__12875 (
            .O(N__74705),
            .I(N__74684));
    InMux I__12874 (
            .O(N__74704),
            .I(N__74684));
    LocalMux I__12873 (
            .O(N__74701),
            .I(N__74681));
    CascadeMux I__12872 (
            .O(N__74700),
            .I(N__74678));
    LocalMux I__12871 (
            .O(N__74697),
            .I(N__74673));
    LocalMux I__12870 (
            .O(N__74692),
            .I(N__74673));
    LocalMux I__12869 (
            .O(N__74689),
            .I(N__74670));
    LocalMux I__12868 (
            .O(N__74684),
            .I(N__74667));
    Sp12to4 I__12867 (
            .O(N__74681),
            .I(N__74664));
    InMux I__12866 (
            .O(N__74678),
            .I(N__74661));
    Span4Mux_v I__12865 (
            .O(N__74673),
            .I(N__74656));
    Span4Mux_v I__12864 (
            .O(N__74670),
            .I(N__74656));
    Span4Mux_v I__12863 (
            .O(N__74667),
            .I(N__74653));
    Span12Mux_v I__12862 (
            .O(N__74664),
            .I(N__74648));
    LocalMux I__12861 (
            .O(N__74661),
            .I(N__74648));
    Span4Mux_v I__12860 (
            .O(N__74656),
            .I(N__74645));
    Odrv4 I__12859 (
            .O(N__74653),
            .I(shift_srl_40Z0Z_15));
    Odrv12 I__12858 (
            .O(N__74648),
            .I(shift_srl_40Z0Z_15));
    Odrv4 I__12857 (
            .O(N__74645),
            .I(shift_srl_40Z0Z_15));
    InMux I__12856 (
            .O(N__74638),
            .I(N__74629));
    InMux I__12855 (
            .O(N__74637),
            .I(N__74629));
    InMux I__12854 (
            .O(N__74636),
            .I(N__74629));
    LocalMux I__12853 (
            .O(N__74629),
            .I(N__74623));
    InMux I__12852 (
            .O(N__74628),
            .I(N__74620));
    InMux I__12851 (
            .O(N__74627),
            .I(N__74617));
    InMux I__12850 (
            .O(N__74626),
            .I(N__74614));
    Span4Mux_h I__12849 (
            .O(N__74623),
            .I(N__74609));
    LocalMux I__12848 (
            .O(N__74620),
            .I(N__74609));
    LocalMux I__12847 (
            .O(N__74617),
            .I(shift_srl_51Z0Z_15));
    LocalMux I__12846 (
            .O(N__74614),
            .I(shift_srl_51Z0Z_15));
    Odrv4 I__12845 (
            .O(N__74609),
            .I(shift_srl_51Z0Z_15));
    CascadeMux I__12844 (
            .O(N__74602),
            .I(shift_srl_47_RNIV3QLZ0Z_15_cascade_));
    IoInMux I__12843 (
            .O(N__74599),
            .I(N__74596));
    LocalMux I__12842 (
            .O(N__74596),
            .I(N__74593));
    Span4Mux_s2_h I__12841 (
            .O(N__74593),
            .I(N__74590));
    Span4Mux_v I__12840 (
            .O(N__74590),
            .I(N__74587));
    Sp12to4 I__12839 (
            .O(N__74587),
            .I(N__74584));
    Odrv12 I__12838 (
            .O(N__74584),
            .I(rco_c_47));
    InMux I__12837 (
            .O(N__74581),
            .I(N__74578));
    LocalMux I__12836 (
            .O(N__74578),
            .I(N__74575));
    Odrv4 I__12835 (
            .O(N__74575),
            .I(shift_srl_50Z0Z_14));
    InMux I__12834 (
            .O(N__74572),
            .I(N__74569));
    LocalMux I__12833 (
            .O(N__74569),
            .I(shift_srl_50Z0Z_11));
    InMux I__12832 (
            .O(N__74566),
            .I(N__74563));
    LocalMux I__12831 (
            .O(N__74563),
            .I(shift_srl_50Z0Z_12));
    InMux I__12830 (
            .O(N__74560),
            .I(N__74557));
    LocalMux I__12829 (
            .O(N__74557),
            .I(N__74554));
    Odrv4 I__12828 (
            .O(N__74554),
            .I(shift_srl_50Z0Z_13));
    InMux I__12827 (
            .O(N__74551),
            .I(N__74548));
    LocalMux I__12826 (
            .O(N__74548),
            .I(shift_srl_52Z0Z_10));
    InMux I__12825 (
            .O(N__74545),
            .I(N__74542));
    LocalMux I__12824 (
            .O(N__74542),
            .I(shift_srl_52Z0Z_11));
    InMux I__12823 (
            .O(N__74539),
            .I(N__74536));
    LocalMux I__12822 (
            .O(N__74536),
            .I(shift_srl_52Z0Z_12));
    InMux I__12821 (
            .O(N__74533),
            .I(N__74530));
    LocalMux I__12820 (
            .O(N__74530),
            .I(shift_srl_49Z0Z_2));
    InMux I__12819 (
            .O(N__74527),
            .I(N__74524));
    LocalMux I__12818 (
            .O(N__74524),
            .I(shift_srl_49Z0Z_3));
    InMux I__12817 (
            .O(N__74521),
            .I(N__74518));
    LocalMux I__12816 (
            .O(N__74518),
            .I(shift_srl_49Z0Z_4));
    InMux I__12815 (
            .O(N__74515),
            .I(N__74512));
    LocalMux I__12814 (
            .O(N__74512),
            .I(shift_srl_49Z0Z_5));
    InMux I__12813 (
            .O(N__74509),
            .I(N__74506));
    LocalMux I__12812 (
            .O(N__74506),
            .I(shift_srl_49Z0Z_6));
    CascadeMux I__12811 (
            .O(N__74503),
            .I(rco_c_44_cascade_));
    InMux I__12810 (
            .O(N__74500),
            .I(N__74491));
    InMux I__12809 (
            .O(N__74499),
            .I(N__74491));
    InMux I__12808 (
            .O(N__74498),
            .I(N__74484));
    InMux I__12807 (
            .O(N__74497),
            .I(N__74484));
    InMux I__12806 (
            .O(N__74496),
            .I(N__74484));
    LocalMux I__12805 (
            .O(N__74491),
            .I(N__74481));
    LocalMux I__12804 (
            .O(N__74484),
            .I(N__74476));
    Span4Mux_v I__12803 (
            .O(N__74481),
            .I(N__74473));
    CascadeMux I__12802 (
            .O(N__74480),
            .I(N__74470));
    InMux I__12801 (
            .O(N__74479),
            .I(N__74466));
    Span4Mux_v I__12800 (
            .O(N__74476),
            .I(N__74463));
    Span4Mux_v I__12799 (
            .O(N__74473),
            .I(N__74460));
    InMux I__12798 (
            .O(N__74470),
            .I(N__74455));
    InMux I__12797 (
            .O(N__74469),
            .I(N__74455));
    LocalMux I__12796 (
            .O(N__74466),
            .I(N__74452));
    Span4Mux_v I__12795 (
            .O(N__74463),
            .I(N__74447));
    Span4Mux_v I__12794 (
            .O(N__74460),
            .I(N__74447));
    LocalMux I__12793 (
            .O(N__74455),
            .I(N__74444));
    Span4Mux_v I__12792 (
            .O(N__74452),
            .I(N__74441));
    Odrv4 I__12791 (
            .O(N__74447),
            .I(rco_int_0_a2_0_a2_0_0_37));
    Odrv4 I__12790 (
            .O(N__74444),
            .I(rco_int_0_a2_0_a2_0_0_37));
    Odrv4 I__12789 (
            .O(N__74441),
            .I(rco_int_0_a2_0_a2_0_0_37));
    CascadeMux I__12788 (
            .O(N__74434),
            .I(clk_en_0_a3_0_a2_sx_49_cascade_));
    CEMux I__12787 (
            .O(N__74431),
            .I(N__74428));
    LocalMux I__12786 (
            .O(N__74428),
            .I(N__74423));
    CEMux I__12785 (
            .O(N__74427),
            .I(N__74420));
    CEMux I__12784 (
            .O(N__74426),
            .I(N__74417));
    Span4Mux_v I__12783 (
            .O(N__74423),
            .I(N__74412));
    LocalMux I__12782 (
            .O(N__74420),
            .I(N__74412));
    LocalMux I__12781 (
            .O(N__74417),
            .I(N__74409));
    Span4Mux_v I__12780 (
            .O(N__74412),
            .I(N__74403));
    Span4Mux_h I__12779 (
            .O(N__74409),
            .I(N__74403));
    CEMux I__12778 (
            .O(N__74408),
            .I(N__74400));
    Span4Mux_h I__12777 (
            .O(N__74403),
            .I(N__74396));
    LocalMux I__12776 (
            .O(N__74400),
            .I(N__74393));
    InMux I__12775 (
            .O(N__74399),
            .I(N__74390));
    Odrv4 I__12774 (
            .O(N__74396),
            .I(clk_en_49));
    Odrv12 I__12773 (
            .O(N__74393),
            .I(clk_en_49));
    LocalMux I__12772 (
            .O(N__74390),
            .I(clk_en_49));
    InMux I__12771 (
            .O(N__74383),
            .I(N__74378));
    InMux I__12770 (
            .O(N__74382),
            .I(N__74373));
    InMux I__12769 (
            .O(N__74381),
            .I(N__74373));
    LocalMux I__12768 (
            .O(N__74378),
            .I(N__74370));
    LocalMux I__12767 (
            .O(N__74373),
            .I(N__74366));
    Span4Mux_h I__12766 (
            .O(N__74370),
            .I(N__74363));
    InMux I__12765 (
            .O(N__74369),
            .I(N__74360));
    Span4Mux_h I__12764 (
            .O(N__74366),
            .I(N__74357));
    Odrv4 I__12763 (
            .O(N__74363),
            .I(shift_srl_46Z0Z_15));
    LocalMux I__12762 (
            .O(N__74360),
            .I(shift_srl_46Z0Z_15));
    Odrv4 I__12761 (
            .O(N__74357),
            .I(shift_srl_46Z0Z_15));
    InMux I__12760 (
            .O(N__74350),
            .I(N__74347));
    LocalMux I__12759 (
            .O(N__74347),
            .I(shift_srl_192Z0Z_13));
    InMux I__12758 (
            .O(N__74344),
            .I(N__74341));
    LocalMux I__12757 (
            .O(N__74341),
            .I(shift_srl_192Z0Z_12));
    InMux I__12756 (
            .O(N__74338),
            .I(N__74335));
    LocalMux I__12755 (
            .O(N__74335),
            .I(shift_srl_192Z0Z_11));
    InMux I__12754 (
            .O(N__74332),
            .I(N__74329));
    LocalMux I__12753 (
            .O(N__74329),
            .I(shift_srl_192Z0Z_10));
    IoInMux I__12752 (
            .O(N__74326),
            .I(N__74323));
    LocalMux I__12751 (
            .O(N__74323),
            .I(N__74320));
    IoSpan4Mux I__12750 (
            .O(N__74320),
            .I(N__74317));
    Span4Mux_s3_v I__12749 (
            .O(N__74317),
            .I(N__74314));
    Sp12to4 I__12748 (
            .O(N__74314),
            .I(N__74311));
    Odrv12 I__12747 (
            .O(N__74311),
            .I(rco_c_46));
    InMux I__12746 (
            .O(N__74308),
            .I(N__74305));
    LocalMux I__12745 (
            .O(N__74305),
            .I(shift_srl_49Z0Z_0));
    InMux I__12744 (
            .O(N__74302),
            .I(N__74299));
    LocalMux I__12743 (
            .O(N__74299),
            .I(shift_srl_49Z0Z_1));
    InMux I__12742 (
            .O(N__74296),
            .I(N__74293));
    LocalMux I__12741 (
            .O(N__74293),
            .I(shift_srl_192Z0Z_1));
    InMux I__12740 (
            .O(N__74290),
            .I(N__74287));
    LocalMux I__12739 (
            .O(N__74287),
            .I(shift_srl_192Z0Z_2));
    InMux I__12738 (
            .O(N__74284),
            .I(N__74281));
    LocalMux I__12737 (
            .O(N__74281),
            .I(shift_srl_192Z0Z_3));
    InMux I__12736 (
            .O(N__74278),
            .I(N__74275));
    LocalMux I__12735 (
            .O(N__74275),
            .I(shift_srl_192Z0Z_4));
    InMux I__12734 (
            .O(N__74272),
            .I(N__74269));
    LocalMux I__12733 (
            .O(N__74269),
            .I(shift_srl_192Z0Z_5));
    InMux I__12732 (
            .O(N__74266),
            .I(N__74263));
    LocalMux I__12731 (
            .O(N__74263),
            .I(shift_srl_192Z0Z_6));
    InMux I__12730 (
            .O(N__74260),
            .I(N__74255));
    CascadeMux I__12729 (
            .O(N__74259),
            .I(N__74252));
    CascadeMux I__12728 (
            .O(N__74258),
            .I(N__74248));
    LocalMux I__12727 (
            .O(N__74255),
            .I(N__74245));
    InMux I__12726 (
            .O(N__74252),
            .I(N__74242));
    InMux I__12725 (
            .O(N__74251),
            .I(N__74237));
    InMux I__12724 (
            .O(N__74248),
            .I(N__74237));
    Span4Mux_v I__12723 (
            .O(N__74245),
            .I(N__74234));
    LocalMux I__12722 (
            .O(N__74242),
            .I(N__74231));
    LocalMux I__12721 (
            .O(N__74237),
            .I(N__74228));
    Span4Mux_h I__12720 (
            .O(N__74234),
            .I(N__74223));
    Span4Mux_v I__12719 (
            .O(N__74231),
            .I(N__74223));
    Odrv12 I__12718 (
            .O(N__74228),
            .I(N_4177));
    Odrv4 I__12717 (
            .O(N__74223),
            .I(N_4177));
    InMux I__12716 (
            .O(N__74218),
            .I(N__74212));
    InMux I__12715 (
            .O(N__74217),
            .I(N__74209));
    InMux I__12714 (
            .O(N__74216),
            .I(N__74204));
    InMux I__12713 (
            .O(N__74215),
            .I(N__74204));
    LocalMux I__12712 (
            .O(N__74212),
            .I(N__74201));
    LocalMux I__12711 (
            .O(N__74209),
            .I(shift_srl_192Z0Z_15));
    LocalMux I__12710 (
            .O(N__74204),
            .I(shift_srl_192Z0Z_15));
    Odrv12 I__12709 (
            .O(N__74201),
            .I(shift_srl_192Z0Z_15));
    IoInMux I__12708 (
            .O(N__74194),
            .I(N__74191));
    LocalMux I__12707 (
            .O(N__74191),
            .I(N__74188));
    Span12Mux_s4_v I__12706 (
            .O(N__74188),
            .I(N__74185));
    Odrv12 I__12705 (
            .O(N__74185),
            .I(rco_c_192));
    InMux I__12704 (
            .O(N__74182),
            .I(N__74179));
    LocalMux I__12703 (
            .O(N__74179),
            .I(shift_srl_192Z0Z_14));
    InMux I__12702 (
            .O(N__74176),
            .I(N__74173));
    LocalMux I__12701 (
            .O(N__74173),
            .I(shift_srl_175Z0Z_10));
    InMux I__12700 (
            .O(N__74170),
            .I(N__74167));
    LocalMux I__12699 (
            .O(N__74167),
            .I(shift_srl_175Z0Z_11));
    InMux I__12698 (
            .O(N__74164),
            .I(N__74161));
    LocalMux I__12697 (
            .O(N__74161),
            .I(shift_srl_175Z0Z_12));
    InMux I__12696 (
            .O(N__74158),
            .I(N__74155));
    LocalMux I__12695 (
            .O(N__74155),
            .I(shift_srl_175Z0Z_13));
    InMux I__12694 (
            .O(N__74152),
            .I(N__74149));
    LocalMux I__12693 (
            .O(N__74149),
            .I(shift_srl_175Z0Z_14));
    InMux I__12692 (
            .O(N__74146),
            .I(N__74143));
    LocalMux I__12691 (
            .O(N__74143),
            .I(shift_srl_175Z0Z_9));
    InMux I__12690 (
            .O(N__74140),
            .I(N__74137));
    LocalMux I__12689 (
            .O(N__74137),
            .I(N__74134));
    Odrv4 I__12688 (
            .O(N__74134),
            .I(shift_srl_175Z0Z_7));
    InMux I__12687 (
            .O(N__74131),
            .I(N__74128));
    LocalMux I__12686 (
            .O(N__74128),
            .I(shift_srl_175Z0Z_8));
    CEMux I__12685 (
            .O(N__74125),
            .I(N__74121));
    CEMux I__12684 (
            .O(N__74124),
            .I(N__74118));
    LocalMux I__12683 (
            .O(N__74121),
            .I(N__74113));
    LocalMux I__12682 (
            .O(N__74118),
            .I(N__74113));
    Odrv4 I__12681 (
            .O(N__74113),
            .I(clk_en_175));
    InMux I__12680 (
            .O(N__74110),
            .I(N__74107));
    LocalMux I__12679 (
            .O(N__74107),
            .I(shift_srl_192Z0Z_0));
    InMux I__12678 (
            .O(N__74104),
            .I(N__74101));
    LocalMux I__12677 (
            .O(N__74101),
            .I(shift_srl_185Z0Z_10));
    InMux I__12676 (
            .O(N__74098),
            .I(N__74095));
    LocalMux I__12675 (
            .O(N__74095),
            .I(shift_srl_185Z0Z_11));
    InMux I__12674 (
            .O(N__74092),
            .I(N__74089));
    LocalMux I__12673 (
            .O(N__74089),
            .I(shift_srl_185Z0Z_12));
    InMux I__12672 (
            .O(N__74086),
            .I(N__74083));
    LocalMux I__12671 (
            .O(N__74083),
            .I(shift_srl_185Z0Z_13));
    InMux I__12670 (
            .O(N__74080),
            .I(N__74077));
    LocalMux I__12669 (
            .O(N__74077),
            .I(shift_srl_185Z0Z_14));
    InMux I__12668 (
            .O(N__74074),
            .I(N__74071));
    LocalMux I__12667 (
            .O(N__74071),
            .I(shift_srl_185Z0Z_9));
    InMux I__12666 (
            .O(N__74068),
            .I(N__74065));
    LocalMux I__12665 (
            .O(N__74065),
            .I(shift_srl_185Z0Z_7));
    InMux I__12664 (
            .O(N__74062),
            .I(N__74059));
    LocalMux I__12663 (
            .O(N__74059),
            .I(shift_srl_185Z0Z_8));
    CEMux I__12662 (
            .O(N__74056),
            .I(N__74052));
    CEMux I__12661 (
            .O(N__74055),
            .I(N__74049));
    LocalMux I__12660 (
            .O(N__74052),
            .I(clk_en_185));
    LocalMux I__12659 (
            .O(N__74049),
            .I(clk_en_185));
    InMux I__12658 (
            .O(N__74044),
            .I(N__74041));
    LocalMux I__12657 (
            .O(N__74041),
            .I(clk_en_0_a2_0_a2_0_sx_192));
    InMux I__12656 (
            .O(N__74038),
            .I(N__74034));
    InMux I__12655 (
            .O(N__74037),
            .I(N__74031));
    LocalMux I__12654 (
            .O(N__74034),
            .I(shift_srl_195Z0Z_15));
    LocalMux I__12653 (
            .O(N__74031),
            .I(shift_srl_195Z0Z_15));
    InMux I__12652 (
            .O(N__74026),
            .I(N__74023));
    LocalMux I__12651 (
            .O(N__74023),
            .I(shift_srl_195Z0Z_0));
    InMux I__12650 (
            .O(N__74020),
            .I(N__74017));
    LocalMux I__12649 (
            .O(N__74017),
            .I(shift_srl_195Z0Z_1));
    InMux I__12648 (
            .O(N__74014),
            .I(N__74011));
    LocalMux I__12647 (
            .O(N__74011),
            .I(shift_srl_195Z0Z_2));
    InMux I__12646 (
            .O(N__74008),
            .I(N__74005));
    LocalMux I__12645 (
            .O(N__74005),
            .I(shift_srl_195Z0Z_3));
    InMux I__12644 (
            .O(N__74002),
            .I(N__73999));
    LocalMux I__12643 (
            .O(N__73999),
            .I(shift_srl_195Z0Z_4));
    InMux I__12642 (
            .O(N__73996),
            .I(N__73993));
    LocalMux I__12641 (
            .O(N__73993),
            .I(shift_srl_195Z0Z_5));
    InMux I__12640 (
            .O(N__73990),
            .I(N__73987));
    LocalMux I__12639 (
            .O(N__73987),
            .I(shift_srl_195Z0Z_6));
    InMux I__12638 (
            .O(N__73984),
            .I(N__73981));
    LocalMux I__12637 (
            .O(N__73981),
            .I(shift_srl_195Z0Z_7));
    CEMux I__12636 (
            .O(N__73978),
            .I(N__73974));
    CEMux I__12635 (
            .O(N__73977),
            .I(N__73971));
    LocalMux I__12634 (
            .O(N__73974),
            .I(N__73966));
    LocalMux I__12633 (
            .O(N__73971),
            .I(N__73966));
    Span4Mux_v I__12632 (
            .O(N__73966),
            .I(N__73963));
    Odrv4 I__12631 (
            .O(N__73963),
            .I(clk_en_195));
    InMux I__12630 (
            .O(N__73960),
            .I(N__73957));
    LocalMux I__12629 (
            .O(N__73957),
            .I(shift_srl_186Z0Z_5));
    InMux I__12628 (
            .O(N__73954),
            .I(N__73951));
    LocalMux I__12627 (
            .O(N__73951),
            .I(shift_srl_186Z0Z_6));
    InMux I__12626 (
            .O(N__73948),
            .I(N__73945));
    LocalMux I__12625 (
            .O(N__73945),
            .I(N__73942));
    Odrv4 I__12624 (
            .O(N__73942),
            .I(shift_srl_184Z0Z_14));
    CEMux I__12623 (
            .O(N__73939),
            .I(N__73936));
    LocalMux I__12622 (
            .O(N__73936),
            .I(N__73931));
    CEMux I__12621 (
            .O(N__73935),
            .I(N__73928));
    CEMux I__12620 (
            .O(N__73934),
            .I(N__73925));
    Span4Mux_h I__12619 (
            .O(N__73931),
            .I(N__73920));
    LocalMux I__12618 (
            .O(N__73928),
            .I(N__73920));
    LocalMux I__12617 (
            .O(N__73925),
            .I(N__73917));
    Span4Mux_v I__12616 (
            .O(N__73920),
            .I(N__73914));
    Odrv4 I__12615 (
            .O(N__73917),
            .I(clk_en_184));
    Odrv4 I__12614 (
            .O(N__73914),
            .I(clk_en_184));
    CascadeMux I__12613 (
            .O(N__73909),
            .I(clk_en_0_a2_0_a2_0_sx_192_cascade_));
    CascadeMux I__12612 (
            .O(N__73906),
            .I(N_4179_cascade_));
    InMux I__12611 (
            .O(N__73903),
            .I(N__73895));
    InMux I__12610 (
            .O(N__73902),
            .I(N__73895));
    InMux I__12609 (
            .O(N__73901),
            .I(N__73892));
    InMux I__12608 (
            .O(N__73900),
            .I(N__73889));
    LocalMux I__12607 (
            .O(N__73895),
            .I(N__73886));
    LocalMux I__12606 (
            .O(N__73892),
            .I(N__73883));
    LocalMux I__12605 (
            .O(N__73889),
            .I(N__73880));
    Span4Mux_v I__12604 (
            .O(N__73886),
            .I(N__73877));
    Span4Mux_h I__12603 (
            .O(N__73883),
            .I(N__73874));
    Span4Mux_h I__12602 (
            .O(N__73880),
            .I(N__73871));
    Odrv4 I__12601 (
            .O(N__73877),
            .I(shift_srl_194Z0Z_15));
    Odrv4 I__12600 (
            .O(N__73874),
            .I(shift_srl_194Z0Z_15));
    Odrv4 I__12599 (
            .O(N__73871),
            .I(shift_srl_194Z0Z_15));
    InMux I__12598 (
            .O(N__73864),
            .I(N__73858));
    InMux I__12597 (
            .O(N__73863),
            .I(N__73858));
    LocalMux I__12596 (
            .O(N__73858),
            .I(N__73854));
    InMux I__12595 (
            .O(N__73857),
            .I(N__73851));
    Span4Mux_v I__12594 (
            .O(N__73854),
            .I(N__73846));
    LocalMux I__12593 (
            .O(N__73851),
            .I(N__73846));
    Span4Mux_h I__12592 (
            .O(N__73846),
            .I(N__73842));
    InMux I__12591 (
            .O(N__73845),
            .I(N__73839));
    Odrv4 I__12590 (
            .O(N__73842),
            .I(N_4179));
    LocalMux I__12589 (
            .O(N__73839),
            .I(N_4179));
    InMux I__12588 (
            .O(N__73834),
            .I(N__73829));
    InMux I__12587 (
            .O(N__73833),
            .I(N__73823));
    InMux I__12586 (
            .O(N__73832),
            .I(N__73823));
    LocalMux I__12585 (
            .O(N__73829),
            .I(N__73819));
    InMux I__12584 (
            .O(N__73828),
            .I(N__73816));
    LocalMux I__12583 (
            .O(N__73823),
            .I(N__73813));
    InMux I__12582 (
            .O(N__73822),
            .I(N__73810));
    Span4Mux_v I__12581 (
            .O(N__73819),
            .I(N__73805));
    LocalMux I__12580 (
            .O(N__73816),
            .I(N__73805));
    Span4Mux_v I__12579 (
            .O(N__73813),
            .I(N__73800));
    LocalMux I__12578 (
            .O(N__73810),
            .I(N__73800));
    Span4Mux_h I__12577 (
            .O(N__73805),
            .I(N__73797));
    Span4Mux_v I__12576 (
            .O(N__73800),
            .I(N__73792));
    Span4Mux_h I__12575 (
            .O(N__73797),
            .I(N__73792));
    Odrv4 I__12574 (
            .O(N__73792),
            .I(N_4181));
    InMux I__12573 (
            .O(N__73789),
            .I(N__73786));
    LocalMux I__12572 (
            .O(N__73786),
            .I(shift_srl_184Z0Z_13));
    InMux I__12571 (
            .O(N__73783),
            .I(N__73780));
    LocalMux I__12570 (
            .O(N__73780),
            .I(shift_srl_184Z0Z_9));
    InMux I__12569 (
            .O(N__73777),
            .I(N__73774));
    LocalMux I__12568 (
            .O(N__73774),
            .I(shift_srl_184Z0Z_7));
    InMux I__12567 (
            .O(N__73771),
            .I(N__73768));
    LocalMux I__12566 (
            .O(N__73768),
            .I(shift_srl_184Z0Z_8));
    InMux I__12565 (
            .O(N__73765),
            .I(N__73762));
    LocalMux I__12564 (
            .O(N__73762),
            .I(shift_srl_186Z0Z_0));
    InMux I__12563 (
            .O(N__73759),
            .I(N__73756));
    LocalMux I__12562 (
            .O(N__73756),
            .I(shift_srl_186Z0Z_1));
    InMux I__12561 (
            .O(N__73753),
            .I(N__73750));
    LocalMux I__12560 (
            .O(N__73750),
            .I(shift_srl_186Z0Z_2));
    InMux I__12559 (
            .O(N__73747),
            .I(N__73744));
    LocalMux I__12558 (
            .O(N__73744),
            .I(shift_srl_186Z0Z_3));
    InMux I__12557 (
            .O(N__73741),
            .I(N__73738));
    LocalMux I__12556 (
            .O(N__73738),
            .I(shift_srl_186Z0Z_4));
    InMux I__12555 (
            .O(N__73735),
            .I(N__73732));
    LocalMux I__12554 (
            .O(N__73732),
            .I(shift_srl_166Z0Z_12));
    InMux I__12553 (
            .O(N__73729),
            .I(N__73726));
    LocalMux I__12552 (
            .O(N__73726),
            .I(shift_srl_166Z0Z_13));
    InMux I__12551 (
            .O(N__73723),
            .I(N__73720));
    LocalMux I__12550 (
            .O(N__73720),
            .I(shift_srl_166Z0Z_14));
    InMux I__12549 (
            .O(N__73717),
            .I(N__73714));
    LocalMux I__12548 (
            .O(N__73714),
            .I(shift_srl_166Z0Z_8));
    InMux I__12547 (
            .O(N__73711),
            .I(N__73708));
    LocalMux I__12546 (
            .O(N__73708),
            .I(shift_srl_166Z0Z_9));
    InMux I__12545 (
            .O(N__73705),
            .I(N__73702));
    LocalMux I__12544 (
            .O(N__73702),
            .I(shift_srl_166Z0Z_0));
    CEMux I__12543 (
            .O(N__73699),
            .I(N__73695));
    CEMux I__12542 (
            .O(N__73698),
            .I(N__73692));
    LocalMux I__12541 (
            .O(N__73695),
            .I(clk_en_166));
    LocalMux I__12540 (
            .O(N__73692),
            .I(clk_en_166));
    InMux I__12539 (
            .O(N__73687),
            .I(N__73684));
    LocalMux I__12538 (
            .O(N__73684),
            .I(shift_srl_184Z0Z_10));
    InMux I__12537 (
            .O(N__73681),
            .I(N__73678));
    LocalMux I__12536 (
            .O(N__73678),
            .I(shift_srl_184Z0Z_11));
    InMux I__12535 (
            .O(N__73675),
            .I(N__73672));
    LocalMux I__12534 (
            .O(N__73672),
            .I(shift_srl_184Z0Z_12));
    InMux I__12533 (
            .O(N__73669),
            .I(N__73666));
    LocalMux I__12532 (
            .O(N__73666),
            .I(shift_srl_166Z0Z_1));
    InMux I__12531 (
            .O(N__73663),
            .I(N__73660));
    LocalMux I__12530 (
            .O(N__73660),
            .I(shift_srl_166Z0Z_2));
    InMux I__12529 (
            .O(N__73657),
            .I(N__73654));
    LocalMux I__12528 (
            .O(N__73654),
            .I(shift_srl_166Z0Z_3));
    InMux I__12527 (
            .O(N__73651),
            .I(N__73648));
    LocalMux I__12526 (
            .O(N__73648),
            .I(shift_srl_166Z0Z_4));
    InMux I__12525 (
            .O(N__73645),
            .I(N__73642));
    LocalMux I__12524 (
            .O(N__73642),
            .I(shift_srl_166Z0Z_5));
    InMux I__12523 (
            .O(N__73639),
            .I(N__73636));
    LocalMux I__12522 (
            .O(N__73636),
            .I(shift_srl_166Z0Z_6));
    InMux I__12521 (
            .O(N__73633),
            .I(N__73630));
    LocalMux I__12520 (
            .O(N__73630),
            .I(shift_srl_166Z0Z_7));
    InMux I__12519 (
            .O(N__73627),
            .I(N__73624));
    LocalMux I__12518 (
            .O(N__73624),
            .I(shift_srl_166Z0Z_10));
    InMux I__12517 (
            .O(N__73621),
            .I(N__73618));
    LocalMux I__12516 (
            .O(N__73618),
            .I(shift_srl_166Z0Z_11));
    InMux I__12515 (
            .O(N__73615),
            .I(N__73612));
    LocalMux I__12514 (
            .O(N__73612),
            .I(shift_srl_174Z0Z_10));
    InMux I__12513 (
            .O(N__73609),
            .I(N__73606));
    LocalMux I__12512 (
            .O(N__73606),
            .I(shift_srl_174Z0Z_11));
    InMux I__12511 (
            .O(N__73603),
            .I(N__73600));
    LocalMux I__12510 (
            .O(N__73600),
            .I(shift_srl_174Z0Z_12));
    InMux I__12509 (
            .O(N__73597),
            .I(N__73594));
    LocalMux I__12508 (
            .O(N__73594),
            .I(shift_srl_174Z0Z_13));
    InMux I__12507 (
            .O(N__73591),
            .I(N__73588));
    LocalMux I__12506 (
            .O(N__73588),
            .I(shift_srl_174Z0Z_14));
    InMux I__12505 (
            .O(N__73585),
            .I(N__73582));
    LocalMux I__12504 (
            .O(N__73582),
            .I(shift_srl_174Z0Z_9));
    InMux I__12503 (
            .O(N__73579),
            .I(N__73576));
    LocalMux I__12502 (
            .O(N__73576),
            .I(shift_srl_174Z0Z_7));
    InMux I__12501 (
            .O(N__73573),
            .I(N__73570));
    LocalMux I__12500 (
            .O(N__73570),
            .I(shift_srl_174Z0Z_8));
    CEMux I__12499 (
            .O(N__73567),
            .I(N__73564));
    LocalMux I__12498 (
            .O(N__73564),
            .I(N__73560));
    CEMux I__12497 (
            .O(N__73563),
            .I(N__73557));
    Span4Mux_v I__12496 (
            .O(N__73560),
            .I(N__73554));
    LocalMux I__12495 (
            .O(N__73557),
            .I(N__73551));
    Odrv4 I__12494 (
            .O(N__73554),
            .I(clk_en_174));
    Odrv12 I__12493 (
            .O(N__73551),
            .I(clk_en_174));
    InMux I__12492 (
            .O(N__73546),
            .I(N__73543));
    LocalMux I__12491 (
            .O(N__73543),
            .I(shift_srl_62Z0Z_10));
    InMux I__12490 (
            .O(N__73540),
            .I(N__73537));
    LocalMux I__12489 (
            .O(N__73537),
            .I(shift_srl_62Z0Z_11));
    InMux I__12488 (
            .O(N__73534),
            .I(N__73531));
    LocalMux I__12487 (
            .O(N__73531),
            .I(shift_srl_62Z0Z_12));
    InMux I__12486 (
            .O(N__73528),
            .I(N__73525));
    LocalMux I__12485 (
            .O(N__73525),
            .I(shift_srl_62Z0Z_13));
    InMux I__12484 (
            .O(N__73522),
            .I(N__73519));
    LocalMux I__12483 (
            .O(N__73519),
            .I(shift_srl_62Z0Z_14));
    InMux I__12482 (
            .O(N__73516),
            .I(N__73512));
    InMux I__12481 (
            .O(N__73515),
            .I(N__73509));
    LocalMux I__12480 (
            .O(N__73512),
            .I(shift_srl_62Z0Z_15));
    LocalMux I__12479 (
            .O(N__73509),
            .I(shift_srl_62Z0Z_15));
    InMux I__12478 (
            .O(N__73504),
            .I(N__73501));
    LocalMux I__12477 (
            .O(N__73501),
            .I(shift_srl_62Z0Z_9));
    InMux I__12476 (
            .O(N__73498),
            .I(N__73495));
    LocalMux I__12475 (
            .O(N__73495),
            .I(shift_srl_62Z0Z_7));
    InMux I__12474 (
            .O(N__73492),
            .I(N__73489));
    LocalMux I__12473 (
            .O(N__73489),
            .I(shift_srl_62Z0Z_8));
    CEMux I__12472 (
            .O(N__73486),
            .I(N__73482));
    CEMux I__12471 (
            .O(N__73485),
            .I(N__73479));
    LocalMux I__12470 (
            .O(N__73482),
            .I(clk_en_62));
    LocalMux I__12469 (
            .O(N__73479),
            .I(clk_en_62));
    InMux I__12468 (
            .O(N__73474),
            .I(N__73471));
    LocalMux I__12467 (
            .O(N__73471),
            .I(shift_srl_61Z0Z_13));
    InMux I__12466 (
            .O(N__73468),
            .I(N__73465));
    LocalMux I__12465 (
            .O(N__73465),
            .I(shift_srl_61Z0Z_14));
    InMux I__12464 (
            .O(N__73462),
            .I(N__73459));
    LocalMux I__12463 (
            .O(N__73459),
            .I(shift_srl_61Z0Z_10));
    InMux I__12462 (
            .O(N__73456),
            .I(N__73453));
    LocalMux I__12461 (
            .O(N__73453),
            .I(shift_srl_61Z0Z_11));
    InMux I__12460 (
            .O(N__73450),
            .I(N__73447));
    LocalMux I__12459 (
            .O(N__73447),
            .I(shift_srl_61Z0Z_8));
    InMux I__12458 (
            .O(N__73444),
            .I(N__73441));
    LocalMux I__12457 (
            .O(N__73441),
            .I(shift_srl_61Z0Z_9));
    CascadeMux I__12456 (
            .O(N__73438),
            .I(shift_srl_61_RNI3LM9Z0Z_15_cascade_));
    InMux I__12455 (
            .O(N__73435),
            .I(N__73430));
    InMux I__12454 (
            .O(N__73434),
            .I(N__73425));
    InMux I__12453 (
            .O(N__73433),
            .I(N__73425));
    LocalMux I__12452 (
            .O(N__73430),
            .I(shift_srl_61Z0Z_15));
    LocalMux I__12451 (
            .O(N__73425),
            .I(shift_srl_61Z0Z_15));
    CascadeMux I__12450 (
            .O(N__73420),
            .I(shift_srl_62_RNIM5RKZ0Z_15_cascade_));
    CEMux I__12449 (
            .O(N__73417),
            .I(N__73413));
    CEMux I__12448 (
            .O(N__73416),
            .I(N__73410));
    LocalMux I__12447 (
            .O(N__73413),
            .I(N__73405));
    LocalMux I__12446 (
            .O(N__73410),
            .I(N__73405));
    Sp12to4 I__12445 (
            .O(N__73405),
            .I(N__73402));
    Odrv12 I__12444 (
            .O(N__73402),
            .I(clk_en_61));
    InMux I__12443 (
            .O(N__73399),
            .I(N__73396));
    LocalMux I__12442 (
            .O(N__73396),
            .I(shift_srl_48Z0Z_13));
    InMux I__12441 (
            .O(N__73393),
            .I(N__73390));
    LocalMux I__12440 (
            .O(N__73390),
            .I(shift_srl_48Z0Z_11));
    InMux I__12439 (
            .O(N__73387),
            .I(N__73384));
    LocalMux I__12438 (
            .O(N__73384),
            .I(shift_srl_48Z0Z_12));
    CEMux I__12437 (
            .O(N__73381),
            .I(N__73376));
    CEMux I__12436 (
            .O(N__73380),
            .I(N__73373));
    CEMux I__12435 (
            .O(N__73379),
            .I(N__73370));
    LocalMux I__12434 (
            .O(N__73376),
            .I(N__73367));
    LocalMux I__12433 (
            .O(N__73373),
            .I(N__73362));
    LocalMux I__12432 (
            .O(N__73370),
            .I(N__73362));
    Span4Mux_h I__12431 (
            .O(N__73367),
            .I(N__73359));
    Span4Mux_h I__12430 (
            .O(N__73362),
            .I(N__73356));
    Odrv4 I__12429 (
            .O(N__73359),
            .I(clk_en_48));
    Odrv4 I__12428 (
            .O(N__73356),
            .I(clk_en_48));
    InMux I__12427 (
            .O(N__73351),
            .I(N__73348));
    LocalMux I__12426 (
            .O(N__73348),
            .I(N__73345));
    Odrv4 I__12425 (
            .O(N__73345),
            .I(shift_srl_55Z0Z_10));
    InMux I__12424 (
            .O(N__73342),
            .I(N__73339));
    LocalMux I__12423 (
            .O(N__73339),
            .I(shift_srl_55Z0Z_9));
    InMux I__12422 (
            .O(N__73336),
            .I(N__73333));
    LocalMux I__12421 (
            .O(N__73333),
            .I(N__73330));
    Odrv4 I__12420 (
            .O(N__73330),
            .I(shift_srl_55Z0Z_7));
    InMux I__12419 (
            .O(N__73327),
            .I(N__73324));
    LocalMux I__12418 (
            .O(N__73324),
            .I(shift_srl_55Z0Z_8));
    InMux I__12417 (
            .O(N__73321),
            .I(N__73318));
    LocalMux I__12416 (
            .O(N__73318),
            .I(shift_srl_61Z0Z_0));
    InMux I__12415 (
            .O(N__73315),
            .I(N__73312));
    LocalMux I__12414 (
            .O(N__73312),
            .I(shift_srl_61Z0Z_12));
    InMux I__12413 (
            .O(N__73309),
            .I(N__73306));
    LocalMux I__12412 (
            .O(N__73306),
            .I(shift_srl_55Z0Z_4));
    InMux I__12411 (
            .O(N__73303),
            .I(N__73300));
    LocalMux I__12410 (
            .O(N__73300),
            .I(shift_srl_55Z0Z_5));
    InMux I__12409 (
            .O(N__73297),
            .I(N__73294));
    LocalMux I__12408 (
            .O(N__73294),
            .I(shift_srl_55Z0Z_6));
    InMux I__12407 (
            .O(N__73291),
            .I(N__73287));
    InMux I__12406 (
            .O(N__73290),
            .I(N__73284));
    LocalMux I__12405 (
            .O(N__73287),
            .I(shift_srl_44Z0Z_15));
    LocalMux I__12404 (
            .O(N__73284),
            .I(shift_srl_44Z0Z_15));
    InMux I__12403 (
            .O(N__73279),
            .I(N__73275));
    InMux I__12402 (
            .O(N__73278),
            .I(N__73272));
    LocalMux I__12401 (
            .O(N__73275),
            .I(N__73268));
    LocalMux I__12400 (
            .O(N__73272),
            .I(N__73265));
    InMux I__12399 (
            .O(N__73271),
            .I(N__73262));
    Span4Mux_v I__12398 (
            .O(N__73268),
            .I(N__73256));
    Span4Mux_h I__12397 (
            .O(N__73265),
            .I(N__73256));
    LocalMux I__12396 (
            .O(N__73262),
            .I(N__73253));
    InMux I__12395 (
            .O(N__73261),
            .I(N__73250));
    Span4Mux_h I__12394 (
            .O(N__73256),
            .I(N__73247));
    Odrv4 I__12393 (
            .O(N__73253),
            .I(shift_srl_43Z0Z_15));
    LocalMux I__12392 (
            .O(N__73250),
            .I(shift_srl_43Z0Z_15));
    Odrv4 I__12391 (
            .O(N__73247),
            .I(shift_srl_43Z0Z_15));
    InMux I__12390 (
            .O(N__73240),
            .I(N__73233));
    InMux I__12389 (
            .O(N__73239),
            .I(N__73233));
    InMux I__12388 (
            .O(N__73238),
            .I(N__73227));
    LocalMux I__12387 (
            .O(N__73233),
            .I(N__73224));
    InMux I__12386 (
            .O(N__73232),
            .I(N__73217));
    InMux I__12385 (
            .O(N__73231),
            .I(N__73217));
    InMux I__12384 (
            .O(N__73230),
            .I(N__73217));
    LocalMux I__12383 (
            .O(N__73227),
            .I(N__73214));
    Span4Mux_v I__12382 (
            .O(N__73224),
            .I(N__73211));
    LocalMux I__12381 (
            .O(N__73217),
            .I(N__73206));
    Span4Mux_h I__12380 (
            .O(N__73214),
            .I(N__73206));
    Odrv4 I__12379 (
            .O(N__73211),
            .I(shift_srl_42Z0Z_15));
    Odrv4 I__12378 (
            .O(N__73206),
            .I(shift_srl_42Z0Z_15));
    CascadeMux I__12377 (
            .O(N__73201),
            .I(rco_int_0_a2_1_a2_0_44_cascade_));
    InMux I__12376 (
            .O(N__73198),
            .I(N__73195));
    LocalMux I__12375 (
            .O(N__73195),
            .I(shift_srl_48Z0Z_14));
    InMux I__12374 (
            .O(N__73192),
            .I(N__73189));
    LocalMux I__12373 (
            .O(N__73189),
            .I(shift_srl_55Z0Z_14));
    InMux I__12372 (
            .O(N__73186),
            .I(N__73183));
    LocalMux I__12371 (
            .O(N__73183),
            .I(shift_srl_55Z0Z_13));
    InMux I__12370 (
            .O(N__73180),
            .I(N__73177));
    LocalMux I__12369 (
            .O(N__73177),
            .I(shift_srl_55Z0Z_12));
    InMux I__12368 (
            .O(N__73174),
            .I(N__73171));
    LocalMux I__12367 (
            .O(N__73171),
            .I(shift_srl_55Z0Z_11));
    InMux I__12366 (
            .O(N__73168),
            .I(N__73165));
    LocalMux I__12365 (
            .O(N__73165),
            .I(shift_srl_55Z0Z_0));
    InMux I__12364 (
            .O(N__73162),
            .I(N__73159));
    LocalMux I__12363 (
            .O(N__73159),
            .I(shift_srl_55Z0Z_1));
    InMux I__12362 (
            .O(N__73156),
            .I(N__73153));
    LocalMux I__12361 (
            .O(N__73153),
            .I(shift_srl_55Z0Z_2));
    InMux I__12360 (
            .O(N__73150),
            .I(N__73147));
    LocalMux I__12359 (
            .O(N__73147),
            .I(shift_srl_55Z0Z_3));
    InMux I__12358 (
            .O(N__73144),
            .I(N__73141));
    LocalMux I__12357 (
            .O(N__73141),
            .I(shift_srl_56Z0Z_11));
    InMux I__12356 (
            .O(N__73138),
            .I(N__73135));
    LocalMux I__12355 (
            .O(N__73135),
            .I(shift_srl_56Z0Z_12));
    InMux I__12354 (
            .O(N__73132),
            .I(N__73129));
    LocalMux I__12353 (
            .O(N__73129),
            .I(shift_srl_56Z0Z_13));
    InMux I__12352 (
            .O(N__73126),
            .I(N__73123));
    LocalMux I__12351 (
            .O(N__73123),
            .I(shift_srl_56Z0Z_14));
    InMux I__12350 (
            .O(N__73120),
            .I(N__73117));
    LocalMux I__12349 (
            .O(N__73117),
            .I(shift_srl_56Z0Z_9));
    CascadeMux I__12348 (
            .O(N__73114),
            .I(shift_srl_58_RNIQMNUZ0Z_15_cascade_));
    CascadeMux I__12347 (
            .O(N__73111),
            .I(shift_srl_54_RNIEAU71Z0Z_15_cascade_));
    CEMux I__12346 (
            .O(N__73108),
            .I(N__73105));
    LocalMux I__12345 (
            .O(N__73105),
            .I(N__73102));
    Span4Mux_h I__12344 (
            .O(N__73102),
            .I(N__73098));
    CEMux I__12343 (
            .O(N__73101),
            .I(N__73095));
    Span4Mux_h I__12342 (
            .O(N__73098),
            .I(N__73090));
    LocalMux I__12341 (
            .O(N__73095),
            .I(N__73090));
    Span4Mux_h I__12340 (
            .O(N__73090),
            .I(N__73086));
    CEMux I__12339 (
            .O(N__73089),
            .I(N__73083));
    Odrv4 I__12338 (
            .O(N__73086),
            .I(clk_en_59));
    LocalMux I__12337 (
            .O(N__73083),
            .I(clk_en_59));
    CascadeMux I__12336 (
            .O(N__73078),
            .I(rco_int_0_a2_0_a2_0_39_cascade_));
    CascadeMux I__12335 (
            .O(N__73075),
            .I(rco_int_0_a2_0_a2_83_m6_0_a2_3_sx_cascade_));
    CascadeMux I__12334 (
            .O(N__73072),
            .I(N__73069));
    InMux I__12333 (
            .O(N__73069),
            .I(N__73065));
    InMux I__12332 (
            .O(N__73068),
            .I(N__73062));
    LocalMux I__12331 (
            .O(N__73065),
            .I(N__73059));
    LocalMux I__12330 (
            .O(N__73062),
            .I(N__73056));
    Span4Mux_v I__12329 (
            .O(N__73059),
            .I(N__73053));
    Span4Mux_h I__12328 (
            .O(N__73056),
            .I(N__73050));
    Span4Mux_h I__12327 (
            .O(N__73053),
            .I(N__73045));
    Span4Mux_h I__12326 (
            .O(N__73050),
            .I(N__73045));
    Odrv4 I__12325 (
            .O(N__73045),
            .I(rco_int_0_a2_0_a2_83_m6_0_a2_3));
    InMux I__12324 (
            .O(N__73042),
            .I(N__73038));
    InMux I__12323 (
            .O(N__73041),
            .I(N__73035));
    LocalMux I__12322 (
            .O(N__73038),
            .I(shift_srl_53Z0Z_15));
    LocalMux I__12321 (
            .O(N__73035),
            .I(shift_srl_53Z0Z_15));
    CascadeMux I__12320 (
            .O(N__73030),
            .I(shift_srl_53_RNI66TQZ0Z_15_cascade_));
    InMux I__12319 (
            .O(N__73027),
            .I(N__73024));
    LocalMux I__12318 (
            .O(N__73024),
            .I(shift_srl_56Z0Z_10));
    InMux I__12317 (
            .O(N__73021),
            .I(N__73018));
    LocalMux I__12316 (
            .O(N__73018),
            .I(shift_srl_51Z0Z_8));
    InMux I__12315 (
            .O(N__73015),
            .I(N__73012));
    LocalMux I__12314 (
            .O(N__73012),
            .I(shift_srl_51Z0Z_9));
    CEMux I__12313 (
            .O(N__73009),
            .I(N__73005));
    CEMux I__12312 (
            .O(N__73008),
            .I(N__73002));
    LocalMux I__12311 (
            .O(N__73005),
            .I(N__72999));
    LocalMux I__12310 (
            .O(N__73002),
            .I(N__72996));
    Span4Mux_v I__12309 (
            .O(N__72999),
            .I(N__72993));
    Span4Mux_v I__12308 (
            .O(N__72996),
            .I(N__72990));
    Odrv4 I__12307 (
            .O(N__72993),
            .I(clk_en_53));
    Odrv4 I__12306 (
            .O(N__72990),
            .I(clk_en_53));
    CascadeMux I__12305 (
            .O(N__72985),
            .I(shift_srl_50_RNI869CZ0Z_15_cascade_));
    CEMux I__12304 (
            .O(N__72982),
            .I(N__72978));
    CEMux I__12303 (
            .O(N__72981),
            .I(N__72975));
    LocalMux I__12302 (
            .O(N__72978),
            .I(clk_en_51));
    LocalMux I__12301 (
            .O(N__72975),
            .I(clk_en_51));
    InMux I__12300 (
            .O(N__72970),
            .I(N__72967));
    LocalMux I__12299 (
            .O(N__72967),
            .I(shift_srl_49Z0Z_14));
    InMux I__12298 (
            .O(N__72964),
            .I(N__72961));
    LocalMux I__12297 (
            .O(N__72961),
            .I(shift_srl_49Z0Z_13));
    InMux I__12296 (
            .O(N__72958),
            .I(N__72955));
    LocalMux I__12295 (
            .O(N__72955),
            .I(shift_srl_49Z0Z_12));
    InMux I__12294 (
            .O(N__72952),
            .I(N__72949));
    LocalMux I__12293 (
            .O(N__72949),
            .I(N__72946));
    Odrv12 I__12292 (
            .O(N__72946),
            .I(shift_srl_49Z0Z_10));
    InMux I__12291 (
            .O(N__72943),
            .I(N__72940));
    LocalMux I__12290 (
            .O(N__72940),
            .I(shift_srl_49Z0Z_11));
    InMux I__12289 (
            .O(N__72937),
            .I(N__72934));
    LocalMux I__12288 (
            .O(N__72934),
            .I(shift_srl_49Z0Z_8));
    InMux I__12287 (
            .O(N__72931),
            .I(N__72928));
    LocalMux I__12286 (
            .O(N__72928),
            .I(shift_srl_49Z0Z_7));
    InMux I__12285 (
            .O(N__72925),
            .I(N__72922));
    LocalMux I__12284 (
            .O(N__72922),
            .I(shift_srl_51Z0Z_0));
    InMux I__12283 (
            .O(N__72919),
            .I(N__72916));
    LocalMux I__12282 (
            .O(N__72916),
            .I(shift_srl_51Z0Z_1));
    InMux I__12281 (
            .O(N__72913),
            .I(N__72910));
    LocalMux I__12280 (
            .O(N__72910),
            .I(shift_srl_51Z0Z_2));
    InMux I__12279 (
            .O(N__72907),
            .I(N__72904));
    LocalMux I__12278 (
            .O(N__72904),
            .I(shift_srl_51Z0Z_3));
    InMux I__12277 (
            .O(N__72901),
            .I(N__72898));
    LocalMux I__12276 (
            .O(N__72898),
            .I(shift_srl_51Z0Z_4));
    InMux I__12275 (
            .O(N__72895),
            .I(N__72892));
    LocalMux I__12274 (
            .O(N__72892),
            .I(shift_srl_51Z0Z_5));
    InMux I__12273 (
            .O(N__72889),
            .I(N__72886));
    LocalMux I__12272 (
            .O(N__72886),
            .I(shift_srl_51Z0Z_7));
    CascadeMux I__12271 (
            .O(N__72883),
            .I(N__72878));
    InMux I__12270 (
            .O(N__72882),
            .I(N__72874));
    InMux I__12269 (
            .O(N__72881),
            .I(N__72868));
    InMux I__12268 (
            .O(N__72878),
            .I(N__72868));
    CascadeMux I__12267 (
            .O(N__72877),
            .I(N__72865));
    LocalMux I__12266 (
            .O(N__72874),
            .I(N__72862));
    InMux I__12265 (
            .O(N__72873),
            .I(N__72859));
    LocalMux I__12264 (
            .O(N__72868),
            .I(N__72856));
    InMux I__12263 (
            .O(N__72865),
            .I(N__72853));
    Span4Mux_v I__12262 (
            .O(N__72862),
            .I(N__72846));
    LocalMux I__12261 (
            .O(N__72859),
            .I(N__72846));
    Span4Mux_v I__12260 (
            .O(N__72856),
            .I(N__72846));
    LocalMux I__12259 (
            .O(N__72853),
            .I(shift_srl_95_RNIHJ49Z0Z_15));
    Odrv4 I__12258 (
            .O(N__72846),
            .I(shift_srl_95_RNIHJ49Z0Z_15));
    IoInMux I__12257 (
            .O(N__72841),
            .I(N__72838));
    LocalMux I__12256 (
            .O(N__72838),
            .I(N__72835));
    IoSpan4Mux I__12255 (
            .O(N__72835),
            .I(N__72832));
    Span4Mux_s3_v I__12254 (
            .O(N__72832),
            .I(N__72829));
    Span4Mux_v I__12253 (
            .O(N__72829),
            .I(N__72826));
    Odrv4 I__12252 (
            .O(N__72826),
            .I(rco_c_95));
    InMux I__12251 (
            .O(N__72823),
            .I(N__72820));
    LocalMux I__12250 (
            .O(N__72820),
            .I(N__72816));
    InMux I__12249 (
            .O(N__72819),
            .I(N__72813));
    Span4Mux_h I__12248 (
            .O(N__72816),
            .I(N__72810));
    LocalMux I__12247 (
            .O(N__72813),
            .I(N__72807));
    Sp12to4 I__12246 (
            .O(N__72810),
            .I(N__72804));
    Span4Mux_v I__12245 (
            .O(N__72807),
            .I(N__72801));
    Odrv12 I__12244 (
            .O(N__72804),
            .I(shift_srl_94_RNI2F961Z0Z_15));
    Odrv4 I__12243 (
            .O(N__72801),
            .I(shift_srl_94_RNI2F961Z0Z_15));
    IoInMux I__12242 (
            .O(N__72796),
            .I(N__72793));
    LocalMux I__12241 (
            .O(N__72793),
            .I(N__72790));
    IoSpan4Mux I__12240 (
            .O(N__72790),
            .I(N__72784));
    InMux I__12239 (
            .O(N__72789),
            .I(N__72777));
    InMux I__12238 (
            .O(N__72788),
            .I(N__72777));
    InMux I__12237 (
            .O(N__72787),
            .I(N__72777));
    IoSpan4Mux I__12236 (
            .O(N__72784),
            .I(N__72773));
    LocalMux I__12235 (
            .O(N__72777),
            .I(N__72770));
    CascadeMux I__12234 (
            .O(N__72776),
            .I(N__72767));
    Span4Mux_s3_v I__12233 (
            .O(N__72773),
            .I(N__72758));
    Span4Mux_h I__12232 (
            .O(N__72770),
            .I(N__72758));
    InMux I__12231 (
            .O(N__72767),
            .I(N__72755));
    InMux I__12230 (
            .O(N__72766),
            .I(N__72750));
    InMux I__12229 (
            .O(N__72765),
            .I(N__72750));
    InMux I__12228 (
            .O(N__72764),
            .I(N__72745));
    InMux I__12227 (
            .O(N__72763),
            .I(N__72745));
    Odrv4 I__12226 (
            .O(N__72758),
            .I(rco_c_93));
    LocalMux I__12225 (
            .O(N__72755),
            .I(rco_c_93));
    LocalMux I__12224 (
            .O(N__72750),
            .I(rco_c_93));
    LocalMux I__12223 (
            .O(N__72745),
            .I(rco_c_93));
    IoInMux I__12222 (
            .O(N__72736),
            .I(N__72733));
    LocalMux I__12221 (
            .O(N__72733),
            .I(N__72730));
    Span12Mux_s3_v I__12220 (
            .O(N__72730),
            .I(N__72727));
    Odrv12 I__12219 (
            .O(N__72727),
            .I(rco_c_98));
    InMux I__12218 (
            .O(N__72724),
            .I(N__72718));
    InMux I__12217 (
            .O(N__72723),
            .I(N__72718));
    LocalMux I__12216 (
            .O(N__72718),
            .I(N__72714));
    InMux I__12215 (
            .O(N__72717),
            .I(N__72709));
    Span4Mux_h I__12214 (
            .O(N__72714),
            .I(N__72706));
    InMux I__12213 (
            .O(N__72713),
            .I(N__72703));
    InMux I__12212 (
            .O(N__72712),
            .I(N__72700));
    LocalMux I__12211 (
            .O(N__72709),
            .I(N__72697));
    Odrv4 I__12210 (
            .O(N__72706),
            .I(shift_srl_94Z0Z_15));
    LocalMux I__12209 (
            .O(N__72703),
            .I(shift_srl_94Z0Z_15));
    LocalMux I__12208 (
            .O(N__72700),
            .I(shift_srl_94Z0Z_15));
    Odrv12 I__12207 (
            .O(N__72697),
            .I(shift_srl_94Z0Z_15));
    InMux I__12206 (
            .O(N__72688),
            .I(N__72685));
    LocalMux I__12205 (
            .O(N__72685),
            .I(shift_srl_94Z0Z_0));
    InMux I__12204 (
            .O(N__72682),
            .I(N__72679));
    LocalMux I__12203 (
            .O(N__72679),
            .I(shift_srl_94Z0Z_1));
    InMux I__12202 (
            .O(N__72676),
            .I(N__72673));
    LocalMux I__12201 (
            .O(N__72673),
            .I(shift_srl_94Z0Z_2));
    InMux I__12200 (
            .O(N__72670),
            .I(N__72667));
    LocalMux I__12199 (
            .O(N__72667),
            .I(shift_srl_94Z0Z_3));
    InMux I__12198 (
            .O(N__72664),
            .I(N__72661));
    LocalMux I__12197 (
            .O(N__72661),
            .I(N__72658));
    Odrv4 I__12196 (
            .O(N__72658),
            .I(shift_srl_94Z0Z_4));
    CEMux I__12195 (
            .O(N__72655),
            .I(N__72651));
    CEMux I__12194 (
            .O(N__72654),
            .I(N__72647));
    LocalMux I__12193 (
            .O(N__72651),
            .I(N__72643));
    CEMux I__12192 (
            .O(N__72650),
            .I(N__72640));
    LocalMux I__12191 (
            .O(N__72647),
            .I(N__72637));
    CEMux I__12190 (
            .O(N__72646),
            .I(N__72634));
    Span4Mux_h I__12189 (
            .O(N__72643),
            .I(N__72631));
    LocalMux I__12188 (
            .O(N__72640),
            .I(N__72628));
    Span4Mux_v I__12187 (
            .O(N__72637),
            .I(N__72623));
    LocalMux I__12186 (
            .O(N__72634),
            .I(N__72623));
    Span4Mux_v I__12185 (
            .O(N__72631),
            .I(N__72620));
    Span4Mux_v I__12184 (
            .O(N__72628),
            .I(N__72617));
    Span4Mux_v I__12183 (
            .O(N__72623),
            .I(N__72614));
    Odrv4 I__12182 (
            .O(N__72620),
            .I(clk_en_94));
    Odrv4 I__12181 (
            .O(N__72617),
            .I(clk_en_94));
    Odrv4 I__12180 (
            .O(N__72614),
            .I(clk_en_94));
    InMux I__12179 (
            .O(N__72607),
            .I(N__72604));
    LocalMux I__12178 (
            .O(N__72604),
            .I(shift_srl_49Z0Z_9));
    InMux I__12177 (
            .O(N__72601),
            .I(N__72598));
    LocalMux I__12176 (
            .O(N__72598),
            .I(shift_srl_182Z0Z_0));
    InMux I__12175 (
            .O(N__72595),
            .I(N__72592));
    LocalMux I__12174 (
            .O(N__72592),
            .I(shift_srl_182Z0Z_1));
    InMux I__12173 (
            .O(N__72589),
            .I(N__72586));
    LocalMux I__12172 (
            .O(N__72586),
            .I(shift_srl_182Z0Z_2));
    InMux I__12171 (
            .O(N__72583),
            .I(N__72580));
    LocalMux I__12170 (
            .O(N__72580),
            .I(shift_srl_182Z0Z_3));
    InMux I__12169 (
            .O(N__72577),
            .I(N__72574));
    LocalMux I__12168 (
            .O(N__72574),
            .I(shift_srl_182Z0Z_4));
    InMux I__12167 (
            .O(N__72571),
            .I(N__72568));
    LocalMux I__12166 (
            .O(N__72568),
            .I(shift_srl_182Z0Z_5));
    InMux I__12165 (
            .O(N__72565),
            .I(N__72562));
    LocalMux I__12164 (
            .O(N__72562),
            .I(shift_srl_182Z0Z_6));
    InMux I__12163 (
            .O(N__72559),
            .I(N__72556));
    LocalMux I__12162 (
            .O(N__72556),
            .I(shift_srl_182Z0Z_7));
    CEMux I__12161 (
            .O(N__72553),
            .I(N__72550));
    LocalMux I__12160 (
            .O(N__72550),
            .I(N__72546));
    CEMux I__12159 (
            .O(N__72549),
            .I(N__72543));
    Span4Mux_s2_v I__12158 (
            .O(N__72546),
            .I(N__72538));
    LocalMux I__12157 (
            .O(N__72543),
            .I(N__72538));
    Span4Mux_v I__12156 (
            .O(N__72538),
            .I(N__72535));
    Odrv4 I__12155 (
            .O(N__72535),
            .I(clk_en_182));
    IoInMux I__12154 (
            .O(N__72532),
            .I(N__72529));
    LocalMux I__12153 (
            .O(N__72529),
            .I(N__72526));
    Span4Mux_s3_v I__12152 (
            .O(N__72526),
            .I(N__72523));
    Span4Mux_h I__12151 (
            .O(N__72523),
            .I(N__72520));
    Odrv4 I__12150 (
            .O(N__72520),
            .I(rco_c_94));
    InMux I__12149 (
            .O(N__72517),
            .I(N__72514));
    LocalMux I__12148 (
            .O(N__72514),
            .I(shift_srl_196Z0Z_10));
    InMux I__12147 (
            .O(N__72511),
            .I(N__72508));
    LocalMux I__12146 (
            .O(N__72508),
            .I(shift_srl_196Z0Z_11));
    CEMux I__12145 (
            .O(N__72505),
            .I(N__72501));
    CEMux I__12144 (
            .O(N__72504),
            .I(N__72498));
    LocalMux I__12143 (
            .O(N__72501),
            .I(N__72494));
    LocalMux I__12142 (
            .O(N__72498),
            .I(N__72491));
    CEMux I__12141 (
            .O(N__72497),
            .I(N__72488));
    Span4Mux_v I__12140 (
            .O(N__72494),
            .I(N__72483));
    Span4Mux_h I__12139 (
            .O(N__72491),
            .I(N__72483));
    LocalMux I__12138 (
            .O(N__72488),
            .I(N__72480));
    Odrv4 I__12137 (
            .O(N__72483),
            .I(clk_en_196));
    Odrv12 I__12136 (
            .O(N__72480),
            .I(clk_en_196));
    InMux I__12135 (
            .O(N__72475),
            .I(N__72472));
    LocalMux I__12134 (
            .O(N__72472),
            .I(shift_srl_182Z0Z_10));
    InMux I__12133 (
            .O(N__72469),
            .I(N__72466));
    LocalMux I__12132 (
            .O(N__72466),
            .I(shift_srl_182Z0Z_11));
    InMux I__12131 (
            .O(N__72463),
            .I(N__72460));
    LocalMux I__12130 (
            .O(N__72460),
            .I(shift_srl_182Z0Z_12));
    InMux I__12129 (
            .O(N__72457),
            .I(N__72454));
    LocalMux I__12128 (
            .O(N__72454),
            .I(shift_srl_182Z0Z_13));
    InMux I__12127 (
            .O(N__72451),
            .I(N__72448));
    LocalMux I__12126 (
            .O(N__72448),
            .I(shift_srl_182Z0Z_14));
    InMux I__12125 (
            .O(N__72445),
            .I(N__72442));
    LocalMux I__12124 (
            .O(N__72442),
            .I(shift_srl_182Z0Z_9));
    InMux I__12123 (
            .O(N__72439),
            .I(N__72436));
    LocalMux I__12122 (
            .O(N__72436),
            .I(shift_srl_182Z0Z_8));
    InMux I__12121 (
            .O(N__72433),
            .I(N__72430));
    LocalMux I__12120 (
            .O(N__72430),
            .I(shift_srl_196Z0Z_6));
    InMux I__12119 (
            .O(N__72427),
            .I(N__72424));
    LocalMux I__12118 (
            .O(N__72424),
            .I(shift_srl_196Z0Z_7));
    InMux I__12117 (
            .O(N__72421),
            .I(N__72418));
    LocalMux I__12116 (
            .O(N__72418),
            .I(shift_srl_196Z0Z_8));
    InMux I__12115 (
            .O(N__72415),
            .I(N__72412));
    LocalMux I__12114 (
            .O(N__72412),
            .I(shift_srl_196Z0Z_9));
    CEMux I__12113 (
            .O(N__72409),
            .I(N__72406));
    LocalMux I__12112 (
            .O(N__72406),
            .I(N__72402));
    CEMux I__12111 (
            .O(N__72405),
            .I(N__72399));
    Span4Mux_s3_v I__12110 (
            .O(N__72402),
            .I(N__72396));
    LocalMux I__12109 (
            .O(N__72399),
            .I(N__72393));
    Span4Mux_h I__12108 (
            .O(N__72396),
            .I(N__72388));
    Span4Mux_v I__12107 (
            .O(N__72393),
            .I(N__72388));
    Odrv4 I__12106 (
            .O(N__72388),
            .I(clk_en_197));
    InMux I__12105 (
            .O(N__72385),
            .I(N__72380));
    InMux I__12104 (
            .O(N__72384),
            .I(N__72377));
    CascadeMux I__12103 (
            .O(N__72383),
            .I(N__72373));
    LocalMux I__12102 (
            .O(N__72380),
            .I(N__72370));
    LocalMux I__12101 (
            .O(N__72377),
            .I(N__72367));
    InMux I__12100 (
            .O(N__72376),
            .I(N__72362));
    InMux I__12099 (
            .O(N__72373),
            .I(N__72362));
    Span12Mux_v I__12098 (
            .O(N__72370),
            .I(N__72359));
    Odrv4 I__12097 (
            .O(N__72367),
            .I(shift_srl_196Z0Z_15));
    LocalMux I__12096 (
            .O(N__72362),
            .I(shift_srl_196Z0Z_15));
    Odrv12 I__12095 (
            .O(N__72359),
            .I(shift_srl_196Z0Z_15));
    IoInMux I__12094 (
            .O(N__72352),
            .I(N__72349));
    LocalMux I__12093 (
            .O(N__72349),
            .I(N__72346));
    Span4Mux_s3_v I__12092 (
            .O(N__72346),
            .I(N__72343));
    Span4Mux_h I__12091 (
            .O(N__72343),
            .I(N__72340));
    Odrv4 I__12090 (
            .O(N__72340),
            .I(rco_c_196));
    InMux I__12089 (
            .O(N__72337),
            .I(N__72334));
    LocalMux I__12088 (
            .O(N__72334),
            .I(shift_srl_196Z0Z_14));
    InMux I__12087 (
            .O(N__72331),
            .I(N__72328));
    LocalMux I__12086 (
            .O(N__72328),
            .I(shift_srl_196Z0Z_13));
    InMux I__12085 (
            .O(N__72325),
            .I(N__72322));
    LocalMux I__12084 (
            .O(N__72322),
            .I(shift_srl_196Z0Z_12));
    InMux I__12083 (
            .O(N__72319),
            .I(N__72316));
    LocalMux I__12082 (
            .O(N__72316),
            .I(shift_srl_196Z0Z_0));
    InMux I__12081 (
            .O(N__72313),
            .I(N__72310));
    LocalMux I__12080 (
            .O(N__72310),
            .I(shift_srl_196Z0Z_1));
    InMux I__12079 (
            .O(N__72307),
            .I(N__72304));
    LocalMux I__12078 (
            .O(N__72304),
            .I(shift_srl_196Z0Z_2));
    InMux I__12077 (
            .O(N__72301),
            .I(N__72298));
    LocalMux I__12076 (
            .O(N__72298),
            .I(shift_srl_196Z0Z_3));
    InMux I__12075 (
            .O(N__72295),
            .I(N__72292));
    LocalMux I__12074 (
            .O(N__72292),
            .I(shift_srl_196Z0Z_4));
    InMux I__12073 (
            .O(N__72289),
            .I(N__72286));
    LocalMux I__12072 (
            .O(N__72286),
            .I(shift_srl_196Z0Z_5));
    InMux I__12071 (
            .O(N__72283),
            .I(N__72280));
    LocalMux I__12070 (
            .O(N__72280),
            .I(shift_srl_185Z0Z_4));
    InMux I__12069 (
            .O(N__72277),
            .I(N__72274));
    LocalMux I__12068 (
            .O(N__72274),
            .I(shift_srl_185Z0Z_5));
    InMux I__12067 (
            .O(N__72271),
            .I(N__72268));
    LocalMux I__12066 (
            .O(N__72268),
            .I(shift_srl_185Z0Z_6));
    CEMux I__12065 (
            .O(N__72265),
            .I(N__72262));
    LocalMux I__12064 (
            .O(N__72262),
            .I(N__72258));
    CEMux I__12063 (
            .O(N__72261),
            .I(N__72255));
    Span4Mux_v I__12062 (
            .O(N__72258),
            .I(N__72249));
    LocalMux I__12061 (
            .O(N__72255),
            .I(N__72249));
    CEMux I__12060 (
            .O(N__72254),
            .I(N__72246));
    Span4Mux_h I__12059 (
            .O(N__72249),
            .I(N__72241));
    LocalMux I__12058 (
            .O(N__72246),
            .I(N__72241));
    Sp12to4 I__12057 (
            .O(N__72241),
            .I(N__72238));
    Odrv12 I__12056 (
            .O(N__72238),
            .I(clk_en_194));
    InMux I__12055 (
            .O(N__72235),
            .I(N__72231));
    InMux I__12054 (
            .O(N__72234),
            .I(N__72228));
    LocalMux I__12053 (
            .O(N__72231),
            .I(N__72225));
    LocalMux I__12052 (
            .O(N__72228),
            .I(N__72222));
    Span4Mux_v I__12051 (
            .O(N__72225),
            .I(N__72217));
    Span4Mux_h I__12050 (
            .O(N__72222),
            .I(N__72217));
    Span4Mux_h I__12049 (
            .O(N__72217),
            .I(N__72213));
    InMux I__12048 (
            .O(N__72216),
            .I(N__72210));
    Odrv4 I__12047 (
            .O(N__72213),
            .I(N_4183));
    LocalMux I__12046 (
            .O(N__72210),
            .I(N_4183));
    CEMux I__12045 (
            .O(N__72205),
            .I(N__72201));
    CEMux I__12044 (
            .O(N__72204),
            .I(N__72197));
    LocalMux I__12043 (
            .O(N__72201),
            .I(N__72194));
    CEMux I__12042 (
            .O(N__72200),
            .I(N__72191));
    LocalMux I__12041 (
            .O(N__72197),
            .I(N__72188));
    Span4Mux_v I__12040 (
            .O(N__72194),
            .I(N__72185));
    LocalMux I__12039 (
            .O(N__72191),
            .I(N__72182));
    Span4Mux_h I__12038 (
            .O(N__72188),
            .I(N__72179));
    Odrv4 I__12037 (
            .O(N__72185),
            .I(clk_en_198));
    Odrv4 I__12036 (
            .O(N__72182),
            .I(clk_en_198));
    Odrv4 I__12035 (
            .O(N__72179),
            .I(clk_en_198));
    CascadeMux I__12034 (
            .O(N__72172),
            .I(rco_c_172_cascade_));
    InMux I__12033 (
            .O(N__72169),
            .I(N__72166));
    LocalMux I__12032 (
            .O(N__72166),
            .I(shift_srl_195Z0Z_12));
    InMux I__12031 (
            .O(N__72163),
            .I(N__72160));
    LocalMux I__12030 (
            .O(N__72160),
            .I(shift_srl_195Z0Z_13));
    InMux I__12029 (
            .O(N__72157),
            .I(N__72154));
    LocalMux I__12028 (
            .O(N__72154),
            .I(shift_srl_195Z0Z_14));
    InMux I__12027 (
            .O(N__72151),
            .I(N__72148));
    LocalMux I__12026 (
            .O(N__72148),
            .I(shift_srl_195Z0Z_9));
    InMux I__12025 (
            .O(N__72145),
            .I(N__72142));
    LocalMux I__12024 (
            .O(N__72142),
            .I(shift_srl_195Z0Z_8));
    InMux I__12023 (
            .O(N__72139),
            .I(N__72136));
    LocalMux I__12022 (
            .O(N__72136),
            .I(shift_srl_185Z0Z_0));
    InMux I__12021 (
            .O(N__72133),
            .I(N__72130));
    LocalMux I__12020 (
            .O(N__72130),
            .I(shift_srl_185Z0Z_1));
    InMux I__12019 (
            .O(N__72127),
            .I(N__72124));
    LocalMux I__12018 (
            .O(N__72124),
            .I(shift_srl_185Z0Z_2));
    InMux I__12017 (
            .O(N__72121),
            .I(N__72118));
    LocalMux I__12016 (
            .O(N__72118),
            .I(shift_srl_185Z0Z_3));
    CascadeMux I__12015 (
            .O(N__72115),
            .I(clk_en_0_a3_0_a2_sx_182_cascade_));
    InMux I__12014 (
            .O(N__72112),
            .I(N__72107));
    InMux I__12013 (
            .O(N__72111),
            .I(N__72104));
    InMux I__12012 (
            .O(N__72110),
            .I(N__72101));
    LocalMux I__12011 (
            .O(N__72107),
            .I(N__72098));
    LocalMux I__12010 (
            .O(N__72104),
            .I(N__72093));
    LocalMux I__12009 (
            .O(N__72101),
            .I(N__72090));
    Span4Mux_v I__12008 (
            .O(N__72098),
            .I(N__72087));
    CascadeMux I__12007 (
            .O(N__72097),
            .I(N__72084));
    CascadeMux I__12006 (
            .O(N__72096),
            .I(N__72081));
    Span4Mux_s3_v I__12005 (
            .O(N__72093),
            .I(N__72078));
    Span4Mux_v I__12004 (
            .O(N__72090),
            .I(N__72075));
    Span4Mux_h I__12003 (
            .O(N__72087),
            .I(N__72072));
    InMux I__12002 (
            .O(N__72084),
            .I(N__72069));
    InMux I__12001 (
            .O(N__72081),
            .I(N__72066));
    Span4Mux_v I__12000 (
            .O(N__72078),
            .I(N__72063));
    Span4Mux_v I__11999 (
            .O(N__72075),
            .I(N__72060));
    Span4Mux_v I__11998 (
            .O(N__72072),
            .I(N__72055));
    LocalMux I__11997 (
            .O(N__72069),
            .I(N__72055));
    LocalMux I__11996 (
            .O(N__72066),
            .I(N__72052));
    Span4Mux_v I__11995 (
            .O(N__72063),
            .I(N__72049));
    Span4Mux_h I__11994 (
            .O(N__72060),
            .I(N__72044));
    Span4Mux_v I__11993 (
            .O(N__72055),
            .I(N__72044));
    Sp12to4 I__11992 (
            .O(N__72052),
            .I(N__72041));
    Odrv4 I__11991 (
            .O(N__72049),
            .I(shift_srl_91_RNI20EN1Z0Z_15));
    Odrv4 I__11990 (
            .O(N__72044),
            .I(shift_srl_91_RNI20EN1Z0Z_15));
    Odrv12 I__11989 (
            .O(N__72041),
            .I(shift_srl_91_RNI20EN1Z0Z_15));
    InMux I__11988 (
            .O(N__72034),
            .I(N__72030));
    InMux I__11987 (
            .O(N__72033),
            .I(N__72025));
    LocalMux I__11986 (
            .O(N__72030),
            .I(N__72022));
    InMux I__11985 (
            .O(N__72029),
            .I(N__72019));
    InMux I__11984 (
            .O(N__72028),
            .I(N__72016));
    LocalMux I__11983 (
            .O(N__72025),
            .I(N__72013));
    Span4Mux_v I__11982 (
            .O(N__72022),
            .I(N__72010));
    LocalMux I__11981 (
            .O(N__72019),
            .I(N__72007));
    LocalMux I__11980 (
            .O(N__72016),
            .I(N__72004));
    Span4Mux_v I__11979 (
            .O(N__72013),
            .I(N__72001));
    Span4Mux_v I__11978 (
            .O(N__72010),
            .I(N__71998));
    Span4Mux_v I__11977 (
            .O(N__72007),
            .I(N__71995));
    Span4Mux_h I__11976 (
            .O(N__72004),
            .I(N__71990));
    Span4Mux_h I__11975 (
            .O(N__72001),
            .I(N__71990));
    Odrv4 I__11974 (
            .O(N__71998),
            .I(rco_int_0_a2_0_a2_99_m6_0_a2_9));
    Odrv4 I__11973 (
            .O(N__71995),
            .I(rco_int_0_a2_0_a2_99_m6_0_a2_9));
    Odrv4 I__11972 (
            .O(N__71990),
            .I(rco_int_0_a2_0_a2_99_m6_0_a2_9));
    InMux I__11971 (
            .O(N__71983),
            .I(N__71980));
    LocalMux I__11970 (
            .O(N__71980),
            .I(N__71977));
    Span4Mux_h I__11969 (
            .O(N__71977),
            .I(N__71973));
    InMux I__11968 (
            .O(N__71976),
            .I(N__71970));
    Span4Mux_v I__11967 (
            .O(N__71973),
            .I(N__71967));
    LocalMux I__11966 (
            .O(N__71970),
            .I(N__71964));
    Span4Mux_v I__11965 (
            .O(N__71967),
            .I(N__71961));
    Odrv12 I__11964 (
            .O(N__71964),
            .I(shift_srl_145_RNIN9307Z0Z_15));
    Odrv4 I__11963 (
            .O(N__71961),
            .I(shift_srl_145_RNIN9307Z0Z_15));
    CascadeMux I__11962 (
            .O(N__71956),
            .I(N__71952));
    InMux I__11961 (
            .O(N__71955),
            .I(N__71949));
    InMux I__11960 (
            .O(N__71952),
            .I(N__71946));
    LocalMux I__11959 (
            .O(N__71949),
            .I(N__71943));
    LocalMux I__11958 (
            .O(N__71946),
            .I(N__71938));
    Span4Mux_v I__11957 (
            .O(N__71943),
            .I(N__71938));
    Sp12to4 I__11956 (
            .O(N__71938),
            .I(N__71935));
    Odrv12 I__11955 (
            .O(N__71935),
            .I(rco_int_0_a2_0_a2_1_1_145));
    CascadeMux I__11954 (
            .O(N__71932),
            .I(rco_int_0_a3_0_a2_sx_183_cascade_));
    InMux I__11953 (
            .O(N__71929),
            .I(N__71926));
    LocalMux I__11952 (
            .O(N__71926),
            .I(shift_srl_195Z0Z_10));
    InMux I__11951 (
            .O(N__71923),
            .I(N__71920));
    LocalMux I__11950 (
            .O(N__71920),
            .I(shift_srl_195Z0Z_11));
    InMux I__11949 (
            .O(N__71917),
            .I(N__71914));
    LocalMux I__11948 (
            .O(N__71914),
            .I(shift_srl_183Z0Z_8));
    InMux I__11947 (
            .O(N__71911),
            .I(N__71908));
    LocalMux I__11946 (
            .O(N__71908),
            .I(shift_srl_183Z0Z_7));
    InMux I__11945 (
            .O(N__71905),
            .I(N__71902));
    LocalMux I__11944 (
            .O(N__71902),
            .I(shift_srl_183Z0Z_1));
    InMux I__11943 (
            .O(N__71899),
            .I(N__71896));
    LocalMux I__11942 (
            .O(N__71896),
            .I(shift_srl_183Z0Z_2));
    InMux I__11941 (
            .O(N__71893),
            .I(N__71890));
    LocalMux I__11940 (
            .O(N__71890),
            .I(shift_srl_183Z0Z_3));
    InMux I__11939 (
            .O(N__71887),
            .I(N__71884));
    LocalMux I__11938 (
            .O(N__71884),
            .I(shift_srl_183Z0Z_4));
    InMux I__11937 (
            .O(N__71881),
            .I(N__71878));
    LocalMux I__11936 (
            .O(N__71878),
            .I(shift_srl_183Z0Z_5));
    InMux I__11935 (
            .O(N__71875),
            .I(N__71872));
    LocalMux I__11934 (
            .O(N__71872),
            .I(shift_srl_183Z0Z_6));
    CEMux I__11933 (
            .O(N__71869),
            .I(N__71866));
    LocalMux I__11932 (
            .O(N__71866),
            .I(N__71861));
    CEMux I__11931 (
            .O(N__71865),
            .I(N__71858));
    CEMux I__11930 (
            .O(N__71864),
            .I(N__71855));
    Span4Mux_h I__11929 (
            .O(N__71861),
            .I(N__71852));
    LocalMux I__11928 (
            .O(N__71858),
            .I(N__71849));
    LocalMux I__11927 (
            .O(N__71855),
            .I(N__71846));
    Odrv4 I__11926 (
            .O(N__71852),
            .I(clk_en_183));
    Odrv4 I__11925 (
            .O(N__71849),
            .I(clk_en_183));
    Odrv12 I__11924 (
            .O(N__71846),
            .I(clk_en_183));
    IoInMux I__11923 (
            .O(N__71839),
            .I(N__71836));
    LocalMux I__11922 (
            .O(N__71836),
            .I(N__71833));
    Span4Mux_s1_v I__11921 (
            .O(N__71833),
            .I(N__71830));
    Span4Mux_v I__11920 (
            .O(N__71830),
            .I(N__71827));
    Span4Mux_v I__11919 (
            .O(N__71827),
            .I(N__71824));
    Odrv4 I__11918 (
            .O(N__71824),
            .I(rco_c_181));
    IoInMux I__11917 (
            .O(N__71821),
            .I(N__71818));
    LocalMux I__11916 (
            .O(N__71818),
            .I(N__71815));
    IoSpan4Mux I__11915 (
            .O(N__71815),
            .I(N__71812));
    Sp12to4 I__11914 (
            .O(N__71812),
            .I(N__71809));
    Odrv12 I__11913 (
            .O(N__71809),
            .I(rco_c_180));
    InMux I__11912 (
            .O(N__71806),
            .I(N__71803));
    LocalMux I__11911 (
            .O(N__71803),
            .I(shift_srl_184Z0Z_4));
    InMux I__11910 (
            .O(N__71800),
            .I(N__71797));
    LocalMux I__11909 (
            .O(N__71797),
            .I(shift_srl_184Z0Z_5));
    InMux I__11908 (
            .O(N__71794),
            .I(N__71791));
    LocalMux I__11907 (
            .O(N__71791),
            .I(shift_srl_184Z0Z_6));
    InMux I__11906 (
            .O(N__71788),
            .I(N__71785));
    LocalMux I__11905 (
            .O(N__71785),
            .I(shift_srl_183Z0Z_10));
    InMux I__11904 (
            .O(N__71782),
            .I(N__71779));
    LocalMux I__11903 (
            .O(N__71779),
            .I(shift_srl_183Z0Z_11));
    InMux I__11902 (
            .O(N__71776),
            .I(N__71773));
    LocalMux I__11901 (
            .O(N__71773),
            .I(shift_srl_183Z0Z_12));
    InMux I__11900 (
            .O(N__71770),
            .I(N__71767));
    LocalMux I__11899 (
            .O(N__71767),
            .I(shift_srl_183Z0Z_13));
    InMux I__11898 (
            .O(N__71764),
            .I(N__71761));
    LocalMux I__11897 (
            .O(N__71761),
            .I(shift_srl_183Z0Z_14));
    InMux I__11896 (
            .O(N__71758),
            .I(N__71755));
    LocalMux I__11895 (
            .O(N__71755),
            .I(shift_srl_183Z0Z_9));
    CascadeMux I__11894 (
            .O(N__71752),
            .I(rco_c_162_cascade_));
    InMux I__11893 (
            .O(N__71749),
            .I(N__71746));
    LocalMux I__11892 (
            .O(N__71746),
            .I(shift_srl_184Z0Z_0));
    InMux I__11891 (
            .O(N__71743),
            .I(N__71740));
    LocalMux I__11890 (
            .O(N__71740),
            .I(shift_srl_184Z0Z_1));
    InMux I__11889 (
            .O(N__71737),
            .I(N__71734));
    LocalMux I__11888 (
            .O(N__71734),
            .I(shift_srl_184Z0Z_2));
    InMux I__11887 (
            .O(N__71731),
            .I(N__71728));
    LocalMux I__11886 (
            .O(N__71728),
            .I(shift_srl_184Z0Z_3));
    InMux I__11885 (
            .O(N__71725),
            .I(N__71722));
    LocalMux I__11884 (
            .O(N__71722),
            .I(shift_srl_174Z0Z_0));
    InMux I__11883 (
            .O(N__71719),
            .I(N__71716));
    LocalMux I__11882 (
            .O(N__71716),
            .I(shift_srl_174Z0Z_1));
    InMux I__11881 (
            .O(N__71713),
            .I(N__71710));
    LocalMux I__11880 (
            .O(N__71710),
            .I(shift_srl_174Z0Z_2));
    InMux I__11879 (
            .O(N__71707),
            .I(N__71704));
    LocalMux I__11878 (
            .O(N__71704),
            .I(shift_srl_174Z0Z_3));
    InMux I__11877 (
            .O(N__71701),
            .I(N__71698));
    LocalMux I__11876 (
            .O(N__71698),
            .I(shift_srl_174Z0Z_4));
    InMux I__11875 (
            .O(N__71695),
            .I(N__71692));
    LocalMux I__11874 (
            .O(N__71692),
            .I(shift_srl_174Z0Z_5));
    InMux I__11873 (
            .O(N__71689),
            .I(N__71686));
    LocalMux I__11872 (
            .O(N__71686),
            .I(shift_srl_174Z0Z_6));
    IoInMux I__11871 (
            .O(N__71683),
            .I(N__71680));
    LocalMux I__11870 (
            .O(N__71680),
            .I(N__71677));
    IoSpan4Mux I__11869 (
            .O(N__71677),
            .I(N__71674));
    Span4Mux_s2_v I__11868 (
            .O(N__71674),
            .I(N__71671));
    Span4Mux_v I__11867 (
            .O(N__71671),
            .I(N__71668));
    Sp12to4 I__11866 (
            .O(N__71668),
            .I(N__71665));
    Span12Mux_h I__11865 (
            .O(N__71665),
            .I(N__71662));
    Span12Mux_v I__11864 (
            .O(N__71662),
            .I(N__71659));
    Odrv12 I__11863 (
            .O(N__71659),
            .I(rco_c_166));
    InMux I__11862 (
            .O(N__71656),
            .I(N__71653));
    LocalMux I__11861 (
            .O(N__71653),
            .I(N__71650));
    Span4Mux_v I__11860 (
            .O(N__71650),
            .I(N__71646));
    InMux I__11859 (
            .O(N__71649),
            .I(N__71643));
    Span4Mux_h I__11858 (
            .O(N__71646),
            .I(N__71638));
    LocalMux I__11857 (
            .O(N__71643),
            .I(N__71638));
    Span4Mux_h I__11856 (
            .O(N__71638),
            .I(N__71635));
    Span4Mux_h I__11855 (
            .O(N__71635),
            .I(N__71631));
    InMux I__11854 (
            .O(N__71634),
            .I(N__71628));
    Odrv4 I__11853 (
            .O(N__71631),
            .I(shift_srl_159_RNIDDRE1Z0Z_15));
    LocalMux I__11852 (
            .O(N__71628),
            .I(shift_srl_159_RNIDDRE1Z0Z_15));
    InMux I__11851 (
            .O(N__71623),
            .I(N__71620));
    LocalMux I__11850 (
            .O(N__71620),
            .I(shift_srl_62Z0Z_0));
    InMux I__11849 (
            .O(N__71617),
            .I(N__71614));
    LocalMux I__11848 (
            .O(N__71614),
            .I(shift_srl_62Z0Z_1));
    InMux I__11847 (
            .O(N__71611),
            .I(N__71608));
    LocalMux I__11846 (
            .O(N__71608),
            .I(shift_srl_62Z0Z_2));
    InMux I__11845 (
            .O(N__71605),
            .I(N__71602));
    LocalMux I__11844 (
            .O(N__71602),
            .I(shift_srl_62Z0Z_3));
    InMux I__11843 (
            .O(N__71599),
            .I(N__71596));
    LocalMux I__11842 (
            .O(N__71596),
            .I(shift_srl_62Z0Z_4));
    InMux I__11841 (
            .O(N__71593),
            .I(N__71590));
    LocalMux I__11840 (
            .O(N__71590),
            .I(shift_srl_62Z0Z_5));
    InMux I__11839 (
            .O(N__71587),
            .I(N__71584));
    LocalMux I__11838 (
            .O(N__71584),
            .I(shift_srl_62Z0Z_6));
    InMux I__11837 (
            .O(N__71581),
            .I(N__71578));
    LocalMux I__11836 (
            .O(N__71578),
            .I(shift_srl_61Z0Z_6));
    InMux I__11835 (
            .O(N__71575),
            .I(N__71572));
    LocalMux I__11834 (
            .O(N__71572),
            .I(shift_srl_61Z0Z_7));
    CascadeMux I__11833 (
            .O(N__71569),
            .I(rco_int_0_a2_0_a2_s_0_0_35_cascade_));
    InMux I__11832 (
            .O(N__71566),
            .I(N__71563));
    LocalMux I__11831 (
            .O(N__71563),
            .I(shift_srl_31_RNI84161_0Z0Z_15));
    InMux I__11830 (
            .O(N__71560),
            .I(N__71557));
    LocalMux I__11829 (
            .O(N__71557),
            .I(shift_srl_37_RNI973EZ0Z_15));
    InMux I__11828 (
            .O(N__71554),
            .I(N__71551));
    LocalMux I__11827 (
            .O(N__71551),
            .I(N__71548));
    Odrv4 I__11826 (
            .O(N__71548),
            .I(rco_int_0_a2_0_a2_99_m6_0_a2_2));
    InMux I__11825 (
            .O(N__71545),
            .I(N__71536));
    InMux I__11824 (
            .O(N__71544),
            .I(N__71536));
    InMux I__11823 (
            .O(N__71543),
            .I(N__71533));
    InMux I__11822 (
            .O(N__71542),
            .I(N__71528));
    InMux I__11821 (
            .O(N__71541),
            .I(N__71528));
    LocalMux I__11820 (
            .O(N__71536),
            .I(N__71523));
    LocalMux I__11819 (
            .O(N__71533),
            .I(N__71518));
    LocalMux I__11818 (
            .O(N__71528),
            .I(N__71518));
    InMux I__11817 (
            .O(N__71527),
            .I(N__71513));
    InMux I__11816 (
            .O(N__71526),
            .I(N__71513));
    Span4Mux_v I__11815 (
            .O(N__71523),
            .I(N__71510));
    Odrv12 I__11814 (
            .O(N__71518),
            .I(shift_srl_26Z0Z_15));
    LocalMux I__11813 (
            .O(N__71513),
            .I(shift_srl_26Z0Z_15));
    Odrv4 I__11812 (
            .O(N__71510),
            .I(shift_srl_26Z0Z_15));
    InMux I__11811 (
            .O(N__71503),
            .I(N__71496));
    CascadeMux I__11810 (
            .O(N__71502),
            .I(N__71493));
    InMux I__11809 (
            .O(N__71501),
            .I(N__71489));
    InMux I__11808 (
            .O(N__71500),
            .I(N__71486));
    InMux I__11807 (
            .O(N__71499),
            .I(N__71483));
    LocalMux I__11806 (
            .O(N__71496),
            .I(N__71480));
    InMux I__11805 (
            .O(N__71493),
            .I(N__71475));
    InMux I__11804 (
            .O(N__71492),
            .I(N__71475));
    LocalMux I__11803 (
            .O(N__71489),
            .I(N__71470));
    LocalMux I__11802 (
            .O(N__71486),
            .I(N__71470));
    LocalMux I__11801 (
            .O(N__71483),
            .I(N__71467));
    Span4Mux_h I__11800 (
            .O(N__71480),
            .I(N__71464));
    LocalMux I__11799 (
            .O(N__71475),
            .I(N__71460));
    Span4Mux_v I__11798 (
            .O(N__71470),
            .I(N__71455));
    Span4Mux_h I__11797 (
            .O(N__71467),
            .I(N__71455));
    Span4Mux_h I__11796 (
            .O(N__71464),
            .I(N__71452));
    InMux I__11795 (
            .O(N__71463),
            .I(N__71449));
    Span12Mux_h I__11794 (
            .O(N__71460),
            .I(N__71446));
    Span4Mux_v I__11793 (
            .O(N__71455),
            .I(N__71443));
    Span4Mux_v I__11792 (
            .O(N__71452),
            .I(N__71440));
    LocalMux I__11791 (
            .O(N__71449),
            .I(shift_srl_25Z0Z_15));
    Odrv12 I__11790 (
            .O(N__71446),
            .I(shift_srl_25Z0Z_15));
    Odrv4 I__11789 (
            .O(N__71443),
            .I(shift_srl_25Z0Z_15));
    Odrv4 I__11788 (
            .O(N__71440),
            .I(shift_srl_25Z0Z_15));
    CascadeMux I__11787 (
            .O(N__71431),
            .I(N__71427));
    CascadeMux I__11786 (
            .O(N__71430),
            .I(N__71423));
    InMux I__11785 (
            .O(N__71427),
            .I(N__71418));
    InMux I__11784 (
            .O(N__71426),
            .I(N__71415));
    InMux I__11783 (
            .O(N__71423),
            .I(N__71410));
    InMux I__11782 (
            .O(N__71422),
            .I(N__71410));
    InMux I__11781 (
            .O(N__71421),
            .I(N__71407));
    LocalMux I__11780 (
            .O(N__71418),
            .I(N__71400));
    LocalMux I__11779 (
            .O(N__71415),
            .I(N__71400));
    LocalMux I__11778 (
            .O(N__71410),
            .I(N__71400));
    LocalMux I__11777 (
            .O(N__71407),
            .I(shift_srl_27Z0Z_15));
    Odrv12 I__11776 (
            .O(N__71400),
            .I(shift_srl_27Z0Z_15));
    InMux I__11775 (
            .O(N__71395),
            .I(N__71392));
    LocalMux I__11774 (
            .O(N__71392),
            .I(shift_srl_27_RNIAA521_0Z0Z_15));
    InMux I__11773 (
            .O(N__71389),
            .I(N__71386));
    LocalMux I__11772 (
            .O(N__71386),
            .I(N__71383));
    Span4Mux_h I__11771 (
            .O(N__71383),
            .I(N__71380));
    Odrv4 I__11770 (
            .O(N__71380),
            .I(rco_int_0_a2_0_a2_99_m6_0_a2_3));
    InMux I__11769 (
            .O(N__71377),
            .I(N__71374));
    LocalMux I__11768 (
            .O(N__71374),
            .I(shift_srl_39Z0Z_10));
    InMux I__11767 (
            .O(N__71371),
            .I(N__71368));
    LocalMux I__11766 (
            .O(N__71368),
            .I(shift_srl_39Z0Z_9));
    InMux I__11765 (
            .O(N__71365),
            .I(N__71362));
    LocalMux I__11764 (
            .O(N__71362),
            .I(shift_srl_61Z0Z_1));
    InMux I__11763 (
            .O(N__71359),
            .I(N__71356));
    LocalMux I__11762 (
            .O(N__71356),
            .I(shift_srl_61Z0Z_2));
    InMux I__11761 (
            .O(N__71353),
            .I(N__71350));
    LocalMux I__11760 (
            .O(N__71350),
            .I(shift_srl_61Z0Z_3));
    InMux I__11759 (
            .O(N__71347),
            .I(N__71344));
    LocalMux I__11758 (
            .O(N__71344),
            .I(shift_srl_61Z0Z_4));
    InMux I__11757 (
            .O(N__71341),
            .I(N__71338));
    LocalMux I__11756 (
            .O(N__71338),
            .I(shift_srl_61Z0Z_5));
    InMux I__11755 (
            .O(N__71335),
            .I(N__71332));
    LocalMux I__11754 (
            .O(N__71332),
            .I(shift_srl_48Z0Z_10));
    InMux I__11753 (
            .O(N__71329),
            .I(N__71326));
    LocalMux I__11752 (
            .O(N__71326),
            .I(shift_srl_48Z0Z_9));
    InMux I__11751 (
            .O(N__71323),
            .I(N__71320));
    LocalMux I__11750 (
            .O(N__71320),
            .I(shift_srl_48Z0Z_8));
    InMux I__11749 (
            .O(N__71317),
            .I(N__71314));
    LocalMux I__11748 (
            .O(N__71314),
            .I(shift_srl_48Z0Z_6));
    InMux I__11747 (
            .O(N__71311),
            .I(N__71308));
    LocalMux I__11746 (
            .O(N__71308),
            .I(shift_srl_48Z0Z_7));
    InMux I__11745 (
            .O(N__71305),
            .I(N__71302));
    LocalMux I__11744 (
            .O(N__71302),
            .I(shift_srl_39_RNIG4I71Z0Z_15));
    InMux I__11743 (
            .O(N__71299),
            .I(N__71296));
    LocalMux I__11742 (
            .O(N__71296),
            .I(shift_srl_39Z0Z_14));
    InMux I__11741 (
            .O(N__71293),
            .I(N__71290));
    LocalMux I__11740 (
            .O(N__71290),
            .I(shift_srl_39Z0Z_13));
    InMux I__11739 (
            .O(N__71287),
            .I(N__71284));
    LocalMux I__11738 (
            .O(N__71284),
            .I(shift_srl_39Z0Z_12));
    InMux I__11737 (
            .O(N__71281),
            .I(N__71278));
    LocalMux I__11736 (
            .O(N__71278),
            .I(shift_srl_39Z0Z_11));
    InMux I__11735 (
            .O(N__71275),
            .I(N__71272));
    LocalMux I__11734 (
            .O(N__71272),
            .I(shift_srl_59Z0Z_6));
    InMux I__11733 (
            .O(N__71269),
            .I(N__71266));
    LocalMux I__11732 (
            .O(N__71266),
            .I(N__71263));
    Odrv12 I__11731 (
            .O(N__71263),
            .I(shift_srl_59Z0Z_7));
    InMux I__11730 (
            .O(N__71260),
            .I(N__71257));
    LocalMux I__11729 (
            .O(N__71257),
            .I(shift_srl_44Z0Z_10));
    InMux I__11728 (
            .O(N__71254),
            .I(N__71251));
    LocalMux I__11727 (
            .O(N__71251),
            .I(shift_srl_44Z0Z_11));
    InMux I__11726 (
            .O(N__71248),
            .I(N__71245));
    LocalMux I__11725 (
            .O(N__71245),
            .I(shift_srl_44Z0Z_12));
    InMux I__11724 (
            .O(N__71242),
            .I(N__71239));
    LocalMux I__11723 (
            .O(N__71239),
            .I(shift_srl_44Z0Z_13));
    InMux I__11722 (
            .O(N__71236),
            .I(N__71233));
    LocalMux I__11721 (
            .O(N__71233),
            .I(shift_srl_44Z0Z_14));
    InMux I__11720 (
            .O(N__71230),
            .I(N__71227));
    LocalMux I__11719 (
            .O(N__71227),
            .I(shift_srl_44Z0Z_9));
    InMux I__11718 (
            .O(N__71224),
            .I(N__71221));
    LocalMux I__11717 (
            .O(N__71221),
            .I(shift_srl_44Z0Z_7));
    InMux I__11716 (
            .O(N__71218),
            .I(N__71215));
    LocalMux I__11715 (
            .O(N__71215),
            .I(shift_srl_44Z0Z_8));
    CEMux I__11714 (
            .O(N__71212),
            .I(N__71208));
    CEMux I__11713 (
            .O(N__71211),
            .I(N__71205));
    LocalMux I__11712 (
            .O(N__71208),
            .I(N__71200));
    LocalMux I__11711 (
            .O(N__71205),
            .I(N__71200));
    Span4Mux_v I__11710 (
            .O(N__71200),
            .I(N__71197));
    Span4Mux_h I__11709 (
            .O(N__71197),
            .I(N__71194));
    Odrv4 I__11708 (
            .O(N__71194),
            .I(clk_en_44));
    InMux I__11707 (
            .O(N__71191),
            .I(N__71188));
    LocalMux I__11706 (
            .O(N__71188),
            .I(shift_srl_41Z0Z_9));
    InMux I__11705 (
            .O(N__71185),
            .I(N__71182));
    LocalMux I__11704 (
            .O(N__71182),
            .I(shift_srl_41Z0Z_8));
    InMux I__11703 (
            .O(N__71179),
            .I(N__71176));
    LocalMux I__11702 (
            .O(N__71176),
            .I(shift_srl_59Z0Z_0));
    InMux I__11701 (
            .O(N__71173),
            .I(N__71170));
    LocalMux I__11700 (
            .O(N__71170),
            .I(shift_srl_59Z0Z_1));
    InMux I__11699 (
            .O(N__71167),
            .I(N__71164));
    LocalMux I__11698 (
            .O(N__71164),
            .I(shift_srl_59Z0Z_2));
    InMux I__11697 (
            .O(N__71161),
            .I(N__71158));
    LocalMux I__11696 (
            .O(N__71158),
            .I(shift_srl_59Z0Z_3));
    InMux I__11695 (
            .O(N__71155),
            .I(N__71152));
    LocalMux I__11694 (
            .O(N__71152),
            .I(shift_srl_59Z0Z_4));
    InMux I__11693 (
            .O(N__71149),
            .I(N__71146));
    LocalMux I__11692 (
            .O(N__71146),
            .I(shift_srl_59Z0Z_5));
    InMux I__11691 (
            .O(N__71143),
            .I(N__71140));
    LocalMux I__11690 (
            .O(N__71140),
            .I(shift_srl_53Z0Z_14));
    InMux I__11689 (
            .O(N__71137),
            .I(N__71134));
    LocalMux I__11688 (
            .O(N__71134),
            .I(shift_srl_53Z0Z_9));
    InMux I__11687 (
            .O(N__71131),
            .I(N__71128));
    LocalMux I__11686 (
            .O(N__71128),
            .I(shift_srl_53Z0Z_7));
    InMux I__11685 (
            .O(N__71125),
            .I(N__71122));
    LocalMux I__11684 (
            .O(N__71122),
            .I(shift_srl_53Z0Z_8));
    InMux I__11683 (
            .O(N__71119),
            .I(N__71116));
    LocalMux I__11682 (
            .O(N__71116),
            .I(shift_srl_41Z0Z_10));
    InMux I__11681 (
            .O(N__71113),
            .I(N__71110));
    LocalMux I__11680 (
            .O(N__71110),
            .I(shift_srl_41Z0Z_11));
    InMux I__11679 (
            .O(N__71107),
            .I(N__71104));
    LocalMux I__11678 (
            .O(N__71104),
            .I(shift_srl_41Z0Z_12));
    InMux I__11677 (
            .O(N__71101),
            .I(N__71098));
    LocalMux I__11676 (
            .O(N__71098),
            .I(shift_srl_41Z0Z_13));
    InMux I__11675 (
            .O(N__71095),
            .I(N__71092));
    LocalMux I__11674 (
            .O(N__71092),
            .I(shift_srl_41Z0Z_14));
    InMux I__11673 (
            .O(N__71089),
            .I(N__71086));
    LocalMux I__11672 (
            .O(N__71086),
            .I(shift_srl_53Z0Z_3));
    InMux I__11671 (
            .O(N__71083),
            .I(N__71080));
    LocalMux I__11670 (
            .O(N__71080),
            .I(shift_srl_53Z0Z_4));
    InMux I__11669 (
            .O(N__71077),
            .I(N__71074));
    LocalMux I__11668 (
            .O(N__71074),
            .I(shift_srl_53Z0Z_5));
    InMux I__11667 (
            .O(N__71071),
            .I(N__71068));
    LocalMux I__11666 (
            .O(N__71068),
            .I(shift_srl_53Z0Z_6));
    InMux I__11665 (
            .O(N__71065),
            .I(N__71062));
    LocalMux I__11664 (
            .O(N__71062),
            .I(shift_srl_53Z0Z_10));
    InMux I__11663 (
            .O(N__71059),
            .I(N__71056));
    LocalMux I__11662 (
            .O(N__71056),
            .I(shift_srl_53Z0Z_11));
    InMux I__11661 (
            .O(N__71053),
            .I(N__71050));
    LocalMux I__11660 (
            .O(N__71050),
            .I(shift_srl_53Z0Z_12));
    InMux I__11659 (
            .O(N__71047),
            .I(N__71044));
    LocalMux I__11658 (
            .O(N__71044),
            .I(shift_srl_53Z0Z_13));
    InMux I__11657 (
            .O(N__71041),
            .I(N__71038));
    LocalMux I__11656 (
            .O(N__71038),
            .I(shift_srl_51Z0Z_11));
    InMux I__11655 (
            .O(N__71035),
            .I(N__71032));
    LocalMux I__11654 (
            .O(N__71032),
            .I(shift_srl_51Z0Z_12));
    InMux I__11653 (
            .O(N__71029),
            .I(N__71026));
    LocalMux I__11652 (
            .O(N__71026),
            .I(shift_srl_51Z0Z_13));
    InMux I__11651 (
            .O(N__71023),
            .I(N__71020));
    LocalMux I__11650 (
            .O(N__71020),
            .I(shift_srl_51Z0Z_14));
    InMux I__11649 (
            .O(N__71017),
            .I(N__71014));
    LocalMux I__11648 (
            .O(N__71014),
            .I(shift_srl_51Z0Z_6));
    InMux I__11647 (
            .O(N__71011),
            .I(N__71008));
    LocalMux I__11646 (
            .O(N__71008),
            .I(shift_srl_53Z0Z_0));
    InMux I__11645 (
            .O(N__71005),
            .I(N__71002));
    LocalMux I__11644 (
            .O(N__71002),
            .I(shift_srl_53Z0Z_1));
    InMux I__11643 (
            .O(N__70999),
            .I(N__70996));
    LocalMux I__11642 (
            .O(N__70996),
            .I(shift_srl_53Z0Z_2));
    InMux I__11641 (
            .O(N__70993),
            .I(N__70990));
    LocalMux I__11640 (
            .O(N__70990),
            .I(shift_srl_97Z0Z_0));
    InMux I__11639 (
            .O(N__70987),
            .I(N__70984));
    LocalMux I__11638 (
            .O(N__70984),
            .I(shift_srl_97Z0Z_1));
    InMux I__11637 (
            .O(N__70981),
            .I(N__70978));
    LocalMux I__11636 (
            .O(N__70978),
            .I(shift_srl_97Z0Z_2));
    InMux I__11635 (
            .O(N__70975),
            .I(N__70972));
    LocalMux I__11634 (
            .O(N__70972),
            .I(shift_srl_97Z0Z_3));
    InMux I__11633 (
            .O(N__70969),
            .I(N__70966));
    LocalMux I__11632 (
            .O(N__70966),
            .I(shift_srl_97Z0Z_4));
    InMux I__11631 (
            .O(N__70963),
            .I(N__70960));
    LocalMux I__11630 (
            .O(N__70960),
            .I(shift_srl_97Z0Z_5));
    InMux I__11629 (
            .O(N__70957),
            .I(N__70954));
    LocalMux I__11628 (
            .O(N__70954),
            .I(shift_srl_97Z0Z_6));
    InMux I__11627 (
            .O(N__70951),
            .I(N__70948));
    LocalMux I__11626 (
            .O(N__70948),
            .I(shift_srl_97Z0Z_7));
    CEMux I__11625 (
            .O(N__70945),
            .I(N__70941));
    CEMux I__11624 (
            .O(N__70944),
            .I(N__70938));
    LocalMux I__11623 (
            .O(N__70941),
            .I(clk_en_97));
    LocalMux I__11622 (
            .O(N__70938),
            .I(clk_en_97));
    InMux I__11621 (
            .O(N__70933),
            .I(N__70930));
    LocalMux I__11620 (
            .O(N__70930),
            .I(shift_srl_51Z0Z_10));
    InMux I__11619 (
            .O(N__70927),
            .I(N__70924));
    LocalMux I__11618 (
            .O(N__70924),
            .I(shift_srl_46Z0Z_7));
    InMux I__11617 (
            .O(N__70921),
            .I(N__70918));
    LocalMux I__11616 (
            .O(N__70918),
            .I(shift_srl_46Z0Z_10));
    InMux I__11615 (
            .O(N__70915),
            .I(N__70912));
    LocalMux I__11614 (
            .O(N__70912),
            .I(shift_srl_46Z0Z_11));
    InMux I__11613 (
            .O(N__70909),
            .I(N__70906));
    LocalMux I__11612 (
            .O(N__70906),
            .I(shift_srl_46Z0Z_12));
    InMux I__11611 (
            .O(N__70903),
            .I(N__70900));
    LocalMux I__11610 (
            .O(N__70900),
            .I(shift_srl_46Z0Z_13));
    InMux I__11609 (
            .O(N__70897),
            .I(N__70894));
    LocalMux I__11608 (
            .O(N__70894),
            .I(shift_srl_46Z0Z_14));
    InMux I__11607 (
            .O(N__70891),
            .I(N__70888));
    LocalMux I__11606 (
            .O(N__70888),
            .I(shift_srl_46Z0Z_6));
    InMux I__11605 (
            .O(N__70885),
            .I(N__70882));
    LocalMux I__11604 (
            .O(N__70882),
            .I(shift_srl_46Z0Z_4));
    InMux I__11603 (
            .O(N__70879),
            .I(N__70876));
    LocalMux I__11602 (
            .O(N__70876),
            .I(shift_srl_46Z0Z_5));
    CEMux I__11601 (
            .O(N__70873),
            .I(N__70869));
    CEMux I__11600 (
            .O(N__70872),
            .I(N__70866));
    LocalMux I__11599 (
            .O(N__70869),
            .I(N__70863));
    LocalMux I__11598 (
            .O(N__70866),
            .I(N__70860));
    Span12Mux_h I__11597 (
            .O(N__70863),
            .I(N__70855));
    Sp12to4 I__11596 (
            .O(N__70860),
            .I(N__70855));
    Odrv12 I__11595 (
            .O(N__70855),
            .I(clk_en_46));
    CascadeMux I__11594 (
            .O(N__70852),
            .I(N__70849));
    InMux I__11593 (
            .O(N__70849),
            .I(N__70844));
    InMux I__11592 (
            .O(N__70848),
            .I(N__70838));
    InMux I__11591 (
            .O(N__70847),
            .I(N__70838));
    LocalMux I__11590 (
            .O(N__70844),
            .I(N__70835));
    InMux I__11589 (
            .O(N__70843),
            .I(N__70832));
    LocalMux I__11588 (
            .O(N__70838),
            .I(N__70829));
    Span12Mux_v I__11587 (
            .O(N__70835),
            .I(N__70826));
    LocalMux I__11586 (
            .O(N__70832),
            .I(shift_srl_97Z0Z_15));
    Odrv4 I__11585 (
            .O(N__70829),
            .I(shift_srl_97Z0Z_15));
    Odrv12 I__11584 (
            .O(N__70826),
            .I(shift_srl_97Z0Z_15));
    InMux I__11583 (
            .O(N__70819),
            .I(N__70816));
    LocalMux I__11582 (
            .O(N__70816),
            .I(shift_srl_92Z0Z_0));
    InMux I__11581 (
            .O(N__70813),
            .I(N__70810));
    LocalMux I__11580 (
            .O(N__70810),
            .I(shift_srl_92Z0Z_1));
    InMux I__11579 (
            .O(N__70807),
            .I(N__70804));
    LocalMux I__11578 (
            .O(N__70804),
            .I(shift_srl_92Z0Z_2));
    InMux I__11577 (
            .O(N__70801),
            .I(N__70798));
    LocalMux I__11576 (
            .O(N__70798),
            .I(shift_srl_92Z0Z_3));
    InMux I__11575 (
            .O(N__70795),
            .I(N__70792));
    LocalMux I__11574 (
            .O(N__70792),
            .I(shift_srl_92Z0Z_4));
    InMux I__11573 (
            .O(N__70789),
            .I(N__70786));
    LocalMux I__11572 (
            .O(N__70786),
            .I(shift_srl_92Z0Z_5));
    InMux I__11571 (
            .O(N__70783),
            .I(N__70780));
    LocalMux I__11570 (
            .O(N__70780),
            .I(shift_srl_92Z0Z_6));
    InMux I__11569 (
            .O(N__70777),
            .I(N__70774));
    LocalMux I__11568 (
            .O(N__70774),
            .I(shift_srl_92Z0Z_7));
    InMux I__11567 (
            .O(N__70771),
            .I(N__70768));
    LocalMux I__11566 (
            .O(N__70768),
            .I(N__70765));
    Odrv4 I__11565 (
            .O(N__70765),
            .I(shift_srl_92Z0Z_8));
    CEMux I__11564 (
            .O(N__70762),
            .I(N__70759));
    LocalMux I__11563 (
            .O(N__70759),
            .I(N__70754));
    CEMux I__11562 (
            .O(N__70758),
            .I(N__70751));
    CEMux I__11561 (
            .O(N__70757),
            .I(N__70748));
    Span4Mux_s2_v I__11560 (
            .O(N__70754),
            .I(N__70743));
    LocalMux I__11559 (
            .O(N__70751),
            .I(N__70743));
    LocalMux I__11558 (
            .O(N__70748),
            .I(N__70740));
    Span4Mux_h I__11557 (
            .O(N__70743),
            .I(N__70737));
    Span4Mux_h I__11556 (
            .O(N__70740),
            .I(N__70734));
    Odrv4 I__11555 (
            .O(N__70737),
            .I(clk_en_92));
    Odrv4 I__11554 (
            .O(N__70734),
            .I(clk_en_92));
    InMux I__11553 (
            .O(N__70729),
            .I(N__70726));
    LocalMux I__11552 (
            .O(N__70726),
            .I(N__70723));
    Span4Mux_v I__11551 (
            .O(N__70723),
            .I(N__70720));
    Span4Mux_v I__11550 (
            .O(N__70720),
            .I(N__70713));
    InMux I__11549 (
            .O(N__70719),
            .I(N__70710));
    CascadeMux I__11548 (
            .O(N__70718),
            .I(N__70707));
    InMux I__11547 (
            .O(N__70717),
            .I(N__70702));
    InMux I__11546 (
            .O(N__70716),
            .I(N__70702));
    Sp12to4 I__11545 (
            .O(N__70713),
            .I(N__70697));
    LocalMux I__11544 (
            .O(N__70710),
            .I(N__70697));
    InMux I__11543 (
            .O(N__70707),
            .I(N__70694));
    LocalMux I__11542 (
            .O(N__70702),
            .I(N__70683));
    Span12Mux_h I__11541 (
            .O(N__70697),
            .I(N__70683));
    LocalMux I__11540 (
            .O(N__70694),
            .I(N__70683));
    InMux I__11539 (
            .O(N__70693),
            .I(N__70674));
    InMux I__11538 (
            .O(N__70692),
            .I(N__70674));
    InMux I__11537 (
            .O(N__70691),
            .I(N__70674));
    InMux I__11536 (
            .O(N__70690),
            .I(N__70674));
    Odrv12 I__11535 (
            .O(N__70683),
            .I(shift_srl_146Z0Z_15));
    LocalMux I__11534 (
            .O(N__70674),
            .I(shift_srl_146Z0Z_15));
    IoInMux I__11533 (
            .O(N__70669),
            .I(N__70666));
    LocalMux I__11532 (
            .O(N__70666),
            .I(N__70663));
    Odrv4 I__11531 (
            .O(N__70663),
            .I(rco_c_146));
    InMux I__11530 (
            .O(N__70660),
            .I(N__70657));
    LocalMux I__11529 (
            .O(N__70657),
            .I(shift_srl_197Z0Z_11));
    InMux I__11528 (
            .O(N__70654),
            .I(N__70651));
    LocalMux I__11527 (
            .O(N__70651),
            .I(shift_srl_197Z0Z_12));
    InMux I__11526 (
            .O(N__70648),
            .I(N__70645));
    LocalMux I__11525 (
            .O(N__70645),
            .I(shift_srl_197Z0Z_13));
    InMux I__11524 (
            .O(N__70642),
            .I(N__70639));
    LocalMux I__11523 (
            .O(N__70639),
            .I(shift_srl_197Z0Z_14));
    InMux I__11522 (
            .O(N__70636),
            .I(N__70633));
    LocalMux I__11521 (
            .O(N__70633),
            .I(N__70630));
    Span4Mux_h I__11520 (
            .O(N__70630),
            .I(N__70626));
    InMux I__11519 (
            .O(N__70629),
            .I(N__70623));
    Span4Mux_v I__11518 (
            .O(N__70626),
            .I(N__70620));
    LocalMux I__11517 (
            .O(N__70623),
            .I(shift_srl_197Z0Z_15));
    Odrv4 I__11516 (
            .O(N__70620),
            .I(shift_srl_197Z0Z_15));
    InMux I__11515 (
            .O(N__70615),
            .I(N__70612));
    LocalMux I__11514 (
            .O(N__70612),
            .I(shift_srl_197Z0Z_9));
    InMux I__11513 (
            .O(N__70609),
            .I(N__70606));
    LocalMux I__11512 (
            .O(N__70606),
            .I(shift_srl_197Z0Z_7));
    InMux I__11511 (
            .O(N__70603),
            .I(N__70600));
    LocalMux I__11510 (
            .O(N__70600),
            .I(shift_srl_197Z0Z_8));
    InMux I__11509 (
            .O(N__70597),
            .I(N__70594));
    LocalMux I__11508 (
            .O(N__70594),
            .I(N__70591));
    Odrv4 I__11507 (
            .O(N__70591),
            .I(shift_srl_93Z0Z_8));
    InMux I__11506 (
            .O(N__70588),
            .I(N__70585));
    LocalMux I__11505 (
            .O(N__70585),
            .I(shift_srl_93Z0Z_6));
    InMux I__11504 (
            .O(N__70582),
            .I(N__70579));
    LocalMux I__11503 (
            .O(N__70579),
            .I(shift_srl_93Z0Z_7));
    CEMux I__11502 (
            .O(N__70576),
            .I(N__70572));
    CEMux I__11501 (
            .O(N__70575),
            .I(N__70568));
    LocalMux I__11500 (
            .O(N__70572),
            .I(N__70565));
    CEMux I__11499 (
            .O(N__70571),
            .I(N__70562));
    LocalMux I__11498 (
            .O(N__70568),
            .I(N__70559));
    Span4Mux_v I__11497 (
            .O(N__70565),
            .I(N__70554));
    LocalMux I__11496 (
            .O(N__70562),
            .I(N__70554));
    Span4Mux_h I__11495 (
            .O(N__70559),
            .I(N__70549));
    Span4Mux_s1_v I__11494 (
            .O(N__70554),
            .I(N__70549));
    Odrv4 I__11493 (
            .O(N__70549),
            .I(clk_en_93));
    InMux I__11492 (
            .O(N__70546),
            .I(N__70543));
    LocalMux I__11491 (
            .O(N__70543),
            .I(shift_srl_197Z0Z_2));
    InMux I__11490 (
            .O(N__70540),
            .I(N__70537));
    LocalMux I__11489 (
            .O(N__70537),
            .I(shift_srl_197Z0Z_3));
    InMux I__11488 (
            .O(N__70534),
            .I(N__70531));
    LocalMux I__11487 (
            .O(N__70531),
            .I(shift_srl_197Z0Z_4));
    InMux I__11486 (
            .O(N__70528),
            .I(N__70525));
    LocalMux I__11485 (
            .O(N__70525),
            .I(shift_srl_197Z0Z_5));
    InMux I__11484 (
            .O(N__70522),
            .I(N__70519));
    LocalMux I__11483 (
            .O(N__70519),
            .I(shift_srl_197Z0Z_6));
    InMux I__11482 (
            .O(N__70516),
            .I(N__70513));
    LocalMux I__11481 (
            .O(N__70513),
            .I(shift_srl_197Z0Z_0));
    InMux I__11480 (
            .O(N__70510),
            .I(N__70507));
    LocalMux I__11479 (
            .O(N__70507),
            .I(shift_srl_197Z0Z_1));
    InMux I__11478 (
            .O(N__70504),
            .I(N__70501));
    LocalMux I__11477 (
            .O(N__70501),
            .I(shift_srl_197Z0Z_10));
    InMux I__11476 (
            .O(N__70498),
            .I(N__70495));
    LocalMux I__11475 (
            .O(N__70495),
            .I(N__70492));
    Odrv4 I__11474 (
            .O(N__70492),
            .I(shift_srl_198Z0Z_7));
    InMux I__11473 (
            .O(N__70489),
            .I(N__70486));
    LocalMux I__11472 (
            .O(N__70486),
            .I(shift_srl_198Z0Z_8));
    IoInMux I__11471 (
            .O(N__70483),
            .I(N__70480));
    LocalMux I__11470 (
            .O(N__70480),
            .I(N__70477));
    IoSpan4Mux I__11469 (
            .O(N__70477),
            .I(N__70474));
    Span4Mux_s3_h I__11468 (
            .O(N__70474),
            .I(N__70471));
    Span4Mux_h I__11467 (
            .O(N__70471),
            .I(N__70468));
    Span4Mux_h I__11466 (
            .O(N__70468),
            .I(N__70465));
    Odrv4 I__11465 (
            .O(N__70465),
            .I(rco_c_197));
    CascadeMux I__11464 (
            .O(N__70462),
            .I(rco_c_197_cascade_));
    IoInMux I__11463 (
            .O(N__70459),
            .I(N__70456));
    LocalMux I__11462 (
            .O(N__70456),
            .I(N__70453));
    Span4Mux_s3_h I__11461 (
            .O(N__70453),
            .I(N__70449));
    InMux I__11460 (
            .O(N__70452),
            .I(N__70446));
    Span4Mux_v I__11459 (
            .O(N__70449),
            .I(N__70443));
    LocalMux I__11458 (
            .O(N__70446),
            .I(N__70440));
    Span4Mux_h I__11457 (
            .O(N__70443),
            .I(N__70437));
    Span4Mux_v I__11456 (
            .O(N__70440),
            .I(N__70434));
    Span4Mux_h I__11455 (
            .O(N__70437),
            .I(N__70429));
    Span4Mux_h I__11454 (
            .O(N__70434),
            .I(N__70429));
    Odrv4 I__11453 (
            .O(N__70429),
            .I(rco_c_198));
    CascadeMux I__11452 (
            .O(N__70426),
            .I(N__70423));
    InMux I__11451 (
            .O(N__70423),
            .I(N__70420));
    LocalMux I__11450 (
            .O(N__70420),
            .I(N__70417));
    Span4Mux_v I__11449 (
            .O(N__70417),
            .I(N__70412));
    InMux I__11448 (
            .O(N__70416),
            .I(N__70407));
    InMux I__11447 (
            .O(N__70415),
            .I(N__70407));
    Span4Mux_h I__11446 (
            .O(N__70412),
            .I(N__70404));
    LocalMux I__11445 (
            .O(N__70407),
            .I(shift_srl_198Z0Z_15));
    Odrv4 I__11444 (
            .O(N__70404),
            .I(shift_srl_198Z0Z_15));
    InMux I__11443 (
            .O(N__70399),
            .I(N__70396));
    LocalMux I__11442 (
            .O(N__70396),
            .I(shift_srl_198Z0Z_0));
    InMux I__11441 (
            .O(N__70393),
            .I(N__70390));
    LocalMux I__11440 (
            .O(N__70390),
            .I(shift_srl_198Z0Z_1));
    InMux I__11439 (
            .O(N__70387),
            .I(N__70384));
    LocalMux I__11438 (
            .O(N__70384),
            .I(shift_srl_198Z0Z_2));
    InMux I__11437 (
            .O(N__70381),
            .I(N__70378));
    LocalMux I__11436 (
            .O(N__70378),
            .I(shift_srl_198Z0Z_3));
    InMux I__11435 (
            .O(N__70375),
            .I(N__70372));
    LocalMux I__11434 (
            .O(N__70372),
            .I(shift_srl_198Z0Z_4));
    InMux I__11433 (
            .O(N__70369),
            .I(N__70366));
    LocalMux I__11432 (
            .O(N__70366),
            .I(N__70363));
    Odrv4 I__11431 (
            .O(N__70363),
            .I(shift_srl_198Z0Z_5));
    InMux I__11430 (
            .O(N__70360),
            .I(N__70357));
    LocalMux I__11429 (
            .O(N__70357),
            .I(shift_srl_175Z0Z_5));
    InMux I__11428 (
            .O(N__70354),
            .I(N__70351));
    LocalMux I__11427 (
            .O(N__70351),
            .I(shift_srl_175Z0Z_6));
    InMux I__11426 (
            .O(N__70348),
            .I(N__70345));
    LocalMux I__11425 (
            .O(N__70345),
            .I(shift_srl_198Z0Z_10));
    InMux I__11424 (
            .O(N__70342),
            .I(N__70339));
    LocalMux I__11423 (
            .O(N__70339),
            .I(shift_srl_198Z0Z_11));
    InMux I__11422 (
            .O(N__70336),
            .I(N__70333));
    LocalMux I__11421 (
            .O(N__70333),
            .I(shift_srl_198Z0Z_12));
    InMux I__11420 (
            .O(N__70330),
            .I(N__70327));
    LocalMux I__11419 (
            .O(N__70327),
            .I(shift_srl_198Z0Z_13));
    InMux I__11418 (
            .O(N__70324),
            .I(N__70321));
    LocalMux I__11417 (
            .O(N__70321),
            .I(shift_srl_198Z0Z_14));
    InMux I__11416 (
            .O(N__70318),
            .I(N__70315));
    LocalMux I__11415 (
            .O(N__70315),
            .I(shift_srl_198Z0Z_9));
    InMux I__11414 (
            .O(N__70312),
            .I(N__70309));
    LocalMux I__11413 (
            .O(N__70309),
            .I(shift_srl_194Z0Z_5));
    InMux I__11412 (
            .O(N__70306),
            .I(N__70303));
    LocalMux I__11411 (
            .O(N__70303),
            .I(shift_srl_194Z0Z_6));
    InMux I__11410 (
            .O(N__70300),
            .I(N__70297));
    LocalMux I__11409 (
            .O(N__70297),
            .I(shift_srl_194Z0Z_7));
    InMux I__11408 (
            .O(N__70294),
            .I(N__70291));
    LocalMux I__11407 (
            .O(N__70291),
            .I(shift_srl_194Z0Z_8));
    InMux I__11406 (
            .O(N__70288),
            .I(N__70285));
    LocalMux I__11405 (
            .O(N__70285),
            .I(shift_srl_175Z0Z_0));
    InMux I__11404 (
            .O(N__70282),
            .I(N__70279));
    LocalMux I__11403 (
            .O(N__70279),
            .I(shift_srl_175Z0Z_1));
    InMux I__11402 (
            .O(N__70276),
            .I(N__70273));
    LocalMux I__11401 (
            .O(N__70273),
            .I(shift_srl_175Z0Z_2));
    InMux I__11400 (
            .O(N__70270),
            .I(N__70267));
    LocalMux I__11399 (
            .O(N__70267),
            .I(shift_srl_175Z0Z_3));
    InMux I__11398 (
            .O(N__70264),
            .I(N__70261));
    LocalMux I__11397 (
            .O(N__70261),
            .I(shift_srl_175Z0Z_4));
    InMux I__11396 (
            .O(N__70258),
            .I(N__70255));
    LocalMux I__11395 (
            .O(N__70255),
            .I(shift_srl_194Z0Z_11));
    InMux I__11394 (
            .O(N__70252),
            .I(N__70249));
    LocalMux I__11393 (
            .O(N__70249),
            .I(shift_srl_194Z0Z_12));
    InMux I__11392 (
            .O(N__70246),
            .I(N__70243));
    LocalMux I__11391 (
            .O(N__70243),
            .I(shift_srl_194Z0Z_13));
    InMux I__11390 (
            .O(N__70240),
            .I(N__70237));
    LocalMux I__11389 (
            .O(N__70237),
            .I(shift_srl_194Z0Z_14));
    InMux I__11388 (
            .O(N__70234),
            .I(N__70231));
    LocalMux I__11387 (
            .O(N__70231),
            .I(shift_srl_194Z0Z_9));
    InMux I__11386 (
            .O(N__70228),
            .I(N__70225));
    LocalMux I__11385 (
            .O(N__70225),
            .I(N__70222));
    Odrv12 I__11384 (
            .O(N__70222),
            .I(shift_srl_194Z0Z_1));
    InMux I__11383 (
            .O(N__70219),
            .I(N__70216));
    LocalMux I__11382 (
            .O(N__70216),
            .I(shift_srl_194Z0Z_2));
    InMux I__11381 (
            .O(N__70213),
            .I(N__70210));
    LocalMux I__11380 (
            .O(N__70210),
            .I(shift_srl_194Z0Z_3));
    InMux I__11379 (
            .O(N__70207),
            .I(N__70204));
    LocalMux I__11378 (
            .O(N__70204),
            .I(shift_srl_194Z0Z_4));
    InMux I__11377 (
            .O(N__70201),
            .I(N__70198));
    LocalMux I__11376 (
            .O(N__70198),
            .I(shift_srl_187Z0Z_10));
    InMux I__11375 (
            .O(N__70195),
            .I(N__70192));
    LocalMux I__11374 (
            .O(N__70192),
            .I(shift_srl_187Z0Z_11));
    InMux I__11373 (
            .O(N__70189),
            .I(N__70186));
    LocalMux I__11372 (
            .O(N__70186),
            .I(shift_srl_187Z0Z_12));
    InMux I__11371 (
            .O(N__70183),
            .I(N__70180));
    LocalMux I__11370 (
            .O(N__70180),
            .I(shift_srl_187Z0Z_13));
    InMux I__11369 (
            .O(N__70177),
            .I(N__70174));
    LocalMux I__11368 (
            .O(N__70174),
            .I(shift_srl_187Z0Z_14));
    InMux I__11367 (
            .O(N__70171),
            .I(N__70168));
    LocalMux I__11366 (
            .O(N__70168),
            .I(shift_srl_187Z0Z_9));
    InMux I__11365 (
            .O(N__70165),
            .I(N__70162));
    LocalMux I__11364 (
            .O(N__70162),
            .I(shift_srl_187Z0Z_7));
    InMux I__11363 (
            .O(N__70159),
            .I(N__70156));
    LocalMux I__11362 (
            .O(N__70156),
            .I(shift_srl_187Z0Z_8));
    CEMux I__11361 (
            .O(N__70153),
            .I(N__70150));
    LocalMux I__11360 (
            .O(N__70150),
            .I(N__70146));
    CEMux I__11359 (
            .O(N__70149),
            .I(N__70143));
    Span4Mux_v I__11358 (
            .O(N__70146),
            .I(N__70140));
    LocalMux I__11357 (
            .O(N__70143),
            .I(N__70137));
    Span4Mux_h I__11356 (
            .O(N__70140),
            .I(N__70134));
    Span4Mux_h I__11355 (
            .O(N__70137),
            .I(N__70131));
    Odrv4 I__11354 (
            .O(N__70134),
            .I(clk_en_187));
    Odrv4 I__11353 (
            .O(N__70131),
            .I(clk_en_187));
    InMux I__11352 (
            .O(N__70126),
            .I(N__70123));
    LocalMux I__11351 (
            .O(N__70123),
            .I(shift_srl_194Z0Z_10));
    InMux I__11350 (
            .O(N__70120),
            .I(N__70117));
    LocalMux I__11349 (
            .O(N__70117),
            .I(shift_srl_156Z0Z_7));
    InMux I__11348 (
            .O(N__70114),
            .I(N__70111));
    LocalMux I__11347 (
            .O(N__70111),
            .I(shift_srl_156Z0Z_8));
    CEMux I__11346 (
            .O(N__70108),
            .I(N__70104));
    CEMux I__11345 (
            .O(N__70107),
            .I(N__70101));
    LocalMux I__11344 (
            .O(N__70104),
            .I(N__70096));
    LocalMux I__11343 (
            .O(N__70101),
            .I(N__70096));
    Odrv4 I__11342 (
            .O(N__70096),
            .I(clk_en_156));
    InMux I__11341 (
            .O(N__70093),
            .I(N__70090));
    LocalMux I__11340 (
            .O(N__70090),
            .I(N__70087));
    Span4Mux_h I__11339 (
            .O(N__70087),
            .I(N__70084));
    Odrv4 I__11338 (
            .O(N__70084),
            .I(g0_15));
    CascadeMux I__11337 (
            .O(N__70081),
            .I(rco_int_0_a3_0_a2_0_183_cascade_));
    CascadeMux I__11336 (
            .O(N__70078),
            .I(clk_en_0_a2_0_a2_1_187_cascade_));
    InMux I__11335 (
            .O(N__70075),
            .I(N__70072));
    LocalMux I__11334 (
            .O(N__70072),
            .I(clk_en_0_a2_0_a2_sx_187));
    CascadeMux I__11333 (
            .O(N__70069),
            .I(N__70066));
    InMux I__11332 (
            .O(N__70066),
            .I(N__70061));
    InMux I__11331 (
            .O(N__70065),
            .I(N__70056));
    InMux I__11330 (
            .O(N__70064),
            .I(N__70056));
    LocalMux I__11329 (
            .O(N__70061),
            .I(shift_srl_183Z0Z_15));
    LocalMux I__11328 (
            .O(N__70056),
            .I(shift_srl_183Z0Z_15));
    InMux I__11327 (
            .O(N__70051),
            .I(N__70048));
    LocalMux I__11326 (
            .O(N__70048),
            .I(shift_srl_183Z0Z_0));
    CEMux I__11325 (
            .O(N__70045),
            .I(N__70041));
    CEMux I__11324 (
            .O(N__70044),
            .I(N__70038));
    LocalMux I__11323 (
            .O(N__70041),
            .I(N__70035));
    LocalMux I__11322 (
            .O(N__70038),
            .I(N__70032));
    Span4Mux_h I__11321 (
            .O(N__70035),
            .I(N__70029));
    Span4Mux_h I__11320 (
            .O(N__70032),
            .I(N__70026));
    Odrv4 I__11319 (
            .O(N__70029),
            .I(clk_en_158));
    Odrv4 I__11318 (
            .O(N__70026),
            .I(clk_en_158));
    InMux I__11317 (
            .O(N__70021),
            .I(N__70018));
    LocalMux I__11316 (
            .O(N__70018),
            .I(shift_srl_156Z0Z_10));
    InMux I__11315 (
            .O(N__70015),
            .I(N__70012));
    LocalMux I__11314 (
            .O(N__70012),
            .I(shift_srl_156Z0Z_11));
    InMux I__11313 (
            .O(N__70009),
            .I(N__70006));
    LocalMux I__11312 (
            .O(N__70006),
            .I(shift_srl_156Z0Z_12));
    InMux I__11311 (
            .O(N__70003),
            .I(N__70000));
    LocalMux I__11310 (
            .O(N__70000),
            .I(shift_srl_156Z0Z_13));
    InMux I__11309 (
            .O(N__69997),
            .I(N__69994));
    LocalMux I__11308 (
            .O(N__69994),
            .I(shift_srl_156Z0Z_14));
    InMux I__11307 (
            .O(N__69991),
            .I(N__69988));
    LocalMux I__11306 (
            .O(N__69988),
            .I(shift_srl_156Z0Z_9));
    InMux I__11305 (
            .O(N__69985),
            .I(N__69982));
    LocalMux I__11304 (
            .O(N__69982),
            .I(shift_srl_158Z0Z_13));
    InMux I__11303 (
            .O(N__69979),
            .I(N__69976));
    LocalMux I__11302 (
            .O(N__69976),
            .I(shift_srl_158Z0Z_14));
    InMux I__11301 (
            .O(N__69973),
            .I(N__69970));
    LocalMux I__11300 (
            .O(N__69970),
            .I(shift_srl_158Z0Z_9));
    InMux I__11299 (
            .O(N__69967),
            .I(N__69964));
    LocalMux I__11298 (
            .O(N__69964),
            .I(shift_srl_158Z0Z_7));
    InMux I__11297 (
            .O(N__69961),
            .I(N__69958));
    LocalMux I__11296 (
            .O(N__69958),
            .I(shift_srl_158Z0Z_8));
    IoInMux I__11295 (
            .O(N__69955),
            .I(N__69952));
    LocalMux I__11294 (
            .O(N__69952),
            .I(N__69949));
    IoSpan4Mux I__11293 (
            .O(N__69949),
            .I(N__69946));
    Span4Mux_s1_h I__11292 (
            .O(N__69946),
            .I(N__69943));
    Sp12to4 I__11291 (
            .O(N__69943),
            .I(N__69940));
    Span12Mux_v I__11290 (
            .O(N__69940),
            .I(N__69937));
    Span12Mux_h I__11289 (
            .O(N__69937),
            .I(N__69934));
    Odrv12 I__11288 (
            .O(N__69934),
            .I(rco_c_158));
    IoInMux I__11287 (
            .O(N__69931),
            .I(N__69928));
    LocalMux I__11286 (
            .O(N__69928),
            .I(N__69925));
    Span4Mux_s0_h I__11285 (
            .O(N__69925),
            .I(N__69922));
    Sp12to4 I__11284 (
            .O(N__69922),
            .I(N__69919));
    Span12Mux_v I__11283 (
            .O(N__69919),
            .I(N__69916));
    Span12Mux_h I__11282 (
            .O(N__69916),
            .I(N__69913));
    Odrv12 I__11281 (
            .O(N__69913),
            .I(rco_c_157));
    InMux I__11280 (
            .O(N__69910),
            .I(N__69907));
    LocalMux I__11279 (
            .O(N__69907),
            .I(N__69904));
    Span4Mux_h I__11278 (
            .O(N__69904),
            .I(N__69901));
    Span4Mux_v I__11277 (
            .O(N__69901),
            .I(N__69898));
    Span4Mux_v I__11276 (
            .O(N__69898),
            .I(N__69895));
    Odrv4 I__11275 (
            .O(N__69895),
            .I(rco_int_0_a2_0_a2_sx_1_153));
    CascadeMux I__11274 (
            .O(N__69892),
            .I(rco_c_153_cascade_));
    CEMux I__11273 (
            .O(N__69889),
            .I(N__69885));
    CEMux I__11272 (
            .O(N__69888),
            .I(N__69882));
    LocalMux I__11271 (
            .O(N__69885),
            .I(N__69879));
    LocalMux I__11270 (
            .O(N__69882),
            .I(N__69876));
    Span4Mux_h I__11269 (
            .O(N__69879),
            .I(N__69873));
    Span4Mux_h I__11268 (
            .O(N__69876),
            .I(N__69870));
    Odrv4 I__11267 (
            .O(N__69873),
            .I(clk_en_162));
    Odrv4 I__11266 (
            .O(N__69870),
            .I(clk_en_162));
    InMux I__11265 (
            .O(N__69865),
            .I(N__69862));
    LocalMux I__11264 (
            .O(N__69862),
            .I(N__69857));
    InMux I__11263 (
            .O(N__69861),
            .I(N__69852));
    InMux I__11262 (
            .O(N__69860),
            .I(N__69852));
    Span4Mux_h I__11261 (
            .O(N__69857),
            .I(N__69849));
    LocalMux I__11260 (
            .O(N__69852),
            .I(N__69846));
    Span4Mux_h I__11259 (
            .O(N__69849),
            .I(N__69843));
    Span12Mux_h I__11258 (
            .O(N__69846),
            .I(N__69839));
    Span4Mux_v I__11257 (
            .O(N__69843),
            .I(N__69836));
    InMux I__11256 (
            .O(N__69842),
            .I(N__69833));
    Odrv12 I__11255 (
            .O(N__69839),
            .I(shift_srl_160_RNIFA2R1Z0Z_15));
    Odrv4 I__11254 (
            .O(N__69836),
            .I(shift_srl_160_RNIFA2R1Z0Z_15));
    LocalMux I__11253 (
            .O(N__69833),
            .I(shift_srl_160_RNIFA2R1Z0Z_15));
    InMux I__11252 (
            .O(N__69826),
            .I(N__69823));
    LocalMux I__11251 (
            .O(N__69823),
            .I(shift_srl_38Z0Z_10));
    InMux I__11250 (
            .O(N__69820),
            .I(N__69817));
    LocalMux I__11249 (
            .O(N__69817),
            .I(shift_srl_38Z0Z_11));
    InMux I__11248 (
            .O(N__69814),
            .I(N__69811));
    LocalMux I__11247 (
            .O(N__69811),
            .I(shift_srl_38Z0Z_12));
    InMux I__11246 (
            .O(N__69808),
            .I(N__69805));
    LocalMux I__11245 (
            .O(N__69805),
            .I(shift_srl_38Z0Z_14));
    InMux I__11244 (
            .O(N__69802),
            .I(N__69799));
    LocalMux I__11243 (
            .O(N__69799),
            .I(shift_srl_38Z0Z_9));
    InMux I__11242 (
            .O(N__69796),
            .I(N__69793));
    LocalMux I__11241 (
            .O(N__69793),
            .I(shift_srl_38Z0Z_7));
    InMux I__11240 (
            .O(N__69790),
            .I(N__69787));
    LocalMux I__11239 (
            .O(N__69787),
            .I(shift_srl_38Z0Z_8));
    CEMux I__11238 (
            .O(N__69784),
            .I(N__69781));
    LocalMux I__11237 (
            .O(N__69781),
            .I(N__69777));
    CEMux I__11236 (
            .O(N__69780),
            .I(N__69774));
    Span4Mux_h I__11235 (
            .O(N__69777),
            .I(N__69768));
    LocalMux I__11234 (
            .O(N__69774),
            .I(N__69768));
    CEMux I__11233 (
            .O(N__69773),
            .I(N__69765));
    Span4Mux_h I__11232 (
            .O(N__69768),
            .I(N__69762));
    LocalMux I__11231 (
            .O(N__69765),
            .I(N__69759));
    Odrv4 I__11230 (
            .O(N__69762),
            .I(clk_en_38));
    Odrv4 I__11229 (
            .O(N__69759),
            .I(clk_en_38));
    InMux I__11228 (
            .O(N__69754),
            .I(N__69751));
    LocalMux I__11227 (
            .O(N__69751),
            .I(shift_srl_158Z0Z_10));
    InMux I__11226 (
            .O(N__69748),
            .I(N__69745));
    LocalMux I__11225 (
            .O(N__69745),
            .I(shift_srl_158Z0Z_11));
    InMux I__11224 (
            .O(N__69742),
            .I(N__69739));
    LocalMux I__11223 (
            .O(N__69739),
            .I(shift_srl_158Z0Z_12));
    InMux I__11222 (
            .O(N__69736),
            .I(N__69733));
    LocalMux I__11221 (
            .O(N__69733),
            .I(shift_srl_38Z0Z_0));
    InMux I__11220 (
            .O(N__69730),
            .I(N__69727));
    LocalMux I__11219 (
            .O(N__69727),
            .I(shift_srl_38Z0Z_1));
    InMux I__11218 (
            .O(N__69724),
            .I(N__69721));
    LocalMux I__11217 (
            .O(N__69721),
            .I(shift_srl_38Z0Z_2));
    InMux I__11216 (
            .O(N__69718),
            .I(N__69715));
    LocalMux I__11215 (
            .O(N__69715),
            .I(shift_srl_38Z0Z_3));
    InMux I__11214 (
            .O(N__69712),
            .I(N__69709));
    LocalMux I__11213 (
            .O(N__69709),
            .I(shift_srl_38Z0Z_4));
    InMux I__11212 (
            .O(N__69706),
            .I(N__69703));
    LocalMux I__11211 (
            .O(N__69703),
            .I(shift_srl_38Z0Z_5));
    InMux I__11210 (
            .O(N__69700),
            .I(N__69697));
    LocalMux I__11209 (
            .O(N__69697),
            .I(shift_srl_38Z0Z_6));
    InMux I__11208 (
            .O(N__69694),
            .I(N__69691));
    LocalMux I__11207 (
            .O(N__69691),
            .I(N__69688));
    Span12Mux_h I__11206 (
            .O(N__69688),
            .I(N__69685));
    Span12Mux_v I__11205 (
            .O(N__69685),
            .I(N__69682));
    Odrv12 I__11204 (
            .O(N__69682),
            .I(shift_srl_40Z0Z_9));
    InMux I__11203 (
            .O(N__69679),
            .I(N__69676));
    LocalMux I__11202 (
            .O(N__69676),
            .I(shift_srl_40Z0Z_10));
    CEMux I__11201 (
            .O(N__69673),
            .I(N__69664));
    CEMux I__11200 (
            .O(N__69672),
            .I(N__69664));
    CEMux I__11199 (
            .O(N__69671),
            .I(N__69664));
    GlobalMux I__11198 (
            .O(N__69664),
            .I(N__69661));
    gio2CtrlBuf I__11197 (
            .O(N__69661),
            .I(clk_en_g_40));
    InMux I__11196 (
            .O(N__69658),
            .I(N__69655));
    LocalMux I__11195 (
            .O(N__69655),
            .I(rco_int_0_a2_0_a2_out_2));
    IoInMux I__11194 (
            .O(N__69652),
            .I(N__69649));
    LocalMux I__11193 (
            .O(N__69649),
            .I(N__69646));
    IoSpan4Mux I__11192 (
            .O(N__69646),
            .I(N__69643));
    Span4Mux_s2_v I__11191 (
            .O(N__69643),
            .I(N__69640));
    Sp12to4 I__11190 (
            .O(N__69640),
            .I(N__69637));
    Span12Mux_s8_v I__11189 (
            .O(N__69637),
            .I(N__69634));
    Odrv12 I__11188 (
            .O(N__69634),
            .I(rco_c_30));
    InMux I__11187 (
            .O(N__69631),
            .I(N__69628));
    LocalMux I__11186 (
            .O(N__69628),
            .I(shift_srl_30Z0Z_0));
    InMux I__11185 (
            .O(N__69625),
            .I(N__69622));
    LocalMux I__11184 (
            .O(N__69622),
            .I(shift_srl_30Z0Z_1));
    InMux I__11183 (
            .O(N__69619),
            .I(N__69616));
    LocalMux I__11182 (
            .O(N__69616),
            .I(shift_srl_30Z0Z_2));
    InMux I__11181 (
            .O(N__69613),
            .I(N__69610));
    LocalMux I__11180 (
            .O(N__69610),
            .I(shift_srl_30Z0Z_3));
    InMux I__11179 (
            .O(N__69607),
            .I(N__69604));
    LocalMux I__11178 (
            .O(N__69604),
            .I(shift_srl_30Z0Z_4));
    InMux I__11177 (
            .O(N__69601),
            .I(N__69598));
    LocalMux I__11176 (
            .O(N__69598),
            .I(shift_srl_30Z0Z_5));
    IoInMux I__11175 (
            .O(N__69595),
            .I(N__69592));
    LocalMux I__11174 (
            .O(N__69592),
            .I(N__69589));
    IoSpan4Mux I__11173 (
            .O(N__69589),
            .I(N__69586));
    IoSpan4Mux I__11172 (
            .O(N__69586),
            .I(N__69583));
    Sp12to4 I__11171 (
            .O(N__69583),
            .I(N__69580));
    Span12Mux_s7_v I__11170 (
            .O(N__69580),
            .I(N__69577));
    Odrv12 I__11169 (
            .O(N__69577),
            .I(rco_c_34));
    InMux I__11168 (
            .O(N__69574),
            .I(N__69571));
    LocalMux I__11167 (
            .O(N__69571),
            .I(N__69568));
    Span4Mux_v I__11166 (
            .O(N__69568),
            .I(N__69565));
    Span4Mux_v I__11165 (
            .O(N__69565),
            .I(N__69562));
    Odrv4 I__11164 (
            .O(N__69562),
            .I(shift_srl_95Z0Z_13));
    InMux I__11163 (
            .O(N__69559),
            .I(N__69556));
    LocalMux I__11162 (
            .O(N__69556),
            .I(shift_srl_95Z0Z_14));
    CEMux I__11161 (
            .O(N__69553),
            .I(N__69549));
    CEMux I__11160 (
            .O(N__69552),
            .I(N__69545));
    LocalMux I__11159 (
            .O(N__69549),
            .I(N__69542));
    CEMux I__11158 (
            .O(N__69548),
            .I(N__69539));
    LocalMux I__11157 (
            .O(N__69545),
            .I(N__69536));
    Span4Mux_v I__11156 (
            .O(N__69542),
            .I(N__69533));
    LocalMux I__11155 (
            .O(N__69539),
            .I(N__69530));
    Span4Mux_v I__11154 (
            .O(N__69536),
            .I(N__69527));
    Odrv4 I__11153 (
            .O(N__69533),
            .I(clk_en_95));
    Odrv4 I__11152 (
            .O(N__69530),
            .I(clk_en_95));
    Odrv4 I__11151 (
            .O(N__69527),
            .I(clk_en_95));
    InMux I__11150 (
            .O(N__69520),
            .I(N__69516));
    InMux I__11149 (
            .O(N__69519),
            .I(N__69513));
    LocalMux I__11148 (
            .O(N__69516),
            .I(N__69510));
    LocalMux I__11147 (
            .O(N__69513),
            .I(N__69505));
    Span12Mux_v I__11146 (
            .O(N__69510),
            .I(N__69505));
    Odrv12 I__11145 (
            .O(N__69505),
            .I(shift_srl_93Z0Z_15));
    InMux I__11144 (
            .O(N__69502),
            .I(N__69499));
    LocalMux I__11143 (
            .O(N__69499),
            .I(shift_srl_40_fastZ0Z_15));
    InMux I__11142 (
            .O(N__69496),
            .I(N__69490));
    InMux I__11141 (
            .O(N__69495),
            .I(N__69490));
    LocalMux I__11140 (
            .O(N__69490),
            .I(shift_srl_40Z0Z_14));
    InMux I__11139 (
            .O(N__69487),
            .I(N__69484));
    LocalMux I__11138 (
            .O(N__69484),
            .I(shift_srl_40Z0Z_13));
    InMux I__11137 (
            .O(N__69481),
            .I(N__69478));
    LocalMux I__11136 (
            .O(N__69478),
            .I(shift_srl_40Z0Z_12));
    InMux I__11135 (
            .O(N__69475),
            .I(N__69472));
    LocalMux I__11134 (
            .O(N__69472),
            .I(shift_srl_40Z0Z_11));
    InMux I__11133 (
            .O(N__69469),
            .I(N__69466));
    LocalMux I__11132 (
            .O(N__69466),
            .I(shift_srl_48Z0Z_4));
    InMux I__11131 (
            .O(N__69463),
            .I(N__69460));
    LocalMux I__11130 (
            .O(N__69460),
            .I(shift_srl_48Z0Z_5));
    CascadeMux I__11129 (
            .O(N__69457),
            .I(shift_srl_94_RNI2F961Z0Z_15_cascade_));
    CascadeMux I__11128 (
            .O(N__69454),
            .I(N__69451));
    InMux I__11127 (
            .O(N__69451),
            .I(N__69441));
    InMux I__11126 (
            .O(N__69450),
            .I(N__69441));
    InMux I__11125 (
            .O(N__69449),
            .I(N__69438));
    InMux I__11124 (
            .O(N__69448),
            .I(N__69435));
    InMux I__11123 (
            .O(N__69447),
            .I(N__69430));
    InMux I__11122 (
            .O(N__69446),
            .I(N__69430));
    LocalMux I__11121 (
            .O(N__69441),
            .I(N__69425));
    LocalMux I__11120 (
            .O(N__69438),
            .I(N__69425));
    LocalMux I__11119 (
            .O(N__69435),
            .I(shift_srl_96Z0Z_15));
    LocalMux I__11118 (
            .O(N__69430),
            .I(shift_srl_96Z0Z_15));
    Odrv12 I__11117 (
            .O(N__69425),
            .I(shift_srl_96Z0Z_15));
    InMux I__11116 (
            .O(N__69418),
            .I(N__69414));
    InMux I__11115 (
            .O(N__69417),
            .I(N__69411));
    LocalMux I__11114 (
            .O(N__69414),
            .I(N__69408));
    LocalMux I__11113 (
            .O(N__69411),
            .I(shift_srl_98Z0Z_15));
    Odrv4 I__11112 (
            .O(N__69408),
            .I(shift_srl_98Z0Z_15));
    InMux I__11111 (
            .O(N__69403),
            .I(N__69400));
    LocalMux I__11110 (
            .O(N__69400),
            .I(shift_srl_98_RNIA7Q31Z0Z_15));
    InMux I__11109 (
            .O(N__69397),
            .I(N__69394));
    LocalMux I__11108 (
            .O(N__69394),
            .I(rco_int_0_a2_0_a2_99_m6_0_a2_1));
    CascadeMux I__11107 (
            .O(N__69391),
            .I(rco_int_0_a2_0_a2_99_m6_0_a2_9_1_cascade_));
    InMux I__11106 (
            .O(N__69388),
            .I(N__69385));
    LocalMux I__11105 (
            .O(N__69385),
            .I(rco_int_0_a2_0_a2_99_m6_0_a2_9_sx));
    InMux I__11104 (
            .O(N__69382),
            .I(N__69378));
    InMux I__11103 (
            .O(N__69381),
            .I(N__69375));
    LocalMux I__11102 (
            .O(N__69378),
            .I(N__69370));
    LocalMux I__11101 (
            .O(N__69375),
            .I(N__69370));
    Span4Mux_v I__11100 (
            .O(N__69370),
            .I(N__69366));
    InMux I__11099 (
            .O(N__69369),
            .I(N__69363));
    Odrv4 I__11098 (
            .O(N__69366),
            .I(shift_srl_95Z0Z_15));
    LocalMux I__11097 (
            .O(N__69363),
            .I(shift_srl_95Z0Z_15));
    InMux I__11096 (
            .O(N__69358),
            .I(N__69355));
    LocalMux I__11095 (
            .O(N__69355),
            .I(shift_srl_44Z0Z_2));
    InMux I__11094 (
            .O(N__69352),
            .I(N__69349));
    LocalMux I__11093 (
            .O(N__69349),
            .I(shift_srl_44Z0Z_3));
    InMux I__11092 (
            .O(N__69346),
            .I(N__69343));
    LocalMux I__11091 (
            .O(N__69343),
            .I(shift_srl_44Z0Z_4));
    InMux I__11090 (
            .O(N__69340),
            .I(N__69337));
    LocalMux I__11089 (
            .O(N__69337),
            .I(shift_srl_44Z0Z_5));
    InMux I__11088 (
            .O(N__69334),
            .I(N__69331));
    LocalMux I__11087 (
            .O(N__69331),
            .I(shift_srl_44Z0Z_6));
    InMux I__11086 (
            .O(N__69328),
            .I(N__69325));
    LocalMux I__11085 (
            .O(N__69325),
            .I(shift_srl_48Z0Z_0));
    InMux I__11084 (
            .O(N__69322),
            .I(N__69319));
    LocalMux I__11083 (
            .O(N__69319),
            .I(shift_srl_48Z0Z_1));
    InMux I__11082 (
            .O(N__69316),
            .I(N__69313));
    LocalMux I__11081 (
            .O(N__69313),
            .I(shift_srl_48Z0Z_2));
    InMux I__11080 (
            .O(N__69310),
            .I(N__69307));
    LocalMux I__11079 (
            .O(N__69307),
            .I(shift_srl_48Z0Z_3));
    InMux I__11078 (
            .O(N__69304),
            .I(N__69301));
    LocalMux I__11077 (
            .O(N__69301),
            .I(N__69298));
    Span4Mux_h I__11076 (
            .O(N__69298),
            .I(N__69295));
    Span4Mux_h I__11075 (
            .O(N__69295),
            .I(N__69291));
    InMux I__11074 (
            .O(N__69294),
            .I(N__69288));
    Span4Mux_h I__11073 (
            .O(N__69291),
            .I(N__69285));
    LocalMux I__11072 (
            .O(N__69288),
            .I(N__69282));
    Odrv4 I__11071 (
            .O(N__69285),
            .I(N_4016_i_0_a2_1));
    Odrv12 I__11070 (
            .O(N__69282),
            .I(N_4016_i_0_a2_1));
    CascadeMux I__11069 (
            .O(N__69277),
            .I(N__69273));
    InMux I__11068 (
            .O(N__69276),
            .I(N__69269));
    InMux I__11067 (
            .O(N__69273),
            .I(N__69266));
    InMux I__11066 (
            .O(N__69272),
            .I(N__69263));
    LocalMux I__11065 (
            .O(N__69269),
            .I(N__69260));
    LocalMux I__11064 (
            .O(N__69266),
            .I(N__69257));
    LocalMux I__11063 (
            .O(N__69263),
            .I(N__69254));
    Span4Mux_h I__11062 (
            .O(N__69260),
            .I(N__69251));
    Span12Mux_h I__11061 (
            .O(N__69257),
            .I(N__69248));
    Span4Mux_v I__11060 (
            .O(N__69254),
            .I(N__69243));
    Span4Mux_v I__11059 (
            .O(N__69251),
            .I(N__69243));
    Odrv12 I__11058 (
            .O(N__69248),
            .I(rco_int_0_a2_21_m6_0_a2_s_7));
    Odrv4 I__11057 (
            .O(N__69243),
            .I(rco_int_0_a2_21_m6_0_a2_s_7));
    InMux I__11056 (
            .O(N__69238),
            .I(N__69235));
    LocalMux I__11055 (
            .O(N__69235),
            .I(N__69232));
    Span4Mux_h I__11054 (
            .O(N__69232),
            .I(N__69228));
    InMux I__11053 (
            .O(N__69231),
            .I(N__69224));
    Span4Mux_h I__11052 (
            .O(N__69228),
            .I(N__69221));
    InMux I__11051 (
            .O(N__69227),
            .I(N__69218));
    LocalMux I__11050 (
            .O(N__69224),
            .I(N__69215));
    Span4Mux_h I__11049 (
            .O(N__69221),
            .I(N__69212));
    LocalMux I__11048 (
            .O(N__69218),
            .I(N__69209));
    Span12Mux_v I__11047 (
            .O(N__69215),
            .I(N__69206));
    Span4Mux_h I__11046 (
            .O(N__69212),
            .I(N__69201));
    Span4Mux_h I__11045 (
            .O(N__69209),
            .I(N__69201));
    Odrv12 I__11044 (
            .O(N__69206),
            .I(rco_int_0_a2_21_m6_0_a2_s_8));
    Odrv4 I__11043 (
            .O(N__69201),
            .I(rco_int_0_a2_21_m6_0_a2_s_8));
    CascadeMux I__11042 (
            .O(N__69196),
            .I(shift_srl_23_RNI0DK37Z0Z_15_cascade_));
    IoInMux I__11041 (
            .O(N__69193),
            .I(N__69189));
    InMux I__11040 (
            .O(N__69192),
            .I(N__69185));
    LocalMux I__11039 (
            .O(N__69189),
            .I(N__69182));
    InMux I__11038 (
            .O(N__69188),
            .I(N__69179));
    LocalMux I__11037 (
            .O(N__69185),
            .I(N__69175));
    Span4Mux_s2_h I__11036 (
            .O(N__69182),
            .I(N__69172));
    LocalMux I__11035 (
            .O(N__69179),
            .I(N__69169));
    InMux I__11034 (
            .O(N__69178),
            .I(N__69166));
    Span4Mux_h I__11033 (
            .O(N__69175),
            .I(N__69163));
    Span4Mux_h I__11032 (
            .O(N__69172),
            .I(N__69160));
    Span4Mux_h I__11031 (
            .O(N__69169),
            .I(N__69157));
    LocalMux I__11030 (
            .O(N__69166),
            .I(N__69154));
    Span4Mux_h I__11029 (
            .O(N__69163),
            .I(N__69151));
    Sp12to4 I__11028 (
            .O(N__69160),
            .I(N__69148));
    Span4Mux_v I__11027 (
            .O(N__69157),
            .I(N__69143));
    Span4Mux_h I__11026 (
            .O(N__69154),
            .I(N__69143));
    Span4Mux_h I__11025 (
            .O(N__69151),
            .I(N__69140));
    Odrv12 I__11024 (
            .O(N__69148),
            .I(rco_c_9));
    Odrv4 I__11023 (
            .O(N__69143),
            .I(rco_c_9));
    Odrv4 I__11022 (
            .O(N__69140),
            .I(rco_c_9));
    CascadeMux I__11021 (
            .O(N__69133),
            .I(rco_c_41_cascade_));
    IoInMux I__11020 (
            .O(N__69130),
            .I(N__69127));
    LocalMux I__11019 (
            .O(N__69127),
            .I(N__69124));
    Span4Mux_s2_h I__11018 (
            .O(N__69124),
            .I(N__69121));
    Span4Mux_h I__11017 (
            .O(N__69121),
            .I(N__69116));
    InMux I__11016 (
            .O(N__69120),
            .I(N__69111));
    InMux I__11015 (
            .O(N__69119),
            .I(N__69111));
    Span4Mux_h I__11014 (
            .O(N__69116),
            .I(N__69106));
    LocalMux I__11013 (
            .O(N__69111),
            .I(N__69103));
    CascadeMux I__11012 (
            .O(N__69110),
            .I(N__69099));
    CascadeMux I__11011 (
            .O(N__69109),
            .I(N__69096));
    Span4Mux_h I__11010 (
            .O(N__69106),
            .I(N__69092));
    Span4Mux_v I__11009 (
            .O(N__69103),
            .I(N__69089));
    InMux I__11008 (
            .O(N__69102),
            .I(N__69080));
    InMux I__11007 (
            .O(N__69099),
            .I(N__69080));
    InMux I__11006 (
            .O(N__69096),
            .I(N__69080));
    InMux I__11005 (
            .O(N__69095),
            .I(N__69080));
    Odrv4 I__11004 (
            .O(N__69092),
            .I(rco_c_41));
    Odrv4 I__11003 (
            .O(N__69089),
            .I(rco_c_41));
    LocalMux I__11002 (
            .O(N__69080),
            .I(rco_c_41));
    CEMux I__11001 (
            .O(N__69073),
            .I(N__69069));
    CEMux I__11000 (
            .O(N__69072),
            .I(N__69066));
    LocalMux I__10999 (
            .O(N__69069),
            .I(N__69061));
    LocalMux I__10998 (
            .O(N__69066),
            .I(N__69061));
    Odrv4 I__10997 (
            .O(N__69061),
            .I(clk_en_45));
    InMux I__10996 (
            .O(N__69058),
            .I(N__69055));
    LocalMux I__10995 (
            .O(N__69055),
            .I(shift_srl_44Z0Z_0));
    InMux I__10994 (
            .O(N__69052),
            .I(N__69049));
    LocalMux I__10993 (
            .O(N__69049),
            .I(shift_srl_44Z0Z_1));
    InMux I__10992 (
            .O(N__69046),
            .I(N__69043));
    LocalMux I__10991 (
            .O(N__69043),
            .I(shift_srl_45Z0Z_10));
    InMux I__10990 (
            .O(N__69040),
            .I(N__69037));
    LocalMux I__10989 (
            .O(N__69037),
            .I(shift_srl_45Z0Z_11));
    InMux I__10988 (
            .O(N__69034),
            .I(N__69031));
    LocalMux I__10987 (
            .O(N__69031),
            .I(shift_srl_45Z0Z_12));
    InMux I__10986 (
            .O(N__69028),
            .I(N__69025));
    LocalMux I__10985 (
            .O(N__69025),
            .I(shift_srl_45Z0Z_13));
    InMux I__10984 (
            .O(N__69022),
            .I(N__69019));
    LocalMux I__10983 (
            .O(N__69019),
            .I(shift_srl_45Z0Z_14));
    InMux I__10982 (
            .O(N__69016),
            .I(N__69013));
    LocalMux I__10981 (
            .O(N__69013),
            .I(shift_srl_45Z0Z_9));
    InMux I__10980 (
            .O(N__69010),
            .I(N__69007));
    LocalMux I__10979 (
            .O(N__69007),
            .I(shift_srl_45Z0Z_7));
    InMux I__10978 (
            .O(N__69004),
            .I(N__69001));
    LocalMux I__10977 (
            .O(N__69001),
            .I(shift_srl_45Z0Z_8));
    CEMux I__10976 (
            .O(N__68998),
            .I(N__68994));
    CEMux I__10975 (
            .O(N__68997),
            .I(N__68991));
    LocalMux I__10974 (
            .O(N__68994),
            .I(N__68987));
    LocalMux I__10973 (
            .O(N__68991),
            .I(N__68984));
    CEMux I__10972 (
            .O(N__68990),
            .I(N__68981));
    Span4Mux_v I__10971 (
            .O(N__68987),
            .I(N__68976));
    Span4Mux_v I__10970 (
            .O(N__68984),
            .I(N__68976));
    LocalMux I__10969 (
            .O(N__68981),
            .I(N__68973));
    Span4Mux_h I__10968 (
            .O(N__68976),
            .I(N__68970));
    Span4Mux_h I__10967 (
            .O(N__68973),
            .I(N__68967));
    Odrv4 I__10966 (
            .O(N__68970),
            .I(clk_en_43));
    Odrv4 I__10965 (
            .O(N__68967),
            .I(clk_en_43));
    InMux I__10964 (
            .O(N__68962),
            .I(N__68959));
    LocalMux I__10963 (
            .O(N__68959),
            .I(shift_srl_96Z0Z_6));
    InMux I__10962 (
            .O(N__68956),
            .I(N__68953));
    LocalMux I__10961 (
            .O(N__68953),
            .I(shift_srl_96Z0Z_4));
    InMux I__10960 (
            .O(N__68950),
            .I(N__68947));
    LocalMux I__10959 (
            .O(N__68947),
            .I(shift_srl_96Z0Z_5));
    InMux I__10958 (
            .O(N__68944),
            .I(N__68941));
    LocalMux I__10957 (
            .O(N__68941),
            .I(shift_srl_96Z0Z_12));
    InMux I__10956 (
            .O(N__68938),
            .I(N__68935));
    LocalMux I__10955 (
            .O(N__68935),
            .I(shift_srl_96Z0Z_13));
    InMux I__10954 (
            .O(N__68932),
            .I(N__68929));
    LocalMux I__10953 (
            .O(N__68929),
            .I(shift_srl_96Z0Z_14));
    InMux I__10952 (
            .O(N__68926),
            .I(N__68923));
    LocalMux I__10951 (
            .O(N__68923),
            .I(shift_srl_96Z0Z_9));
    InMux I__10950 (
            .O(N__68920),
            .I(N__68917));
    LocalMux I__10949 (
            .O(N__68917),
            .I(shift_srl_96Z0Z_7));
    InMux I__10948 (
            .O(N__68914),
            .I(N__68911));
    LocalMux I__10947 (
            .O(N__68911),
            .I(shift_srl_96Z0Z_8));
    CEMux I__10946 (
            .O(N__68908),
            .I(N__68904));
    CEMux I__10945 (
            .O(N__68907),
            .I(N__68901));
    LocalMux I__10944 (
            .O(N__68904),
            .I(N__68898));
    LocalMux I__10943 (
            .O(N__68901),
            .I(N__68895));
    Odrv4 I__10942 (
            .O(N__68898),
            .I(clk_en_96));
    Odrv4 I__10941 (
            .O(N__68895),
            .I(clk_en_96));
    InMux I__10940 (
            .O(N__68890),
            .I(N__68887));
    LocalMux I__10939 (
            .O(N__68887),
            .I(N__68884));
    Span4Mux_v I__10938 (
            .O(N__68884),
            .I(N__68881));
    Odrv4 I__10937 (
            .O(N__68881),
            .I(shift_srl_94Z0Z_10));
    InMux I__10936 (
            .O(N__68878),
            .I(N__68875));
    LocalMux I__10935 (
            .O(N__68875),
            .I(shift_srl_94Z0Z_11));
    InMux I__10934 (
            .O(N__68872),
            .I(N__68869));
    LocalMux I__10933 (
            .O(N__68869),
            .I(shift_srl_96Z0Z_1));
    InMux I__10932 (
            .O(N__68866),
            .I(N__68863));
    LocalMux I__10931 (
            .O(N__68863),
            .I(shift_srl_96Z0Z_2));
    InMux I__10930 (
            .O(N__68860),
            .I(N__68857));
    LocalMux I__10929 (
            .O(N__68857),
            .I(shift_srl_96Z0Z_3));
    InMux I__10928 (
            .O(N__68854),
            .I(N__68851));
    LocalMux I__10927 (
            .O(N__68851),
            .I(shift_srl_96Z0Z_0));
    InMux I__10926 (
            .O(N__68848),
            .I(N__68845));
    LocalMux I__10925 (
            .O(N__68845),
            .I(shift_srl_96Z0Z_10));
    InMux I__10924 (
            .O(N__68842),
            .I(N__68839));
    LocalMux I__10923 (
            .O(N__68839),
            .I(shift_srl_96Z0Z_11));
    InMux I__10922 (
            .O(N__68836),
            .I(N__68833));
    LocalMux I__10921 (
            .O(N__68833),
            .I(shift_srl_97Z0Z_14));
    InMux I__10920 (
            .O(N__68830),
            .I(N__68827));
    LocalMux I__10919 (
            .O(N__68827),
            .I(shift_srl_97Z0Z_9));
    InMux I__10918 (
            .O(N__68824),
            .I(N__68821));
    LocalMux I__10917 (
            .O(N__68821),
            .I(shift_srl_97Z0Z_8));
    CascadeMux I__10916 (
            .O(N__68818),
            .I(shift_srl_95_RNIHJ49Z0Z_15_cascade_));
    IoInMux I__10915 (
            .O(N__68815),
            .I(N__68812));
    LocalMux I__10914 (
            .O(N__68812),
            .I(N__68809));
    IoSpan4Mux I__10913 (
            .O(N__68809),
            .I(N__68806));
    Span4Mux_s2_v I__10912 (
            .O(N__68806),
            .I(N__68803));
    Odrv4 I__10911 (
            .O(N__68803),
            .I(rco_c_96));
    InMux I__10910 (
            .O(N__68800),
            .I(N__68797));
    LocalMux I__10909 (
            .O(N__68797),
            .I(shift_srl_94Z0Z_14));
    InMux I__10908 (
            .O(N__68794),
            .I(N__68791));
    LocalMux I__10907 (
            .O(N__68791),
            .I(shift_srl_94Z0Z_13));
    InMux I__10906 (
            .O(N__68788),
            .I(N__68785));
    LocalMux I__10905 (
            .O(N__68785),
            .I(shift_srl_94Z0Z_12));
    InMux I__10904 (
            .O(N__68782),
            .I(N__68779));
    LocalMux I__10903 (
            .O(N__68779),
            .I(shift_srl_46Z0Z_3));
    InMux I__10902 (
            .O(N__68776),
            .I(N__68773));
    LocalMux I__10901 (
            .O(N__68773),
            .I(shift_srl_46Z0Z_8));
    InMux I__10900 (
            .O(N__68770),
            .I(N__68767));
    LocalMux I__10899 (
            .O(N__68767),
            .I(shift_srl_46Z0Z_9));
    InMux I__10898 (
            .O(N__68764),
            .I(N__68761));
    LocalMux I__10897 (
            .O(N__68761),
            .I(shift_srl_46Z0Z_1));
    InMux I__10896 (
            .O(N__68758),
            .I(N__68755));
    LocalMux I__10895 (
            .O(N__68755),
            .I(shift_srl_46Z0Z_2));
    InMux I__10894 (
            .O(N__68752),
            .I(N__68749));
    LocalMux I__10893 (
            .O(N__68749),
            .I(shift_srl_97Z0Z_10));
    InMux I__10892 (
            .O(N__68746),
            .I(N__68743));
    LocalMux I__10891 (
            .O(N__68743),
            .I(shift_srl_97Z0Z_11));
    InMux I__10890 (
            .O(N__68740),
            .I(N__68737));
    LocalMux I__10889 (
            .O(N__68737),
            .I(shift_srl_97Z0Z_12));
    InMux I__10888 (
            .O(N__68734),
            .I(N__68731));
    LocalMux I__10887 (
            .O(N__68731),
            .I(shift_srl_97Z0Z_13));
    InMux I__10886 (
            .O(N__68728),
            .I(N__68725));
    LocalMux I__10885 (
            .O(N__68725),
            .I(shift_srl_93Z0Z_11));
    InMux I__10884 (
            .O(N__68722),
            .I(N__68719));
    LocalMux I__10883 (
            .O(N__68719),
            .I(shift_srl_93Z0Z_12));
    InMux I__10882 (
            .O(N__68716),
            .I(N__68713));
    LocalMux I__10881 (
            .O(N__68713),
            .I(shift_srl_93Z0Z_13));
    InMux I__10880 (
            .O(N__68710),
            .I(N__68707));
    LocalMux I__10879 (
            .O(N__68707),
            .I(shift_srl_93Z0Z_14));
    InMux I__10878 (
            .O(N__68704),
            .I(N__68701));
    LocalMux I__10877 (
            .O(N__68701),
            .I(shift_srl_93Z0Z_9));
    InMux I__10876 (
            .O(N__68698),
            .I(N__68695));
    LocalMux I__10875 (
            .O(N__68695),
            .I(shift_srl_46Z0Z_0));
    InMux I__10874 (
            .O(N__68692),
            .I(N__68689));
    LocalMux I__10873 (
            .O(N__68689),
            .I(shift_srl_93Z0Z_5));
    InMux I__10872 (
            .O(N__68686),
            .I(N__68683));
    LocalMux I__10871 (
            .O(N__68683),
            .I(N__68677));
    InMux I__10870 (
            .O(N__68682),
            .I(N__68672));
    InMux I__10869 (
            .O(N__68681),
            .I(N__68672));
    InMux I__10868 (
            .O(N__68680),
            .I(N__68668));
    Span4Mux_h I__10867 (
            .O(N__68677),
            .I(N__68665));
    LocalMux I__10866 (
            .O(N__68672),
            .I(N__68662));
    InMux I__10865 (
            .O(N__68671),
            .I(N__68659));
    LocalMux I__10864 (
            .O(N__68668),
            .I(N__68656));
    Span4Mux_v I__10863 (
            .O(N__68665),
            .I(N__68648));
    Span4Mux_h I__10862 (
            .O(N__68662),
            .I(N__68648));
    LocalMux I__10861 (
            .O(N__68659),
            .I(N__68648));
    Span12Mux_s10_v I__10860 (
            .O(N__68656),
            .I(N__68644));
    InMux I__10859 (
            .O(N__68655),
            .I(N__68641));
    Span4Mux_v I__10858 (
            .O(N__68648),
            .I(N__68638));
    InMux I__10857 (
            .O(N__68647),
            .I(N__68635));
    Odrv12 I__10856 (
            .O(N__68644),
            .I(shift_srl_84Z0Z_15));
    LocalMux I__10855 (
            .O(N__68641),
            .I(shift_srl_84Z0Z_15));
    Odrv4 I__10854 (
            .O(N__68638),
            .I(shift_srl_84Z0Z_15));
    LocalMux I__10853 (
            .O(N__68635),
            .I(shift_srl_84Z0Z_15));
    IoInMux I__10852 (
            .O(N__68626),
            .I(N__68623));
    LocalMux I__10851 (
            .O(N__68623),
            .I(N__68620));
    IoSpan4Mux I__10850 (
            .O(N__68620),
            .I(N__68617));
    Span4Mux_s2_v I__10849 (
            .O(N__68617),
            .I(N__68614));
    Odrv4 I__10848 (
            .O(N__68614),
            .I(rco_c_84));
    InMux I__10847 (
            .O(N__68611),
            .I(N__68605));
    InMux I__10846 (
            .O(N__68610),
            .I(N__68602));
    InMux I__10845 (
            .O(N__68609),
            .I(N__68597));
    InMux I__10844 (
            .O(N__68608),
            .I(N__68597));
    LocalMux I__10843 (
            .O(N__68605),
            .I(N__68594));
    LocalMux I__10842 (
            .O(N__68602),
            .I(N__68591));
    LocalMux I__10841 (
            .O(N__68597),
            .I(N__68588));
    Span4Mux_v I__10840 (
            .O(N__68594),
            .I(N__68585));
    Span4Mux_v I__10839 (
            .O(N__68591),
            .I(N__68582));
    Span4Mux_v I__10838 (
            .O(N__68588),
            .I(N__68579));
    Odrv4 I__10837 (
            .O(N__68585),
            .I(shift_srl_89_RNIPCQF1Z0Z_15));
    Odrv4 I__10836 (
            .O(N__68582),
            .I(shift_srl_89_RNIPCQF1Z0Z_15));
    Odrv4 I__10835 (
            .O(N__68579),
            .I(shift_srl_89_RNIPCQF1Z0Z_15));
    IoInMux I__10834 (
            .O(N__68572),
            .I(N__68569));
    LocalMux I__10833 (
            .O(N__68569),
            .I(N__68566));
    Span4Mux_s2_v I__10832 (
            .O(N__68566),
            .I(N__68563));
    Odrv4 I__10831 (
            .O(N__68563),
            .I(rco_c_89));
    InMux I__10830 (
            .O(N__68560),
            .I(N__68554));
    InMux I__10829 (
            .O(N__68559),
            .I(N__68554));
    LocalMux I__10828 (
            .O(N__68554),
            .I(N__68551));
    Span4Mux_s3_v I__10827 (
            .O(N__68551),
            .I(N__68546));
    InMux I__10826 (
            .O(N__68550),
            .I(N__68543));
    InMux I__10825 (
            .O(N__68549),
            .I(N__68540));
    Odrv4 I__10824 (
            .O(N__68546),
            .I(shift_srl_91_RNIOVG12Z0Z_15));
    LocalMux I__10823 (
            .O(N__68543),
            .I(shift_srl_91_RNIOVG12Z0Z_15));
    LocalMux I__10822 (
            .O(N__68540),
            .I(shift_srl_91_RNIOVG12Z0Z_15));
    IoInMux I__10821 (
            .O(N__68533),
            .I(N__68530));
    LocalMux I__10820 (
            .O(N__68530),
            .I(N__68526));
    InMux I__10819 (
            .O(N__68529),
            .I(N__68523));
    IoSpan4Mux I__10818 (
            .O(N__68526),
            .I(N__68510));
    LocalMux I__10817 (
            .O(N__68523),
            .I(N__68510));
    InMux I__10816 (
            .O(N__68522),
            .I(N__68506));
    InMux I__10815 (
            .O(N__68521),
            .I(N__68502));
    InMux I__10814 (
            .O(N__68520),
            .I(N__68497));
    InMux I__10813 (
            .O(N__68519),
            .I(N__68497));
    InMux I__10812 (
            .O(N__68518),
            .I(N__68488));
    InMux I__10811 (
            .O(N__68517),
            .I(N__68488));
    InMux I__10810 (
            .O(N__68516),
            .I(N__68488));
    InMux I__10809 (
            .O(N__68515),
            .I(N__68488));
    Span4Mux_s2_v I__10808 (
            .O(N__68510),
            .I(N__68485));
    CascadeMux I__10807 (
            .O(N__68509),
            .I(N__68482));
    LocalMux I__10806 (
            .O(N__68506),
            .I(N__68474));
    InMux I__10805 (
            .O(N__68505),
            .I(N__68471));
    LocalMux I__10804 (
            .O(N__68502),
            .I(N__68464));
    LocalMux I__10803 (
            .O(N__68497),
            .I(N__68464));
    LocalMux I__10802 (
            .O(N__68488),
            .I(N__68464));
    Span4Mux_v I__10801 (
            .O(N__68485),
            .I(N__68461));
    InMux I__10800 (
            .O(N__68482),
            .I(N__68452));
    InMux I__10799 (
            .O(N__68481),
            .I(N__68452));
    InMux I__10798 (
            .O(N__68480),
            .I(N__68452));
    InMux I__10797 (
            .O(N__68479),
            .I(N__68452));
    InMux I__10796 (
            .O(N__68478),
            .I(N__68447));
    InMux I__10795 (
            .O(N__68477),
            .I(N__68447));
    Span4Mux_h I__10794 (
            .O(N__68474),
            .I(N__68440));
    LocalMux I__10793 (
            .O(N__68471),
            .I(N__68440));
    Span4Mux_h I__10792 (
            .O(N__68464),
            .I(N__68440));
    Odrv4 I__10791 (
            .O(N__68461),
            .I(rco_c_83));
    LocalMux I__10790 (
            .O(N__68452),
            .I(rco_c_83));
    LocalMux I__10789 (
            .O(N__68447),
            .I(rco_c_83));
    Odrv4 I__10788 (
            .O(N__68440),
            .I(rco_c_83));
    IoInMux I__10787 (
            .O(N__68431),
            .I(N__68428));
    LocalMux I__10786 (
            .O(N__68428),
            .I(N__68425));
    Span4Mux_s2_v I__10785 (
            .O(N__68425),
            .I(N__68422));
    Odrv4 I__10784 (
            .O(N__68422),
            .I(rco_c_92));
    InMux I__10783 (
            .O(N__68419),
            .I(N__68415));
    InMux I__10782 (
            .O(N__68418),
            .I(N__68412));
    LocalMux I__10781 (
            .O(N__68415),
            .I(N__68408));
    LocalMux I__10780 (
            .O(N__68412),
            .I(N__68405));
    InMux I__10779 (
            .O(N__68411),
            .I(N__68402));
    Sp12to4 I__10778 (
            .O(N__68408),
            .I(N__68397));
    Span12Mux_v I__10777 (
            .O(N__68405),
            .I(N__68397));
    LocalMux I__10776 (
            .O(N__68402),
            .I(shift_srl_92Z0Z_15));
    Odrv12 I__10775 (
            .O(N__68397),
            .I(shift_srl_92Z0Z_15));
    InMux I__10774 (
            .O(N__68392),
            .I(N__68389));
    LocalMux I__10773 (
            .O(N__68389),
            .I(shift_srl_93Z0Z_10));
    InMux I__10772 (
            .O(N__68386),
            .I(N__68383));
    LocalMux I__10771 (
            .O(N__68383),
            .I(shift_srl_40Z0Z_6));
    IoInMux I__10770 (
            .O(N__68380),
            .I(N__68377));
    LocalMux I__10769 (
            .O(N__68377),
            .I(N__68374));
    IoSpan4Mux I__10768 (
            .O(N__68374),
            .I(N__68371));
    Span4Mux_s3_v I__10767 (
            .O(N__68371),
            .I(N__68368));
    Span4Mux_h I__10766 (
            .O(N__68368),
            .I(N__68365));
    Odrv4 I__10765 (
            .O(N__68365),
            .I(rco_c_54));
    InMux I__10764 (
            .O(N__68362),
            .I(N__68359));
    LocalMux I__10763 (
            .O(N__68359),
            .I(shift_srl_198Z0Z_6));
    InMux I__10762 (
            .O(N__68356),
            .I(N__68353));
    LocalMux I__10761 (
            .O(N__68353),
            .I(shift_srl_93Z0Z_0));
    InMux I__10760 (
            .O(N__68350),
            .I(N__68347));
    LocalMux I__10759 (
            .O(N__68347),
            .I(shift_srl_93Z0Z_1));
    InMux I__10758 (
            .O(N__68344),
            .I(N__68341));
    LocalMux I__10757 (
            .O(N__68341),
            .I(shift_srl_93Z0Z_2));
    InMux I__10756 (
            .O(N__68338),
            .I(N__68335));
    LocalMux I__10755 (
            .O(N__68335),
            .I(shift_srl_93Z0Z_3));
    InMux I__10754 (
            .O(N__68332),
            .I(N__68329));
    LocalMux I__10753 (
            .O(N__68329),
            .I(shift_srl_93Z0Z_4));
    InMux I__10752 (
            .O(N__68326),
            .I(N__68323));
    LocalMux I__10751 (
            .O(N__68323),
            .I(shift_srl_119Z0Z_5));
    InMux I__10750 (
            .O(N__68320),
            .I(N__68317));
    LocalMux I__10749 (
            .O(N__68317),
            .I(shift_srl_119Z0Z_6));
    InMux I__10748 (
            .O(N__68314),
            .I(N__68311));
    LocalMux I__10747 (
            .O(N__68311),
            .I(shift_srl_119Z0Z_11));
    InMux I__10746 (
            .O(N__68308),
            .I(N__68305));
    LocalMux I__10745 (
            .O(N__68305),
            .I(shift_srl_119Z0Z_12));
    CEMux I__10744 (
            .O(N__68302),
            .I(N__68298));
    CEMux I__10743 (
            .O(N__68301),
            .I(N__68295));
    LocalMux I__10742 (
            .O(N__68298),
            .I(N__68289));
    LocalMux I__10741 (
            .O(N__68295),
            .I(N__68289));
    CEMux I__10740 (
            .O(N__68294),
            .I(N__68286));
    Span4Mux_v I__10739 (
            .O(N__68289),
            .I(N__68280));
    LocalMux I__10738 (
            .O(N__68286),
            .I(N__68280));
    CEMux I__10737 (
            .O(N__68285),
            .I(N__68277));
    Span4Mux_h I__10736 (
            .O(N__68280),
            .I(N__68274));
    LocalMux I__10735 (
            .O(N__68277),
            .I(N__68271));
    Span4Mux_h I__10734 (
            .O(N__68274),
            .I(N__68268));
    Odrv4 I__10733 (
            .O(N__68271),
            .I(clk_en_119));
    Odrv4 I__10732 (
            .O(N__68268),
            .I(clk_en_119));
    InMux I__10731 (
            .O(N__68263),
            .I(N__68260));
    LocalMux I__10730 (
            .O(N__68260),
            .I(shift_srl_40Z0Z_0));
    InMux I__10729 (
            .O(N__68257),
            .I(N__68254));
    LocalMux I__10728 (
            .O(N__68254),
            .I(shift_srl_40Z0Z_1));
    InMux I__10727 (
            .O(N__68251),
            .I(N__68248));
    LocalMux I__10726 (
            .O(N__68248),
            .I(shift_srl_40Z0Z_2));
    InMux I__10725 (
            .O(N__68245),
            .I(N__68242));
    LocalMux I__10724 (
            .O(N__68242),
            .I(shift_srl_40Z0Z_3));
    InMux I__10723 (
            .O(N__68239),
            .I(N__68236));
    LocalMux I__10722 (
            .O(N__68236),
            .I(shift_srl_40Z0Z_4));
    InMux I__10721 (
            .O(N__68233),
            .I(N__68230));
    LocalMux I__10720 (
            .O(N__68230),
            .I(shift_srl_40Z0Z_5));
    InMux I__10719 (
            .O(N__68227),
            .I(N__68224));
    LocalMux I__10718 (
            .O(N__68224),
            .I(shift_srl_127Z0Z_6));
    InMux I__10717 (
            .O(N__68221),
            .I(N__68218));
    LocalMux I__10716 (
            .O(N__68218),
            .I(shift_srl_127Z0Z_7));
    CEMux I__10715 (
            .O(N__68215),
            .I(N__68211));
    CEMux I__10714 (
            .O(N__68214),
            .I(N__68208));
    LocalMux I__10713 (
            .O(N__68211),
            .I(N__68205));
    LocalMux I__10712 (
            .O(N__68208),
            .I(N__68202));
    Odrv12 I__10711 (
            .O(N__68205),
            .I(clk_en_127));
    Odrv12 I__10710 (
            .O(N__68202),
            .I(clk_en_127));
    InMux I__10709 (
            .O(N__68197),
            .I(N__68194));
    LocalMux I__10708 (
            .O(N__68194),
            .I(shift_srl_173Z0Z_0));
    InMux I__10707 (
            .O(N__68191),
            .I(N__68188));
    LocalMux I__10706 (
            .O(N__68188),
            .I(shift_srl_173Z0Z_1));
    InMux I__10705 (
            .O(N__68185),
            .I(N__68182));
    LocalMux I__10704 (
            .O(N__68182),
            .I(shift_srl_173Z0Z_2));
    InMux I__10703 (
            .O(N__68179),
            .I(N__68176));
    LocalMux I__10702 (
            .O(N__68176),
            .I(shift_srl_173Z0Z_3));
    InMux I__10701 (
            .O(N__68173),
            .I(N__68170));
    LocalMux I__10700 (
            .O(N__68170),
            .I(shift_srl_173Z0Z_4));
    InMux I__10699 (
            .O(N__68167),
            .I(N__68164));
    LocalMux I__10698 (
            .O(N__68164),
            .I(shift_srl_173Z0Z_5));
    InMux I__10697 (
            .O(N__68161),
            .I(N__68158));
    LocalMux I__10696 (
            .O(N__68158),
            .I(shift_srl_173Z0Z_6));
    InMux I__10695 (
            .O(N__68155),
            .I(N__68152));
    LocalMux I__10694 (
            .O(N__68152),
            .I(shift_srl_119Z0Z_7));
    InMux I__10693 (
            .O(N__68149),
            .I(N__68146));
    LocalMux I__10692 (
            .O(N__68146),
            .I(shift_srl_111Z0Z_9));
    InMux I__10691 (
            .O(N__68143),
            .I(N__68140));
    LocalMux I__10690 (
            .O(N__68140),
            .I(N__68137));
    Span4Mux_h I__10689 (
            .O(N__68137),
            .I(N__68134));
    Odrv4 I__10688 (
            .O(N__68134),
            .I(shift_srl_111Z0Z_7));
    InMux I__10687 (
            .O(N__68131),
            .I(N__68128));
    LocalMux I__10686 (
            .O(N__68128),
            .I(shift_srl_111Z0Z_8));
    CEMux I__10685 (
            .O(N__68125),
            .I(N__68121));
    CEMux I__10684 (
            .O(N__68124),
            .I(N__68118));
    LocalMux I__10683 (
            .O(N__68121),
            .I(N__68115));
    LocalMux I__10682 (
            .O(N__68118),
            .I(N__68111));
    Span4Mux_v I__10681 (
            .O(N__68115),
            .I(N__68108));
    CEMux I__10680 (
            .O(N__68114),
            .I(N__68105));
    Span4Mux_v I__10679 (
            .O(N__68111),
            .I(N__68098));
    Span4Mux_h I__10678 (
            .O(N__68108),
            .I(N__68098));
    LocalMux I__10677 (
            .O(N__68105),
            .I(N__68098));
    Span4Mux_h I__10676 (
            .O(N__68098),
            .I(N__68095));
    Odrv4 I__10675 (
            .O(N__68095),
            .I(clk_en_111));
    CascadeMux I__10674 (
            .O(N__68092),
            .I(N__68089));
    InMux I__10673 (
            .O(N__68089),
            .I(N__68086));
    LocalMux I__10672 (
            .O(N__68086),
            .I(N__68083));
    Span4Mux_h I__10671 (
            .O(N__68083),
            .I(N__68079));
    InMux I__10670 (
            .O(N__68082),
            .I(N__68076));
    Span4Mux_h I__10669 (
            .O(N__68079),
            .I(N__68073));
    LocalMux I__10668 (
            .O(N__68076),
            .I(shift_srl_127Z0Z_15));
    Odrv4 I__10667 (
            .O(N__68073),
            .I(shift_srl_127Z0Z_15));
    InMux I__10666 (
            .O(N__68068),
            .I(N__68065));
    LocalMux I__10665 (
            .O(N__68065),
            .I(shift_srl_127Z0Z_0));
    InMux I__10664 (
            .O(N__68062),
            .I(N__68059));
    LocalMux I__10663 (
            .O(N__68059),
            .I(shift_srl_127Z0Z_1));
    InMux I__10662 (
            .O(N__68056),
            .I(N__68053));
    LocalMux I__10661 (
            .O(N__68053),
            .I(shift_srl_127Z0Z_2));
    InMux I__10660 (
            .O(N__68050),
            .I(N__68047));
    LocalMux I__10659 (
            .O(N__68047),
            .I(shift_srl_127Z0Z_3));
    InMux I__10658 (
            .O(N__68044),
            .I(N__68041));
    LocalMux I__10657 (
            .O(N__68041),
            .I(shift_srl_127Z0Z_4));
    InMux I__10656 (
            .O(N__68038),
            .I(N__68035));
    LocalMux I__10655 (
            .O(N__68035),
            .I(shift_srl_127Z0Z_5));
    InMux I__10654 (
            .O(N__68032),
            .I(N__68029));
    LocalMux I__10653 (
            .O(N__68029),
            .I(shift_srl_187Z0Z_1));
    InMux I__10652 (
            .O(N__68026),
            .I(N__68023));
    LocalMux I__10651 (
            .O(N__68023),
            .I(shift_srl_187Z0Z_2));
    InMux I__10650 (
            .O(N__68020),
            .I(N__68017));
    LocalMux I__10649 (
            .O(N__68017),
            .I(shift_srl_187Z0Z_3));
    InMux I__10648 (
            .O(N__68014),
            .I(N__68011));
    LocalMux I__10647 (
            .O(N__68011),
            .I(shift_srl_187Z0Z_4));
    InMux I__10646 (
            .O(N__68008),
            .I(N__68005));
    LocalMux I__10645 (
            .O(N__68005),
            .I(shift_srl_187Z0Z_5));
    InMux I__10644 (
            .O(N__68002),
            .I(N__67999));
    LocalMux I__10643 (
            .O(N__67999),
            .I(shift_srl_187Z0Z_6));
    InMux I__10642 (
            .O(N__67996),
            .I(N__67993));
    LocalMux I__10641 (
            .O(N__67993),
            .I(shift_srl_111Z0Z_10));
    InMux I__10640 (
            .O(N__67990),
            .I(N__67987));
    LocalMux I__10639 (
            .O(N__67987),
            .I(shift_srl_111Z0Z_11));
    InMux I__10638 (
            .O(N__67984),
            .I(N__67981));
    LocalMux I__10637 (
            .O(N__67981),
            .I(N__67978));
    Span4Mux_h I__10636 (
            .O(N__67978),
            .I(N__67975));
    Odrv4 I__10635 (
            .O(N__67975),
            .I(shift_srl_111Z0Z_12));
    InMux I__10634 (
            .O(N__67972),
            .I(N__67969));
    LocalMux I__10633 (
            .O(N__67969),
            .I(shift_srl_156Z0Z_0));
    InMux I__10632 (
            .O(N__67966),
            .I(N__67963));
    LocalMux I__10631 (
            .O(N__67963),
            .I(shift_srl_156Z0Z_1));
    InMux I__10630 (
            .O(N__67960),
            .I(N__67957));
    LocalMux I__10629 (
            .O(N__67957),
            .I(shift_srl_156Z0Z_2));
    InMux I__10628 (
            .O(N__67954),
            .I(N__67951));
    LocalMux I__10627 (
            .O(N__67951),
            .I(shift_srl_156Z0Z_3));
    InMux I__10626 (
            .O(N__67948),
            .I(N__67945));
    LocalMux I__10625 (
            .O(N__67945),
            .I(shift_srl_156Z0Z_4));
    InMux I__10624 (
            .O(N__67942),
            .I(N__67939));
    LocalMux I__10623 (
            .O(N__67939),
            .I(shift_srl_156Z0Z_5));
    InMux I__10622 (
            .O(N__67936),
            .I(N__67933));
    LocalMux I__10621 (
            .O(N__67933),
            .I(shift_srl_156Z0Z_6));
    InMux I__10620 (
            .O(N__67930),
            .I(N__67927));
    LocalMux I__10619 (
            .O(N__67927),
            .I(shift_srl_187Z0Z_0));
    InMux I__10618 (
            .O(N__67924),
            .I(N__67921));
    LocalMux I__10617 (
            .O(N__67921),
            .I(shift_srl_162Z0Z_0));
    InMux I__10616 (
            .O(N__67918),
            .I(N__67915));
    LocalMux I__10615 (
            .O(N__67915),
            .I(shift_srl_162Z0Z_1));
    InMux I__10614 (
            .O(N__67912),
            .I(N__67909));
    LocalMux I__10613 (
            .O(N__67909),
            .I(shift_srl_162Z0Z_2));
    InMux I__10612 (
            .O(N__67906),
            .I(N__67903));
    LocalMux I__10611 (
            .O(N__67903),
            .I(shift_srl_162Z0Z_3));
    InMux I__10610 (
            .O(N__67900),
            .I(N__67897));
    LocalMux I__10609 (
            .O(N__67897),
            .I(shift_srl_162Z0Z_4));
    InMux I__10608 (
            .O(N__67894),
            .I(N__67891));
    LocalMux I__10607 (
            .O(N__67891),
            .I(shift_srl_162Z0Z_5));
    InMux I__10606 (
            .O(N__67888),
            .I(N__67885));
    LocalMux I__10605 (
            .O(N__67885),
            .I(shift_srl_162Z0Z_11));
    InMux I__10604 (
            .O(N__67882),
            .I(N__67879));
    LocalMux I__10603 (
            .O(N__67879),
            .I(shift_srl_162Z0Z_12));
    InMux I__10602 (
            .O(N__67876),
            .I(N__67873));
    LocalMux I__10601 (
            .O(N__67873),
            .I(shift_srl_162Z0Z_13));
    InMux I__10600 (
            .O(N__67870),
            .I(N__67867));
    LocalMux I__10599 (
            .O(N__67867),
            .I(shift_srl_38Z0Z_13));
    InMux I__10598 (
            .O(N__67864),
            .I(N__67861));
    LocalMux I__10597 (
            .O(N__67861),
            .I(shift_srl_158Z0Z_0));
    InMux I__10596 (
            .O(N__67858),
            .I(N__67855));
    LocalMux I__10595 (
            .O(N__67855),
            .I(shift_srl_158Z0Z_1));
    InMux I__10594 (
            .O(N__67852),
            .I(N__67849));
    LocalMux I__10593 (
            .O(N__67849),
            .I(shift_srl_158Z0Z_2));
    InMux I__10592 (
            .O(N__67846),
            .I(N__67843));
    LocalMux I__10591 (
            .O(N__67843),
            .I(shift_srl_158Z0Z_3));
    InMux I__10590 (
            .O(N__67840),
            .I(N__67837));
    LocalMux I__10589 (
            .O(N__67837),
            .I(shift_srl_158Z0Z_4));
    InMux I__10588 (
            .O(N__67834),
            .I(N__67831));
    LocalMux I__10587 (
            .O(N__67831),
            .I(shift_srl_158Z0Z_5));
    InMux I__10586 (
            .O(N__67828),
            .I(N__67825));
    LocalMux I__10585 (
            .O(N__67825),
            .I(shift_srl_158Z0Z_6));
    InMux I__10584 (
            .O(N__67822),
            .I(N__67819));
    LocalMux I__10583 (
            .O(N__67819),
            .I(N__67816));
    Odrv4 I__10582 (
            .O(N__67816),
            .I(shift_srl_29Z0Z_9));
    InMux I__10581 (
            .O(N__67813),
            .I(N__67810));
    LocalMux I__10580 (
            .O(N__67810),
            .I(shift_srl_29Z0Z_10));
    InMux I__10579 (
            .O(N__67807),
            .I(N__67804));
    LocalMux I__10578 (
            .O(N__67804),
            .I(shift_srl_29Z0Z_11));
    InMux I__10577 (
            .O(N__67801),
            .I(N__67798));
    LocalMux I__10576 (
            .O(N__67798),
            .I(shift_srl_29Z0Z_12));
    InMux I__10575 (
            .O(N__67795),
            .I(N__67792));
    LocalMux I__10574 (
            .O(N__67792),
            .I(N__67789));
    Odrv4 I__10573 (
            .O(N__67789),
            .I(shift_srl_29Z0Z_1));
    InMux I__10572 (
            .O(N__67786),
            .I(N__67783));
    LocalMux I__10571 (
            .O(N__67783),
            .I(shift_srl_29Z0Z_0));
    InMux I__10570 (
            .O(N__67780),
            .I(N__67777));
    LocalMux I__10569 (
            .O(N__67777),
            .I(shift_srl_29Z0Z_13));
    InMux I__10568 (
            .O(N__67774),
            .I(N__67771));
    LocalMux I__10567 (
            .O(N__67771),
            .I(shift_srl_29Z0Z_14));
    CEMux I__10566 (
            .O(N__67768),
            .I(N__67765));
    LocalMux I__10565 (
            .O(N__67765),
            .I(N__67762));
    Span4Mux_v I__10564 (
            .O(N__67762),
            .I(N__67758));
    CEMux I__10563 (
            .O(N__67761),
            .I(N__67755));
    Span4Mux_h I__10562 (
            .O(N__67758),
            .I(N__67752));
    LocalMux I__10561 (
            .O(N__67755),
            .I(N__67749));
    Odrv4 I__10560 (
            .O(N__67752),
            .I(clk_en_29));
    Odrv12 I__10559 (
            .O(N__67749),
            .I(clk_en_29));
    InMux I__10558 (
            .O(N__67744),
            .I(N__67741));
    LocalMux I__10557 (
            .O(N__67741),
            .I(shift_srl_29Z0Z_7));
    InMux I__10556 (
            .O(N__67738),
            .I(N__67735));
    LocalMux I__10555 (
            .O(N__67735),
            .I(shift_srl_29Z0Z_8));
    IoInMux I__10554 (
            .O(N__67732),
            .I(N__67729));
    LocalMux I__10553 (
            .O(N__67729),
            .I(N__67726));
    Span12Mux_s11_h I__10552 (
            .O(N__67726),
            .I(N__67723));
    Odrv12 I__10551 (
            .O(N__67723),
            .I(rco_c_27));
    CascadeMux I__10550 (
            .O(N__67720),
            .I(rco_c_27_cascade_));
    CEMux I__10549 (
            .O(N__67717),
            .I(N__67713));
    CEMux I__10548 (
            .O(N__67716),
            .I(N__67710));
    LocalMux I__10547 (
            .O(N__67713),
            .I(clk_en_28));
    LocalMux I__10546 (
            .O(N__67710),
            .I(clk_en_28));
    InMux I__10545 (
            .O(N__67705),
            .I(N__67699));
    InMux I__10544 (
            .O(N__67704),
            .I(N__67699));
    LocalMux I__10543 (
            .O(N__67699),
            .I(rco_int_0_a2_0_a2_out_1));
    IoInMux I__10542 (
            .O(N__67696),
            .I(N__67693));
    LocalMux I__10541 (
            .O(N__67693),
            .I(N__67690));
    Span12Mux_s9_h I__10540 (
            .O(N__67690),
            .I(N__67687));
    Odrv12 I__10539 (
            .O(N__67687),
            .I(rco_c_28));
    CascadeMux I__10538 (
            .O(N__67684),
            .I(rco_c_28_cascade_));
    CascadeMux I__10537 (
            .O(N__67681),
            .I(shift_srl_27_RNIP5TNZ0Z_15_cascade_));
    CascadeMux I__10536 (
            .O(N__67678),
            .I(rco_int_0_a2_0_a2_out_2_cascade_));
    InMux I__10535 (
            .O(N__67675),
            .I(N__67672));
    LocalMux I__10534 (
            .O(N__67672),
            .I(shift_srl_99Z0Z_3));
    InMux I__10533 (
            .O(N__67669),
            .I(N__67666));
    LocalMux I__10532 (
            .O(N__67666),
            .I(shift_srl_99Z0Z_4));
    InMux I__10531 (
            .O(N__67663),
            .I(N__67660));
    LocalMux I__10530 (
            .O(N__67660),
            .I(N__67657));
    Span4Mux_h I__10529 (
            .O(N__67657),
            .I(N__67654));
    Odrv4 I__10528 (
            .O(N__67654),
            .I(shift_srl_99Z0Z_5));
    CEMux I__10527 (
            .O(N__67651),
            .I(N__67647));
    CEMux I__10526 (
            .O(N__67650),
            .I(N__67644));
    LocalMux I__10525 (
            .O(N__67647),
            .I(N__67641));
    LocalMux I__10524 (
            .O(N__67644),
            .I(N__67637));
    Span4Mux_v I__10523 (
            .O(N__67641),
            .I(N__67634));
    CEMux I__10522 (
            .O(N__67640),
            .I(N__67631));
    Span4Mux_v I__10521 (
            .O(N__67637),
            .I(N__67628));
    Span4Mux_h I__10520 (
            .O(N__67634),
            .I(N__67625));
    LocalMux I__10519 (
            .O(N__67631),
            .I(N__67622));
    Odrv4 I__10518 (
            .O(N__67628),
            .I(clk_en_99));
    Odrv4 I__10517 (
            .O(N__67625),
            .I(clk_en_99));
    Odrv12 I__10516 (
            .O(N__67622),
            .I(clk_en_99));
    InMux I__10515 (
            .O(N__67615),
            .I(N__67612));
    LocalMux I__10514 (
            .O(N__67612),
            .I(shift_srl_29Z0Z_2));
    InMux I__10513 (
            .O(N__67609),
            .I(N__67606));
    LocalMux I__10512 (
            .O(N__67606),
            .I(shift_srl_29Z0Z_3));
    InMux I__10511 (
            .O(N__67603),
            .I(N__67600));
    LocalMux I__10510 (
            .O(N__67600),
            .I(shift_srl_29Z0Z_4));
    InMux I__10509 (
            .O(N__67597),
            .I(N__67594));
    LocalMux I__10508 (
            .O(N__67594),
            .I(shift_srl_29Z0Z_5));
    InMux I__10507 (
            .O(N__67591),
            .I(N__67588));
    LocalMux I__10506 (
            .O(N__67588),
            .I(shift_srl_29Z0Z_6));
    InMux I__10505 (
            .O(N__67585),
            .I(N__67582));
    LocalMux I__10504 (
            .O(N__67582),
            .I(shift_srl_98Z0Z_14));
    InMux I__10503 (
            .O(N__67579),
            .I(N__67576));
    LocalMux I__10502 (
            .O(N__67576),
            .I(shift_srl_98Z0Z_9));
    InMux I__10501 (
            .O(N__67573),
            .I(N__67570));
    LocalMux I__10500 (
            .O(N__67570),
            .I(shift_srl_98Z0Z_7));
    InMux I__10499 (
            .O(N__67567),
            .I(N__67564));
    LocalMux I__10498 (
            .O(N__67564),
            .I(shift_srl_98Z0Z_8));
    CEMux I__10497 (
            .O(N__67561),
            .I(N__67558));
    LocalMux I__10496 (
            .O(N__67558),
            .I(N__67555));
    Span4Mux_v I__10495 (
            .O(N__67555),
            .I(N__67551));
    CEMux I__10494 (
            .O(N__67554),
            .I(N__67548));
    Span4Mux_v I__10493 (
            .O(N__67551),
            .I(N__67543));
    LocalMux I__10492 (
            .O(N__67548),
            .I(N__67543));
    Span4Mux_v I__10491 (
            .O(N__67543),
            .I(N__67540));
    Odrv4 I__10490 (
            .O(N__67540),
            .I(clk_en_98));
    InMux I__10489 (
            .O(N__67537),
            .I(N__67534));
    LocalMux I__10488 (
            .O(N__67534),
            .I(N__67531));
    Span4Mux_v I__10487 (
            .O(N__67531),
            .I(N__67528));
    Odrv4 I__10486 (
            .O(N__67528),
            .I(shift_srl_99Z0Z_14));
    InMux I__10485 (
            .O(N__67525),
            .I(N__67519));
    InMux I__10484 (
            .O(N__67524),
            .I(N__67519));
    LocalMux I__10483 (
            .O(N__67519),
            .I(shift_srl_99Z0Z_15));
    InMux I__10482 (
            .O(N__67516),
            .I(N__67513));
    LocalMux I__10481 (
            .O(N__67513),
            .I(shift_srl_99Z0Z_0));
    InMux I__10480 (
            .O(N__67510),
            .I(N__67507));
    LocalMux I__10479 (
            .O(N__67507),
            .I(shift_srl_99Z0Z_1));
    InMux I__10478 (
            .O(N__67504),
            .I(N__67501));
    LocalMux I__10477 (
            .O(N__67501),
            .I(shift_srl_99Z0Z_2));
    InMux I__10476 (
            .O(N__67498),
            .I(N__67495));
    LocalMux I__10475 (
            .O(N__67495),
            .I(shift_srl_98Z0Z_3));
    InMux I__10474 (
            .O(N__67492),
            .I(N__67489));
    LocalMux I__10473 (
            .O(N__67489),
            .I(shift_srl_98Z0Z_4));
    InMux I__10472 (
            .O(N__67486),
            .I(N__67483));
    LocalMux I__10471 (
            .O(N__67483),
            .I(shift_srl_98Z0Z_5));
    InMux I__10470 (
            .O(N__67480),
            .I(N__67477));
    LocalMux I__10469 (
            .O(N__67477),
            .I(shift_srl_98Z0Z_6));
    InMux I__10468 (
            .O(N__67474),
            .I(N__67471));
    LocalMux I__10467 (
            .O(N__67471),
            .I(shift_srl_98Z0Z_10));
    InMux I__10466 (
            .O(N__67468),
            .I(N__67465));
    LocalMux I__10465 (
            .O(N__67465),
            .I(shift_srl_98Z0Z_11));
    InMux I__10464 (
            .O(N__67462),
            .I(N__67459));
    LocalMux I__10463 (
            .O(N__67459),
            .I(shift_srl_98Z0Z_12));
    InMux I__10462 (
            .O(N__67456),
            .I(N__67453));
    LocalMux I__10461 (
            .O(N__67453),
            .I(shift_srl_98Z0Z_13));
    InMux I__10460 (
            .O(N__67450),
            .I(N__67447));
    LocalMux I__10459 (
            .O(N__67447),
            .I(shift_srl_59Z0Z_13));
    InMux I__10458 (
            .O(N__67444),
            .I(N__67441));
    LocalMux I__10457 (
            .O(N__67441),
            .I(shift_srl_59Z0Z_12));
    InMux I__10456 (
            .O(N__67438),
            .I(N__67435));
    LocalMux I__10455 (
            .O(N__67435),
            .I(shift_srl_59Z0Z_11));
    InMux I__10454 (
            .O(N__67432),
            .I(N__67429));
    LocalMux I__10453 (
            .O(N__67429),
            .I(shift_srl_59Z0Z_10));
    InMux I__10452 (
            .O(N__67426),
            .I(N__67423));
    LocalMux I__10451 (
            .O(N__67423),
            .I(shift_srl_59Z0Z_8));
    InMux I__10450 (
            .O(N__67420),
            .I(N__67417));
    LocalMux I__10449 (
            .O(N__67417),
            .I(shift_srl_59Z0Z_9));
    InMux I__10448 (
            .O(N__67414),
            .I(N__67411));
    LocalMux I__10447 (
            .O(N__67411),
            .I(shift_srl_98Z0Z_0));
    InMux I__10446 (
            .O(N__67408),
            .I(N__67405));
    LocalMux I__10445 (
            .O(N__67405),
            .I(shift_srl_98Z0Z_1));
    InMux I__10444 (
            .O(N__67402),
            .I(N__67399));
    LocalMux I__10443 (
            .O(N__67399),
            .I(shift_srl_98Z0Z_2));
    InMux I__10442 (
            .O(N__67396),
            .I(N__67393));
    LocalMux I__10441 (
            .O(N__67393),
            .I(shift_srl_45Z0Z_0));
    InMux I__10440 (
            .O(N__67390),
            .I(N__67387));
    LocalMux I__10439 (
            .O(N__67387),
            .I(shift_srl_45Z0Z_1));
    InMux I__10438 (
            .O(N__67384),
            .I(N__67381));
    LocalMux I__10437 (
            .O(N__67381),
            .I(shift_srl_45Z0Z_2));
    InMux I__10436 (
            .O(N__67378),
            .I(N__67375));
    LocalMux I__10435 (
            .O(N__67375),
            .I(shift_srl_45Z0Z_3));
    InMux I__10434 (
            .O(N__67372),
            .I(N__67369));
    LocalMux I__10433 (
            .O(N__67369),
            .I(shift_srl_45Z0Z_4));
    InMux I__10432 (
            .O(N__67366),
            .I(N__67363));
    LocalMux I__10431 (
            .O(N__67363),
            .I(shift_srl_45Z0Z_5));
    InMux I__10430 (
            .O(N__67360),
            .I(N__67357));
    LocalMux I__10429 (
            .O(N__67357),
            .I(shift_srl_45Z0Z_6));
    InMux I__10428 (
            .O(N__67354),
            .I(N__67350));
    InMux I__10427 (
            .O(N__67353),
            .I(N__67347));
    LocalMux I__10426 (
            .O(N__67350),
            .I(N__67344));
    LocalMux I__10425 (
            .O(N__67347),
            .I(N__67341));
    Span4Mux_h I__10424 (
            .O(N__67344),
            .I(N__67338));
    Span4Mux_h I__10423 (
            .O(N__67341),
            .I(N__67335));
    Odrv4 I__10422 (
            .O(N__67338),
            .I(rco_int_0_a2_0_a2_83_m6_0_a2_sx));
    Odrv4 I__10421 (
            .O(N__67335),
            .I(rco_int_0_a2_0_a2_83_m6_0_a2_sx));
    InMux I__10420 (
            .O(N__67330),
            .I(N__67327));
    LocalMux I__10419 (
            .O(N__67327),
            .I(shift_srl_59Z0Z_14));
    IoInMux I__10418 (
            .O(N__67324),
            .I(N__67321));
    LocalMux I__10417 (
            .O(N__67321),
            .I(N__67318));
    Span4Mux_s0_v I__10416 (
            .O(N__67318),
            .I(N__67315));
    Span4Mux_v I__10415 (
            .O(N__67315),
            .I(N__67312));
    Span4Mux_v I__10414 (
            .O(N__67312),
            .I(N__67309));
    Span4Mux_h I__10413 (
            .O(N__67309),
            .I(N__67306));
    Odrv4 I__10412 (
            .O(N__67306),
            .I(rco_c_40));
    CEMux I__10411 (
            .O(N__67303),
            .I(N__67299));
    CEMux I__10410 (
            .O(N__67302),
            .I(N__67296));
    LocalMux I__10409 (
            .O(N__67299),
            .I(N__67292));
    LocalMux I__10408 (
            .O(N__67296),
            .I(N__67289));
    CEMux I__10407 (
            .O(N__67295),
            .I(N__67286));
    Span4Mux_v I__10406 (
            .O(N__67292),
            .I(N__67283));
    Span4Mux_h I__10405 (
            .O(N__67289),
            .I(N__67280));
    LocalMux I__10404 (
            .O(N__67286),
            .I(N__67277));
    Odrv4 I__10403 (
            .O(N__67283),
            .I(clk_en_42));
    Odrv4 I__10402 (
            .O(N__67280),
            .I(clk_en_42));
    Odrv4 I__10401 (
            .O(N__67277),
            .I(clk_en_42));
    CascadeMux I__10400 (
            .O(N__67270),
            .I(rco_c_39_cascade_));
    IoInMux I__10399 (
            .O(N__67267),
            .I(N__67264));
    LocalMux I__10398 (
            .O(N__67264),
            .I(N__67261));
    Span12Mux_s11_v I__10397 (
            .O(N__67261),
            .I(N__67258));
    Span12Mux_v I__10396 (
            .O(N__67258),
            .I(N__67255));
    Odrv12 I__10395 (
            .O(N__67255),
            .I(clk_en_40));
    IoInMux I__10394 (
            .O(N__67252),
            .I(N__67249));
    LocalMux I__10393 (
            .O(N__67249),
            .I(N__67246));
    Span4Mux_s0_v I__10392 (
            .O(N__67246),
            .I(N__67243));
    Span4Mux_v I__10391 (
            .O(N__67243),
            .I(N__67240));
    Span4Mux_v I__10390 (
            .O(N__67240),
            .I(N__67237));
    Span4Mux_h I__10389 (
            .O(N__67237),
            .I(N__67232));
    InMux I__10388 (
            .O(N__67236),
            .I(N__67229));
    InMux I__10387 (
            .O(N__67235),
            .I(N__67226));
    Odrv4 I__10386 (
            .O(N__67232),
            .I(rco_c_39));
    LocalMux I__10385 (
            .O(N__67229),
            .I(rco_c_39));
    LocalMux I__10384 (
            .O(N__67226),
            .I(rco_c_39));
    CascadeMux I__10383 (
            .O(N__67219),
            .I(clk_en_0_a3_0_a2_sx_98_cascade_));
    IoInMux I__10382 (
            .O(N__67216),
            .I(N__67213));
    LocalMux I__10381 (
            .O(N__67213),
            .I(N__67210));
    IoSpan4Mux I__10380 (
            .O(N__67210),
            .I(N__67207));
    Span4Mux_s3_v I__10379 (
            .O(N__67207),
            .I(N__67204));
    Span4Mux_v I__10378 (
            .O(N__67204),
            .I(N__67201));
    Span4Mux_h I__10377 (
            .O(N__67201),
            .I(N__67198));
    Odrv4 I__10376 (
            .O(N__67198),
            .I(rco_c_97));
    InMux I__10375 (
            .O(N__67195),
            .I(N__67192));
    LocalMux I__10374 (
            .O(N__67192),
            .I(shift_srl_95Z0Z_6));
    InMux I__10373 (
            .O(N__67189),
            .I(N__67186));
    LocalMux I__10372 (
            .O(N__67186),
            .I(shift_srl_95Z0Z_7));
    InMux I__10371 (
            .O(N__67183),
            .I(N__67180));
    LocalMux I__10370 (
            .O(N__67180),
            .I(N__67177));
    Odrv12 I__10369 (
            .O(N__67177),
            .I(shift_srl_86Z0Z_14));
    CEMux I__10368 (
            .O(N__67174),
            .I(N__67171));
    LocalMux I__10367 (
            .O(N__67171),
            .I(N__67166));
    CEMux I__10366 (
            .O(N__67170),
            .I(N__67163));
    CEMux I__10365 (
            .O(N__67169),
            .I(N__67160));
    Span4Mux_h I__10364 (
            .O(N__67166),
            .I(N__67157));
    LocalMux I__10363 (
            .O(N__67163),
            .I(N__67154));
    LocalMux I__10362 (
            .O(N__67160),
            .I(N__67151));
    Odrv4 I__10361 (
            .O(N__67157),
            .I(clk_en_86));
    Odrv4 I__10360 (
            .O(N__67154),
            .I(clk_en_86));
    Odrv4 I__10359 (
            .O(N__67151),
            .I(clk_en_86));
    InMux I__10358 (
            .O(N__67144),
            .I(N__67140));
    InMux I__10357 (
            .O(N__67143),
            .I(N__67137));
    LocalMux I__10356 (
            .O(N__67140),
            .I(N__67133));
    LocalMux I__10355 (
            .O(N__67137),
            .I(N__67130));
    InMux I__10354 (
            .O(N__67136),
            .I(N__67127));
    Span4Mux_v I__10353 (
            .O(N__67133),
            .I(N__67124));
    Odrv12 I__10352 (
            .O(N__67130),
            .I(shift_srl_86Z0Z_15));
    LocalMux I__10351 (
            .O(N__67127),
            .I(shift_srl_86Z0Z_15));
    Odrv4 I__10350 (
            .O(N__67124),
            .I(shift_srl_86Z0Z_15));
    CascadeMux I__10349 (
            .O(N__67117),
            .I(N__67114));
    InMux I__10348 (
            .O(N__67114),
            .I(N__67111));
    LocalMux I__10347 (
            .O(N__67111),
            .I(N__67107));
    InMux I__10346 (
            .O(N__67110),
            .I(N__67101));
    Span4Mux_v I__10345 (
            .O(N__67107),
            .I(N__67096));
    InMux I__10344 (
            .O(N__67106),
            .I(N__67093));
    InMux I__10343 (
            .O(N__67105),
            .I(N__67088));
    InMux I__10342 (
            .O(N__67104),
            .I(N__67088));
    LocalMux I__10341 (
            .O(N__67101),
            .I(N__67085));
    InMux I__10340 (
            .O(N__67100),
            .I(N__67080));
    InMux I__10339 (
            .O(N__67099),
            .I(N__67080));
    Span4Mux_h I__10338 (
            .O(N__67096),
            .I(N__67077));
    LocalMux I__10337 (
            .O(N__67093),
            .I(N__67072));
    LocalMux I__10336 (
            .O(N__67088),
            .I(N__67072));
    Odrv12 I__10335 (
            .O(N__67085),
            .I(shift_srl_87Z0Z_15));
    LocalMux I__10334 (
            .O(N__67080),
            .I(shift_srl_87Z0Z_15));
    Odrv4 I__10333 (
            .O(N__67077),
            .I(shift_srl_87Z0Z_15));
    Odrv12 I__10332 (
            .O(N__67072),
            .I(shift_srl_87Z0Z_15));
    InMux I__10331 (
            .O(N__67063),
            .I(N__67058));
    InMux I__10330 (
            .O(N__67062),
            .I(N__67054));
    InMux I__10329 (
            .O(N__67061),
            .I(N__67051));
    LocalMux I__10328 (
            .O(N__67058),
            .I(N__67048));
    InMux I__10327 (
            .O(N__67057),
            .I(N__67044));
    LocalMux I__10326 (
            .O(N__67054),
            .I(N__67041));
    LocalMux I__10325 (
            .O(N__67051),
            .I(N__67038));
    Span4Mux_v I__10324 (
            .O(N__67048),
            .I(N__67035));
    InMux I__10323 (
            .O(N__67047),
            .I(N__67032));
    LocalMux I__10322 (
            .O(N__67044),
            .I(N__67025));
    Span4Mux_h I__10321 (
            .O(N__67041),
            .I(N__67025));
    Span4Mux_v I__10320 (
            .O(N__67038),
            .I(N__67025));
    Odrv4 I__10319 (
            .O(N__67035),
            .I(shift_srl_85Z0Z_15));
    LocalMux I__10318 (
            .O(N__67032),
            .I(shift_srl_85Z0Z_15));
    Odrv4 I__10317 (
            .O(N__67025),
            .I(shift_srl_85Z0Z_15));
    InMux I__10316 (
            .O(N__67018),
            .I(N__67015));
    LocalMux I__10315 (
            .O(N__67015),
            .I(N__67012));
    Span4Mux_h I__10314 (
            .O(N__67012),
            .I(N__67008));
    InMux I__10313 (
            .O(N__67011),
            .I(N__67004));
    Span4Mux_v I__10312 (
            .O(N__67008),
            .I(N__67001));
    InMux I__10311 (
            .O(N__67007),
            .I(N__66998));
    LocalMux I__10310 (
            .O(N__67004),
            .I(shift_srl_89Z0Z_15));
    Odrv4 I__10309 (
            .O(N__67001),
            .I(shift_srl_89Z0Z_15));
    LocalMux I__10308 (
            .O(N__66998),
            .I(shift_srl_89Z0Z_15));
    CascadeMux I__10307 (
            .O(N__66991),
            .I(rco_int_0_a2_0_a2_0_sx_89_cascade_));
    InMux I__10306 (
            .O(N__66988),
            .I(N__66982));
    InMux I__10305 (
            .O(N__66987),
            .I(N__66977));
    InMux I__10304 (
            .O(N__66986),
            .I(N__66977));
    InMux I__10303 (
            .O(N__66985),
            .I(N__66974));
    LocalMux I__10302 (
            .O(N__66982),
            .I(N__66970));
    LocalMux I__10301 (
            .O(N__66977),
            .I(N__66967));
    LocalMux I__10300 (
            .O(N__66974),
            .I(N__66964));
    InMux I__10299 (
            .O(N__66973),
            .I(N__66961));
    Span4Mux_h I__10298 (
            .O(N__66970),
            .I(N__66958));
    Span12Mux_v I__10297 (
            .O(N__66967),
            .I(N__66955));
    Odrv4 I__10296 (
            .O(N__66964),
            .I(shift_srl_88Z0Z_15));
    LocalMux I__10295 (
            .O(N__66961),
            .I(shift_srl_88Z0Z_15));
    Odrv4 I__10294 (
            .O(N__66958),
            .I(shift_srl_88Z0Z_15));
    Odrv12 I__10293 (
            .O(N__66955),
            .I(shift_srl_88Z0Z_15));
    InMux I__10292 (
            .O(N__66946),
            .I(N__66942));
    InMux I__10291 (
            .O(N__66945),
            .I(N__66939));
    LocalMux I__10290 (
            .O(N__66942),
            .I(N__66935));
    LocalMux I__10289 (
            .O(N__66939),
            .I(N__66932));
    InMux I__10288 (
            .O(N__66938),
            .I(N__66929));
    Span4Mux_h I__10287 (
            .O(N__66935),
            .I(N__66926));
    Span4Mux_v I__10286 (
            .O(N__66932),
            .I(N__66923));
    LocalMux I__10285 (
            .O(N__66929),
            .I(shift_srl_91Z0Z_15));
    Odrv4 I__10284 (
            .O(N__66926),
            .I(shift_srl_91Z0Z_15));
    Odrv4 I__10283 (
            .O(N__66923),
            .I(shift_srl_91Z0Z_15));
    InMux I__10282 (
            .O(N__66916),
            .I(N__66911));
    CascadeMux I__10281 (
            .O(N__66915),
            .I(N__66908));
    InMux I__10280 (
            .O(N__66914),
            .I(N__66905));
    LocalMux I__10279 (
            .O(N__66911),
            .I(N__66901));
    InMux I__10278 (
            .O(N__66908),
            .I(N__66898));
    LocalMux I__10277 (
            .O(N__66905),
            .I(N__66895));
    CascadeMux I__10276 (
            .O(N__66904),
            .I(N__66891));
    Span4Mux_h I__10275 (
            .O(N__66901),
            .I(N__66886));
    LocalMux I__10274 (
            .O(N__66898),
            .I(N__66886));
    Span4Mux_v I__10273 (
            .O(N__66895),
            .I(N__66883));
    InMux I__10272 (
            .O(N__66894),
            .I(N__66880));
    InMux I__10271 (
            .O(N__66891),
            .I(N__66877));
    Span4Mux_v I__10270 (
            .O(N__66886),
            .I(N__66874));
    Odrv4 I__10269 (
            .O(N__66883),
            .I(shift_srl_90Z0Z_15));
    LocalMux I__10268 (
            .O(N__66880),
            .I(shift_srl_90Z0Z_15));
    LocalMux I__10267 (
            .O(N__66877),
            .I(shift_srl_90Z0Z_15));
    Odrv4 I__10266 (
            .O(N__66874),
            .I(shift_srl_90Z0Z_15));
    CascadeMux I__10265 (
            .O(N__66865),
            .I(shift_srl_89_RNIPCQF1Z0Z_15_cascade_));
    CascadeMux I__10264 (
            .O(N__66862),
            .I(shift_srl_91_RNIOVG12Z0Z_15_cascade_));
    CascadeMux I__10263 (
            .O(N__66859),
            .I(rco_c_93_cascade_));
    InMux I__10262 (
            .O(N__66856),
            .I(N__66853));
    LocalMux I__10261 (
            .O(N__66853),
            .I(shift_srl_95Z0Z_9));
    InMux I__10260 (
            .O(N__66850),
            .I(N__66847));
    LocalMux I__10259 (
            .O(N__66847),
            .I(shift_srl_95Z0Z_8));
    InMux I__10258 (
            .O(N__66844),
            .I(N__66841));
    LocalMux I__10257 (
            .O(N__66841),
            .I(shift_srl_95Z0Z_0));
    InMux I__10256 (
            .O(N__66838),
            .I(N__66835));
    LocalMux I__10255 (
            .O(N__66835),
            .I(shift_srl_95Z0Z_1));
    InMux I__10254 (
            .O(N__66832),
            .I(N__66829));
    LocalMux I__10253 (
            .O(N__66829),
            .I(shift_srl_95Z0Z_2));
    InMux I__10252 (
            .O(N__66826),
            .I(N__66823));
    LocalMux I__10251 (
            .O(N__66823),
            .I(shift_srl_95Z0Z_3));
    InMux I__10250 (
            .O(N__66820),
            .I(N__66817));
    LocalMux I__10249 (
            .O(N__66817),
            .I(shift_srl_95Z0Z_4));
    InMux I__10248 (
            .O(N__66814),
            .I(N__66811));
    LocalMux I__10247 (
            .O(N__66811),
            .I(shift_srl_95Z0Z_5));
    CascadeMux I__10246 (
            .O(N__66808),
            .I(N__66801));
    InMux I__10245 (
            .O(N__66807),
            .I(N__66797));
    InMux I__10244 (
            .O(N__66806),
            .I(N__66794));
    InMux I__10243 (
            .O(N__66805),
            .I(N__66791));
    InMux I__10242 (
            .O(N__66804),
            .I(N__66784));
    InMux I__10241 (
            .O(N__66801),
            .I(N__66784));
    InMux I__10240 (
            .O(N__66800),
            .I(N__66784));
    LocalMux I__10239 (
            .O(N__66797),
            .I(N__66779));
    LocalMux I__10238 (
            .O(N__66794),
            .I(N__66779));
    LocalMux I__10237 (
            .O(N__66791),
            .I(N__66776));
    LocalMux I__10236 (
            .O(N__66784),
            .I(N__66773));
    Span12Mux_h I__10235 (
            .O(N__66779),
            .I(N__66770));
    Span4Mux_v I__10234 (
            .O(N__66776),
            .I(N__66767));
    Span4Mux_h I__10233 (
            .O(N__66773),
            .I(N__66764));
    Span12Mux_v I__10232 (
            .O(N__66770),
            .I(N__66761));
    Span4Mux_v I__10231 (
            .O(N__66767),
            .I(N__66756));
    Span4Mux_h I__10230 (
            .O(N__66764),
            .I(N__66756));
    Odrv12 I__10229 (
            .O(N__66761),
            .I(shift_srl_146_RNIVSUTZ0Z_15));
    Odrv4 I__10228 (
            .O(N__66756),
            .I(shift_srl_146_RNIVSUTZ0Z_15));
    IoInMux I__10227 (
            .O(N__66751),
            .I(N__66748));
    LocalMux I__10226 (
            .O(N__66748),
            .I(N__66745));
    Span12Mux_s3_v I__10225 (
            .O(N__66745),
            .I(N__66742));
    Odrv12 I__10224 (
            .O(N__66742),
            .I(rco_c_150));
    IoInMux I__10223 (
            .O(N__66739),
            .I(N__66736));
    LocalMux I__10222 (
            .O(N__66736),
            .I(N__66733));
    IoSpan4Mux I__10221 (
            .O(N__66733),
            .I(N__66730));
    Span4Mux_s3_v I__10220 (
            .O(N__66730),
            .I(N__66727));
    Odrv4 I__10219 (
            .O(N__66727),
            .I(rco_c_173));
    IoInMux I__10218 (
            .O(N__66724),
            .I(N__66721));
    LocalMux I__10217 (
            .O(N__66721),
            .I(N__66718));
    Span12Mux_s4_v I__10216 (
            .O(N__66718),
            .I(N__66715));
    Odrv12 I__10215 (
            .O(N__66715),
            .I(rco_c_176));
    IoInMux I__10214 (
            .O(N__66712),
            .I(N__66709));
    LocalMux I__10213 (
            .O(N__66709),
            .I(N__66706));
    Span12Mux_s4_v I__10212 (
            .O(N__66706),
            .I(N__66703));
    Odrv12 I__10211 (
            .O(N__66703),
            .I(rco_c_179));
    IoInMux I__10210 (
            .O(N__66700),
            .I(N__66697));
    LocalMux I__10209 (
            .O(N__66697),
            .I(N__66694));
    Span4Mux_s0_v I__10208 (
            .O(N__66694),
            .I(N__66691));
    Span4Mux_v I__10207 (
            .O(N__66691),
            .I(N__66688));
    Odrv4 I__10206 (
            .O(N__66688),
            .I(rco_c_182));
    InMux I__10205 (
            .O(N__66685),
            .I(N__66682));
    LocalMux I__10204 (
            .O(N__66682),
            .I(shift_srl_95Z0Z_10));
    InMux I__10203 (
            .O(N__66679),
            .I(N__66676));
    LocalMux I__10202 (
            .O(N__66676),
            .I(shift_srl_95Z0Z_11));
    InMux I__10201 (
            .O(N__66673),
            .I(N__66670));
    LocalMux I__10200 (
            .O(N__66670),
            .I(shift_srl_95Z0Z_12));
    InMux I__10199 (
            .O(N__66667),
            .I(N__66664));
    LocalMux I__10198 (
            .O(N__66664),
            .I(shift_srl_92Z0Z_14));
    InMux I__10197 (
            .O(N__66661),
            .I(N__66658));
    LocalMux I__10196 (
            .O(N__66658),
            .I(shift_srl_92Z0Z_9));
    InMux I__10195 (
            .O(N__66655),
            .I(N__66652));
    LocalMux I__10194 (
            .O(N__66652),
            .I(shift_srl_94Z0Z_8));
    InMux I__10193 (
            .O(N__66649),
            .I(N__66646));
    LocalMux I__10192 (
            .O(N__66646),
            .I(shift_srl_94Z0Z_9));
    InMux I__10191 (
            .O(N__66643),
            .I(N__66640));
    LocalMux I__10190 (
            .O(N__66640),
            .I(shift_srl_94Z0Z_7));
    InMux I__10189 (
            .O(N__66637),
            .I(N__66634));
    LocalMux I__10188 (
            .O(N__66634),
            .I(shift_srl_94Z0Z_6));
    InMux I__10187 (
            .O(N__66631),
            .I(N__66628));
    LocalMux I__10186 (
            .O(N__66628),
            .I(shift_srl_94Z0Z_5));
    InMux I__10185 (
            .O(N__66625),
            .I(N__66622));
    LocalMux I__10184 (
            .O(N__66622),
            .I(N__66618));
    InMux I__10183 (
            .O(N__66621),
            .I(N__66615));
    Span4Mux_h I__10182 (
            .O(N__66618),
            .I(N__66612));
    LocalMux I__10181 (
            .O(N__66615),
            .I(N__66608));
    Span4Mux_v I__10180 (
            .O(N__66612),
            .I(N__66604));
    InMux I__10179 (
            .O(N__66611),
            .I(N__66597));
    Span4Mux_v I__10178 (
            .O(N__66608),
            .I(N__66594));
    InMux I__10177 (
            .O(N__66607),
            .I(N__66591));
    Sp12to4 I__10176 (
            .O(N__66604),
            .I(N__66588));
    InMux I__10175 (
            .O(N__66603),
            .I(N__66579));
    InMux I__10174 (
            .O(N__66602),
            .I(N__66579));
    InMux I__10173 (
            .O(N__66601),
            .I(N__66579));
    InMux I__10172 (
            .O(N__66600),
            .I(N__66579));
    LocalMux I__10171 (
            .O(N__66597),
            .I(N__66576));
    Span4Mux_h I__10170 (
            .O(N__66594),
            .I(N__66571));
    LocalMux I__10169 (
            .O(N__66591),
            .I(N__66571));
    Odrv12 I__10168 (
            .O(N__66588),
            .I(shift_srl_141_RNI9SAMZ0Z_15));
    LocalMux I__10167 (
            .O(N__66579),
            .I(shift_srl_141_RNI9SAMZ0Z_15));
    Odrv4 I__10166 (
            .O(N__66576),
            .I(shift_srl_141_RNI9SAMZ0Z_15));
    Odrv4 I__10165 (
            .O(N__66571),
            .I(shift_srl_141_RNI9SAMZ0Z_15));
    IoInMux I__10164 (
            .O(N__66562),
            .I(N__66559));
    LocalMux I__10163 (
            .O(N__66559),
            .I(N__66556));
    Span4Mux_s0_v I__10162 (
            .O(N__66556),
            .I(N__66553));
    Span4Mux_v I__10161 (
            .O(N__66553),
            .I(N__66550));
    Odrv4 I__10160 (
            .O(N__66550),
            .I(rco_c_141));
    InMux I__10159 (
            .O(N__66547),
            .I(N__66544));
    LocalMux I__10158 (
            .O(N__66544),
            .I(N__66541));
    Span4Mux_h I__10157 (
            .O(N__66541),
            .I(N__66537));
    InMux I__10156 (
            .O(N__66540),
            .I(N__66533));
    Sp12to4 I__10155 (
            .O(N__66537),
            .I(N__66530));
    InMux I__10154 (
            .O(N__66536),
            .I(N__66527));
    LocalMux I__10153 (
            .O(N__66533),
            .I(N__66524));
    Span12Mux_v I__10152 (
            .O(N__66530),
            .I(N__66521));
    LocalMux I__10151 (
            .O(N__66527),
            .I(N__66516));
    Span4Mux_v I__10150 (
            .O(N__66524),
            .I(N__66516));
    Odrv12 I__10149 (
            .O(N__66521),
            .I(shift_srl_144_RNIIPPI1Z0Z_15));
    Odrv4 I__10148 (
            .O(N__66516),
            .I(shift_srl_144_RNIIPPI1Z0Z_15));
    IoInMux I__10147 (
            .O(N__66511),
            .I(N__66508));
    LocalMux I__10146 (
            .O(N__66508),
            .I(N__66505));
    Span4Mux_s0_v I__10145 (
            .O(N__66505),
            .I(N__66502));
    Span4Mux_v I__10144 (
            .O(N__66502),
            .I(N__66499));
    Odrv4 I__10143 (
            .O(N__66499),
            .I(rco_c_144));
    IoInMux I__10142 (
            .O(N__66496),
            .I(N__66492));
    InMux I__10141 (
            .O(N__66495),
            .I(N__66489));
    LocalMux I__10140 (
            .O(N__66492),
            .I(N__66486));
    LocalMux I__10139 (
            .O(N__66489),
            .I(N__66483));
    Span12Mux_s9_v I__10138 (
            .O(N__66486),
            .I(N__66480));
    Span4Mux_v I__10137 (
            .O(N__66483),
            .I(N__66477));
    Span12Mux_h I__10136 (
            .O(N__66480),
            .I(N__66474));
    Span4Mux_v I__10135 (
            .O(N__66477),
            .I(N__66471));
    Odrv12 I__10134 (
            .O(N__66474),
            .I(rco_c_116));
    Odrv4 I__10133 (
            .O(N__66471),
            .I(rco_c_116));
    InMux I__10132 (
            .O(N__66466),
            .I(N__66463));
    LocalMux I__10131 (
            .O(N__66463),
            .I(N__66457));
    CascadeMux I__10130 (
            .O(N__66462),
            .I(N__66451));
    InMux I__10129 (
            .O(N__66461),
            .I(N__66448));
    CascadeMux I__10128 (
            .O(N__66460),
            .I(N__66444));
    Span4Mux_v I__10127 (
            .O(N__66457),
            .I(N__66438));
    InMux I__10126 (
            .O(N__66456),
            .I(N__66433));
    InMux I__10125 (
            .O(N__66455),
            .I(N__66433));
    InMux I__10124 (
            .O(N__66454),
            .I(N__66430));
    InMux I__10123 (
            .O(N__66451),
            .I(N__66427));
    LocalMux I__10122 (
            .O(N__66448),
            .I(N__66424));
    InMux I__10121 (
            .O(N__66447),
            .I(N__66419));
    InMux I__10120 (
            .O(N__66444),
            .I(N__66419));
    InMux I__10119 (
            .O(N__66443),
            .I(N__66416));
    InMux I__10118 (
            .O(N__66442),
            .I(N__66412));
    InMux I__10117 (
            .O(N__66441),
            .I(N__66409));
    Span4Mux_h I__10116 (
            .O(N__66438),
            .I(N__66406));
    LocalMux I__10115 (
            .O(N__66433),
            .I(N__66403));
    LocalMux I__10114 (
            .O(N__66430),
            .I(N__66398));
    LocalMux I__10113 (
            .O(N__66427),
            .I(N__66398));
    Span4Mux_v I__10112 (
            .O(N__66424),
            .I(N__66393));
    LocalMux I__10111 (
            .O(N__66419),
            .I(N__66393));
    LocalMux I__10110 (
            .O(N__66416),
            .I(N__66388));
    InMux I__10109 (
            .O(N__66415),
            .I(N__66383));
    LocalMux I__10108 (
            .O(N__66412),
            .I(N__66380));
    LocalMux I__10107 (
            .O(N__66409),
            .I(N__66377));
    Span4Mux_v I__10106 (
            .O(N__66406),
            .I(N__66372));
    Span4Mux_h I__10105 (
            .O(N__66403),
            .I(N__66372));
    Span12Mux_s11_h I__10104 (
            .O(N__66398),
            .I(N__66369));
    Span4Mux_h I__10103 (
            .O(N__66393),
            .I(N__66366));
    InMux I__10102 (
            .O(N__66392),
            .I(N__66361));
    InMux I__10101 (
            .O(N__66391),
            .I(N__66361));
    Span12Mux_s11_h I__10100 (
            .O(N__66388),
            .I(N__66358));
    InMux I__10099 (
            .O(N__66387),
            .I(N__66353));
    InMux I__10098 (
            .O(N__66386),
            .I(N__66353));
    LocalMux I__10097 (
            .O(N__66383),
            .I(shift_srl_117Z0Z_15));
    Odrv4 I__10096 (
            .O(N__66380),
            .I(shift_srl_117Z0Z_15));
    Odrv4 I__10095 (
            .O(N__66377),
            .I(shift_srl_117Z0Z_15));
    Odrv4 I__10094 (
            .O(N__66372),
            .I(shift_srl_117Z0Z_15));
    Odrv12 I__10093 (
            .O(N__66369),
            .I(shift_srl_117Z0Z_15));
    Odrv4 I__10092 (
            .O(N__66366),
            .I(shift_srl_117Z0Z_15));
    LocalMux I__10091 (
            .O(N__66361),
            .I(shift_srl_117Z0Z_15));
    Odrv12 I__10090 (
            .O(N__66358),
            .I(shift_srl_117Z0Z_15));
    LocalMux I__10089 (
            .O(N__66353),
            .I(shift_srl_117Z0Z_15));
    IoInMux I__10088 (
            .O(N__66334),
            .I(N__66331));
    LocalMux I__10087 (
            .O(N__66331),
            .I(N__66328));
    IoSpan4Mux I__10086 (
            .O(N__66328),
            .I(N__66325));
    Span4Mux_s3_v I__10085 (
            .O(N__66325),
            .I(N__66322));
    Span4Mux_h I__10084 (
            .O(N__66322),
            .I(N__66319));
    Odrv4 I__10083 (
            .O(N__66319),
            .I(rco_c_117));
    IoInMux I__10082 (
            .O(N__66316),
            .I(N__66313));
    LocalMux I__10081 (
            .O(N__66313),
            .I(N__66310));
    IoSpan4Mux I__10080 (
            .O(N__66310),
            .I(N__66306));
    InMux I__10079 (
            .O(N__66309),
            .I(N__66303));
    Span4Mux_s3_v I__10078 (
            .O(N__66306),
            .I(N__66296));
    LocalMux I__10077 (
            .O(N__66303),
            .I(N__66293));
    InMux I__10076 (
            .O(N__66302),
            .I(N__66286));
    InMux I__10075 (
            .O(N__66301),
            .I(N__66286));
    InMux I__10074 (
            .O(N__66300),
            .I(N__66286));
    InMux I__10073 (
            .O(N__66299),
            .I(N__66283));
    Span4Mux_h I__10072 (
            .O(N__66296),
            .I(N__66278));
    Span4Mux_s3_v I__10071 (
            .O(N__66293),
            .I(N__66278));
    LocalMux I__10070 (
            .O(N__66286),
            .I(N__66273));
    LocalMux I__10069 (
            .O(N__66283),
            .I(N__66273));
    Span4Mux_h I__10068 (
            .O(N__66278),
            .I(N__66270));
    Span4Mux_v I__10067 (
            .O(N__66273),
            .I(N__66267));
    Span4Mux_v I__10066 (
            .O(N__66270),
            .I(N__66262));
    Span4Mux_h I__10065 (
            .O(N__66267),
            .I(N__66262));
    Odrv4 I__10064 (
            .O(N__66262),
            .I(rco_c_132));
    InMux I__10063 (
            .O(N__66259),
            .I(N__66254));
    InMux I__10062 (
            .O(N__66258),
            .I(N__66251));
    CascadeMux I__10061 (
            .O(N__66257),
            .I(N__66248));
    LocalMux I__10060 (
            .O(N__66254),
            .I(N__66245));
    LocalMux I__10059 (
            .O(N__66251),
            .I(N__66238));
    InMux I__10058 (
            .O(N__66248),
            .I(N__66234));
    Span4Mux_v I__10057 (
            .O(N__66245),
            .I(N__66231));
    InMux I__10056 (
            .O(N__66244),
            .I(N__66226));
    InMux I__10055 (
            .O(N__66243),
            .I(N__66226));
    InMux I__10054 (
            .O(N__66242),
            .I(N__66223));
    InMux I__10053 (
            .O(N__66241),
            .I(N__66220));
    Span12Mux_v I__10052 (
            .O(N__66238),
            .I(N__66217));
    CascadeMux I__10051 (
            .O(N__66237),
            .I(N__66214));
    LocalMux I__10050 (
            .O(N__66234),
            .I(N__66211));
    Span4Mux_h I__10049 (
            .O(N__66231),
            .I(N__66202));
    LocalMux I__10048 (
            .O(N__66226),
            .I(N__66202));
    LocalMux I__10047 (
            .O(N__66223),
            .I(N__66202));
    LocalMux I__10046 (
            .O(N__66220),
            .I(N__66202));
    Span12Mux_h I__10045 (
            .O(N__66217),
            .I(N__66199));
    InMux I__10044 (
            .O(N__66214),
            .I(N__66196));
    Span4Mux_h I__10043 (
            .O(N__66211),
            .I(N__66191));
    Span4Mux_v I__10042 (
            .O(N__66202),
            .I(N__66191));
    Odrv12 I__10041 (
            .O(N__66199),
            .I(shift_srl_133Z0Z_15));
    LocalMux I__10040 (
            .O(N__66196),
            .I(shift_srl_133Z0Z_15));
    Odrv4 I__10039 (
            .O(N__66191),
            .I(shift_srl_133Z0Z_15));
    IoInMux I__10038 (
            .O(N__66184),
            .I(N__66181));
    LocalMux I__10037 (
            .O(N__66181),
            .I(N__66178));
    Span4Mux_s2_v I__10036 (
            .O(N__66178),
            .I(N__66175));
    Span4Mux_h I__10035 (
            .O(N__66175),
            .I(N__66172));
    Odrv4 I__10034 (
            .O(N__66172),
            .I(rco_c_133));
    IoInMux I__10033 (
            .O(N__66169),
            .I(N__66166));
    LocalMux I__10032 (
            .O(N__66166),
            .I(N__66163));
    IoSpan4Mux I__10031 (
            .O(N__66163),
            .I(N__66160));
    Odrv4 I__10030 (
            .O(N__66160),
            .I(rco_c_58));
    IoInMux I__10029 (
            .O(N__66157),
            .I(N__66154));
    LocalMux I__10028 (
            .O(N__66154),
            .I(N__66151));
    Span4Mux_s1_v I__10027 (
            .O(N__66151),
            .I(N__66148));
    Span4Mux_h I__10026 (
            .O(N__66148),
            .I(N__66145));
    Odrv4 I__10025 (
            .O(N__66145),
            .I(rco_c_85));
    InMux I__10024 (
            .O(N__66142),
            .I(N__66139));
    LocalMux I__10023 (
            .O(N__66139),
            .I(shift_srl_92Z0Z_10));
    InMux I__10022 (
            .O(N__66136),
            .I(N__66133));
    LocalMux I__10021 (
            .O(N__66133),
            .I(shift_srl_92Z0Z_11));
    InMux I__10020 (
            .O(N__66130),
            .I(N__66127));
    LocalMux I__10019 (
            .O(N__66127),
            .I(shift_srl_92Z0Z_12));
    InMux I__10018 (
            .O(N__66124),
            .I(N__66121));
    LocalMux I__10017 (
            .O(N__66121),
            .I(shift_srl_92Z0Z_13));
    InMux I__10016 (
            .O(N__66118),
            .I(N__66115));
    LocalMux I__10015 (
            .O(N__66115),
            .I(shift_srl_119Z0Z_10));
    InMux I__10014 (
            .O(N__66112),
            .I(N__66109));
    LocalMux I__10013 (
            .O(N__66109),
            .I(N__66106));
    Odrv4 I__10012 (
            .O(N__66106),
            .I(shift_srl_119Z0Z_13));
    InMux I__10011 (
            .O(N__66103),
            .I(N__66100));
    LocalMux I__10010 (
            .O(N__66100),
            .I(shift_srl_119Z0Z_9));
    InMux I__10009 (
            .O(N__66097),
            .I(N__66094));
    LocalMux I__10008 (
            .O(N__66094),
            .I(shift_srl_119Z0Z_8));
    InMux I__10007 (
            .O(N__66091),
            .I(N__66088));
    LocalMux I__10006 (
            .O(N__66088),
            .I(shift_srl_119Z0Z_4));
    InMux I__10005 (
            .O(N__66085),
            .I(N__66082));
    LocalMux I__10004 (
            .O(N__66082),
            .I(shift_srl_40Z0Z_8));
    InMux I__10003 (
            .O(N__66079),
            .I(N__66076));
    LocalMux I__10002 (
            .O(N__66076),
            .I(shift_srl_40Z0Z_7));
    InMux I__10001 (
            .O(N__66073),
            .I(N__66070));
    LocalMux I__10000 (
            .O(N__66070),
            .I(N__66067));
    Span4Mux_h I__9999 (
            .O(N__66067),
            .I(N__66064));
    Span4Mux_h I__9998 (
            .O(N__66064),
            .I(N__66058));
    InMux I__9997 (
            .O(N__66063),
            .I(N__66053));
    InMux I__9996 (
            .O(N__66062),
            .I(N__66053));
    InMux I__9995 (
            .O(N__66061),
            .I(N__66050));
    Span4Mux_v I__9994 (
            .O(N__66058),
            .I(N__66047));
    LocalMux I__9993 (
            .O(N__66053),
            .I(N__66044));
    LocalMux I__9992 (
            .O(N__66050),
            .I(shift_srl_126Z0Z_15));
    Odrv4 I__9991 (
            .O(N__66047),
            .I(shift_srl_126Z0Z_15));
    Odrv4 I__9990 (
            .O(N__66044),
            .I(shift_srl_126Z0Z_15));
    InMux I__9989 (
            .O(N__66037),
            .I(N__66033));
    InMux I__9988 (
            .O(N__66036),
            .I(N__66030));
    LocalMux I__9987 (
            .O(N__66033),
            .I(N__66025));
    LocalMux I__9986 (
            .O(N__66030),
            .I(N__66022));
    CascadeMux I__9985 (
            .O(N__66029),
            .I(N__66019));
    CascadeMux I__9984 (
            .O(N__66028),
            .I(N__66016));
    Span4Mux_h I__9983 (
            .O(N__66025),
            .I(N__66011));
    Span4Mux_h I__9982 (
            .O(N__66022),
            .I(N__66008));
    InMux I__9981 (
            .O(N__66019),
            .I(N__66005));
    InMux I__9980 (
            .O(N__66016),
            .I(N__66000));
    InMux I__9979 (
            .O(N__66015),
            .I(N__66000));
    InMux I__9978 (
            .O(N__66014),
            .I(N__65997));
    Span4Mux_h I__9977 (
            .O(N__66011),
            .I(N__65992));
    Span4Mux_h I__9976 (
            .O(N__66008),
            .I(N__65992));
    LocalMux I__9975 (
            .O(N__66005),
            .I(N__65987));
    LocalMux I__9974 (
            .O(N__66000),
            .I(N__65987));
    LocalMux I__9973 (
            .O(N__65997),
            .I(shift_srl_125Z0Z_15));
    Odrv4 I__9972 (
            .O(N__65992),
            .I(shift_srl_125Z0Z_15));
    Odrv4 I__9971 (
            .O(N__65987),
            .I(shift_srl_125Z0Z_15));
    CascadeMux I__9970 (
            .O(N__65980),
            .I(clk_en_0_a3_0_a2_1_127_cascade_));
    IoInMux I__9969 (
            .O(N__65977),
            .I(N__65974));
    LocalMux I__9968 (
            .O(N__65974),
            .I(N__65967));
    InMux I__9967 (
            .O(N__65973),
            .I(N__65962));
    InMux I__9966 (
            .O(N__65972),
            .I(N__65962));
    InMux I__9965 (
            .O(N__65971),
            .I(N__65957));
    InMux I__9964 (
            .O(N__65970),
            .I(N__65957));
    Span12Mux_s8_h I__9963 (
            .O(N__65967),
            .I(N__65954));
    LocalMux I__9962 (
            .O(N__65962),
            .I(N__65949));
    LocalMux I__9961 (
            .O(N__65957),
            .I(N__65949));
    Span12Mux_h I__9960 (
            .O(N__65954),
            .I(N__65944));
    Span4Mux_v I__9959 (
            .O(N__65949),
            .I(N__65941));
    InMux I__9958 (
            .O(N__65948),
            .I(N__65936));
    InMux I__9957 (
            .O(N__65947),
            .I(N__65936));
    Odrv12 I__9956 (
            .O(N__65944),
            .I(rco_c_118));
    Odrv4 I__9955 (
            .O(N__65941),
            .I(rco_c_118));
    LocalMux I__9954 (
            .O(N__65936),
            .I(rco_c_118));
    InMux I__9953 (
            .O(N__65929),
            .I(N__65926));
    LocalMux I__9952 (
            .O(N__65926),
            .I(shift_srl_119Z0Z_14));
    InMux I__9951 (
            .O(N__65923),
            .I(N__65920));
    LocalMux I__9950 (
            .O(N__65920),
            .I(N__65917));
    Span4Mux_h I__9949 (
            .O(N__65917),
            .I(N__65914));
    Odrv4 I__9948 (
            .O(N__65914),
            .I(clk_en_0_a3_0_a2_sx_119));
    InMux I__9947 (
            .O(N__65911),
            .I(N__65908));
    LocalMux I__9946 (
            .O(N__65908),
            .I(N__65905));
    Span4Mux_v I__9945 (
            .O(N__65905),
            .I(N__65899));
    InMux I__9944 (
            .O(N__65904),
            .I(N__65896));
    InMux I__9943 (
            .O(N__65903),
            .I(N__65891));
    InMux I__9942 (
            .O(N__65902),
            .I(N__65891));
    Span4Mux_h I__9941 (
            .O(N__65899),
            .I(N__65883));
    LocalMux I__9940 (
            .O(N__65896),
            .I(N__65883));
    LocalMux I__9939 (
            .O(N__65891),
            .I(N__65883));
    CascadeMux I__9938 (
            .O(N__65890),
            .I(N__65879));
    Span4Mux_v I__9937 (
            .O(N__65883),
            .I(N__65876));
    InMux I__9936 (
            .O(N__65882),
            .I(N__65871));
    InMux I__9935 (
            .O(N__65879),
            .I(N__65871));
    Odrv4 I__9934 (
            .O(N__65876),
            .I(rco_int_0_a2_1_a2_0_0_116));
    LocalMux I__9933 (
            .O(N__65871),
            .I(rco_int_0_a2_1_a2_0_0_116));
    InMux I__9932 (
            .O(N__65866),
            .I(N__65863));
    LocalMux I__9931 (
            .O(N__65863),
            .I(N__65860));
    Span4Mux_s3_h I__9930 (
            .O(N__65860),
            .I(N__65856));
    CascadeMux I__9929 (
            .O(N__65859),
            .I(N__65852));
    Span4Mux_h I__9928 (
            .O(N__65856),
            .I(N__65848));
    InMux I__9927 (
            .O(N__65855),
            .I(N__65845));
    InMux I__9926 (
            .O(N__65852),
            .I(N__65838));
    InMux I__9925 (
            .O(N__65851),
            .I(N__65838));
    Span4Mux_h I__9924 (
            .O(N__65848),
            .I(N__65833));
    LocalMux I__9923 (
            .O(N__65845),
            .I(N__65833));
    InMux I__9922 (
            .O(N__65844),
            .I(N__65830));
    InMux I__9921 (
            .O(N__65843),
            .I(N__65827));
    LocalMux I__9920 (
            .O(N__65838),
            .I(N__65822));
    Span4Mux_h I__9919 (
            .O(N__65833),
            .I(N__65822));
    LocalMux I__9918 (
            .O(N__65830),
            .I(shift_srl_119Z0Z_15));
    LocalMux I__9917 (
            .O(N__65827),
            .I(shift_srl_119Z0Z_15));
    Odrv4 I__9916 (
            .O(N__65822),
            .I(shift_srl_119Z0Z_15));
    InMux I__9915 (
            .O(N__65815),
            .I(N__65812));
    LocalMux I__9914 (
            .O(N__65812),
            .I(shift_srl_119Z0Z_0));
    InMux I__9913 (
            .O(N__65809),
            .I(N__65806));
    LocalMux I__9912 (
            .O(N__65806),
            .I(shift_srl_119Z0Z_1));
    InMux I__9911 (
            .O(N__65803),
            .I(N__65800));
    LocalMux I__9910 (
            .O(N__65800),
            .I(shift_srl_119Z0Z_2));
    InMux I__9909 (
            .O(N__65797),
            .I(N__65794));
    LocalMux I__9908 (
            .O(N__65794),
            .I(shift_srl_119Z0Z_3));
    InMux I__9907 (
            .O(N__65791),
            .I(N__65788));
    LocalMux I__9906 (
            .O(N__65788),
            .I(shift_srl_127Z0Z_11));
    InMux I__9905 (
            .O(N__65785),
            .I(N__65782));
    LocalMux I__9904 (
            .O(N__65782),
            .I(shift_srl_127Z0Z_12));
    InMux I__9903 (
            .O(N__65779),
            .I(N__65776));
    LocalMux I__9902 (
            .O(N__65776),
            .I(shift_srl_127Z0Z_13));
    InMux I__9901 (
            .O(N__65773),
            .I(N__65770));
    LocalMux I__9900 (
            .O(N__65770),
            .I(shift_srl_127Z0Z_14));
    InMux I__9899 (
            .O(N__65767),
            .I(N__65764));
    LocalMux I__9898 (
            .O(N__65764),
            .I(shift_srl_127Z0Z_9));
    InMux I__9897 (
            .O(N__65761),
            .I(N__65758));
    LocalMux I__9896 (
            .O(N__65758),
            .I(shift_srl_127Z0Z_8));
    CascadeMux I__9895 (
            .O(N__65755),
            .I(N__65747));
    CascadeMux I__9894 (
            .O(N__65754),
            .I(N__65743));
    InMux I__9893 (
            .O(N__65753),
            .I(N__65734));
    InMux I__9892 (
            .O(N__65752),
            .I(N__65734));
    InMux I__9891 (
            .O(N__65751),
            .I(N__65729));
    InMux I__9890 (
            .O(N__65750),
            .I(N__65729));
    InMux I__9889 (
            .O(N__65747),
            .I(N__65725));
    InMux I__9888 (
            .O(N__65746),
            .I(N__65718));
    InMux I__9887 (
            .O(N__65743),
            .I(N__65718));
    InMux I__9886 (
            .O(N__65742),
            .I(N__65718));
    InMux I__9885 (
            .O(N__65741),
            .I(N__65713));
    InMux I__9884 (
            .O(N__65740),
            .I(N__65710));
    InMux I__9883 (
            .O(N__65739),
            .I(N__65706));
    LocalMux I__9882 (
            .O(N__65734),
            .I(N__65703));
    LocalMux I__9881 (
            .O(N__65729),
            .I(N__65700));
    InMux I__9880 (
            .O(N__65728),
            .I(N__65697));
    LocalMux I__9879 (
            .O(N__65725),
            .I(N__65692));
    LocalMux I__9878 (
            .O(N__65718),
            .I(N__65692));
    InMux I__9877 (
            .O(N__65717),
            .I(N__65689));
    InMux I__9876 (
            .O(N__65716),
            .I(N__65686));
    LocalMux I__9875 (
            .O(N__65713),
            .I(N__65683));
    LocalMux I__9874 (
            .O(N__65710),
            .I(N__65680));
    InMux I__9873 (
            .O(N__65709),
            .I(N__65677));
    LocalMux I__9872 (
            .O(N__65706),
            .I(N__65674));
    Span4Mux_v I__9871 (
            .O(N__65703),
            .I(N__65669));
    Span4Mux_s2_h I__9870 (
            .O(N__65700),
            .I(N__65669));
    LocalMux I__9869 (
            .O(N__65697),
            .I(N__65662));
    Span4Mux_h I__9868 (
            .O(N__65692),
            .I(N__65662));
    LocalMux I__9867 (
            .O(N__65689),
            .I(N__65662));
    LocalMux I__9866 (
            .O(N__65686),
            .I(N__65659));
    Span4Mux_h I__9865 (
            .O(N__65683),
            .I(N__65655));
    Span4Mux_h I__9864 (
            .O(N__65680),
            .I(N__65652));
    LocalMux I__9863 (
            .O(N__65677),
            .I(N__65649));
    Span4Mux_v I__9862 (
            .O(N__65674),
            .I(N__65646));
    Span4Mux_h I__9861 (
            .O(N__65669),
            .I(N__65641));
    Span4Mux_v I__9860 (
            .O(N__65662),
            .I(N__65641));
    Span12Mux_h I__9859 (
            .O(N__65659),
            .I(N__65638));
    InMux I__9858 (
            .O(N__65658),
            .I(N__65635));
    Span4Mux_v I__9857 (
            .O(N__65655),
            .I(N__65630));
    Span4Mux_h I__9856 (
            .O(N__65652),
            .I(N__65630));
    Span4Mux_v I__9855 (
            .O(N__65649),
            .I(N__65623));
    Span4Mux_v I__9854 (
            .O(N__65646),
            .I(N__65623));
    Span4Mux_h I__9853 (
            .O(N__65641),
            .I(N__65623));
    Odrv12 I__9852 (
            .O(N__65638),
            .I(rco_int_0_a2_1_a2_0_127));
    LocalMux I__9851 (
            .O(N__65635),
            .I(rco_int_0_a2_1_a2_0_127));
    Odrv4 I__9850 (
            .O(N__65630),
            .I(rco_int_0_a2_1_a2_0_127));
    Odrv4 I__9849 (
            .O(N__65623),
            .I(rco_int_0_a2_1_a2_0_127));
    InMux I__9848 (
            .O(N__65614),
            .I(N__65611));
    LocalMux I__9847 (
            .O(N__65611),
            .I(N__65608));
    Span4Mux_h I__9846 (
            .O(N__65608),
            .I(N__65605));
    Span4Mux_h I__9845 (
            .O(N__65605),
            .I(N__65599));
    InMux I__9844 (
            .O(N__65604),
            .I(N__65596));
    CascadeMux I__9843 (
            .O(N__65603),
            .I(N__65593));
    InMux I__9842 (
            .O(N__65602),
            .I(N__65590));
    Span4Mux_h I__9841 (
            .O(N__65599),
            .I(N__65587));
    LocalMux I__9840 (
            .O(N__65596),
            .I(N__65584));
    InMux I__9839 (
            .O(N__65593),
            .I(N__65581));
    LocalMux I__9838 (
            .O(N__65590),
            .I(shift_srl_120Z0Z_15));
    Odrv4 I__9837 (
            .O(N__65587),
            .I(shift_srl_120Z0Z_15));
    Odrv4 I__9836 (
            .O(N__65584),
            .I(shift_srl_120Z0Z_15));
    LocalMux I__9835 (
            .O(N__65581),
            .I(shift_srl_120Z0Z_15));
    CascadeMux I__9834 (
            .O(N__65572),
            .I(N__65569));
    InMux I__9833 (
            .O(N__65569),
            .I(N__65563));
    InMux I__9832 (
            .O(N__65568),
            .I(N__65560));
    InMux I__9831 (
            .O(N__65567),
            .I(N__65557));
    CascadeMux I__9830 (
            .O(N__65566),
            .I(N__65554));
    LocalMux I__9829 (
            .O(N__65563),
            .I(N__65547));
    LocalMux I__9828 (
            .O(N__65560),
            .I(N__65544));
    LocalMux I__9827 (
            .O(N__65557),
            .I(N__65541));
    InMux I__9826 (
            .O(N__65554),
            .I(N__65538));
    InMux I__9825 (
            .O(N__65553),
            .I(N__65533));
    InMux I__9824 (
            .O(N__65552),
            .I(N__65533));
    InMux I__9823 (
            .O(N__65551),
            .I(N__65530));
    CascadeMux I__9822 (
            .O(N__65550),
            .I(N__65527));
    Span4Mux_v I__9821 (
            .O(N__65547),
            .I(N__65524));
    Span4Mux_v I__9820 (
            .O(N__65544),
            .I(N__65518));
    Span4Mux_v I__9819 (
            .O(N__65541),
            .I(N__65518));
    LocalMux I__9818 (
            .O(N__65538),
            .I(N__65515));
    LocalMux I__9817 (
            .O(N__65533),
            .I(N__65511));
    LocalMux I__9816 (
            .O(N__65530),
            .I(N__65508));
    InMux I__9815 (
            .O(N__65527),
            .I(N__65505));
    Span4Mux_h I__9814 (
            .O(N__65524),
            .I(N__65502));
    InMux I__9813 (
            .O(N__65523),
            .I(N__65499));
    Sp12to4 I__9812 (
            .O(N__65518),
            .I(N__65496));
    Span12Mux_v I__9811 (
            .O(N__65515),
            .I(N__65493));
    InMux I__9810 (
            .O(N__65514),
            .I(N__65490));
    Span4Mux_h I__9809 (
            .O(N__65511),
            .I(N__65485));
    Span4Mux_h I__9808 (
            .O(N__65508),
            .I(N__65485));
    LocalMux I__9807 (
            .O(N__65505),
            .I(N__65482));
    Span4Mux_h I__9806 (
            .O(N__65502),
            .I(N__65477));
    LocalMux I__9805 (
            .O(N__65499),
            .I(N__65477));
    Span12Mux_h I__9804 (
            .O(N__65496),
            .I(N__65474));
    Span12Mux_h I__9803 (
            .O(N__65493),
            .I(N__65471));
    LocalMux I__9802 (
            .O(N__65490),
            .I(rco_int_0_a2_1_a2_0_120));
    Odrv4 I__9801 (
            .O(N__65485),
            .I(rco_int_0_a2_1_a2_0_120));
    Odrv12 I__9800 (
            .O(N__65482),
            .I(rco_int_0_a2_1_a2_0_120));
    Odrv4 I__9799 (
            .O(N__65477),
            .I(rco_int_0_a2_1_a2_0_120));
    Odrv12 I__9798 (
            .O(N__65474),
            .I(rco_int_0_a2_1_a2_0_120));
    Odrv12 I__9797 (
            .O(N__65471),
            .I(rco_int_0_a2_1_a2_0_120));
    InMux I__9796 (
            .O(N__65458),
            .I(N__65454));
    InMux I__9795 (
            .O(N__65457),
            .I(N__65450));
    LocalMux I__9794 (
            .O(N__65454),
            .I(N__65447));
    InMux I__9793 (
            .O(N__65453),
            .I(N__65444));
    LocalMux I__9792 (
            .O(N__65450),
            .I(N__65441));
    Span4Mux_v I__9791 (
            .O(N__65447),
            .I(N__65436));
    LocalMux I__9790 (
            .O(N__65444),
            .I(N__65433));
    Span4Mux_v I__9789 (
            .O(N__65441),
            .I(N__65430));
    InMux I__9788 (
            .O(N__65440),
            .I(N__65427));
    InMux I__9787 (
            .O(N__65439),
            .I(N__65424));
    Span4Mux_h I__9786 (
            .O(N__65436),
            .I(N__65421));
    Span4Mux_v I__9785 (
            .O(N__65433),
            .I(N__65418));
    Span4Mux_h I__9784 (
            .O(N__65430),
            .I(N__65413));
    LocalMux I__9783 (
            .O(N__65427),
            .I(N__65413));
    LocalMux I__9782 (
            .O(N__65424),
            .I(N__65407));
    Span4Mux_h I__9781 (
            .O(N__65421),
            .I(N__65402));
    Span4Mux_h I__9780 (
            .O(N__65418),
            .I(N__65402));
    Span4Mux_v I__9779 (
            .O(N__65413),
            .I(N__65399));
    InMux I__9778 (
            .O(N__65412),
            .I(N__65392));
    InMux I__9777 (
            .O(N__65411),
            .I(N__65392));
    InMux I__9776 (
            .O(N__65410),
            .I(N__65392));
    Odrv4 I__9775 (
            .O(N__65407),
            .I(shift_srl_124Z0Z_15));
    Odrv4 I__9774 (
            .O(N__65402),
            .I(shift_srl_124Z0Z_15));
    Odrv4 I__9773 (
            .O(N__65399),
            .I(shift_srl_124Z0Z_15));
    LocalMux I__9772 (
            .O(N__65392),
            .I(shift_srl_124Z0Z_15));
    CascadeMux I__9771 (
            .O(N__65383),
            .I(rco_int_0_a2_1_a2_0_120_cascade_));
    CascadeMux I__9770 (
            .O(N__65380),
            .I(N__65376));
    CascadeMux I__9769 (
            .O(N__65379),
            .I(N__65371));
    InMux I__9768 (
            .O(N__65376),
            .I(N__65365));
    InMux I__9767 (
            .O(N__65375),
            .I(N__65365));
    InMux I__9766 (
            .O(N__65374),
            .I(N__65359));
    InMux I__9765 (
            .O(N__65371),
            .I(N__65355));
    InMux I__9764 (
            .O(N__65370),
            .I(N__65352));
    LocalMux I__9763 (
            .O(N__65365),
            .I(N__65349));
    InMux I__9762 (
            .O(N__65364),
            .I(N__65345));
    InMux I__9761 (
            .O(N__65363),
            .I(N__65342));
    InMux I__9760 (
            .O(N__65362),
            .I(N__65338));
    LocalMux I__9759 (
            .O(N__65359),
            .I(N__65335));
    InMux I__9758 (
            .O(N__65358),
            .I(N__65332));
    LocalMux I__9757 (
            .O(N__65355),
            .I(N__65329));
    LocalMux I__9756 (
            .O(N__65352),
            .I(N__65326));
    Span4Mux_h I__9755 (
            .O(N__65349),
            .I(N__65323));
    InMux I__9754 (
            .O(N__65348),
            .I(N__65320));
    LocalMux I__9753 (
            .O(N__65345),
            .I(N__65317));
    LocalMux I__9752 (
            .O(N__65342),
            .I(N__65314));
    InMux I__9751 (
            .O(N__65341),
            .I(N__65311));
    LocalMux I__9750 (
            .O(N__65338),
            .I(N__65307));
    Span4Mux_v I__9749 (
            .O(N__65335),
            .I(N__65302));
    LocalMux I__9748 (
            .O(N__65332),
            .I(N__65302));
    Span4Mux_v I__9747 (
            .O(N__65329),
            .I(N__65294));
    Span4Mux_h I__9746 (
            .O(N__65326),
            .I(N__65294));
    Span4Mux_h I__9745 (
            .O(N__65323),
            .I(N__65294));
    LocalMux I__9744 (
            .O(N__65320),
            .I(N__65291));
    Span4Mux_v I__9743 (
            .O(N__65317),
            .I(N__65286));
    Span4Mux_s2_h I__9742 (
            .O(N__65314),
            .I(N__65286));
    LocalMux I__9741 (
            .O(N__65311),
            .I(N__65283));
    InMux I__9740 (
            .O(N__65310),
            .I(N__65280));
    Span4Mux_v I__9739 (
            .O(N__65307),
            .I(N__65277));
    Span4Mux_v I__9738 (
            .O(N__65302),
            .I(N__65274));
    InMux I__9737 (
            .O(N__65301),
            .I(N__65271));
    Span4Mux_v I__9736 (
            .O(N__65294),
            .I(N__65268));
    Span4Mux_v I__9735 (
            .O(N__65291),
            .I(N__65261));
    Span4Mux_h I__9734 (
            .O(N__65286),
            .I(N__65261));
    Span4Mux_h I__9733 (
            .O(N__65283),
            .I(N__65261));
    LocalMux I__9732 (
            .O(N__65280),
            .I(N__65254));
    Span4Mux_h I__9731 (
            .O(N__65277),
            .I(N__65254));
    Span4Mux_h I__9730 (
            .O(N__65274),
            .I(N__65254));
    LocalMux I__9729 (
            .O(N__65271),
            .I(rco_int_0_a2_1_a2_0_123));
    Odrv4 I__9728 (
            .O(N__65268),
            .I(rco_int_0_a2_1_a2_0_123));
    Odrv4 I__9727 (
            .O(N__65261),
            .I(rco_int_0_a2_1_a2_0_123));
    Odrv4 I__9726 (
            .O(N__65254),
            .I(rco_int_0_a2_1_a2_0_123));
    InMux I__9725 (
            .O(N__65245),
            .I(N__65242));
    LocalMux I__9724 (
            .O(N__65242),
            .I(shift_srl_120Z0Z_5));
    InMux I__9723 (
            .O(N__65239),
            .I(N__65236));
    LocalMux I__9722 (
            .O(N__65236),
            .I(shift_srl_120Z0Z_3));
    InMux I__9721 (
            .O(N__65233),
            .I(N__65230));
    LocalMux I__9720 (
            .O(N__65230),
            .I(shift_srl_120Z0Z_4));
    IoInMux I__9719 (
            .O(N__65227),
            .I(N__65224));
    LocalMux I__9718 (
            .O(N__65224),
            .I(N__65221));
    IoSpan4Mux I__9717 (
            .O(N__65221),
            .I(N__65218));
    Sp12to4 I__9716 (
            .O(N__65218),
            .I(N__65215));
    Span12Mux_s9_h I__9715 (
            .O(N__65215),
            .I(N__65212));
    Odrv12 I__9714 (
            .O(N__65212),
            .I(rco_c_119));
    InMux I__9713 (
            .O(N__65209),
            .I(N__65206));
    LocalMux I__9712 (
            .O(N__65206),
            .I(shift_srl_120Z0Z_0));
    InMux I__9711 (
            .O(N__65203),
            .I(N__65200));
    LocalMux I__9710 (
            .O(N__65200),
            .I(shift_srl_120Z0Z_1));
    InMux I__9709 (
            .O(N__65197),
            .I(N__65194));
    LocalMux I__9708 (
            .O(N__65194),
            .I(shift_srl_120Z0Z_2));
    CEMux I__9707 (
            .O(N__65191),
            .I(N__65187));
    CEMux I__9706 (
            .O(N__65190),
            .I(N__65183));
    LocalMux I__9705 (
            .O(N__65187),
            .I(N__65180));
    CEMux I__9704 (
            .O(N__65186),
            .I(N__65177));
    LocalMux I__9703 (
            .O(N__65183),
            .I(N__65174));
    Span4Mux_v I__9702 (
            .O(N__65180),
            .I(N__65171));
    LocalMux I__9701 (
            .O(N__65177),
            .I(N__65168));
    Odrv12 I__9700 (
            .O(N__65174),
            .I(clk_en_120));
    Odrv4 I__9699 (
            .O(N__65171),
            .I(clk_en_120));
    Odrv4 I__9698 (
            .O(N__65168),
            .I(clk_en_120));
    InMux I__9697 (
            .O(N__65161),
            .I(N__65158));
    LocalMux I__9696 (
            .O(N__65158),
            .I(shift_srl_127Z0Z_10));
    InMux I__9695 (
            .O(N__65155),
            .I(N__65152));
    LocalMux I__9694 (
            .O(N__65152),
            .I(shift_srl_162Z0Z_10));
    InMux I__9693 (
            .O(N__65149),
            .I(N__65146));
    LocalMux I__9692 (
            .O(N__65146),
            .I(shift_srl_162Z0Z_6));
    InMux I__9691 (
            .O(N__65143),
            .I(N__65140));
    LocalMux I__9690 (
            .O(N__65140),
            .I(shift_srl_162Z0Z_14));
    InMux I__9689 (
            .O(N__65137),
            .I(N__65134));
    LocalMux I__9688 (
            .O(N__65134),
            .I(shift_srl_162Z0Z_9));
    InMux I__9687 (
            .O(N__65131),
            .I(N__65128));
    LocalMux I__9686 (
            .O(N__65128),
            .I(shift_srl_162Z0Z_7));
    InMux I__9685 (
            .O(N__65125),
            .I(N__65122));
    LocalMux I__9684 (
            .O(N__65122),
            .I(shift_srl_162Z0Z_8));
    InMux I__9683 (
            .O(N__65119),
            .I(N__65116));
    LocalMux I__9682 (
            .O(N__65116),
            .I(shift_srl_120Z0Z_6));
    InMux I__9681 (
            .O(N__65113),
            .I(N__65110));
    LocalMux I__9680 (
            .O(N__65110),
            .I(shift_srl_120Z0Z_7));
    InMux I__9679 (
            .O(N__65107),
            .I(N__65104));
    LocalMux I__9678 (
            .O(N__65104),
            .I(shift_srl_28Z0Z_7));
    InMux I__9677 (
            .O(N__65101),
            .I(N__65098));
    LocalMux I__9676 (
            .O(N__65098),
            .I(N__65095));
    Span4Mux_h I__9675 (
            .O(N__65095),
            .I(N__65092));
    Odrv4 I__9674 (
            .O(N__65092),
            .I(shift_srl_117Z0Z_7));
    InMux I__9673 (
            .O(N__65089),
            .I(N__65086));
    LocalMux I__9672 (
            .O(N__65086),
            .I(shift_srl_117Z0Z_8));
    InMux I__9671 (
            .O(N__65083),
            .I(N__65080));
    LocalMux I__9670 (
            .O(N__65080),
            .I(N__65077));
    Span4Mux_v I__9669 (
            .O(N__65077),
            .I(N__65074));
    Span4Mux_h I__9668 (
            .O(N__65074),
            .I(N__65071));
    Odrv4 I__9667 (
            .O(N__65071),
            .I(shift_srl_117Z0Z_9));
    CEMux I__9666 (
            .O(N__65068),
            .I(N__65065));
    LocalMux I__9665 (
            .O(N__65065),
            .I(N__65061));
    CEMux I__9664 (
            .O(N__65064),
            .I(N__65057));
    Span4Mux_v I__9663 (
            .O(N__65061),
            .I(N__65054));
    CEMux I__9662 (
            .O(N__65060),
            .I(N__65051));
    LocalMux I__9661 (
            .O(N__65057),
            .I(N__65048));
    Span4Mux_h I__9660 (
            .O(N__65054),
            .I(N__65043));
    LocalMux I__9659 (
            .O(N__65051),
            .I(N__65043));
    Span4Mux_v I__9658 (
            .O(N__65048),
            .I(N__65040));
    Span4Mux_h I__9657 (
            .O(N__65043),
            .I(N__65037));
    Odrv4 I__9656 (
            .O(N__65040),
            .I(clk_en_117));
    Odrv4 I__9655 (
            .O(N__65037),
            .I(clk_en_117));
    InMux I__9654 (
            .O(N__65032),
            .I(N__65029));
    LocalMux I__9653 (
            .O(N__65029),
            .I(N__65024));
    InMux I__9652 (
            .O(N__65028),
            .I(N__65017));
    InMux I__9651 (
            .O(N__65027),
            .I(N__65014));
    Span4Mux_v I__9650 (
            .O(N__65024),
            .I(N__65011));
    InMux I__9649 (
            .O(N__65023),
            .I(N__65002));
    InMux I__9648 (
            .O(N__65022),
            .I(N__65002));
    InMux I__9647 (
            .O(N__65021),
            .I(N__65002));
    InMux I__9646 (
            .O(N__65020),
            .I(N__65002));
    LocalMux I__9645 (
            .O(N__65017),
            .I(N__64997));
    LocalMux I__9644 (
            .O(N__65014),
            .I(N__64997));
    Odrv4 I__9643 (
            .O(N__65011),
            .I(rco_int_0_a3_0_a2_138_m6_0_a2_7));
    LocalMux I__9642 (
            .O(N__65002),
            .I(rco_int_0_a3_0_a2_138_m6_0_a2_7));
    Odrv4 I__9641 (
            .O(N__64997),
            .I(rco_int_0_a3_0_a2_138_m6_0_a2_7));
    InMux I__9640 (
            .O(N__64990),
            .I(N__64987));
    LocalMux I__9639 (
            .O(N__64987),
            .I(N__64980));
    InMux I__9638 (
            .O(N__64986),
            .I(N__64968));
    InMux I__9637 (
            .O(N__64985),
            .I(N__64968));
    InMux I__9636 (
            .O(N__64984),
            .I(N__64968));
    InMux I__9635 (
            .O(N__64983),
            .I(N__64965));
    Span4Mux_h I__9634 (
            .O(N__64980),
            .I(N__64962));
    InMux I__9633 (
            .O(N__64979),
            .I(N__64955));
    InMux I__9632 (
            .O(N__64978),
            .I(N__64955));
    InMux I__9631 (
            .O(N__64977),
            .I(N__64955));
    InMux I__9630 (
            .O(N__64976),
            .I(N__64952));
    InMux I__9629 (
            .O(N__64975),
            .I(N__64940));
    LocalMux I__9628 (
            .O(N__64968),
            .I(N__64937));
    LocalMux I__9627 (
            .O(N__64965),
            .I(N__64934));
    Span4Mux_h I__9626 (
            .O(N__64962),
            .I(N__64927));
    LocalMux I__9625 (
            .O(N__64955),
            .I(N__64927));
    LocalMux I__9624 (
            .O(N__64952),
            .I(N__64927));
    InMux I__9623 (
            .O(N__64951),
            .I(N__64924));
    InMux I__9622 (
            .O(N__64950),
            .I(N__64921));
    InMux I__9621 (
            .O(N__64949),
            .I(N__64918));
    InMux I__9620 (
            .O(N__64948),
            .I(N__64909));
    InMux I__9619 (
            .O(N__64947),
            .I(N__64909));
    InMux I__9618 (
            .O(N__64946),
            .I(N__64909));
    InMux I__9617 (
            .O(N__64945),
            .I(N__64909));
    InMux I__9616 (
            .O(N__64944),
            .I(N__64904));
    InMux I__9615 (
            .O(N__64943),
            .I(N__64904));
    LocalMux I__9614 (
            .O(N__64940),
            .I(N__64899));
    Span4Mux_h I__9613 (
            .O(N__64937),
            .I(N__64899));
    Span4Mux_h I__9612 (
            .O(N__64934),
            .I(N__64894));
    Span4Mux_h I__9611 (
            .O(N__64927),
            .I(N__64894));
    LocalMux I__9610 (
            .O(N__64924),
            .I(rco_int_0_a2_0_a2_out_5));
    LocalMux I__9609 (
            .O(N__64921),
            .I(rco_int_0_a2_0_a2_out_5));
    LocalMux I__9608 (
            .O(N__64918),
            .I(rco_int_0_a2_0_a2_out_5));
    LocalMux I__9607 (
            .O(N__64909),
            .I(rco_int_0_a2_0_a2_out_5));
    LocalMux I__9606 (
            .O(N__64904),
            .I(rco_int_0_a2_0_a2_out_5));
    Odrv4 I__9605 (
            .O(N__64899),
            .I(rco_int_0_a2_0_a2_out_5));
    Odrv4 I__9604 (
            .O(N__64894),
            .I(rco_int_0_a2_0_a2_out_5));
    InMux I__9603 (
            .O(N__64879),
            .I(N__64873));
    InMux I__9602 (
            .O(N__64878),
            .I(N__64870));
    InMux I__9601 (
            .O(N__64877),
            .I(N__64867));
    InMux I__9600 (
            .O(N__64876),
            .I(N__64864));
    LocalMux I__9599 (
            .O(N__64873),
            .I(shift_srl_140Z0Z_15));
    LocalMux I__9598 (
            .O(N__64870),
            .I(shift_srl_140Z0Z_15));
    LocalMux I__9597 (
            .O(N__64867),
            .I(shift_srl_140Z0Z_15));
    LocalMux I__9596 (
            .O(N__64864),
            .I(shift_srl_140Z0Z_15));
    InMux I__9595 (
            .O(N__64855),
            .I(N__64852));
    LocalMux I__9594 (
            .O(N__64852),
            .I(shift_srl_139Z0Z_14));
    InMux I__9593 (
            .O(N__64849),
            .I(N__64846));
    LocalMux I__9592 (
            .O(N__64846),
            .I(N__64843));
    Span4Mux_v I__9591 (
            .O(N__64843),
            .I(N__64840));
    Span4Mux_v I__9590 (
            .O(N__64840),
            .I(N__64837));
    Odrv4 I__9589 (
            .O(N__64837),
            .I(shift_srl_139Z0Z_12));
    InMux I__9588 (
            .O(N__64834),
            .I(N__64831));
    LocalMux I__9587 (
            .O(N__64831),
            .I(shift_srl_139Z0Z_13));
    CEMux I__9586 (
            .O(N__64828),
            .I(N__64824));
    CEMux I__9585 (
            .O(N__64827),
            .I(N__64821));
    LocalMux I__9584 (
            .O(N__64824),
            .I(N__64815));
    LocalMux I__9583 (
            .O(N__64821),
            .I(N__64815));
    CEMux I__9582 (
            .O(N__64820),
            .I(N__64812));
    Span4Mux_v I__9581 (
            .O(N__64815),
            .I(N__64808));
    LocalMux I__9580 (
            .O(N__64812),
            .I(N__64805));
    CEMux I__9579 (
            .O(N__64811),
            .I(N__64802));
    Span4Mux_h I__9578 (
            .O(N__64808),
            .I(N__64796));
    Span4Mux_h I__9577 (
            .O(N__64805),
            .I(N__64796));
    LocalMux I__9576 (
            .O(N__64802),
            .I(N__64793));
    CEMux I__9575 (
            .O(N__64801),
            .I(N__64790));
    Span4Mux_v I__9574 (
            .O(N__64796),
            .I(N__64787));
    Span4Mux_v I__9573 (
            .O(N__64793),
            .I(N__64784));
    LocalMux I__9572 (
            .O(N__64790),
            .I(N__64781));
    Odrv4 I__9571 (
            .O(N__64787),
            .I(clk_en_139));
    Odrv4 I__9570 (
            .O(N__64784),
            .I(clk_en_139));
    Odrv12 I__9569 (
            .O(N__64781),
            .I(clk_en_139));
    InMux I__9568 (
            .O(N__64774),
            .I(N__64771));
    LocalMux I__9567 (
            .O(N__64771),
            .I(shift_srl_28Z0Z_1));
    InMux I__9566 (
            .O(N__64768),
            .I(N__64765));
    LocalMux I__9565 (
            .O(N__64765),
            .I(shift_srl_28Z0Z_2));
    InMux I__9564 (
            .O(N__64762),
            .I(N__64759));
    LocalMux I__9563 (
            .O(N__64759),
            .I(shift_srl_28Z0Z_3));
    InMux I__9562 (
            .O(N__64756),
            .I(N__64753));
    LocalMux I__9561 (
            .O(N__64753),
            .I(shift_srl_28Z0Z_11));
    InMux I__9560 (
            .O(N__64750),
            .I(N__64747));
    LocalMux I__9559 (
            .O(N__64747),
            .I(shift_srl_28Z0Z_8));
    InMux I__9558 (
            .O(N__64744),
            .I(N__64741));
    LocalMux I__9557 (
            .O(N__64741),
            .I(shift_srl_28Z0Z_12));
    InMux I__9556 (
            .O(N__64738),
            .I(N__64735));
    LocalMux I__9555 (
            .O(N__64735),
            .I(shift_srl_28Z0Z_13));
    InMux I__9554 (
            .O(N__64732),
            .I(N__64729));
    LocalMux I__9553 (
            .O(N__64729),
            .I(shift_srl_28Z0Z_14));
    InMux I__9552 (
            .O(N__64726),
            .I(N__64723));
    LocalMux I__9551 (
            .O(N__64723),
            .I(shift_srl_28Z0Z_4));
    InMux I__9550 (
            .O(N__64720),
            .I(N__64717));
    LocalMux I__9549 (
            .O(N__64717),
            .I(shift_srl_28Z0Z_5));
    InMux I__9548 (
            .O(N__64714),
            .I(N__64711));
    LocalMux I__9547 (
            .O(N__64711),
            .I(shift_srl_28Z0Z_6));
    InMux I__9546 (
            .O(N__64708),
            .I(N__64705));
    LocalMux I__9545 (
            .O(N__64705),
            .I(shift_srl_26Z0Z_14));
    InMux I__9544 (
            .O(N__64702),
            .I(N__64699));
    LocalMux I__9543 (
            .O(N__64699),
            .I(shift_srl_26Z0Z_9));
    InMux I__9542 (
            .O(N__64696),
            .I(N__64693));
    LocalMux I__9541 (
            .O(N__64693),
            .I(N__64690));
    Odrv12 I__9540 (
            .O(N__64690),
            .I(shift_srl_26Z0Z_7));
    InMux I__9539 (
            .O(N__64687),
            .I(N__64684));
    LocalMux I__9538 (
            .O(N__64684),
            .I(shift_srl_26Z0Z_8));
    CEMux I__9537 (
            .O(N__64681),
            .I(N__64678));
    LocalMux I__9536 (
            .O(N__64678),
            .I(N__64674));
    CEMux I__9535 (
            .O(N__64677),
            .I(N__64671));
    Span4Mux_h I__9534 (
            .O(N__64674),
            .I(N__64666));
    LocalMux I__9533 (
            .O(N__64671),
            .I(N__64666));
    Span4Mux_h I__9532 (
            .O(N__64666),
            .I(N__64663));
    Odrv4 I__9531 (
            .O(N__64663),
            .I(clk_en_26));
    InMux I__9530 (
            .O(N__64660),
            .I(N__64657));
    LocalMux I__9529 (
            .O(N__64657),
            .I(shift_srl_28Z0Z_0));
    InMux I__9528 (
            .O(N__64654),
            .I(N__64651));
    LocalMux I__9527 (
            .O(N__64651),
            .I(shift_srl_28Z0Z_10));
    InMux I__9526 (
            .O(N__64648),
            .I(N__64645));
    LocalMux I__9525 (
            .O(N__64645),
            .I(shift_srl_28Z0Z_9));
    InMux I__9524 (
            .O(N__64642),
            .I(N__64639));
    LocalMux I__9523 (
            .O(N__64639),
            .I(shift_srl_42Z0Z_0));
    InMux I__9522 (
            .O(N__64636),
            .I(N__64633));
    LocalMux I__9521 (
            .O(N__64633),
            .I(shift_srl_42Z0Z_1));
    InMux I__9520 (
            .O(N__64630),
            .I(N__64627));
    LocalMux I__9519 (
            .O(N__64627),
            .I(shift_srl_42Z0Z_2));
    InMux I__9518 (
            .O(N__64624),
            .I(N__64621));
    LocalMux I__9517 (
            .O(N__64621),
            .I(shift_srl_42Z0Z_3));
    InMux I__9516 (
            .O(N__64618),
            .I(N__64615));
    LocalMux I__9515 (
            .O(N__64615),
            .I(N__64612));
    Odrv12 I__9514 (
            .O(N__64612),
            .I(shift_srl_42Z0Z_4));
    InMux I__9513 (
            .O(N__64609),
            .I(N__64606));
    LocalMux I__9512 (
            .O(N__64606),
            .I(shift_srl_26Z0Z_10));
    InMux I__9511 (
            .O(N__64603),
            .I(N__64600));
    LocalMux I__9510 (
            .O(N__64600),
            .I(shift_srl_26Z0Z_11));
    InMux I__9509 (
            .O(N__64597),
            .I(N__64594));
    LocalMux I__9508 (
            .O(N__64594),
            .I(shift_srl_26Z0Z_12));
    InMux I__9507 (
            .O(N__64591),
            .I(N__64588));
    LocalMux I__9506 (
            .O(N__64588),
            .I(shift_srl_26Z0Z_13));
    InMux I__9505 (
            .O(N__64585),
            .I(N__64582));
    LocalMux I__9504 (
            .O(N__64582),
            .I(shift_srl_42Z0Z_12));
    InMux I__9503 (
            .O(N__64579),
            .I(N__64576));
    LocalMux I__9502 (
            .O(N__64576),
            .I(shift_srl_42Z0Z_13));
    InMux I__9501 (
            .O(N__64573),
            .I(N__64570));
    LocalMux I__9500 (
            .O(N__64570),
            .I(shift_srl_42Z0Z_14));
    InMux I__9499 (
            .O(N__64567),
            .I(N__64564));
    LocalMux I__9498 (
            .O(N__64564),
            .I(shift_srl_42Z0Z_9));
    InMux I__9497 (
            .O(N__64561),
            .I(N__64558));
    LocalMux I__9496 (
            .O(N__64558),
            .I(shift_srl_42Z0Z_7));
    InMux I__9495 (
            .O(N__64555),
            .I(N__64552));
    LocalMux I__9494 (
            .O(N__64552),
            .I(shift_srl_42Z0Z_8));
    IoInMux I__9493 (
            .O(N__64549),
            .I(N__64546));
    LocalMux I__9492 (
            .O(N__64546),
            .I(N__64543));
    Span4Mux_s0_v I__9491 (
            .O(N__64543),
            .I(N__64540));
    Sp12to4 I__9490 (
            .O(N__64540),
            .I(N__64537));
    Span12Mux_h I__9489 (
            .O(N__64537),
            .I(N__64534));
    Span12Mux_v I__9488 (
            .O(N__64534),
            .I(N__64531));
    Odrv12 I__9487 (
            .O(N__64531),
            .I(rco_c_43));
    IoInMux I__9486 (
            .O(N__64528),
            .I(N__64525));
    LocalMux I__9485 (
            .O(N__64525),
            .I(N__64522));
    IoSpan4Mux I__9484 (
            .O(N__64522),
            .I(N__64519));
    Span4Mux_s0_v I__9483 (
            .O(N__64519),
            .I(N__64516));
    Sp12to4 I__9482 (
            .O(N__64516),
            .I(N__64513));
    Span12Mux_s11_v I__9481 (
            .O(N__64513),
            .I(N__64510));
    Span12Mux_h I__9480 (
            .O(N__64510),
            .I(N__64507));
    Odrv12 I__9479 (
            .O(N__64507),
            .I(rco_c_42));
    InMux I__9478 (
            .O(N__64504),
            .I(N__64501));
    LocalMux I__9477 (
            .O(N__64501),
            .I(shift_srl_99Z0Z_9));
    InMux I__9476 (
            .O(N__64498),
            .I(N__64495));
    LocalMux I__9475 (
            .O(N__64495),
            .I(shift_srl_99Z0Z_8));
    InMux I__9474 (
            .O(N__64492),
            .I(N__64489));
    LocalMux I__9473 (
            .O(N__64489),
            .I(N__64486));
    Span4Mux_h I__9472 (
            .O(N__64486),
            .I(N__64483));
    Odrv4 I__9471 (
            .O(N__64483),
            .I(shift_srl_99Z0Z_6));
    InMux I__9470 (
            .O(N__64480),
            .I(N__64477));
    LocalMux I__9469 (
            .O(N__64477),
            .I(shift_srl_99Z0Z_7));
    InMux I__9468 (
            .O(N__64474),
            .I(N__64471));
    LocalMux I__9467 (
            .O(N__64471),
            .I(shift_srl_42Z0Z_6));
    InMux I__9466 (
            .O(N__64468),
            .I(N__64465));
    LocalMux I__9465 (
            .O(N__64465),
            .I(shift_srl_42Z0Z_5));
    InMux I__9464 (
            .O(N__64462),
            .I(N__64459));
    LocalMux I__9463 (
            .O(N__64459),
            .I(shift_srl_42Z0Z_10));
    InMux I__9462 (
            .O(N__64456),
            .I(N__64453));
    LocalMux I__9461 (
            .O(N__64453),
            .I(shift_srl_42Z0Z_11));
    InMux I__9460 (
            .O(N__64450),
            .I(N__64447));
    LocalMux I__9459 (
            .O(N__64447),
            .I(shift_srl_87Z0Z_2));
    InMux I__9458 (
            .O(N__64444),
            .I(N__64441));
    LocalMux I__9457 (
            .O(N__64441),
            .I(shift_srl_87Z0Z_3));
    InMux I__9456 (
            .O(N__64438),
            .I(N__64435));
    LocalMux I__9455 (
            .O(N__64435),
            .I(shift_srl_87Z0Z_4));
    InMux I__9454 (
            .O(N__64432),
            .I(N__64429));
    LocalMux I__9453 (
            .O(N__64429),
            .I(shift_srl_87Z0Z_5));
    InMux I__9452 (
            .O(N__64426),
            .I(N__64423));
    LocalMux I__9451 (
            .O(N__64423),
            .I(shift_srl_87Z0Z_6));
    InMux I__9450 (
            .O(N__64420),
            .I(N__64417));
    LocalMux I__9449 (
            .O(N__64417),
            .I(N__64414));
    Odrv4 I__9448 (
            .O(N__64414),
            .I(shift_srl_87Z0Z_7));
    CEMux I__9447 (
            .O(N__64411),
            .I(N__64407));
    CEMux I__9446 (
            .O(N__64410),
            .I(N__64404));
    LocalMux I__9445 (
            .O(N__64407),
            .I(N__64401));
    LocalMux I__9444 (
            .O(N__64404),
            .I(N__64398));
    Odrv4 I__9443 (
            .O(N__64401),
            .I(clk_en_87));
    Odrv4 I__9442 (
            .O(N__64398),
            .I(clk_en_87));
    InMux I__9441 (
            .O(N__64393),
            .I(N__64390));
    LocalMux I__9440 (
            .O(N__64390),
            .I(shift_srl_99Z0Z_10));
    InMux I__9439 (
            .O(N__64387),
            .I(N__64384));
    LocalMux I__9438 (
            .O(N__64384),
            .I(shift_srl_99Z0Z_11));
    InMux I__9437 (
            .O(N__64381),
            .I(N__64378));
    LocalMux I__9436 (
            .O(N__64378),
            .I(shift_srl_99Z0Z_12));
    InMux I__9435 (
            .O(N__64375),
            .I(N__64372));
    LocalMux I__9434 (
            .O(N__64372),
            .I(shift_srl_99Z0Z_13));
    InMux I__9433 (
            .O(N__64369),
            .I(N__64366));
    LocalMux I__9432 (
            .O(N__64366),
            .I(shift_srl_88Z0Z_1));
    InMux I__9431 (
            .O(N__64363),
            .I(N__64360));
    LocalMux I__9430 (
            .O(N__64360),
            .I(shift_srl_88Z0Z_2));
    InMux I__9429 (
            .O(N__64357),
            .I(N__64354));
    LocalMux I__9428 (
            .O(N__64354),
            .I(shift_srl_88Z0Z_3));
    InMux I__9427 (
            .O(N__64351),
            .I(N__64348));
    LocalMux I__9426 (
            .O(N__64348),
            .I(shift_srl_88Z0Z_4));
    InMux I__9425 (
            .O(N__64345),
            .I(N__64342));
    LocalMux I__9424 (
            .O(N__64342),
            .I(shift_srl_88Z0Z_5));
    InMux I__9423 (
            .O(N__64339),
            .I(N__64336));
    LocalMux I__9422 (
            .O(N__64336),
            .I(shift_srl_88Z0Z_6));
    InMux I__9421 (
            .O(N__64333),
            .I(N__64330));
    LocalMux I__9420 (
            .O(N__64330),
            .I(shift_srl_88Z0Z_7));
    CEMux I__9419 (
            .O(N__64327),
            .I(N__64323));
    CEMux I__9418 (
            .O(N__64326),
            .I(N__64320));
    LocalMux I__9417 (
            .O(N__64323),
            .I(N__64317));
    LocalMux I__9416 (
            .O(N__64320),
            .I(N__64314));
    Span4Mux_v I__9415 (
            .O(N__64317),
            .I(N__64311));
    Span4Mux_h I__9414 (
            .O(N__64314),
            .I(N__64308));
    Odrv4 I__9413 (
            .O(N__64311),
            .I(clk_en_88));
    Odrv4 I__9412 (
            .O(N__64308),
            .I(clk_en_88));
    InMux I__9411 (
            .O(N__64303),
            .I(N__64300));
    LocalMux I__9410 (
            .O(N__64300),
            .I(shift_srl_87Z0Z_0));
    InMux I__9409 (
            .O(N__64297),
            .I(N__64294));
    LocalMux I__9408 (
            .O(N__64294),
            .I(shift_srl_87Z0Z_1));
    InMux I__9407 (
            .O(N__64291),
            .I(N__64288));
    LocalMux I__9406 (
            .O(N__64288),
            .I(shift_srl_85Z0Z_0));
    InMux I__9405 (
            .O(N__64285),
            .I(N__64282));
    LocalMux I__9404 (
            .O(N__64282),
            .I(shift_srl_85Z0Z_1));
    InMux I__9403 (
            .O(N__64279),
            .I(N__64276));
    LocalMux I__9402 (
            .O(N__64276),
            .I(shift_srl_85Z0Z_2));
    InMux I__9401 (
            .O(N__64273),
            .I(N__64270));
    LocalMux I__9400 (
            .O(N__64270),
            .I(shift_srl_85Z0Z_3));
    InMux I__9399 (
            .O(N__64267),
            .I(N__64264));
    LocalMux I__9398 (
            .O(N__64264),
            .I(shift_srl_85Z0Z_4));
    InMux I__9397 (
            .O(N__64261),
            .I(N__64258));
    LocalMux I__9396 (
            .O(N__64258),
            .I(shift_srl_85Z0Z_5));
    InMux I__9395 (
            .O(N__64255),
            .I(N__64252));
    LocalMux I__9394 (
            .O(N__64252),
            .I(shift_srl_85Z0Z_6));
    InMux I__9393 (
            .O(N__64249),
            .I(N__64246));
    LocalMux I__9392 (
            .O(N__64246),
            .I(shift_srl_85Z0Z_7));
    CEMux I__9391 (
            .O(N__64243),
            .I(N__64240));
    LocalMux I__9390 (
            .O(N__64240),
            .I(N__64236));
    CEMux I__9389 (
            .O(N__64239),
            .I(N__64233));
    Span4Mux_v I__9388 (
            .O(N__64236),
            .I(N__64230));
    LocalMux I__9387 (
            .O(N__64233),
            .I(N__64227));
    Odrv4 I__9386 (
            .O(N__64230),
            .I(clk_en_85));
    Odrv4 I__9385 (
            .O(N__64227),
            .I(clk_en_85));
    InMux I__9384 (
            .O(N__64222),
            .I(N__64219));
    LocalMux I__9383 (
            .O(N__64219),
            .I(shift_srl_88Z0Z_0));
    IoInMux I__9382 (
            .O(N__64216),
            .I(N__64213));
    LocalMux I__9381 (
            .O(N__64213),
            .I(N__64210));
    IoSpan4Mux I__9380 (
            .O(N__64210),
            .I(N__64207));
    Span4Mux_s1_h I__9379 (
            .O(N__64207),
            .I(N__64204));
    Sp12to4 I__9378 (
            .O(N__64204),
            .I(N__64201));
    Span12Mux_h I__9377 (
            .O(N__64201),
            .I(N__64198));
    Span12Mux_v I__9376 (
            .O(N__64198),
            .I(N__64195));
    Odrv12 I__9375 (
            .O(N__64195),
            .I(rco_c_191));
    IoInMux I__9374 (
            .O(N__64192),
            .I(N__64189));
    LocalMux I__9373 (
            .O(N__64189),
            .I(N__64186));
    Span12Mux_s2_h I__9372 (
            .O(N__64186),
            .I(N__64183));
    Span12Mux_h I__9371 (
            .O(N__64183),
            .I(N__64180));
    Span12Mux_v I__9370 (
            .O(N__64180),
            .I(N__64177));
    Odrv12 I__9369 (
            .O(N__64177),
            .I(rco_c_195));
    InMux I__9368 (
            .O(N__64174),
            .I(N__64171));
    LocalMux I__9367 (
            .O(N__64171),
            .I(shift_srl_194Z0Z_0));
    InMux I__9366 (
            .O(N__64168),
            .I(N__64165));
    LocalMux I__9365 (
            .O(N__64165),
            .I(shift_srl_139Z0Z_11));
    IoInMux I__9364 (
            .O(N__64162),
            .I(N__64159));
    LocalMux I__9363 (
            .O(N__64159),
            .I(N__64156));
    Span4Mux_s2_v I__9362 (
            .O(N__64156),
            .I(N__64153));
    Odrv4 I__9361 (
            .O(N__64153),
            .I(rco_c_90));
    IoInMux I__9360 (
            .O(N__64150),
            .I(N__64147));
    LocalMux I__9359 (
            .O(N__64147),
            .I(N__64144));
    Span4Mux_s1_v I__9358 (
            .O(N__64144),
            .I(N__64141));
    Span4Mux_h I__9357 (
            .O(N__64141),
            .I(N__64138));
    Odrv4 I__9356 (
            .O(N__64138),
            .I(rco_c_91));
    InMux I__9355 (
            .O(N__64135),
            .I(N__64132));
    LocalMux I__9354 (
            .O(N__64132),
            .I(shift_srl_115Z0Z_12));
    InMux I__9353 (
            .O(N__64129),
            .I(N__64126));
    LocalMux I__9352 (
            .O(N__64126),
            .I(shift_srl_115Z0Z_13));
    InMux I__9351 (
            .O(N__64123),
            .I(N__64120));
    LocalMux I__9350 (
            .O(N__64120),
            .I(N__64117));
    Span4Mux_v I__9349 (
            .O(N__64117),
            .I(N__64114));
    Sp12to4 I__9348 (
            .O(N__64114),
            .I(N__64111));
    Odrv12 I__9347 (
            .O(N__64111),
            .I(shift_srl_115Z0Z_14));
    InMux I__9346 (
            .O(N__64108),
            .I(N__64105));
    LocalMux I__9345 (
            .O(N__64105),
            .I(shift_srl_115Z0Z_9));
    InMux I__9344 (
            .O(N__64102),
            .I(N__64099));
    LocalMux I__9343 (
            .O(N__64099),
            .I(shift_srl_115Z0Z_8));
    InMux I__9342 (
            .O(N__64096),
            .I(N__64093));
    LocalMux I__9341 (
            .O(N__64093),
            .I(shift_srl_115Z0Z_6));
    InMux I__9340 (
            .O(N__64090),
            .I(N__64087));
    LocalMux I__9339 (
            .O(N__64087),
            .I(shift_srl_115Z0Z_7));
    CEMux I__9338 (
            .O(N__64084),
            .I(N__64081));
    LocalMux I__9337 (
            .O(N__64081),
            .I(N__64077));
    CEMux I__9336 (
            .O(N__64080),
            .I(N__64074));
    Span4Mux_h I__9335 (
            .O(N__64077),
            .I(N__64070));
    LocalMux I__9334 (
            .O(N__64074),
            .I(N__64067));
    CEMux I__9333 (
            .O(N__64073),
            .I(N__64064));
    Span4Mux_h I__9332 (
            .O(N__64070),
            .I(N__64061));
    Span4Mux_h I__9331 (
            .O(N__64067),
            .I(N__64058));
    LocalMux I__9330 (
            .O(N__64064),
            .I(N__64055));
    Odrv4 I__9329 (
            .O(N__64061),
            .I(clk_en_115));
    Odrv4 I__9328 (
            .O(N__64058),
            .I(clk_en_115));
    Odrv12 I__9327 (
            .O(N__64055),
            .I(clk_en_115));
    IoInMux I__9326 (
            .O(N__64048),
            .I(N__64045));
    LocalMux I__9325 (
            .O(N__64045),
            .I(N__64042));
    Span4Mux_s2_h I__9324 (
            .O(N__64042),
            .I(N__64039));
    Sp12to4 I__9323 (
            .O(N__64039),
            .I(N__64036));
    Span12Mux_v I__9322 (
            .O(N__64036),
            .I(N__64033));
    Span12Mux_h I__9321 (
            .O(N__64033),
            .I(N__64030));
    Odrv12 I__9320 (
            .O(N__64030),
            .I(rco_c_194));
    IoInMux I__9319 (
            .O(N__64027),
            .I(N__64024));
    LocalMux I__9318 (
            .O(N__64024),
            .I(N__64021));
    Span4Mux_s2_h I__9317 (
            .O(N__64021),
            .I(N__64018));
    Sp12to4 I__9316 (
            .O(N__64018),
            .I(N__64015));
    Span12Mux_v I__9315 (
            .O(N__64015),
            .I(N__64012));
    Span12Mux_h I__9314 (
            .O(N__64012),
            .I(N__64009));
    Odrv12 I__9313 (
            .O(N__64009),
            .I(rco_c_193));
    IoInMux I__9312 (
            .O(N__64006),
            .I(N__64003));
    LocalMux I__9311 (
            .O(N__64003),
            .I(N__64000));
    Span12Mux_s2_h I__9310 (
            .O(N__64000),
            .I(N__63997));
    Span12Mux_h I__9309 (
            .O(N__63997),
            .I(N__63994));
    Span12Mux_v I__9308 (
            .O(N__63994),
            .I(N__63991));
    Odrv12 I__9307 (
            .O(N__63991),
            .I(rco_c_184));
    IoInMux I__9306 (
            .O(N__63988),
            .I(N__63985));
    LocalMux I__9305 (
            .O(N__63985),
            .I(N__63982));
    Span12Mux_s2_h I__9304 (
            .O(N__63982),
            .I(N__63979));
    Span12Mux_h I__9303 (
            .O(N__63979),
            .I(N__63976));
    Span12Mux_v I__9302 (
            .O(N__63976),
            .I(N__63973));
    Odrv12 I__9301 (
            .O(N__63973),
            .I(rco_c_187));
    InMux I__9300 (
            .O(N__63970),
            .I(N__63967));
    LocalMux I__9299 (
            .O(N__63967),
            .I(shift_srl_115Z0Z_0));
    InMux I__9298 (
            .O(N__63964),
            .I(N__63961));
    LocalMux I__9297 (
            .O(N__63961),
            .I(shift_srl_115Z0Z_1));
    InMux I__9296 (
            .O(N__63958),
            .I(N__63955));
    LocalMux I__9295 (
            .O(N__63955),
            .I(shift_srl_115Z0Z_2));
    InMux I__9294 (
            .O(N__63952),
            .I(N__63949));
    LocalMux I__9293 (
            .O(N__63949),
            .I(shift_srl_115Z0Z_3));
    InMux I__9292 (
            .O(N__63946),
            .I(N__63943));
    LocalMux I__9291 (
            .O(N__63943),
            .I(shift_srl_115Z0Z_4));
    InMux I__9290 (
            .O(N__63940),
            .I(N__63937));
    LocalMux I__9289 (
            .O(N__63937),
            .I(shift_srl_115Z0Z_5));
    InMux I__9288 (
            .O(N__63934),
            .I(N__63931));
    LocalMux I__9287 (
            .O(N__63931),
            .I(shift_srl_115Z0Z_10));
    InMux I__9286 (
            .O(N__63928),
            .I(N__63925));
    LocalMux I__9285 (
            .O(N__63925),
            .I(shift_srl_115Z0Z_11));
    InMux I__9284 (
            .O(N__63922),
            .I(N__63919));
    LocalMux I__9283 (
            .O(N__63919),
            .I(shift_srl_120Z0Z_10));
    InMux I__9282 (
            .O(N__63916),
            .I(N__63913));
    LocalMux I__9281 (
            .O(N__63913),
            .I(shift_srl_120Z0Z_11));
    InMux I__9280 (
            .O(N__63910),
            .I(N__63907));
    LocalMux I__9279 (
            .O(N__63907),
            .I(shift_srl_120Z0Z_12));
    InMux I__9278 (
            .O(N__63904),
            .I(N__63901));
    LocalMux I__9277 (
            .O(N__63901),
            .I(shift_srl_120Z0Z_13));
    InMux I__9276 (
            .O(N__63898),
            .I(N__63895));
    LocalMux I__9275 (
            .O(N__63895),
            .I(shift_srl_120Z0Z_14));
    InMux I__9274 (
            .O(N__63892),
            .I(N__63889));
    LocalMux I__9273 (
            .O(N__63889),
            .I(shift_srl_120Z0Z_9));
    InMux I__9272 (
            .O(N__63886),
            .I(N__63883));
    LocalMux I__9271 (
            .O(N__63883),
            .I(shift_srl_120Z0Z_8));
    IoInMux I__9270 (
            .O(N__63880),
            .I(N__63877));
    LocalMux I__9269 (
            .O(N__63877),
            .I(N__63874));
    Span12Mux_s6_h I__9268 (
            .O(N__63874),
            .I(N__63870));
    InMux I__9267 (
            .O(N__63873),
            .I(N__63867));
    Span12Mux_h I__9266 (
            .O(N__63870),
            .I(N__63864));
    LocalMux I__9265 (
            .O(N__63867),
            .I(N__63861));
    Odrv12 I__9264 (
            .O(N__63864),
            .I(N_162));
    Odrv4 I__9263 (
            .O(N__63861),
            .I(N_162));
    IoInMux I__9262 (
            .O(N__63856),
            .I(N__63853));
    LocalMux I__9261 (
            .O(N__63853),
            .I(N__63850));
    IoSpan4Mux I__9260 (
            .O(N__63850),
            .I(N__63847));
    Span4Mux_s2_h I__9259 (
            .O(N__63847),
            .I(N__63844));
    Sp12to4 I__9258 (
            .O(N__63844),
            .I(N__63841));
    Span12Mux_s9_h I__9257 (
            .O(N__63841),
            .I(N__63838));
    Odrv12 I__9256 (
            .O(N__63838),
            .I(rco_c_115));
    InMux I__9255 (
            .O(N__63835),
            .I(N__63827));
    InMux I__9254 (
            .O(N__63834),
            .I(N__63827));
    InMux I__9253 (
            .O(N__63833),
            .I(N__63822));
    InMux I__9252 (
            .O(N__63832),
            .I(N__63822));
    LocalMux I__9251 (
            .O(N__63827),
            .I(N__63819));
    LocalMux I__9250 (
            .O(N__63822),
            .I(N__63815));
    Span4Mux_v I__9249 (
            .O(N__63819),
            .I(N__63806));
    InMux I__9248 (
            .O(N__63818),
            .I(N__63803));
    Span4Mux_v I__9247 (
            .O(N__63815),
            .I(N__63800));
    InMux I__9246 (
            .O(N__63814),
            .I(N__63797));
    InMux I__9245 (
            .O(N__63813),
            .I(N__63794));
    InMux I__9244 (
            .O(N__63812),
            .I(N__63791));
    InMux I__9243 (
            .O(N__63811),
            .I(N__63784));
    InMux I__9242 (
            .O(N__63810),
            .I(N__63784));
    InMux I__9241 (
            .O(N__63809),
            .I(N__63784));
    Sp12to4 I__9240 (
            .O(N__63806),
            .I(N__63775));
    LocalMux I__9239 (
            .O(N__63803),
            .I(N__63775));
    Sp12to4 I__9238 (
            .O(N__63800),
            .I(N__63775));
    LocalMux I__9237 (
            .O(N__63797),
            .I(N__63775));
    LocalMux I__9236 (
            .O(N__63794),
            .I(shift_srl_115Z0Z_15));
    LocalMux I__9235 (
            .O(N__63791),
            .I(shift_srl_115Z0Z_15));
    LocalMux I__9234 (
            .O(N__63784),
            .I(shift_srl_115Z0Z_15));
    Odrv12 I__9233 (
            .O(N__63775),
            .I(shift_srl_115Z0Z_15));
    CascadeMux I__9232 (
            .O(N__63766),
            .I(N__63758));
    CascadeMux I__9231 (
            .O(N__63765),
            .I(N__63755));
    InMux I__9230 (
            .O(N__63764),
            .I(N__63749));
    InMux I__9229 (
            .O(N__63763),
            .I(N__63749));
    InMux I__9228 (
            .O(N__63762),
            .I(N__63745));
    InMux I__9227 (
            .O(N__63761),
            .I(N__63738));
    InMux I__9226 (
            .O(N__63758),
            .I(N__63738));
    InMux I__9225 (
            .O(N__63755),
            .I(N__63738));
    InMux I__9224 (
            .O(N__63754),
            .I(N__63735));
    LocalMux I__9223 (
            .O(N__63749),
            .I(N__63732));
    InMux I__9222 (
            .O(N__63748),
            .I(N__63729));
    LocalMux I__9221 (
            .O(N__63745),
            .I(N__63722));
    LocalMux I__9220 (
            .O(N__63738),
            .I(N__63722));
    LocalMux I__9219 (
            .O(N__63735),
            .I(N__63722));
    Span4Mux_h I__9218 (
            .O(N__63732),
            .I(N__63719));
    LocalMux I__9217 (
            .O(N__63729),
            .I(N__63716));
    Span4Mux_h I__9216 (
            .O(N__63722),
            .I(N__63711));
    Span4Mux_h I__9215 (
            .O(N__63719),
            .I(N__63711));
    Odrv4 I__9214 (
            .O(N__63716),
            .I(shift_srl_142Z0Z_15));
    Odrv4 I__9213 (
            .O(N__63711),
            .I(shift_srl_142Z0Z_15));
    InMux I__9212 (
            .O(N__63706),
            .I(N__63703));
    LocalMux I__9211 (
            .O(N__63703),
            .I(shift_srl_142Z0Z_0));
    InMux I__9210 (
            .O(N__63700),
            .I(N__63697));
    LocalMux I__9209 (
            .O(N__63697),
            .I(shift_srl_142Z0Z_1));
    InMux I__9208 (
            .O(N__63694),
            .I(N__63691));
    LocalMux I__9207 (
            .O(N__63691),
            .I(shift_srl_142Z0Z_2));
    InMux I__9206 (
            .O(N__63688),
            .I(N__63685));
    LocalMux I__9205 (
            .O(N__63685),
            .I(shift_srl_142Z0Z_3));
    InMux I__9204 (
            .O(N__63682),
            .I(N__63679));
    LocalMux I__9203 (
            .O(N__63679),
            .I(shift_srl_142Z0Z_4));
    InMux I__9202 (
            .O(N__63676),
            .I(N__63673));
    LocalMux I__9201 (
            .O(N__63673),
            .I(shift_srl_142Z0Z_5));
    InMux I__9200 (
            .O(N__63670),
            .I(N__63667));
    LocalMux I__9199 (
            .O(N__63667),
            .I(shift_srl_142Z0Z_6));
    InMux I__9198 (
            .O(N__63664),
            .I(N__63661));
    LocalMux I__9197 (
            .O(N__63661),
            .I(N__63658));
    Odrv4 I__9196 (
            .O(N__63658),
            .I(shift_srl_142Z0Z_7));
    CEMux I__9195 (
            .O(N__63655),
            .I(N__63651));
    CEMux I__9194 (
            .O(N__63654),
            .I(N__63648));
    LocalMux I__9193 (
            .O(N__63651),
            .I(N__63645));
    LocalMux I__9192 (
            .O(N__63648),
            .I(N__63642));
    Span4Mux_h I__9191 (
            .O(N__63645),
            .I(N__63639));
    Odrv12 I__9190 (
            .O(N__63642),
            .I(clk_en_142));
    Odrv4 I__9189 (
            .O(N__63639),
            .I(clk_en_142));
    InMux I__9188 (
            .O(N__63634),
            .I(N__63631));
    LocalMux I__9187 (
            .O(N__63631),
            .I(shift_srl_140Z0Z_6));
    InMux I__9186 (
            .O(N__63628),
            .I(N__63625));
    LocalMux I__9185 (
            .O(N__63625),
            .I(shift_srl_140Z0Z_7));
    CEMux I__9184 (
            .O(N__63622),
            .I(N__63618));
    CEMux I__9183 (
            .O(N__63621),
            .I(N__63615));
    LocalMux I__9182 (
            .O(N__63618),
            .I(N__63612));
    LocalMux I__9181 (
            .O(N__63615),
            .I(N__63609));
    Span4Mux_v I__9180 (
            .O(N__63612),
            .I(N__63606));
    Span12Mux_h I__9179 (
            .O(N__63609),
            .I(N__63603));
    Odrv4 I__9178 (
            .O(N__63606),
            .I(N_124_i));
    Odrv12 I__9177 (
            .O(N__63603),
            .I(N_124_i));
    InMux I__9176 (
            .O(N__63598),
            .I(N__63595));
    LocalMux I__9175 (
            .O(N__63595),
            .I(N__63592));
    Span4Mux_v I__9174 (
            .O(N__63592),
            .I(N__63587));
    InMux I__9173 (
            .O(N__63591),
            .I(N__63584));
    InMux I__9172 (
            .O(N__63590),
            .I(N__63580));
    Span4Mux_h I__9171 (
            .O(N__63587),
            .I(N__63575));
    LocalMux I__9170 (
            .O(N__63584),
            .I(N__63575));
    InMux I__9169 (
            .O(N__63583),
            .I(N__63572));
    LocalMux I__9168 (
            .O(N__63580),
            .I(N__63567));
    Span4Mux_h I__9167 (
            .O(N__63575),
            .I(N__63567));
    LocalMux I__9166 (
            .O(N__63572),
            .I(shift_srl_145Z0Z_15));
    Odrv4 I__9165 (
            .O(N__63567),
            .I(shift_srl_145Z0Z_15));
    InMux I__9164 (
            .O(N__63562),
            .I(N__63559));
    LocalMux I__9163 (
            .O(N__63559),
            .I(shift_srl_145Z0Z_0));
    InMux I__9162 (
            .O(N__63556),
            .I(N__63553));
    LocalMux I__9161 (
            .O(N__63553),
            .I(shift_srl_145Z0Z_1));
    InMux I__9160 (
            .O(N__63550),
            .I(N__63547));
    LocalMux I__9159 (
            .O(N__63547),
            .I(shift_srl_145Z0Z_2));
    InMux I__9158 (
            .O(N__63544),
            .I(N__63541));
    LocalMux I__9157 (
            .O(N__63541),
            .I(shift_srl_145Z0Z_3));
    InMux I__9156 (
            .O(N__63538),
            .I(N__63535));
    LocalMux I__9155 (
            .O(N__63535),
            .I(shift_srl_145Z0Z_4));
    InMux I__9154 (
            .O(N__63532),
            .I(N__63529));
    LocalMux I__9153 (
            .O(N__63529),
            .I(shift_srl_145Z0Z_5));
    InMux I__9152 (
            .O(N__63526),
            .I(N__63523));
    LocalMux I__9151 (
            .O(N__63523),
            .I(shift_srl_145Z0Z_6));
    InMux I__9150 (
            .O(N__63520),
            .I(N__63517));
    LocalMux I__9149 (
            .O(N__63517),
            .I(shift_srl_145Z0Z_7));
    CEMux I__9148 (
            .O(N__63514),
            .I(N__63510));
    CEMux I__9147 (
            .O(N__63513),
            .I(N__63507));
    LocalMux I__9146 (
            .O(N__63510),
            .I(N__63504));
    LocalMux I__9145 (
            .O(N__63507),
            .I(N__63501));
    Span4Mux_h I__9144 (
            .O(N__63504),
            .I(N__63496));
    Span4Mux_h I__9143 (
            .O(N__63501),
            .I(N__63496));
    Odrv4 I__9142 (
            .O(N__63496),
            .I(clk_en_145));
    InMux I__9141 (
            .O(N__63493),
            .I(N__63490));
    LocalMux I__9140 (
            .O(N__63490),
            .I(shift_srl_140Z0Z_14));
    InMux I__9139 (
            .O(N__63487),
            .I(N__63484));
    LocalMux I__9138 (
            .O(N__63484),
            .I(shift_srl_140Z0Z_9));
    InMux I__9137 (
            .O(N__63481),
            .I(N__63478));
    LocalMux I__9136 (
            .O(N__63478),
            .I(shift_srl_140Z0Z_8));
    InMux I__9135 (
            .O(N__63475),
            .I(N__63472));
    LocalMux I__9134 (
            .O(N__63472),
            .I(shift_srl_140Z0Z_0));
    InMux I__9133 (
            .O(N__63469),
            .I(N__63466));
    LocalMux I__9132 (
            .O(N__63466),
            .I(shift_srl_140Z0Z_1));
    InMux I__9131 (
            .O(N__63463),
            .I(N__63460));
    LocalMux I__9130 (
            .O(N__63460),
            .I(shift_srl_140Z0Z_2));
    InMux I__9129 (
            .O(N__63457),
            .I(N__63454));
    LocalMux I__9128 (
            .O(N__63454),
            .I(shift_srl_140Z0Z_3));
    InMux I__9127 (
            .O(N__63451),
            .I(N__63448));
    LocalMux I__9126 (
            .O(N__63448),
            .I(shift_srl_140Z0Z_4));
    InMux I__9125 (
            .O(N__63445),
            .I(N__63442));
    LocalMux I__9124 (
            .O(N__63442),
            .I(shift_srl_140Z0Z_5));
    InMux I__9123 (
            .O(N__63439),
            .I(N__63436));
    LocalMux I__9122 (
            .O(N__63436),
            .I(shift_srl_151Z0Z_13));
    InMux I__9121 (
            .O(N__63433),
            .I(N__63430));
    LocalMux I__9120 (
            .O(N__63430),
            .I(shift_srl_151Z0Z_14));
    InMux I__9119 (
            .O(N__63427),
            .I(N__63424));
    LocalMux I__9118 (
            .O(N__63424),
            .I(N__63420));
    InMux I__9117 (
            .O(N__63423),
            .I(N__63417));
    Span4Mux_h I__9116 (
            .O(N__63420),
            .I(N__63412));
    LocalMux I__9115 (
            .O(N__63417),
            .I(N__63412));
    Span4Mux_v I__9114 (
            .O(N__63412),
            .I(N__63409));
    Span4Mux_v I__9113 (
            .O(N__63409),
            .I(N__63402));
    InMux I__9112 (
            .O(N__63408),
            .I(N__63397));
    InMux I__9111 (
            .O(N__63407),
            .I(N__63397));
    InMux I__9110 (
            .O(N__63406),
            .I(N__63394));
    InMux I__9109 (
            .O(N__63405),
            .I(N__63391));
    Span4Mux_h I__9108 (
            .O(N__63402),
            .I(N__63386));
    LocalMux I__9107 (
            .O(N__63397),
            .I(N__63386));
    LocalMux I__9106 (
            .O(N__63394),
            .I(N__63383));
    LocalMux I__9105 (
            .O(N__63391),
            .I(shift_srl_151Z0Z_15));
    Odrv4 I__9104 (
            .O(N__63386),
            .I(shift_srl_151Z0Z_15));
    Odrv12 I__9103 (
            .O(N__63383),
            .I(shift_srl_151Z0Z_15));
    InMux I__9102 (
            .O(N__63376),
            .I(N__63373));
    LocalMux I__9101 (
            .O(N__63373),
            .I(shift_srl_151Z0Z_9));
    InMux I__9100 (
            .O(N__63370),
            .I(N__63367));
    LocalMux I__9099 (
            .O(N__63367),
            .I(shift_srl_151Z0Z_7));
    InMux I__9098 (
            .O(N__63364),
            .I(N__63361));
    LocalMux I__9097 (
            .O(N__63361),
            .I(shift_srl_151Z0Z_8));
    CEMux I__9096 (
            .O(N__63358),
            .I(N__63354));
    CEMux I__9095 (
            .O(N__63357),
            .I(N__63351));
    LocalMux I__9094 (
            .O(N__63354),
            .I(N__63348));
    LocalMux I__9093 (
            .O(N__63351),
            .I(N__63345));
    Span4Mux_v I__9092 (
            .O(N__63348),
            .I(N__63342));
    Span4Mux_h I__9091 (
            .O(N__63345),
            .I(N__63339));
    Span4Mux_h I__9090 (
            .O(N__63342),
            .I(N__63336));
    Odrv4 I__9089 (
            .O(N__63339),
            .I(clk_en_151));
    Odrv4 I__9088 (
            .O(N__63336),
            .I(clk_en_151));
    InMux I__9087 (
            .O(N__63331),
            .I(N__63328));
    LocalMux I__9086 (
            .O(N__63328),
            .I(shift_srl_140Z0Z_10));
    InMux I__9085 (
            .O(N__63325),
            .I(N__63322));
    LocalMux I__9084 (
            .O(N__63322),
            .I(shift_srl_140Z0Z_11));
    InMux I__9083 (
            .O(N__63319),
            .I(N__63316));
    LocalMux I__9082 (
            .O(N__63316),
            .I(shift_srl_140Z0Z_12));
    InMux I__9081 (
            .O(N__63313),
            .I(N__63310));
    LocalMux I__9080 (
            .O(N__63310),
            .I(shift_srl_140Z0Z_13));
    InMux I__9079 (
            .O(N__63307),
            .I(N__63304));
    LocalMux I__9078 (
            .O(N__63304),
            .I(shift_srl_151Z0Z_2));
    InMux I__9077 (
            .O(N__63301),
            .I(N__63298));
    LocalMux I__9076 (
            .O(N__63298),
            .I(shift_srl_151Z0Z_3));
    InMux I__9075 (
            .O(N__63295),
            .I(N__63292));
    LocalMux I__9074 (
            .O(N__63292),
            .I(shift_srl_151Z0Z_4));
    InMux I__9073 (
            .O(N__63289),
            .I(N__63286));
    LocalMux I__9072 (
            .O(N__63286),
            .I(shift_srl_151Z0Z_5));
    InMux I__9071 (
            .O(N__63283),
            .I(N__63280));
    LocalMux I__9070 (
            .O(N__63280),
            .I(shift_srl_151Z0Z_6));
    InMux I__9069 (
            .O(N__63277),
            .I(N__63274));
    LocalMux I__9068 (
            .O(N__63274),
            .I(shift_srl_151Z0Z_10));
    InMux I__9067 (
            .O(N__63271),
            .I(N__63268));
    LocalMux I__9066 (
            .O(N__63268),
            .I(shift_srl_151Z0Z_11));
    InMux I__9065 (
            .O(N__63265),
            .I(N__63262));
    LocalMux I__9064 (
            .O(N__63262),
            .I(shift_srl_151Z0Z_12));
    CascadeMux I__9063 (
            .O(N__63259),
            .I(N__63256));
    InMux I__9062 (
            .O(N__63256),
            .I(N__63253));
    LocalMux I__9061 (
            .O(N__63253),
            .I(N__63249));
    InMux I__9060 (
            .O(N__63252),
            .I(N__63245));
    Span4Mux_h I__9059 (
            .O(N__63249),
            .I(N__63242));
    CascadeMux I__9058 (
            .O(N__63248),
            .I(N__63238));
    LocalMux I__9057 (
            .O(N__63245),
            .I(N__63235));
    Span4Mux_v I__9056 (
            .O(N__63242),
            .I(N__63232));
    InMux I__9055 (
            .O(N__63241),
            .I(N__63229));
    InMux I__9054 (
            .O(N__63238),
            .I(N__63226));
    Span4Mux_h I__9053 (
            .O(N__63235),
            .I(N__63223));
    Odrv4 I__9052 (
            .O(N__63232),
            .I(shift_srl_152Z0Z_15));
    LocalMux I__9051 (
            .O(N__63229),
            .I(shift_srl_152Z0Z_15));
    LocalMux I__9050 (
            .O(N__63226),
            .I(shift_srl_152Z0Z_15));
    Odrv4 I__9049 (
            .O(N__63223),
            .I(shift_srl_152Z0Z_15));
    CascadeMux I__9048 (
            .O(N__63214),
            .I(clk_en_0_a3_0_a2_sx_153_cascade_));
    CEMux I__9047 (
            .O(N__63211),
            .I(N__63207));
    CEMux I__9046 (
            .O(N__63210),
            .I(N__63204));
    LocalMux I__9045 (
            .O(N__63207),
            .I(clk_en_153));
    LocalMux I__9044 (
            .O(N__63204),
            .I(clk_en_153));
    CascadeMux I__9043 (
            .O(N__63199),
            .I(shift_srl_91_RNIUH4HPZ0Z_15_cascade_));
    CascadeMux I__9042 (
            .O(N__63196),
            .I(rco_c_145_cascade_));
    CEMux I__9041 (
            .O(N__63193),
            .I(N__63189));
    CEMux I__9040 (
            .O(N__63192),
            .I(N__63186));
    LocalMux I__9039 (
            .O(N__63189),
            .I(N__63181));
    LocalMux I__9038 (
            .O(N__63186),
            .I(N__63181));
    Odrv4 I__9037 (
            .O(N__63181),
            .I(clk_en_152));
    InMux I__9036 (
            .O(N__63178),
            .I(N__63175));
    LocalMux I__9035 (
            .O(N__63175),
            .I(shift_srl_151Z0Z_0));
    InMux I__9034 (
            .O(N__63172),
            .I(N__63169));
    LocalMux I__9033 (
            .O(N__63169),
            .I(shift_srl_151Z0Z_1));
    InMux I__9032 (
            .O(N__63166),
            .I(N__63163));
    LocalMux I__9031 (
            .O(N__63163),
            .I(shift_srl_24Z0Z_8));
    InMux I__9030 (
            .O(N__63160),
            .I(N__63157));
    LocalMux I__9029 (
            .O(N__63157),
            .I(shift_srl_24Z0Z_9));
    CEMux I__9028 (
            .O(N__63154),
            .I(N__63151));
    LocalMux I__9027 (
            .O(N__63151),
            .I(N__63146));
    CEMux I__9026 (
            .O(N__63150),
            .I(N__63143));
    CEMux I__9025 (
            .O(N__63149),
            .I(N__63140));
    Span4Mux_h I__9024 (
            .O(N__63146),
            .I(N__63135));
    LocalMux I__9023 (
            .O(N__63143),
            .I(N__63135));
    LocalMux I__9022 (
            .O(N__63140),
            .I(N__63132));
    Span4Mux_h I__9021 (
            .O(N__63135),
            .I(N__63129));
    Odrv12 I__9020 (
            .O(N__63132),
            .I(clk_en_24));
    Odrv4 I__9019 (
            .O(N__63129),
            .I(clk_en_24));
    InMux I__9018 (
            .O(N__63124),
            .I(N__63121));
    LocalMux I__9017 (
            .O(N__63121),
            .I(shift_srl_152Z0Z_0));
    InMux I__9016 (
            .O(N__63118),
            .I(N__63115));
    LocalMux I__9015 (
            .O(N__63115),
            .I(shift_srl_152Z0Z_1));
    InMux I__9014 (
            .O(N__63112),
            .I(N__63109));
    LocalMux I__9013 (
            .O(N__63109),
            .I(shift_srl_152Z0Z_2));
    InMux I__9012 (
            .O(N__63106),
            .I(N__63103));
    LocalMux I__9011 (
            .O(N__63103),
            .I(shift_srl_152Z0Z_3));
    InMux I__9010 (
            .O(N__63100),
            .I(N__63097));
    LocalMux I__9009 (
            .O(N__63097),
            .I(shift_srl_152Z0Z_4));
    InMux I__9008 (
            .O(N__63094),
            .I(N__63091));
    LocalMux I__9007 (
            .O(N__63091),
            .I(shift_srl_152Z0Z_5));
    InMux I__9006 (
            .O(N__63088),
            .I(N__63085));
    LocalMux I__9005 (
            .O(N__63085),
            .I(shift_srl_152Z0Z_6));
    InMux I__9004 (
            .O(N__63082),
            .I(N__63079));
    LocalMux I__9003 (
            .O(N__63079),
            .I(shift_srl_152Z0Z_7));
    InMux I__9002 (
            .O(N__63076),
            .I(N__63073));
    LocalMux I__9001 (
            .O(N__63073),
            .I(shift_srl_43Z0Z_0));
    InMux I__9000 (
            .O(N__63070),
            .I(N__63067));
    LocalMux I__8999 (
            .O(N__63067),
            .I(shift_srl_43Z0Z_1));
    InMux I__8998 (
            .O(N__63064),
            .I(N__63061));
    LocalMux I__8997 (
            .O(N__63061),
            .I(shift_srl_43Z0Z_6));
    InMux I__8996 (
            .O(N__63058),
            .I(N__63055));
    LocalMux I__8995 (
            .O(N__63055),
            .I(shift_srl_43Z0Z_7));
    InMux I__8994 (
            .O(N__63052),
            .I(N__63049));
    LocalMux I__8993 (
            .O(N__63049),
            .I(shift_srl_24Z0Z_10));
    InMux I__8992 (
            .O(N__63046),
            .I(N__63043));
    LocalMux I__8991 (
            .O(N__63043),
            .I(shift_srl_24Z0Z_11));
    InMux I__8990 (
            .O(N__63040),
            .I(N__63037));
    LocalMux I__8989 (
            .O(N__63037),
            .I(shift_srl_24Z0Z_12));
    InMux I__8988 (
            .O(N__63034),
            .I(N__63031));
    LocalMux I__8987 (
            .O(N__63031),
            .I(shift_srl_24Z0Z_13));
    InMux I__8986 (
            .O(N__63028),
            .I(N__63025));
    LocalMux I__8985 (
            .O(N__63025),
            .I(shift_srl_24Z0Z_14));
    InMux I__8984 (
            .O(N__63022),
            .I(N__63019));
    LocalMux I__8983 (
            .O(N__63019),
            .I(shift_srl_43Z0Z_13));
    InMux I__8982 (
            .O(N__63016),
            .I(N__63013));
    LocalMux I__8981 (
            .O(N__63013),
            .I(shift_srl_43Z0Z_14));
    InMux I__8980 (
            .O(N__63010),
            .I(N__63007));
    LocalMux I__8979 (
            .O(N__63007),
            .I(shift_srl_43Z0Z_9));
    InMux I__8978 (
            .O(N__63004),
            .I(N__63001));
    LocalMux I__8977 (
            .O(N__63001),
            .I(shift_srl_43Z0Z_8));
    InMux I__8976 (
            .O(N__62998),
            .I(N__62995));
    LocalMux I__8975 (
            .O(N__62995),
            .I(shift_srl_43Z0Z_2));
    InMux I__8974 (
            .O(N__62992),
            .I(N__62989));
    LocalMux I__8973 (
            .O(N__62989),
            .I(shift_srl_43Z0Z_3));
    InMux I__8972 (
            .O(N__62986),
            .I(N__62983));
    LocalMux I__8971 (
            .O(N__62983),
            .I(shift_srl_43Z0Z_4));
    InMux I__8970 (
            .O(N__62980),
            .I(N__62977));
    LocalMux I__8969 (
            .O(N__62977),
            .I(shift_srl_43Z0Z_5));
    InMux I__8968 (
            .O(N__62974),
            .I(N__62971));
    LocalMux I__8967 (
            .O(N__62971),
            .I(shift_srl_86Z0Z_5));
    InMux I__8966 (
            .O(N__62968),
            .I(N__62965));
    LocalMux I__8965 (
            .O(N__62965),
            .I(shift_srl_86Z0Z_6));
    InMux I__8964 (
            .O(N__62962),
            .I(N__62959));
    LocalMux I__8963 (
            .O(N__62959),
            .I(shift_srl_86Z0Z_12));
    InMux I__8962 (
            .O(N__62956),
            .I(N__62953));
    LocalMux I__8961 (
            .O(N__62953),
            .I(shift_srl_86Z0Z_13));
    InMux I__8960 (
            .O(N__62950),
            .I(N__62947));
    LocalMux I__8959 (
            .O(N__62947),
            .I(shift_srl_86Z0Z_9));
    InMux I__8958 (
            .O(N__62944),
            .I(N__62941));
    LocalMux I__8957 (
            .O(N__62941),
            .I(shift_srl_86Z0Z_7));
    InMux I__8956 (
            .O(N__62938),
            .I(N__62935));
    LocalMux I__8955 (
            .O(N__62935),
            .I(shift_srl_86Z0Z_8));
    InMux I__8954 (
            .O(N__62932),
            .I(N__62929));
    LocalMux I__8953 (
            .O(N__62929),
            .I(shift_srl_43Z0Z_11));
    InMux I__8952 (
            .O(N__62926),
            .I(N__62923));
    LocalMux I__8951 (
            .O(N__62923),
            .I(shift_srl_43Z0Z_10));
    InMux I__8950 (
            .O(N__62920),
            .I(N__62917));
    LocalMux I__8949 (
            .O(N__62917),
            .I(shift_srl_43Z0Z_12));
    InMux I__8948 (
            .O(N__62914),
            .I(N__62911));
    LocalMux I__8947 (
            .O(N__62911),
            .I(shift_srl_88Z0Z_8));
    IoInMux I__8946 (
            .O(N__62908),
            .I(N__62905));
    LocalMux I__8945 (
            .O(N__62905),
            .I(N__62902));
    Span4Mux_s3_v I__8944 (
            .O(N__62902),
            .I(N__62899));
    Span4Mux_h I__8943 (
            .O(N__62899),
            .I(N__62896));
    Odrv4 I__8942 (
            .O(N__62896),
            .I(rco_c_88));
    CascadeMux I__8941 (
            .O(N__62893),
            .I(rco_c_83_cascade_));
    InMux I__8940 (
            .O(N__62890),
            .I(N__62885));
    InMux I__8939 (
            .O(N__62889),
            .I(N__62882));
    CascadeMux I__8938 (
            .O(N__62888),
            .I(N__62878));
    LocalMux I__8937 (
            .O(N__62885),
            .I(N__62872));
    LocalMux I__8936 (
            .O(N__62882),
            .I(N__62872));
    InMux I__8935 (
            .O(N__62881),
            .I(N__62865));
    InMux I__8934 (
            .O(N__62878),
            .I(N__62865));
    InMux I__8933 (
            .O(N__62877),
            .I(N__62865));
    Span4Mux_v I__8932 (
            .O(N__62872),
            .I(N__62860));
    LocalMux I__8931 (
            .O(N__62865),
            .I(N__62860));
    Span4Mux_v I__8930 (
            .O(N__62860),
            .I(N__62855));
    InMux I__8929 (
            .O(N__62859),
            .I(N__62850));
    InMux I__8928 (
            .O(N__62858),
            .I(N__62850));
    Odrv4 I__8927 (
            .O(N__62855),
            .I(shift_srl_86_RNI8K1LZ0Z_15));
    LocalMux I__8926 (
            .O(N__62850),
            .I(shift_srl_86_RNI8K1LZ0Z_15));
    InMux I__8925 (
            .O(N__62845),
            .I(N__62842));
    LocalMux I__8924 (
            .O(N__62842),
            .I(shift_srl_86Z0Z_10));
    InMux I__8923 (
            .O(N__62839),
            .I(N__62836));
    LocalMux I__8922 (
            .O(N__62836),
            .I(shift_srl_85Z0Z_9));
    InMux I__8921 (
            .O(N__62833),
            .I(N__62830));
    LocalMux I__8920 (
            .O(N__62830),
            .I(shift_srl_85Z0Z_8));
    InMux I__8919 (
            .O(N__62827),
            .I(N__62824));
    LocalMux I__8918 (
            .O(N__62824),
            .I(shift_srl_88Z0Z_10));
    InMux I__8917 (
            .O(N__62821),
            .I(N__62818));
    LocalMux I__8916 (
            .O(N__62818),
            .I(shift_srl_88Z0Z_11));
    InMux I__8915 (
            .O(N__62815),
            .I(N__62812));
    LocalMux I__8914 (
            .O(N__62812),
            .I(shift_srl_88Z0Z_12));
    InMux I__8913 (
            .O(N__62809),
            .I(N__62806));
    LocalMux I__8912 (
            .O(N__62806),
            .I(shift_srl_88Z0Z_13));
    InMux I__8911 (
            .O(N__62803),
            .I(N__62800));
    LocalMux I__8910 (
            .O(N__62800),
            .I(shift_srl_88Z0Z_14));
    InMux I__8909 (
            .O(N__62797),
            .I(N__62794));
    LocalMux I__8908 (
            .O(N__62794),
            .I(shift_srl_88Z0Z_9));
    InMux I__8907 (
            .O(N__62791),
            .I(N__62788));
    LocalMux I__8906 (
            .O(N__62788),
            .I(N__62785));
    Span4Mux_v I__8905 (
            .O(N__62785),
            .I(N__62782));
    Odrv4 I__8904 (
            .O(N__62782),
            .I(shift_srl_139Z0Z_7));
    InMux I__8903 (
            .O(N__62779),
            .I(N__62776));
    LocalMux I__8902 (
            .O(N__62776),
            .I(shift_srl_139Z0Z_8));
    InMux I__8901 (
            .O(N__62773),
            .I(N__62770));
    LocalMux I__8900 (
            .O(N__62770),
            .I(shift_srl_139Z0Z_9));
    InMux I__8899 (
            .O(N__62767),
            .I(N__62764));
    LocalMux I__8898 (
            .O(N__62764),
            .I(shift_srl_139Z0Z_10));
    InMux I__8897 (
            .O(N__62761),
            .I(N__62758));
    LocalMux I__8896 (
            .O(N__62758),
            .I(shift_srl_85Z0Z_10));
    InMux I__8895 (
            .O(N__62755),
            .I(N__62752));
    LocalMux I__8894 (
            .O(N__62752),
            .I(shift_srl_85Z0Z_11));
    InMux I__8893 (
            .O(N__62749),
            .I(N__62746));
    LocalMux I__8892 (
            .O(N__62746),
            .I(shift_srl_85Z0Z_12));
    InMux I__8891 (
            .O(N__62743),
            .I(N__62740));
    LocalMux I__8890 (
            .O(N__62740),
            .I(shift_srl_85Z0Z_13));
    InMux I__8889 (
            .O(N__62737),
            .I(N__62734));
    LocalMux I__8888 (
            .O(N__62734),
            .I(shift_srl_85Z0Z_14));
    CEMux I__8887 (
            .O(N__62731),
            .I(N__62728));
    LocalMux I__8886 (
            .O(N__62728),
            .I(N__62725));
    Span4Mux_h I__8885 (
            .O(N__62725),
            .I(N__62722));
    Span4Mux_h I__8884 (
            .O(N__62722),
            .I(N__62717));
    CEMux I__8883 (
            .O(N__62721),
            .I(N__62714));
    CEMux I__8882 (
            .O(N__62720),
            .I(N__62711));
    Odrv4 I__8881 (
            .O(N__62717),
            .I(clk_en_199));
    LocalMux I__8880 (
            .O(N__62714),
            .I(clk_en_199));
    LocalMux I__8879 (
            .O(N__62711),
            .I(clk_en_199));
    InMux I__8878 (
            .O(N__62704),
            .I(N__62699));
    InMux I__8877 (
            .O(N__62703),
            .I(N__62693));
    InMux I__8876 (
            .O(N__62702),
            .I(N__62690));
    LocalMux I__8875 (
            .O(N__62699),
            .I(N__62687));
    InMux I__8874 (
            .O(N__62698),
            .I(N__62680));
    InMux I__8873 (
            .O(N__62697),
            .I(N__62680));
    InMux I__8872 (
            .O(N__62696),
            .I(N__62680));
    LocalMux I__8871 (
            .O(N__62693),
            .I(shift_srl_102Z0Z_15));
    LocalMux I__8870 (
            .O(N__62690),
            .I(shift_srl_102Z0Z_15));
    Odrv4 I__8869 (
            .O(N__62687),
            .I(shift_srl_102Z0Z_15));
    LocalMux I__8868 (
            .O(N__62680),
            .I(shift_srl_102Z0Z_15));
    InMux I__8867 (
            .O(N__62671),
            .I(N__62668));
    LocalMux I__8866 (
            .O(N__62668),
            .I(shift_srl_102Z0Z_0));
    InMux I__8865 (
            .O(N__62665),
            .I(N__62662));
    LocalMux I__8864 (
            .O(N__62662),
            .I(shift_srl_102Z0Z_1));
    InMux I__8863 (
            .O(N__62659),
            .I(N__62656));
    LocalMux I__8862 (
            .O(N__62656),
            .I(shift_srl_102Z0Z_2));
    InMux I__8861 (
            .O(N__62653),
            .I(N__62650));
    LocalMux I__8860 (
            .O(N__62650),
            .I(shift_srl_102Z0Z_3));
    InMux I__8859 (
            .O(N__62647),
            .I(N__62644));
    LocalMux I__8858 (
            .O(N__62644),
            .I(shift_srl_102Z0Z_4));
    InMux I__8857 (
            .O(N__62641),
            .I(N__62638));
    LocalMux I__8856 (
            .O(N__62638),
            .I(shift_srl_102Z0Z_5));
    InMux I__8855 (
            .O(N__62635),
            .I(N__62632));
    LocalMux I__8854 (
            .O(N__62632),
            .I(shift_srl_102Z0Z_6));
    InMux I__8853 (
            .O(N__62629),
            .I(N__62626));
    LocalMux I__8852 (
            .O(N__62626),
            .I(shift_srl_102Z0Z_8));
    InMux I__8851 (
            .O(N__62623),
            .I(N__62620));
    LocalMux I__8850 (
            .O(N__62620),
            .I(shift_srl_102Z0Z_9));
    CEMux I__8849 (
            .O(N__62617),
            .I(N__62614));
    LocalMux I__8848 (
            .O(N__62614),
            .I(N__62611));
    Span4Mux_v I__8847 (
            .O(N__62611),
            .I(N__62607));
    CEMux I__8846 (
            .O(N__62610),
            .I(N__62604));
    Span4Mux_h I__8845 (
            .O(N__62607),
            .I(N__62601));
    LocalMux I__8844 (
            .O(N__62604),
            .I(N__62598));
    Odrv4 I__8843 (
            .O(N__62601),
            .I(clk_en_102));
    Odrv12 I__8842 (
            .O(N__62598),
            .I(clk_en_102));
    CascadeMux I__8841 (
            .O(N__62593),
            .I(N__62590));
    InMux I__8840 (
            .O(N__62590),
            .I(N__62582));
    InMux I__8839 (
            .O(N__62589),
            .I(N__62577));
    InMux I__8838 (
            .O(N__62588),
            .I(N__62577));
    InMux I__8837 (
            .O(N__62587),
            .I(N__62574));
    InMux I__8836 (
            .O(N__62586),
            .I(N__62569));
    InMux I__8835 (
            .O(N__62585),
            .I(N__62569));
    LocalMux I__8834 (
            .O(N__62582),
            .I(N__62566));
    LocalMux I__8833 (
            .O(N__62577),
            .I(N__62561));
    LocalMux I__8832 (
            .O(N__62574),
            .I(N__62561));
    LocalMux I__8831 (
            .O(N__62569),
            .I(N__62558));
    Span4Mux_h I__8830 (
            .O(N__62566),
            .I(N__62555));
    Span4Mux_v I__8829 (
            .O(N__62561),
            .I(N__62552));
    Span12Mux_h I__8828 (
            .O(N__62558),
            .I(N__62549));
    Odrv4 I__8827 (
            .O(N__62555),
            .I(rco_int_0_a2_1_a2_out_0));
    Odrv4 I__8826 (
            .O(N__62552),
            .I(rco_int_0_a2_1_a2_out_0));
    Odrv12 I__8825 (
            .O(N__62549),
            .I(rco_int_0_a2_1_a2_out_0));
    InMux I__8824 (
            .O(N__62542),
            .I(N__62539));
    LocalMux I__8823 (
            .O(N__62539),
            .I(g0_8));
    InMux I__8822 (
            .O(N__62536),
            .I(N__62533));
    LocalMux I__8821 (
            .O(N__62533),
            .I(shift_srl_199Z0Z_10));
    InMux I__8820 (
            .O(N__62530),
            .I(N__62527));
    LocalMux I__8819 (
            .O(N__62527),
            .I(shift_srl_199Z0Z_11));
    InMux I__8818 (
            .O(N__62524),
            .I(N__62521));
    LocalMux I__8817 (
            .O(N__62521),
            .I(shift_srl_199Z0Z_12));
    InMux I__8816 (
            .O(N__62518),
            .I(N__62515));
    LocalMux I__8815 (
            .O(N__62515),
            .I(shift_srl_199Z0Z_13));
    InMux I__8814 (
            .O(N__62512),
            .I(N__62509));
    LocalMux I__8813 (
            .O(N__62509),
            .I(shift_srl_199Z0Z_14));
    InMux I__8812 (
            .O(N__62506),
            .I(N__62500));
    InMux I__8811 (
            .O(N__62505),
            .I(N__62500));
    LocalMux I__8810 (
            .O(N__62500),
            .I(shift_srl_199Z0Z_15));
    InMux I__8809 (
            .O(N__62497),
            .I(N__62494));
    LocalMux I__8808 (
            .O(N__62494),
            .I(shift_srl_199Z0Z_9));
    InMux I__8807 (
            .O(N__62491),
            .I(N__62488));
    LocalMux I__8806 (
            .O(N__62488),
            .I(N__62485));
    Span4Mux_h I__8805 (
            .O(N__62485),
            .I(N__62482));
    Span4Mux_h I__8804 (
            .O(N__62482),
            .I(N__62479));
    Odrv4 I__8803 (
            .O(N__62479),
            .I(shift_srl_199Z0Z_7));
    InMux I__8802 (
            .O(N__62476),
            .I(N__62473));
    LocalMux I__8801 (
            .O(N__62473),
            .I(shift_srl_199Z0Z_8));
    InMux I__8800 (
            .O(N__62470),
            .I(N__62467));
    LocalMux I__8799 (
            .O(N__62467),
            .I(N__62464));
    Span4Mux_h I__8798 (
            .O(N__62464),
            .I(N__62461));
    Span4Mux_h I__8797 (
            .O(N__62461),
            .I(N__62458));
    Odrv4 I__8796 (
            .O(N__62458),
            .I(shift_srl_110Z0Z_14));
    CEMux I__8795 (
            .O(N__62455),
            .I(N__62452));
    LocalMux I__8794 (
            .O(N__62452),
            .I(N__62449));
    Span4Mux_h I__8793 (
            .O(N__62449),
            .I(N__62444));
    CEMux I__8792 (
            .O(N__62448),
            .I(N__62441));
    CEMux I__8791 (
            .O(N__62447),
            .I(N__62438));
    Odrv4 I__8790 (
            .O(N__62444),
            .I(clk_en_110));
    LocalMux I__8789 (
            .O(N__62441),
            .I(clk_en_110));
    LocalMux I__8788 (
            .O(N__62438),
            .I(clk_en_110));
    InMux I__8787 (
            .O(N__62431),
            .I(N__62428));
    LocalMux I__8786 (
            .O(N__62428),
            .I(N__62425));
    Span4Mux_v I__8785 (
            .O(N__62425),
            .I(N__62420));
    InMux I__8784 (
            .O(N__62424),
            .I(N__62415));
    InMux I__8783 (
            .O(N__62423),
            .I(N__62415));
    Odrv4 I__8782 (
            .O(N__62420),
            .I(shift_srl_110Z0Z_15));
    LocalMux I__8781 (
            .O(N__62415),
            .I(shift_srl_110Z0Z_15));
    InMux I__8780 (
            .O(N__62410),
            .I(N__62407));
    LocalMux I__8779 (
            .O(N__62407),
            .I(N__62404));
    Sp12to4 I__8778 (
            .O(N__62404),
            .I(N__62397));
    InMux I__8777 (
            .O(N__62403),
            .I(N__62392));
    InMux I__8776 (
            .O(N__62402),
            .I(N__62392));
    InMux I__8775 (
            .O(N__62401),
            .I(N__62389));
    InMux I__8774 (
            .O(N__62400),
            .I(N__62386));
    Span12Mux_s9_v I__8773 (
            .O(N__62397),
            .I(N__62381));
    LocalMux I__8772 (
            .O(N__62392),
            .I(N__62381));
    LocalMux I__8771 (
            .O(N__62389),
            .I(shift_srl_109Z0Z_15));
    LocalMux I__8770 (
            .O(N__62386),
            .I(shift_srl_109Z0Z_15));
    Odrv12 I__8769 (
            .O(N__62381),
            .I(shift_srl_109Z0Z_15));
    CascadeMux I__8768 (
            .O(N__62374),
            .I(N__62367));
    InMux I__8767 (
            .O(N__62373),
            .I(N__62362));
    InMux I__8766 (
            .O(N__62372),
            .I(N__62362));
    InMux I__8765 (
            .O(N__62371),
            .I(N__62359));
    InMux I__8764 (
            .O(N__62370),
            .I(N__62355));
    InMux I__8763 (
            .O(N__62367),
            .I(N__62352));
    LocalMux I__8762 (
            .O(N__62362),
            .I(N__62349));
    LocalMux I__8761 (
            .O(N__62359),
            .I(N__62346));
    InMux I__8760 (
            .O(N__62358),
            .I(N__62341));
    LocalMux I__8759 (
            .O(N__62355),
            .I(N__62336));
    LocalMux I__8758 (
            .O(N__62352),
            .I(N__62336));
    Span12Mux_s7_v I__8757 (
            .O(N__62349),
            .I(N__62333));
    Span4Mux_v I__8756 (
            .O(N__62346),
            .I(N__62330));
    InMux I__8755 (
            .O(N__62345),
            .I(N__62325));
    InMux I__8754 (
            .O(N__62344),
            .I(N__62325));
    LocalMux I__8753 (
            .O(N__62341),
            .I(N__62322));
    Span4Mux_h I__8752 (
            .O(N__62336),
            .I(N__62319));
    Odrv12 I__8751 (
            .O(N__62333),
            .I(shift_srl_107Z0Z_15));
    Odrv4 I__8750 (
            .O(N__62330),
            .I(shift_srl_107Z0Z_15));
    LocalMux I__8749 (
            .O(N__62325),
            .I(shift_srl_107Z0Z_15));
    Odrv4 I__8748 (
            .O(N__62322),
            .I(shift_srl_107Z0Z_15));
    Odrv4 I__8747 (
            .O(N__62319),
            .I(shift_srl_107Z0Z_15));
    InMux I__8746 (
            .O(N__62308),
            .I(N__62305));
    LocalMux I__8745 (
            .O(N__62305),
            .I(N__62299));
    InMux I__8744 (
            .O(N__62304),
            .I(N__62296));
    InMux I__8743 (
            .O(N__62303),
            .I(N__62289));
    InMux I__8742 (
            .O(N__62302),
            .I(N__62289));
    Span12Mux_s9_h I__8741 (
            .O(N__62299),
            .I(N__62284));
    LocalMux I__8740 (
            .O(N__62296),
            .I(N__62284));
    InMux I__8739 (
            .O(N__62295),
            .I(N__62279));
    InMux I__8738 (
            .O(N__62294),
            .I(N__62279));
    LocalMux I__8737 (
            .O(N__62289),
            .I(N__62276));
    Odrv12 I__8736 (
            .O(N__62284),
            .I(shift_srl_108Z0Z_15));
    LocalMux I__8735 (
            .O(N__62279),
            .I(shift_srl_108Z0Z_15));
    Odrv12 I__8734 (
            .O(N__62276),
            .I(shift_srl_108Z0Z_15));
    InMux I__8733 (
            .O(N__62269),
            .I(N__62263));
    InMux I__8732 (
            .O(N__62268),
            .I(N__62263));
    LocalMux I__8731 (
            .O(N__62263),
            .I(N__62260));
    Span4Mux_h I__8730 (
            .O(N__62260),
            .I(N__62257));
    Odrv4 I__8729 (
            .O(N__62257),
            .I(rco_int_0_a3_0_a2_s_0_1_104));
    CascadeMux I__8728 (
            .O(N__62254),
            .I(shift_srl_110_RNI91581Z0Z_15_cascade_));
    InMux I__8727 (
            .O(N__62251),
            .I(N__62245));
    InMux I__8726 (
            .O(N__62250),
            .I(N__62245));
    LocalMux I__8725 (
            .O(N__62245),
            .I(N__62242));
    Span4Mux_h I__8724 (
            .O(N__62242),
            .I(N__62239));
    Odrv4 I__8723 (
            .O(N__62239),
            .I(rco_int_0_a2_0_a2_s_0_sx_110));
    InMux I__8722 (
            .O(N__62236),
            .I(N__62232));
    InMux I__8721 (
            .O(N__62235),
            .I(N__62229));
    LocalMux I__8720 (
            .O(N__62232),
            .I(N__62226));
    LocalMux I__8719 (
            .O(N__62229),
            .I(N__62221));
    Span4Mux_h I__8718 (
            .O(N__62226),
            .I(N__62221));
    Odrv4 I__8717 (
            .O(N__62221),
            .I(rco_int_0_a3_0_a2_138_m6_0_a2_7_4));
    CascadeMux I__8716 (
            .O(N__62218),
            .I(shift_srl_110_RNI4QDG2Z0Z_15_cascade_));
    InMux I__8715 (
            .O(N__62215),
            .I(N__62212));
    LocalMux I__8714 (
            .O(N__62212),
            .I(N__62209));
    Span4Mux_h I__8713 (
            .O(N__62209),
            .I(N__62206));
    Span4Mux_h I__8712 (
            .O(N__62206),
            .I(N__62203));
    Odrv4 I__8711 (
            .O(N__62203),
            .I(g0_4));
    InMux I__8710 (
            .O(N__62200),
            .I(N__62197));
    LocalMux I__8709 (
            .O(N__62197),
            .I(N__62194));
    Span4Mux_h I__8708 (
            .O(N__62194),
            .I(N__62191));
    Span4Mux_h I__8707 (
            .O(N__62191),
            .I(N__62188));
    Span4Mux_h I__8706 (
            .O(N__62188),
            .I(N__62185));
    Odrv4 I__8705 (
            .O(N__62185),
            .I(g0_0));
    InMux I__8704 (
            .O(N__62182),
            .I(N__62177));
    InMux I__8703 (
            .O(N__62181),
            .I(N__62174));
    InMux I__8702 (
            .O(N__62180),
            .I(N__62171));
    LocalMux I__8701 (
            .O(N__62177),
            .I(N__62168));
    LocalMux I__8700 (
            .O(N__62174),
            .I(N__62165));
    LocalMux I__8699 (
            .O(N__62171),
            .I(N__62162));
    Span4Mux_v I__8698 (
            .O(N__62168),
            .I(N__62157));
    Span4Mux_v I__8697 (
            .O(N__62165),
            .I(N__62157));
    Span4Mux_v I__8696 (
            .O(N__62162),
            .I(N__62152));
    Span4Mux_h I__8695 (
            .O(N__62157),
            .I(N__62152));
    Span4Mux_h I__8694 (
            .O(N__62152),
            .I(N__62148));
    InMux I__8693 (
            .O(N__62151),
            .I(N__62145));
    Odrv4 I__8692 (
            .O(N__62148),
            .I(rco_int_0_a3_0_a2_0_132));
    LocalMux I__8691 (
            .O(N__62145),
            .I(rco_int_0_a3_0_a2_0_132));
    CascadeMux I__8690 (
            .O(N__62140),
            .I(g0_9_cascade_));
    CascadeMux I__8689 (
            .O(N__62137),
            .I(g0_16_cascade_));
    InMux I__8688 (
            .O(N__62134),
            .I(N__62131));
    LocalMux I__8687 (
            .O(N__62131),
            .I(N__62126));
    InMux I__8686 (
            .O(N__62130),
            .I(N__62122));
    InMux I__8685 (
            .O(N__62129),
            .I(N__62119));
    Span4Mux_v I__8684 (
            .O(N__62126),
            .I(N__62116));
    InMux I__8683 (
            .O(N__62125),
            .I(N__62113));
    LocalMux I__8682 (
            .O(N__62122),
            .I(N__62110));
    LocalMux I__8681 (
            .O(N__62119),
            .I(N__62107));
    Sp12to4 I__8680 (
            .O(N__62116),
            .I(N__62102));
    LocalMux I__8679 (
            .O(N__62113),
            .I(N__62102));
    Span4Mux_v I__8678 (
            .O(N__62110),
            .I(N__62097));
    Span4Mux_h I__8677 (
            .O(N__62107),
            .I(N__62097));
    Span12Mux_h I__8676 (
            .O(N__62102),
            .I(N__62094));
    Span4Mux_h I__8675 (
            .O(N__62097),
            .I(N__62091));
    Odrv12 I__8674 (
            .O(N__62094),
            .I(rco_int_0_a3_0_a2_0_138));
    Odrv4 I__8673 (
            .O(N__62091),
            .I(rco_int_0_a3_0_a2_0_138));
    InMux I__8672 (
            .O(N__62086),
            .I(N__62083));
    LocalMux I__8671 (
            .O(N__62083),
            .I(g0_12));
    InMux I__8670 (
            .O(N__62080),
            .I(N__62077));
    LocalMux I__8669 (
            .O(N__62077),
            .I(shift_srl_139Z0Z_2));
    InMux I__8668 (
            .O(N__62074),
            .I(N__62071));
    LocalMux I__8667 (
            .O(N__62071),
            .I(shift_srl_139Z0Z_3));
    InMux I__8666 (
            .O(N__62068),
            .I(N__62065));
    LocalMux I__8665 (
            .O(N__62065),
            .I(shift_srl_139Z0Z_4));
    InMux I__8664 (
            .O(N__62062),
            .I(N__62059));
    LocalMux I__8663 (
            .O(N__62059),
            .I(shift_srl_139Z0Z_5));
    InMux I__8662 (
            .O(N__62056),
            .I(N__62053));
    LocalMux I__8661 (
            .O(N__62053),
            .I(shift_srl_139Z0Z_6));
    CascadeMux I__8660 (
            .O(N__62050),
            .I(rco_int_0_a2_0_a2_s_0_1_110_cascade_));
    CascadeMux I__8659 (
            .O(N__62047),
            .I(rco_int_0_a2_0_a2_out_5_cascade_));
    CascadeMux I__8658 (
            .O(N__62044),
            .I(rco_int_0_a3_0_a2_138_m6_0_a2_7_cascade_));
    CEMux I__8657 (
            .O(N__62041),
            .I(N__62038));
    LocalMux I__8656 (
            .O(N__62038),
            .I(N__62033));
    CEMux I__8655 (
            .O(N__62037),
            .I(N__62030));
    CEMux I__8654 (
            .O(N__62036),
            .I(N__62027));
    Span4Mux_h I__8653 (
            .O(N__62033),
            .I(N__62022));
    LocalMux I__8652 (
            .O(N__62030),
            .I(N__62022));
    LocalMux I__8651 (
            .O(N__62027),
            .I(N__62019));
    Span4Mux_v I__8650 (
            .O(N__62022),
            .I(N__62016));
    Odrv4 I__8649 (
            .O(N__62019),
            .I(N_122_i));
    Odrv4 I__8648 (
            .O(N__62016),
            .I(N_122_i));
    IoInMux I__8647 (
            .O(N__62011),
            .I(N__62008));
    LocalMux I__8646 (
            .O(N__62008),
            .I(N__62005));
    Span4Mux_s3_h I__8645 (
            .O(N__62005),
            .I(N__62001));
    InMux I__8644 (
            .O(N__62004),
            .I(N__61995));
    Span4Mux_h I__8643 (
            .O(N__62001),
            .I(N__61992));
    InMux I__8642 (
            .O(N__62000),
            .I(N__61986));
    InMux I__8641 (
            .O(N__61999),
            .I(N__61986));
    InMux I__8640 (
            .O(N__61998),
            .I(N__61983));
    LocalMux I__8639 (
            .O(N__61995),
            .I(N__61980));
    Span4Mux_h I__8638 (
            .O(N__61992),
            .I(N__61977));
    InMux I__8637 (
            .O(N__61991),
            .I(N__61968));
    LocalMux I__8636 (
            .O(N__61986),
            .I(N__61965));
    LocalMux I__8635 (
            .O(N__61983),
            .I(N__61960));
    Span4Mux_h I__8634 (
            .O(N__61980),
            .I(N__61960));
    Span4Mux_h I__8633 (
            .O(N__61977),
            .I(N__61957));
    InMux I__8632 (
            .O(N__61976),
            .I(N__61952));
    InMux I__8631 (
            .O(N__61975),
            .I(N__61952));
    InMux I__8630 (
            .O(N__61974),
            .I(N__61943));
    InMux I__8629 (
            .O(N__61973),
            .I(N__61943));
    InMux I__8628 (
            .O(N__61972),
            .I(N__61943));
    InMux I__8627 (
            .O(N__61971),
            .I(N__61943));
    LocalMux I__8626 (
            .O(N__61968),
            .I(N__61940));
    Span4Mux_h I__8625 (
            .O(N__61965),
            .I(N__61935));
    Span4Mux_h I__8624 (
            .O(N__61960),
            .I(N__61935));
    Span4Mux_h I__8623 (
            .O(N__61957),
            .I(N__61932));
    LocalMux I__8622 (
            .O(N__61952),
            .I(N__61929));
    LocalMux I__8621 (
            .O(N__61943),
            .I(N__61924));
    Span4Mux_h I__8620 (
            .O(N__61940),
            .I(N__61924));
    Span4Mux_h I__8619 (
            .O(N__61935),
            .I(N__61921));
    Odrv4 I__8618 (
            .O(N__61932),
            .I(rco_c_110));
    Odrv12 I__8617 (
            .O(N__61929),
            .I(rco_c_110));
    Odrv4 I__8616 (
            .O(N__61924),
            .I(rco_c_110));
    Odrv4 I__8615 (
            .O(N__61921),
            .I(rco_c_110));
    InMux I__8614 (
            .O(N__61912),
            .I(N__61909));
    LocalMux I__8613 (
            .O(N__61909),
            .I(rco_int_0_a3_0_a2_138_m6_0_a2_7_4_1));
    InMux I__8612 (
            .O(N__61906),
            .I(N__61903));
    LocalMux I__8611 (
            .O(N__61903),
            .I(N__61900));
    Odrv4 I__8610 (
            .O(N__61900),
            .I(rco_int_0_a3_0_a2_138_m6_0_a2_7_0));
    InMux I__8609 (
            .O(N__61897),
            .I(N__61894));
    LocalMux I__8608 (
            .O(N__61894),
            .I(shift_srl_120_RNIG17D2Z0Z_15));
    InMux I__8607 (
            .O(N__61891),
            .I(N__61888));
    LocalMux I__8606 (
            .O(N__61888),
            .I(shift_srl_139Z0Z_0));
    InMux I__8605 (
            .O(N__61885),
            .I(N__61882));
    LocalMux I__8604 (
            .O(N__61882),
            .I(shift_srl_139Z0Z_1));
    InMux I__8603 (
            .O(N__61879),
            .I(N__61876));
    LocalMux I__8602 (
            .O(N__61876),
            .I(shift_srl_145Z0Z_10));
    InMux I__8601 (
            .O(N__61873),
            .I(N__61870));
    LocalMux I__8600 (
            .O(N__61870),
            .I(shift_srl_145Z0Z_11));
    InMux I__8599 (
            .O(N__61867),
            .I(N__61864));
    LocalMux I__8598 (
            .O(N__61864),
            .I(shift_srl_145Z0Z_12));
    InMux I__8597 (
            .O(N__61861),
            .I(N__61858));
    LocalMux I__8596 (
            .O(N__61858),
            .I(shift_srl_145Z0Z_13));
    InMux I__8595 (
            .O(N__61855),
            .I(N__61852));
    LocalMux I__8594 (
            .O(N__61852),
            .I(shift_srl_145Z0Z_14));
    InMux I__8593 (
            .O(N__61849),
            .I(N__61846));
    LocalMux I__8592 (
            .O(N__61846),
            .I(shift_srl_145Z0Z_9));
    InMux I__8591 (
            .O(N__61843),
            .I(N__61840));
    LocalMux I__8590 (
            .O(N__61840),
            .I(shift_srl_145Z0Z_8));
    CascadeMux I__8589 (
            .O(N__61837),
            .I(rco_int_0_a3_0_a2_138_m6_0_a2_7_4_cascade_));
    InMux I__8588 (
            .O(N__61834),
            .I(N__61831));
    LocalMux I__8587 (
            .O(N__61831),
            .I(shift_srl_141Z0Z_3));
    InMux I__8586 (
            .O(N__61828),
            .I(N__61825));
    LocalMux I__8585 (
            .O(N__61825),
            .I(shift_srl_141Z0Z_13));
    InMux I__8584 (
            .O(N__61822),
            .I(N__61816));
    InMux I__8583 (
            .O(N__61821),
            .I(N__61811));
    InMux I__8582 (
            .O(N__61820),
            .I(N__61811));
    InMux I__8581 (
            .O(N__61819),
            .I(N__61808));
    LocalMux I__8580 (
            .O(N__61816),
            .I(N__61805));
    LocalMux I__8579 (
            .O(N__61811),
            .I(N__61802));
    LocalMux I__8578 (
            .O(N__61808),
            .I(shift_srl_144Z0Z_15));
    Odrv4 I__8577 (
            .O(N__61805),
            .I(shift_srl_144Z0Z_15));
    Odrv12 I__8576 (
            .O(N__61802),
            .I(shift_srl_144Z0Z_15));
    CascadeMux I__8575 (
            .O(N__61795),
            .I(rco_int_0_a2_0_a2_0_sx_144_cascade_));
    CascadeMux I__8574 (
            .O(N__61792),
            .I(N__61789));
    InMux I__8573 (
            .O(N__61789),
            .I(N__61782));
    InMux I__8572 (
            .O(N__61788),
            .I(N__61782));
    CascadeMux I__8571 (
            .O(N__61787),
            .I(N__61778));
    LocalMux I__8570 (
            .O(N__61782),
            .I(N__61773));
    InMux I__8569 (
            .O(N__61781),
            .I(N__61770));
    InMux I__8568 (
            .O(N__61778),
            .I(N__61765));
    InMux I__8567 (
            .O(N__61777),
            .I(N__61765));
    InMux I__8566 (
            .O(N__61776),
            .I(N__61762));
    Span4Mux_h I__8565 (
            .O(N__61773),
            .I(N__61759));
    LocalMux I__8564 (
            .O(N__61770),
            .I(N__61756));
    LocalMux I__8563 (
            .O(N__61765),
            .I(N__61751));
    LocalMux I__8562 (
            .O(N__61762),
            .I(N__61751));
    Span4Mux_h I__8561 (
            .O(N__61759),
            .I(N__61748));
    Odrv4 I__8560 (
            .O(N__61756),
            .I(shift_srl_143Z0Z_15));
    Odrv4 I__8559 (
            .O(N__61751),
            .I(shift_srl_143Z0Z_15));
    Odrv4 I__8558 (
            .O(N__61748),
            .I(shift_srl_143Z0Z_15));
    InMux I__8557 (
            .O(N__61741),
            .I(N__61738));
    LocalMux I__8556 (
            .O(N__61738),
            .I(shift_srl_141Z0Z_14));
    CascadeMux I__8555 (
            .O(N__61735),
            .I(N__61732));
    InMux I__8554 (
            .O(N__61732),
            .I(N__61727));
    InMux I__8553 (
            .O(N__61731),
            .I(N__61722));
    InMux I__8552 (
            .O(N__61730),
            .I(N__61722));
    LocalMux I__8551 (
            .O(N__61727),
            .I(shift_srl_141Z0Z_15));
    LocalMux I__8550 (
            .O(N__61722),
            .I(shift_srl_141Z0Z_15));
    InMux I__8549 (
            .O(N__61717),
            .I(N__61714));
    LocalMux I__8548 (
            .O(N__61714),
            .I(shift_srl_141Z0Z_0));
    InMux I__8547 (
            .O(N__61711),
            .I(N__61708));
    LocalMux I__8546 (
            .O(N__61708),
            .I(shift_srl_141Z0Z_1));
    InMux I__8545 (
            .O(N__61705),
            .I(N__61702));
    LocalMux I__8544 (
            .O(N__61702),
            .I(shift_srl_141Z0Z_2));
    InMux I__8543 (
            .O(N__61699),
            .I(N__61696));
    LocalMux I__8542 (
            .O(N__61696),
            .I(shift_srl_141Z0Z_10));
    InMux I__8541 (
            .O(N__61693),
            .I(N__61690));
    LocalMux I__8540 (
            .O(N__61690),
            .I(shift_srl_141Z0Z_11));
    InMux I__8539 (
            .O(N__61687),
            .I(N__61684));
    LocalMux I__8538 (
            .O(N__61684),
            .I(shift_srl_141Z0Z_12));
    InMux I__8537 (
            .O(N__61681),
            .I(N__61678));
    LocalMux I__8536 (
            .O(N__61678),
            .I(shift_srl_141Z0Z_9));
    InMux I__8535 (
            .O(N__61675),
            .I(N__61672));
    LocalMux I__8534 (
            .O(N__61672),
            .I(shift_srl_141Z0Z_7));
    InMux I__8533 (
            .O(N__61669),
            .I(N__61666));
    LocalMux I__8532 (
            .O(N__61666),
            .I(shift_srl_141Z0Z_8));
    InMux I__8531 (
            .O(N__61663),
            .I(N__61660));
    LocalMux I__8530 (
            .O(N__61660),
            .I(shift_srl_141Z0Z_4));
    InMux I__8529 (
            .O(N__61657),
            .I(N__61654));
    LocalMux I__8528 (
            .O(N__61654),
            .I(shift_srl_141Z0Z_5));
    InMux I__8527 (
            .O(N__61651),
            .I(N__61648));
    LocalMux I__8526 (
            .O(N__61648),
            .I(shift_srl_141Z0Z_6));
    InMux I__8525 (
            .O(N__61645),
            .I(N__61642));
    LocalMux I__8524 (
            .O(N__61642),
            .I(N__61638));
    InMux I__8523 (
            .O(N__61641),
            .I(N__61635));
    Span4Mux_h I__8522 (
            .O(N__61638),
            .I(N__61632));
    LocalMux I__8521 (
            .O(N__61635),
            .I(shift_srl_153Z0Z_15));
    Odrv4 I__8520 (
            .O(N__61632),
            .I(shift_srl_153Z0Z_15));
    InMux I__8519 (
            .O(N__61627),
            .I(N__61624));
    LocalMux I__8518 (
            .O(N__61624),
            .I(shift_srl_153Z0Z_0));
    InMux I__8517 (
            .O(N__61621),
            .I(N__61618));
    LocalMux I__8516 (
            .O(N__61618),
            .I(shift_srl_153Z0Z_1));
    InMux I__8515 (
            .O(N__61615),
            .I(N__61612));
    LocalMux I__8514 (
            .O(N__61612),
            .I(shift_srl_153Z0Z_2));
    InMux I__8513 (
            .O(N__61609),
            .I(N__61606));
    LocalMux I__8512 (
            .O(N__61606),
            .I(shift_srl_153Z0Z_3));
    InMux I__8511 (
            .O(N__61603),
            .I(N__61600));
    LocalMux I__8510 (
            .O(N__61600),
            .I(shift_srl_153Z0Z_4));
    InMux I__8509 (
            .O(N__61597),
            .I(N__61594));
    LocalMux I__8508 (
            .O(N__61594),
            .I(shift_srl_153Z0Z_5));
    InMux I__8507 (
            .O(N__61591),
            .I(N__61588));
    LocalMux I__8506 (
            .O(N__61588),
            .I(shift_srl_153Z0Z_6));
    InMux I__8505 (
            .O(N__61585),
            .I(N__61582));
    LocalMux I__8504 (
            .O(N__61582),
            .I(shift_srl_153Z0Z_7));
    InMux I__8503 (
            .O(N__61579),
            .I(N__61576));
    LocalMux I__8502 (
            .O(N__61576),
            .I(shift_srl_152Z0Z_8));
    InMux I__8501 (
            .O(N__61573),
            .I(N__61570));
    LocalMux I__8500 (
            .O(N__61570),
            .I(shift_srl_153Z0Z_10));
    InMux I__8499 (
            .O(N__61567),
            .I(N__61564));
    LocalMux I__8498 (
            .O(N__61564),
            .I(shift_srl_153Z0Z_11));
    InMux I__8497 (
            .O(N__61561),
            .I(N__61558));
    LocalMux I__8496 (
            .O(N__61558),
            .I(shift_srl_153Z0Z_12));
    InMux I__8495 (
            .O(N__61555),
            .I(N__61552));
    LocalMux I__8494 (
            .O(N__61552),
            .I(shift_srl_153Z0Z_13));
    InMux I__8493 (
            .O(N__61549),
            .I(N__61546));
    LocalMux I__8492 (
            .O(N__61546),
            .I(shift_srl_153Z0Z_14));
    InMux I__8491 (
            .O(N__61543),
            .I(N__61540));
    LocalMux I__8490 (
            .O(N__61540),
            .I(shift_srl_153Z0Z_9));
    InMux I__8489 (
            .O(N__61537),
            .I(N__61534));
    LocalMux I__8488 (
            .O(N__61534),
            .I(shift_srl_153Z0Z_8));
    InMux I__8487 (
            .O(N__61531),
            .I(N__61528));
    LocalMux I__8486 (
            .O(N__61528),
            .I(shift_srl_24Z0Z_3));
    InMux I__8485 (
            .O(N__61525),
            .I(N__61522));
    LocalMux I__8484 (
            .O(N__61522),
            .I(shift_srl_24Z0Z_4));
    InMux I__8483 (
            .O(N__61519),
            .I(N__61516));
    LocalMux I__8482 (
            .O(N__61516),
            .I(shift_srl_24Z0Z_7));
    InMux I__8481 (
            .O(N__61513),
            .I(N__61510));
    LocalMux I__8480 (
            .O(N__61510),
            .I(shift_srl_24Z0Z_5));
    InMux I__8479 (
            .O(N__61507),
            .I(N__61504));
    LocalMux I__8478 (
            .O(N__61504),
            .I(shift_srl_24Z0Z_6));
    InMux I__8477 (
            .O(N__61501),
            .I(N__61498));
    LocalMux I__8476 (
            .O(N__61498),
            .I(shift_srl_152Z0Z_10));
    InMux I__8475 (
            .O(N__61495),
            .I(N__61492));
    LocalMux I__8474 (
            .O(N__61492),
            .I(shift_srl_152Z0Z_11));
    InMux I__8473 (
            .O(N__61489),
            .I(N__61486));
    LocalMux I__8472 (
            .O(N__61486),
            .I(shift_srl_152Z0Z_12));
    InMux I__8471 (
            .O(N__61483),
            .I(N__61480));
    LocalMux I__8470 (
            .O(N__61480),
            .I(shift_srl_152Z0Z_13));
    InMux I__8469 (
            .O(N__61477),
            .I(N__61474));
    LocalMux I__8468 (
            .O(N__61474),
            .I(shift_srl_152Z0Z_14));
    InMux I__8467 (
            .O(N__61471),
            .I(N__61468));
    LocalMux I__8466 (
            .O(N__61468),
            .I(shift_srl_152Z0Z_9));
    CascadeMux I__8465 (
            .O(N__61465),
            .I(rco_int_0_a2_0_a2_0_sx_91_cascade_));
    CascadeMux I__8464 (
            .O(N__61462),
            .I(shift_srl_91_RNI20EN1Z0Z_15_cascade_));
    CascadeMux I__8463 (
            .O(N__61459),
            .I(shift_srl_83_RNIKTI68Z0Z_15_cascade_));
    CEMux I__8462 (
            .O(N__61456),
            .I(N__61452));
    CEMux I__8461 (
            .O(N__61455),
            .I(N__61449));
    LocalMux I__8460 (
            .O(N__61452),
            .I(N__61446));
    LocalMux I__8459 (
            .O(N__61449),
            .I(N__61443));
    Odrv4 I__8458 (
            .O(N__61446),
            .I(clk_en_84));
    Odrv12 I__8457 (
            .O(N__61443),
            .I(clk_en_84));
    CascadeMux I__8456 (
            .O(N__61438),
            .I(clk_en_84_cascade_));
    InMux I__8455 (
            .O(N__61435),
            .I(N__61432));
    LocalMux I__8454 (
            .O(N__61432),
            .I(shift_srl_89Z0Z_14));
    CEMux I__8453 (
            .O(N__61429),
            .I(N__61425));
    CEMux I__8452 (
            .O(N__61428),
            .I(N__61421));
    LocalMux I__8451 (
            .O(N__61425),
            .I(N__61418));
    CEMux I__8450 (
            .O(N__61424),
            .I(N__61415));
    LocalMux I__8449 (
            .O(N__61421),
            .I(N__61412));
    Span4Mux_h I__8448 (
            .O(N__61418),
            .I(N__61407));
    LocalMux I__8447 (
            .O(N__61415),
            .I(N__61407));
    Odrv4 I__8446 (
            .O(N__61412),
            .I(clk_en_89));
    Odrv4 I__8445 (
            .O(N__61407),
            .I(clk_en_89));
    InMux I__8444 (
            .O(N__61402),
            .I(N__61399));
    LocalMux I__8443 (
            .O(N__61399),
            .I(shift_srl_84Z0Z_10));
    InMux I__8442 (
            .O(N__61396),
            .I(N__61393));
    LocalMux I__8441 (
            .O(N__61393),
            .I(shift_srl_84Z0Z_11));
    InMux I__8440 (
            .O(N__61390),
            .I(N__61387));
    LocalMux I__8439 (
            .O(N__61387),
            .I(shift_srl_84Z0Z_12));
    InMux I__8438 (
            .O(N__61384),
            .I(N__61381));
    LocalMux I__8437 (
            .O(N__61381),
            .I(shift_srl_84Z0Z_13));
    InMux I__8436 (
            .O(N__61378),
            .I(N__61375));
    LocalMux I__8435 (
            .O(N__61375),
            .I(shift_srl_84Z0Z_14));
    InMux I__8434 (
            .O(N__61372),
            .I(N__61369));
    LocalMux I__8433 (
            .O(N__61369),
            .I(shift_srl_84Z0Z_9));
    InMux I__8432 (
            .O(N__61366),
            .I(N__61363));
    LocalMux I__8431 (
            .O(N__61363),
            .I(shift_srl_84Z0Z_7));
    InMux I__8430 (
            .O(N__61360),
            .I(N__61357));
    LocalMux I__8429 (
            .O(N__61357),
            .I(shift_srl_84Z0Z_8));
    InMux I__8428 (
            .O(N__61354),
            .I(N__61351));
    LocalMux I__8427 (
            .O(N__61351),
            .I(shift_srl_86Z0Z_11));
    InMux I__8426 (
            .O(N__61348),
            .I(N__61345));
    LocalMux I__8425 (
            .O(N__61345),
            .I(shift_srl_84Z0Z_0));
    InMux I__8424 (
            .O(N__61342),
            .I(N__61339));
    LocalMux I__8423 (
            .O(N__61339),
            .I(shift_srl_84Z0Z_1));
    InMux I__8422 (
            .O(N__61336),
            .I(N__61333));
    LocalMux I__8421 (
            .O(N__61333),
            .I(shift_srl_84Z0Z_2));
    InMux I__8420 (
            .O(N__61330),
            .I(N__61327));
    LocalMux I__8419 (
            .O(N__61327),
            .I(shift_srl_84Z0Z_3));
    InMux I__8418 (
            .O(N__61324),
            .I(N__61321));
    LocalMux I__8417 (
            .O(N__61321),
            .I(shift_srl_84Z0Z_4));
    InMux I__8416 (
            .O(N__61318),
            .I(N__61315));
    LocalMux I__8415 (
            .O(N__61315),
            .I(shift_srl_84Z0Z_5));
    InMux I__8414 (
            .O(N__61312),
            .I(N__61309));
    LocalMux I__8413 (
            .O(N__61309),
            .I(shift_srl_84Z0Z_6));
    InMux I__8412 (
            .O(N__61306),
            .I(N__61303));
    LocalMux I__8411 (
            .O(N__61303),
            .I(shift_srl_87Z0Z_14));
    InMux I__8410 (
            .O(N__61300),
            .I(N__61297));
    LocalMux I__8409 (
            .O(N__61297),
            .I(shift_srl_87Z0Z_9));
    InMux I__8408 (
            .O(N__61294),
            .I(N__61291));
    LocalMux I__8407 (
            .O(N__61291),
            .I(shift_srl_87Z0Z_8));
    InMux I__8406 (
            .O(N__61288),
            .I(N__61285));
    LocalMux I__8405 (
            .O(N__61285),
            .I(shift_srl_86Z0Z_0));
    InMux I__8404 (
            .O(N__61282),
            .I(N__61279));
    LocalMux I__8403 (
            .O(N__61279),
            .I(shift_srl_86Z0Z_1));
    InMux I__8402 (
            .O(N__61276),
            .I(N__61273));
    LocalMux I__8401 (
            .O(N__61273),
            .I(shift_srl_86Z0Z_2));
    InMux I__8400 (
            .O(N__61270),
            .I(N__61267));
    LocalMux I__8399 (
            .O(N__61267),
            .I(shift_srl_86Z0Z_3));
    InMux I__8398 (
            .O(N__61264),
            .I(N__61261));
    LocalMux I__8397 (
            .O(N__61261),
            .I(shift_srl_86Z0Z_4));
    InMux I__8396 (
            .O(N__61258),
            .I(N__61255));
    LocalMux I__8395 (
            .O(N__61255),
            .I(shift_srl_90Z0Z_14));
    InMux I__8394 (
            .O(N__61252),
            .I(N__61249));
    LocalMux I__8393 (
            .O(N__61249),
            .I(shift_srl_90Z0Z_13));
    InMux I__8392 (
            .O(N__61246),
            .I(N__61243));
    LocalMux I__8391 (
            .O(N__61243),
            .I(shift_srl_90Z0Z_12));
    InMux I__8390 (
            .O(N__61240),
            .I(N__61237));
    LocalMux I__8389 (
            .O(N__61237),
            .I(shift_srl_90Z0Z_10));
    InMux I__8388 (
            .O(N__61234),
            .I(N__61231));
    LocalMux I__8387 (
            .O(N__61231),
            .I(shift_srl_90Z0Z_11));
    CEMux I__8386 (
            .O(N__61228),
            .I(N__61223));
    CEMux I__8385 (
            .O(N__61227),
            .I(N__61220));
    CEMux I__8384 (
            .O(N__61226),
            .I(N__61217));
    LocalMux I__8383 (
            .O(N__61223),
            .I(clk_en_90));
    LocalMux I__8382 (
            .O(N__61220),
            .I(clk_en_90));
    LocalMux I__8381 (
            .O(N__61217),
            .I(clk_en_90));
    InMux I__8380 (
            .O(N__61210),
            .I(N__61207));
    LocalMux I__8379 (
            .O(N__61207),
            .I(shift_srl_87Z0Z_10));
    InMux I__8378 (
            .O(N__61204),
            .I(N__61201));
    LocalMux I__8377 (
            .O(N__61201),
            .I(shift_srl_87Z0Z_11));
    InMux I__8376 (
            .O(N__61198),
            .I(N__61195));
    LocalMux I__8375 (
            .O(N__61195),
            .I(shift_srl_87Z0Z_12));
    InMux I__8374 (
            .O(N__61192),
            .I(N__61189));
    LocalMux I__8373 (
            .O(N__61189),
            .I(shift_srl_87Z0Z_13));
    InMux I__8372 (
            .O(N__61186),
            .I(N__61183));
    LocalMux I__8371 (
            .O(N__61183),
            .I(shift_srl_90Z0Z_0));
    InMux I__8370 (
            .O(N__61180),
            .I(N__61177));
    LocalMux I__8369 (
            .O(N__61177),
            .I(shift_srl_90Z0Z_1));
    InMux I__8368 (
            .O(N__61174),
            .I(N__61171));
    LocalMux I__8367 (
            .O(N__61171),
            .I(shift_srl_90Z0Z_2));
    InMux I__8366 (
            .O(N__61168),
            .I(N__61165));
    LocalMux I__8365 (
            .O(N__61165),
            .I(shift_srl_90Z0Z_3));
    InMux I__8364 (
            .O(N__61162),
            .I(N__61159));
    LocalMux I__8363 (
            .O(N__61159),
            .I(shift_srl_90Z0Z_4));
    InMux I__8362 (
            .O(N__61156),
            .I(N__61153));
    LocalMux I__8361 (
            .O(N__61153),
            .I(shift_srl_90Z0Z_5));
    CEMux I__8360 (
            .O(N__61150),
            .I(N__61147));
    LocalMux I__8359 (
            .O(N__61147),
            .I(N__61143));
    CEMux I__8358 (
            .O(N__61146),
            .I(N__61140));
    Span4Mux_v I__8357 (
            .O(N__61143),
            .I(N__61137));
    LocalMux I__8356 (
            .O(N__61140),
            .I(N__61134));
    Span4Mux_h I__8355 (
            .O(N__61137),
            .I(N__61129));
    Span4Mux_v I__8354 (
            .O(N__61134),
            .I(N__61129));
    Odrv4 I__8353 (
            .O(N__61129),
            .I(clk_en_91));
    InMux I__8352 (
            .O(N__61126),
            .I(N__61123));
    LocalMux I__8351 (
            .O(N__61123),
            .I(shift_srl_103Z0Z_10));
    InMux I__8350 (
            .O(N__61120),
            .I(N__61117));
    LocalMux I__8349 (
            .O(N__61117),
            .I(shift_srl_103Z0Z_11));
    InMux I__8348 (
            .O(N__61114),
            .I(N__61111));
    LocalMux I__8347 (
            .O(N__61111),
            .I(shift_srl_103Z0Z_12));
    InMux I__8346 (
            .O(N__61108),
            .I(N__61105));
    LocalMux I__8345 (
            .O(N__61105),
            .I(shift_srl_103Z0Z_13));
    InMux I__8344 (
            .O(N__61102),
            .I(N__61099));
    LocalMux I__8343 (
            .O(N__61099),
            .I(shift_srl_103Z0Z_14));
    CascadeMux I__8342 (
            .O(N__61096),
            .I(N__61090));
    InMux I__8341 (
            .O(N__61095),
            .I(N__61084));
    InMux I__8340 (
            .O(N__61094),
            .I(N__61084));
    InMux I__8339 (
            .O(N__61093),
            .I(N__61081));
    InMux I__8338 (
            .O(N__61090),
            .I(N__61076));
    InMux I__8337 (
            .O(N__61089),
            .I(N__61076));
    LocalMux I__8336 (
            .O(N__61084),
            .I(shift_srl_103Z0Z_15));
    LocalMux I__8335 (
            .O(N__61081),
            .I(shift_srl_103Z0Z_15));
    LocalMux I__8334 (
            .O(N__61076),
            .I(shift_srl_103Z0Z_15));
    InMux I__8333 (
            .O(N__61069),
            .I(N__61066));
    LocalMux I__8332 (
            .O(N__61066),
            .I(shift_srl_103Z0Z_9));
    InMux I__8331 (
            .O(N__61063),
            .I(N__61060));
    LocalMux I__8330 (
            .O(N__61060),
            .I(N__61057));
    Odrv4 I__8329 (
            .O(N__61057),
            .I(shift_srl_103Z0Z_7));
    InMux I__8328 (
            .O(N__61054),
            .I(N__61051));
    LocalMux I__8327 (
            .O(N__61051),
            .I(shift_srl_103Z0Z_8));
    CEMux I__8326 (
            .O(N__61048),
            .I(N__61043));
    CEMux I__8325 (
            .O(N__61047),
            .I(N__61040));
    CEMux I__8324 (
            .O(N__61046),
            .I(N__61037));
    LocalMux I__8323 (
            .O(N__61043),
            .I(N__61034));
    LocalMux I__8322 (
            .O(N__61040),
            .I(N__61029));
    LocalMux I__8321 (
            .O(N__61037),
            .I(N__61029));
    Odrv4 I__8320 (
            .O(N__61034),
            .I(clk_en_103));
    Odrv4 I__8319 (
            .O(N__61029),
            .I(clk_en_103));
    IoInMux I__8318 (
            .O(N__61024),
            .I(N__61021));
    LocalMux I__8317 (
            .O(N__61021),
            .I(N__61018));
    Span4Mux_s2_v I__8316 (
            .O(N__61018),
            .I(N__61015));
    Odrv4 I__8315 (
            .O(N__61015),
            .I(rco_c_87));
    IoInMux I__8314 (
            .O(N__61012),
            .I(N__61009));
    LocalMux I__8313 (
            .O(N__61009),
            .I(N__61006));
    Span12Mux_s3_v I__8312 (
            .O(N__61006),
            .I(N__61003));
    Odrv12 I__8311 (
            .O(N__61003),
            .I(rco_c_86));
    InMux I__8310 (
            .O(N__61000),
            .I(N__60995));
    InMux I__8309 (
            .O(N__60999),
            .I(N__60990));
    InMux I__8308 (
            .O(N__60998),
            .I(N__60990));
    LocalMux I__8307 (
            .O(N__60995),
            .I(shift_srl_104Z0Z_15));
    LocalMux I__8306 (
            .O(N__60990),
            .I(shift_srl_104Z0Z_15));
    InMux I__8305 (
            .O(N__60985),
            .I(N__60978));
    InMux I__8304 (
            .O(N__60984),
            .I(N__60978));
    CascadeMux I__8303 (
            .O(N__60983),
            .I(N__60975));
    LocalMux I__8302 (
            .O(N__60978),
            .I(N__60970));
    InMux I__8301 (
            .O(N__60975),
            .I(N__60967));
    InMux I__8300 (
            .O(N__60974),
            .I(N__60962));
    InMux I__8299 (
            .O(N__60973),
            .I(N__60962));
    Span4Mux_v I__8298 (
            .O(N__60970),
            .I(N__60952));
    LocalMux I__8297 (
            .O(N__60967),
            .I(N__60952));
    LocalMux I__8296 (
            .O(N__60962),
            .I(N__60952));
    InMux I__8295 (
            .O(N__60961),
            .I(N__60945));
    InMux I__8294 (
            .O(N__60960),
            .I(N__60945));
    InMux I__8293 (
            .O(N__60959),
            .I(N__60945));
    Odrv4 I__8292 (
            .O(N__60952),
            .I(shift_srl_101Z0Z_15));
    LocalMux I__8291 (
            .O(N__60945),
            .I(shift_srl_101Z0Z_15));
    InMux I__8290 (
            .O(N__60940),
            .I(N__60937));
    LocalMux I__8289 (
            .O(N__60937),
            .I(N__60934));
    Span4Mux_h I__8288 (
            .O(N__60934),
            .I(N__60931));
    Odrv4 I__8287 (
            .O(N__60931),
            .I(rco_int_0_a3_0_a2_s_0_sx_104));
    InMux I__8286 (
            .O(N__60928),
            .I(N__60925));
    LocalMux I__8285 (
            .O(N__60925),
            .I(shift_srl_100Z0Z_14));
    InMux I__8284 (
            .O(N__60922),
            .I(N__60919));
    LocalMux I__8283 (
            .O(N__60919),
            .I(shift_srl_100Z0Z_13));
    InMux I__8282 (
            .O(N__60916),
            .I(N__60913));
    LocalMux I__8281 (
            .O(N__60913),
            .I(shift_srl_100Z0Z_12));
    InMux I__8280 (
            .O(N__60910),
            .I(N__60907));
    LocalMux I__8279 (
            .O(N__60907),
            .I(N__60904));
    Odrv4 I__8278 (
            .O(N__60904),
            .I(shift_srl_100Z0Z_10));
    InMux I__8277 (
            .O(N__60901),
            .I(N__60898));
    LocalMux I__8276 (
            .O(N__60898),
            .I(shift_srl_100Z0Z_11));
    CEMux I__8275 (
            .O(N__60895),
            .I(N__60892));
    LocalMux I__8274 (
            .O(N__60892),
            .I(N__60887));
    CEMux I__8273 (
            .O(N__60891),
            .I(N__60884));
    CEMux I__8272 (
            .O(N__60890),
            .I(N__60881));
    Span4Mux_v I__8271 (
            .O(N__60887),
            .I(N__60874));
    LocalMux I__8270 (
            .O(N__60884),
            .I(N__60874));
    LocalMux I__8269 (
            .O(N__60881),
            .I(N__60874));
    Span4Mux_v I__8268 (
            .O(N__60874),
            .I(N__60871));
    Odrv4 I__8267 (
            .O(N__60871),
            .I(clk_en_100));
    InMux I__8266 (
            .O(N__60868),
            .I(N__60865));
    LocalMux I__8265 (
            .O(N__60865),
            .I(shift_srl_199Z0Z_5));
    InMux I__8264 (
            .O(N__60862),
            .I(N__60859));
    LocalMux I__8263 (
            .O(N__60859),
            .I(N__60856));
    Span4Mux_h I__8262 (
            .O(N__60856),
            .I(N__60853));
    Span4Mux_h I__8261 (
            .O(N__60853),
            .I(N__60850));
    Odrv4 I__8260 (
            .O(N__60850),
            .I(shift_srl_199Z0Z_6));
    InMux I__8259 (
            .O(N__60847),
            .I(N__60844));
    LocalMux I__8258 (
            .O(N__60844),
            .I(shift_srl_102Z0Z_10));
    InMux I__8257 (
            .O(N__60841),
            .I(N__60838));
    LocalMux I__8256 (
            .O(N__60838),
            .I(shift_srl_102Z0Z_11));
    InMux I__8255 (
            .O(N__60835),
            .I(N__60832));
    LocalMux I__8254 (
            .O(N__60832),
            .I(shift_srl_102Z0Z_12));
    InMux I__8253 (
            .O(N__60829),
            .I(N__60826));
    LocalMux I__8252 (
            .O(N__60826),
            .I(shift_srl_102Z0Z_13));
    InMux I__8251 (
            .O(N__60823),
            .I(N__60820));
    LocalMux I__8250 (
            .O(N__60820),
            .I(shift_srl_102Z0Z_14));
    InMux I__8249 (
            .O(N__60817),
            .I(N__60814));
    LocalMux I__8248 (
            .O(N__60814),
            .I(shift_srl_102Z0Z_7));
    CEMux I__8247 (
            .O(N__60811),
            .I(N__60807));
    CEMux I__8246 (
            .O(N__60810),
            .I(N__60804));
    LocalMux I__8245 (
            .O(N__60807),
            .I(N__60801));
    LocalMux I__8244 (
            .O(N__60804),
            .I(N__60797));
    Span4Mux_v I__8243 (
            .O(N__60801),
            .I(N__60794));
    CEMux I__8242 (
            .O(N__60800),
            .I(N__60791));
    Span4Mux_h I__8241 (
            .O(N__60797),
            .I(N__60788));
    Span4Mux_h I__8240 (
            .O(N__60794),
            .I(N__60783));
    LocalMux I__8239 (
            .O(N__60791),
            .I(N__60783));
    Odrv4 I__8238 (
            .O(N__60788),
            .I(clk_en_118));
    Odrv4 I__8237 (
            .O(N__60783),
            .I(clk_en_118));
    CascadeMux I__8236 (
            .O(N__60778),
            .I(N__60772));
    InMux I__8235 (
            .O(N__60777),
            .I(N__60769));
    CascadeMux I__8234 (
            .O(N__60776),
            .I(N__60766));
    CascadeMux I__8233 (
            .O(N__60775),
            .I(N__60762));
    InMux I__8232 (
            .O(N__60772),
            .I(N__60759));
    LocalMux I__8231 (
            .O(N__60769),
            .I(N__60756));
    InMux I__8230 (
            .O(N__60766),
            .I(N__60748));
    InMux I__8229 (
            .O(N__60765),
            .I(N__60748));
    InMux I__8228 (
            .O(N__60762),
            .I(N__60745));
    LocalMux I__8227 (
            .O(N__60759),
            .I(N__60742));
    Span4Mux_v I__8226 (
            .O(N__60756),
            .I(N__60739));
    CascadeMux I__8225 (
            .O(N__60755),
            .I(N__60736));
    CascadeMux I__8224 (
            .O(N__60754),
            .I(N__60733));
    CascadeMux I__8223 (
            .O(N__60753),
            .I(N__60727));
    LocalMux I__8222 (
            .O(N__60748),
            .I(N__60724));
    LocalMux I__8221 (
            .O(N__60745),
            .I(N__60719));
    Span4Mux_v I__8220 (
            .O(N__60742),
            .I(N__60719));
    Span4Mux_h I__8219 (
            .O(N__60739),
            .I(N__60716));
    InMux I__8218 (
            .O(N__60736),
            .I(N__60709));
    InMux I__8217 (
            .O(N__60733),
            .I(N__60709));
    InMux I__8216 (
            .O(N__60732),
            .I(N__60709));
    CascadeMux I__8215 (
            .O(N__60731),
            .I(N__60706));
    InMux I__8214 (
            .O(N__60730),
            .I(N__60702));
    InMux I__8213 (
            .O(N__60727),
            .I(N__60699));
    Span4Mux_h I__8212 (
            .O(N__60724),
            .I(N__60696));
    Span4Mux_h I__8211 (
            .O(N__60719),
            .I(N__60693));
    Sp12to4 I__8210 (
            .O(N__60716),
            .I(N__60688));
    LocalMux I__8209 (
            .O(N__60709),
            .I(N__60688));
    InMux I__8208 (
            .O(N__60706),
            .I(N__60683));
    InMux I__8207 (
            .O(N__60705),
            .I(N__60683));
    LocalMux I__8206 (
            .O(N__60702),
            .I(shift_srl_111Z0Z_15));
    LocalMux I__8205 (
            .O(N__60699),
            .I(shift_srl_111Z0Z_15));
    Odrv4 I__8204 (
            .O(N__60696),
            .I(shift_srl_111Z0Z_15));
    Odrv4 I__8203 (
            .O(N__60693),
            .I(shift_srl_111Z0Z_15));
    Odrv12 I__8202 (
            .O(N__60688),
            .I(shift_srl_111Z0Z_15));
    LocalMux I__8201 (
            .O(N__60683),
            .I(shift_srl_111Z0Z_15));
    IoInMux I__8200 (
            .O(N__60670),
            .I(N__60667));
    LocalMux I__8199 (
            .O(N__60667),
            .I(N__60664));
    Span4Mux_s2_v I__8198 (
            .O(N__60664),
            .I(N__60661));
    Sp12to4 I__8197 (
            .O(N__60661),
            .I(N__60658));
    Span12Mux_h I__8196 (
            .O(N__60658),
            .I(N__60655));
    Odrv12 I__8195 (
            .O(N__60655),
            .I(rco_c_111));
    InMux I__8194 (
            .O(N__60652),
            .I(N__60644));
    InMux I__8193 (
            .O(N__60651),
            .I(N__60644));
    InMux I__8192 (
            .O(N__60650),
            .I(N__60641));
    InMux I__8191 (
            .O(N__60649),
            .I(N__60638));
    LocalMux I__8190 (
            .O(N__60644),
            .I(N__60635));
    LocalMux I__8189 (
            .O(N__60641),
            .I(N__60632));
    LocalMux I__8188 (
            .O(N__60638),
            .I(N__60627));
    Span4Mux_h I__8187 (
            .O(N__60635),
            .I(N__60627));
    Span12Mux_h I__8186 (
            .O(N__60632),
            .I(N__60624));
    Span4Mux_v I__8185 (
            .O(N__60627),
            .I(N__60621));
    Odrv12 I__8184 (
            .O(N__60624),
            .I(rco_int_0_a2_1_a2_1_120));
    Odrv4 I__8183 (
            .O(N__60621),
            .I(rco_int_0_a2_1_a2_1_120));
    IoInMux I__8182 (
            .O(N__60616),
            .I(N__60613));
    LocalMux I__8181 (
            .O(N__60613),
            .I(N__60610));
    Span4Mux_s3_v I__8180 (
            .O(N__60610),
            .I(N__60607));
    Span4Mux_h I__8179 (
            .O(N__60607),
            .I(N__60604));
    Span4Mux_h I__8178 (
            .O(N__60604),
            .I(N__60601));
    Span4Mux_v I__8177 (
            .O(N__60601),
            .I(N__60598));
    Odrv4 I__8176 (
            .O(N__60598),
            .I(rco_c_199));
    InMux I__8175 (
            .O(N__60595),
            .I(N__60592));
    LocalMux I__8174 (
            .O(N__60592),
            .I(shift_srl_199Z0Z_0));
    InMux I__8173 (
            .O(N__60589),
            .I(N__60586));
    LocalMux I__8172 (
            .O(N__60586),
            .I(shift_srl_199Z0Z_1));
    InMux I__8171 (
            .O(N__60583),
            .I(N__60580));
    LocalMux I__8170 (
            .O(N__60580),
            .I(shift_srl_199Z0Z_2));
    InMux I__8169 (
            .O(N__60577),
            .I(N__60574));
    LocalMux I__8168 (
            .O(N__60574),
            .I(shift_srl_199Z0Z_3));
    InMux I__8167 (
            .O(N__60571),
            .I(N__60568));
    LocalMux I__8166 (
            .O(N__60568),
            .I(shift_srl_199Z0Z_4));
    InMux I__8165 (
            .O(N__60565),
            .I(N__60562));
    LocalMux I__8164 (
            .O(N__60562),
            .I(shift_srl_111Z0Z_2));
    InMux I__8163 (
            .O(N__60559),
            .I(N__60556));
    LocalMux I__8162 (
            .O(N__60556),
            .I(shift_srl_111Z0Z_3));
    InMux I__8161 (
            .O(N__60553),
            .I(N__60550));
    LocalMux I__8160 (
            .O(N__60550),
            .I(shift_srl_111Z0Z_4));
    InMux I__8159 (
            .O(N__60547),
            .I(N__60544));
    LocalMux I__8158 (
            .O(N__60544),
            .I(shift_srl_111Z0Z_5));
    InMux I__8157 (
            .O(N__60541),
            .I(N__60538));
    LocalMux I__8156 (
            .O(N__60538),
            .I(shift_srl_111Z0Z_6));
    CascadeMux I__8155 (
            .O(N__60535),
            .I(N__60531));
    InMux I__8154 (
            .O(N__60534),
            .I(N__60525));
    InMux I__8153 (
            .O(N__60531),
            .I(N__60522));
    InMux I__8152 (
            .O(N__60530),
            .I(N__60519));
    InMux I__8151 (
            .O(N__60529),
            .I(N__60516));
    InMux I__8150 (
            .O(N__60528),
            .I(N__60512));
    LocalMux I__8149 (
            .O(N__60525),
            .I(N__60509));
    LocalMux I__8148 (
            .O(N__60522),
            .I(N__60506));
    LocalMux I__8147 (
            .O(N__60519),
            .I(N__60501));
    LocalMux I__8146 (
            .O(N__60516),
            .I(N__60498));
    CascadeMux I__8145 (
            .O(N__60515),
            .I(N__60493));
    LocalMux I__8144 (
            .O(N__60512),
            .I(N__60488));
    Span4Mux_v I__8143 (
            .O(N__60509),
            .I(N__60488));
    Span4Mux_v I__8142 (
            .O(N__60506),
            .I(N__60485));
    InMux I__8141 (
            .O(N__60505),
            .I(N__60480));
    InMux I__8140 (
            .O(N__60504),
            .I(N__60480));
    Span4Mux_h I__8139 (
            .O(N__60501),
            .I(N__60477));
    Span4Mux_v I__8138 (
            .O(N__60498),
            .I(N__60474));
    InMux I__8137 (
            .O(N__60497),
            .I(N__60467));
    InMux I__8136 (
            .O(N__60496),
            .I(N__60467));
    InMux I__8135 (
            .O(N__60493),
            .I(N__60467));
    Sp12to4 I__8134 (
            .O(N__60488),
            .I(N__60460));
    Sp12to4 I__8133 (
            .O(N__60485),
            .I(N__60460));
    LocalMux I__8132 (
            .O(N__60480),
            .I(N__60460));
    Odrv4 I__8131 (
            .O(N__60477),
            .I(shift_srl_112Z0Z_15));
    Odrv4 I__8130 (
            .O(N__60474),
            .I(shift_srl_112Z0Z_15));
    LocalMux I__8129 (
            .O(N__60467),
            .I(shift_srl_112Z0Z_15));
    Odrv12 I__8128 (
            .O(N__60460),
            .I(shift_srl_112Z0Z_15));
    InMux I__8127 (
            .O(N__60451),
            .I(N__60445));
    InMux I__8126 (
            .O(N__60450),
            .I(N__60442));
    InMux I__8125 (
            .O(N__60449),
            .I(N__60439));
    InMux I__8124 (
            .O(N__60448),
            .I(N__60436));
    LocalMux I__8123 (
            .O(N__60445),
            .I(N__60433));
    LocalMux I__8122 (
            .O(N__60442),
            .I(N__60430));
    LocalMux I__8121 (
            .O(N__60439),
            .I(N__60427));
    LocalMux I__8120 (
            .O(N__60436),
            .I(N__60424));
    Span4Mux_v I__8119 (
            .O(N__60433),
            .I(N__60419));
    Span4Mux_v I__8118 (
            .O(N__60430),
            .I(N__60419));
    Span4Mux_v I__8117 (
            .O(N__60427),
            .I(N__60409));
    Span4Mux_v I__8116 (
            .O(N__60424),
            .I(N__60409));
    Span4Mux_h I__8115 (
            .O(N__60419),
            .I(N__60406));
    InMux I__8114 (
            .O(N__60418),
            .I(N__60397));
    InMux I__8113 (
            .O(N__60417),
            .I(N__60397));
    InMux I__8112 (
            .O(N__60416),
            .I(N__60397));
    InMux I__8111 (
            .O(N__60415),
            .I(N__60397));
    InMux I__8110 (
            .O(N__60414),
            .I(N__60394));
    Odrv4 I__8109 (
            .O(N__60409),
            .I(shift_srl_113Z0Z_15));
    Odrv4 I__8108 (
            .O(N__60406),
            .I(shift_srl_113Z0Z_15));
    LocalMux I__8107 (
            .O(N__60397),
            .I(shift_srl_113Z0Z_15));
    LocalMux I__8106 (
            .O(N__60394),
            .I(shift_srl_113Z0Z_15));
    CascadeMux I__8105 (
            .O(N__60385),
            .I(shift_srl_112_RNIV16I3Z0Z_15_cascade_));
    CEMux I__8104 (
            .O(N__60382),
            .I(N__60379));
    LocalMux I__8103 (
            .O(N__60379),
            .I(N__60376));
    Span4Mux_v I__8102 (
            .O(N__60376),
            .I(N__60372));
    CEMux I__8101 (
            .O(N__60375),
            .I(N__60369));
    Odrv4 I__8100 (
            .O(N__60372),
            .I(clk_en_114));
    LocalMux I__8099 (
            .O(N__60369),
            .I(clk_en_114));
    IoInMux I__8098 (
            .O(N__60364),
            .I(N__60361));
    LocalMux I__8097 (
            .O(N__60361),
            .I(N__60358));
    IoSpan4Mux I__8096 (
            .O(N__60358),
            .I(N__60355));
    Span4Mux_s0_h I__8095 (
            .O(N__60355),
            .I(N__60351));
    InMux I__8094 (
            .O(N__60354),
            .I(N__60348));
    Sp12to4 I__8093 (
            .O(N__60351),
            .I(N__60345));
    LocalMux I__8092 (
            .O(N__60348),
            .I(N__60342));
    Span12Mux_h I__8091 (
            .O(N__60345),
            .I(N__60337));
    Span12Mux_s10_v I__8090 (
            .O(N__60342),
            .I(N__60337));
    Odrv12 I__8089 (
            .O(N__60337),
            .I(N_91));
    CascadeMux I__8088 (
            .O(N__60334),
            .I(N__60329));
    CascadeMux I__8087 (
            .O(N__60333),
            .I(N__60324));
    InMux I__8086 (
            .O(N__60332),
            .I(N__60316));
    InMux I__8085 (
            .O(N__60329),
            .I(N__60311));
    InMux I__8084 (
            .O(N__60328),
            .I(N__60308));
    InMux I__8083 (
            .O(N__60327),
            .I(N__60303));
    InMux I__8082 (
            .O(N__60324),
            .I(N__60303));
    CascadeMux I__8081 (
            .O(N__60323),
            .I(N__60299));
    InMux I__8080 (
            .O(N__60322),
            .I(N__60295));
    InMux I__8079 (
            .O(N__60321),
            .I(N__60288));
    InMux I__8078 (
            .O(N__60320),
            .I(N__60288));
    InMux I__8077 (
            .O(N__60319),
            .I(N__60288));
    LocalMux I__8076 (
            .O(N__60316),
            .I(N__60285));
    InMux I__8075 (
            .O(N__60315),
            .I(N__60282));
    InMux I__8074 (
            .O(N__60314),
            .I(N__60279));
    LocalMux I__8073 (
            .O(N__60311),
            .I(N__60272));
    LocalMux I__8072 (
            .O(N__60308),
            .I(N__60272));
    LocalMux I__8071 (
            .O(N__60303),
            .I(N__60272));
    InMux I__8070 (
            .O(N__60302),
            .I(N__60269));
    InMux I__8069 (
            .O(N__60299),
            .I(N__60264));
    InMux I__8068 (
            .O(N__60298),
            .I(N__60264));
    LocalMux I__8067 (
            .O(N__60295),
            .I(N__60261));
    LocalMux I__8066 (
            .O(N__60288),
            .I(N__60258));
    Span4Mux_h I__8065 (
            .O(N__60285),
            .I(N__60255));
    LocalMux I__8064 (
            .O(N__60282),
            .I(N__60248));
    LocalMux I__8063 (
            .O(N__60279),
            .I(N__60248));
    Span4Mux_v I__8062 (
            .O(N__60272),
            .I(N__60248));
    LocalMux I__8061 (
            .O(N__60269),
            .I(shift_srl_118Z0Z_15));
    LocalMux I__8060 (
            .O(N__60264),
            .I(shift_srl_118Z0Z_15));
    Odrv4 I__8059 (
            .O(N__60261),
            .I(shift_srl_118Z0Z_15));
    Odrv4 I__8058 (
            .O(N__60258),
            .I(shift_srl_118Z0Z_15));
    Odrv4 I__8057 (
            .O(N__60255),
            .I(shift_srl_118Z0Z_15));
    Odrv4 I__8056 (
            .O(N__60248),
            .I(shift_srl_118Z0Z_15));
    InMux I__8055 (
            .O(N__60235),
            .I(N__60232));
    LocalMux I__8054 (
            .O(N__60232),
            .I(shift_srl_111Z0Z_14));
    InMux I__8053 (
            .O(N__60229),
            .I(N__60226));
    LocalMux I__8052 (
            .O(N__60226),
            .I(shift_srl_111Z0Z_13));
    InMux I__8051 (
            .O(N__60223),
            .I(N__60220));
    LocalMux I__8050 (
            .O(N__60220),
            .I(shift_srl_111Z0Z_0));
    InMux I__8049 (
            .O(N__60217),
            .I(N__60214));
    LocalMux I__8048 (
            .O(N__60214),
            .I(shift_srl_111Z0Z_1));
    InMux I__8047 (
            .O(N__60211),
            .I(N__60208));
    LocalMux I__8046 (
            .O(N__60208),
            .I(shift_srl_142Z0Z_10));
    InMux I__8045 (
            .O(N__60205),
            .I(N__60202));
    LocalMux I__8044 (
            .O(N__60202),
            .I(shift_srl_142Z0Z_11));
    InMux I__8043 (
            .O(N__60199),
            .I(N__60196));
    LocalMux I__8042 (
            .O(N__60196),
            .I(shift_srl_142Z0Z_12));
    InMux I__8041 (
            .O(N__60193),
            .I(N__60190));
    LocalMux I__8040 (
            .O(N__60190),
            .I(shift_srl_142Z0Z_13));
    InMux I__8039 (
            .O(N__60187),
            .I(N__60184));
    LocalMux I__8038 (
            .O(N__60184),
            .I(shift_srl_142Z0Z_14));
    InMux I__8037 (
            .O(N__60181),
            .I(N__60178));
    LocalMux I__8036 (
            .O(N__60178),
            .I(shift_srl_142Z0Z_9));
    InMux I__8035 (
            .O(N__60175),
            .I(N__60172));
    LocalMux I__8034 (
            .O(N__60172),
            .I(shift_srl_142Z0Z_8));
    CEMux I__8033 (
            .O(N__60169),
            .I(N__60166));
    LocalMux I__8032 (
            .O(N__60166),
            .I(N__60161));
    CEMux I__8031 (
            .O(N__60165),
            .I(N__60158));
    CEMux I__8030 (
            .O(N__60164),
            .I(N__60155));
    Span4Mux_h I__8029 (
            .O(N__60161),
            .I(N__60150));
    LocalMux I__8028 (
            .O(N__60158),
            .I(N__60150));
    LocalMux I__8027 (
            .O(N__60155),
            .I(N__60147));
    Span4Mux_h I__8026 (
            .O(N__60150),
            .I(N__60144));
    Odrv12 I__8025 (
            .O(N__60147),
            .I(clk_en_112));
    Odrv4 I__8024 (
            .O(N__60144),
            .I(clk_en_112));
    CascadeMux I__8023 (
            .O(N__60139),
            .I(rco_c_99_cascade_));
    InMux I__8022 (
            .O(N__60136),
            .I(N__60133));
    LocalMux I__8021 (
            .O(N__60133),
            .I(N__60128));
    InMux I__8020 (
            .O(N__60132),
            .I(N__60125));
    InMux I__8019 (
            .O(N__60131),
            .I(N__60122));
    Span12Mux_s10_h I__8018 (
            .O(N__60128),
            .I(N__60118));
    LocalMux I__8017 (
            .O(N__60125),
            .I(N__60113));
    LocalMux I__8016 (
            .O(N__60122),
            .I(N__60113));
    InMux I__8015 (
            .O(N__60121),
            .I(N__60110));
    Odrv12 I__8014 (
            .O(N__60118),
            .I(shift_srl_122Z0Z_15));
    Odrv12 I__8013 (
            .O(N__60113),
            .I(shift_srl_122Z0Z_15));
    LocalMux I__8012 (
            .O(N__60110),
            .I(shift_srl_122Z0Z_15));
    InMux I__8011 (
            .O(N__60103),
            .I(N__60100));
    LocalMux I__8010 (
            .O(N__60100),
            .I(shift_srl_122Z0Z_0));
    InMux I__8009 (
            .O(N__60097),
            .I(N__60094));
    LocalMux I__8008 (
            .O(N__60094),
            .I(shift_srl_122Z0Z_1));
    InMux I__8007 (
            .O(N__60091),
            .I(N__60088));
    LocalMux I__8006 (
            .O(N__60088),
            .I(shift_srl_122Z0Z_2));
    InMux I__8005 (
            .O(N__60085),
            .I(N__60082));
    LocalMux I__8004 (
            .O(N__60082),
            .I(shift_srl_122Z0Z_3));
    InMux I__8003 (
            .O(N__60079),
            .I(N__60076));
    LocalMux I__8002 (
            .O(N__60076),
            .I(shift_srl_122Z0Z_4));
    InMux I__8001 (
            .O(N__60073),
            .I(N__60070));
    LocalMux I__8000 (
            .O(N__60070),
            .I(shift_srl_122Z0Z_5));
    InMux I__7999 (
            .O(N__60067),
            .I(N__60064));
    LocalMux I__7998 (
            .O(N__60064),
            .I(shift_srl_122Z0Z_6));
    InMux I__7997 (
            .O(N__60061),
            .I(N__60058));
    LocalMux I__7996 (
            .O(N__60058),
            .I(N__60055));
    Odrv4 I__7995 (
            .O(N__60055),
            .I(shift_srl_122Z0Z_7));
    CEMux I__7994 (
            .O(N__60052),
            .I(N__60048));
    CEMux I__7993 (
            .O(N__60051),
            .I(N__60045));
    LocalMux I__7992 (
            .O(N__60048),
            .I(N__60040));
    LocalMux I__7991 (
            .O(N__60045),
            .I(N__60040));
    Odrv4 I__7990 (
            .O(N__60040),
            .I(clk_en_122));
    InMux I__7989 (
            .O(N__60037),
            .I(N__60034));
    LocalMux I__7988 (
            .O(N__60034),
            .I(shift_srl_117Z0Z_5));
    InMux I__7987 (
            .O(N__60031),
            .I(N__60028));
    LocalMux I__7986 (
            .O(N__60028),
            .I(shift_srl_117Z0Z_6));
    IoInMux I__7985 (
            .O(N__60025),
            .I(N__60022));
    LocalMux I__7984 (
            .O(N__60022),
            .I(N__60019));
    Span12Mux_s11_h I__7983 (
            .O(N__60019),
            .I(N__60016));
    Odrv12 I__7982 (
            .O(N__60016),
            .I(rco_c_143));
    IoInMux I__7981 (
            .O(N__60013),
            .I(N__60010));
    LocalMux I__7980 (
            .O(N__60010),
            .I(N__60007));
    Span4Mux_s3_h I__7979 (
            .O(N__60007),
            .I(N__60004));
    Span4Mux_h I__7978 (
            .O(N__60004),
            .I(N__60001));
    Span4Mux_h I__7977 (
            .O(N__60001),
            .I(N__59998));
    Span4Mux_h I__7976 (
            .O(N__59998),
            .I(N__59995));
    Odrv4 I__7975 (
            .O(N__59995),
            .I(rco_c_142));
    CascadeMux I__7974 (
            .O(N__59992),
            .I(clk_en_0_a3_0_a2_sx_144_cascade_));
    CEMux I__7973 (
            .O(N__59989),
            .I(N__59985));
    CEMux I__7972 (
            .O(N__59988),
            .I(N__59982));
    LocalMux I__7971 (
            .O(N__59985),
            .I(clk_en_144));
    LocalMux I__7970 (
            .O(N__59982),
            .I(clk_en_144));
    CascadeMux I__7969 (
            .O(N__59977),
            .I(clk_en_0_a3_0_a2_sx_143_cascade_));
    CEMux I__7968 (
            .O(N__59974),
            .I(N__59971));
    LocalMux I__7967 (
            .O(N__59971),
            .I(N__59967));
    CEMux I__7966 (
            .O(N__59970),
            .I(N__59964));
    Span4Mux_v I__7965 (
            .O(N__59967),
            .I(N__59959));
    LocalMux I__7964 (
            .O(N__59964),
            .I(N__59959));
    Odrv4 I__7963 (
            .O(N__59959),
            .I(clk_en_143));
    InMux I__7962 (
            .O(N__59956),
            .I(N__59953));
    LocalMux I__7961 (
            .O(N__59953),
            .I(shift_srl_143Z0Z_14));
    InMux I__7960 (
            .O(N__59950),
            .I(N__59947));
    LocalMux I__7959 (
            .O(N__59947),
            .I(shift_srl_143Z0Z_9));
    InMux I__7958 (
            .O(N__59944),
            .I(N__59941));
    LocalMux I__7957 (
            .O(N__59941),
            .I(N__59938));
    Odrv4 I__7956 (
            .O(N__59938),
            .I(shift_srl_143Z0Z_7));
    InMux I__7955 (
            .O(N__59935),
            .I(N__59932));
    LocalMux I__7954 (
            .O(N__59932),
            .I(shift_srl_143Z0Z_8));
    InMux I__7953 (
            .O(N__59929),
            .I(N__59926));
    LocalMux I__7952 (
            .O(N__59926),
            .I(shift_srl_117Z0Z_0));
    InMux I__7951 (
            .O(N__59923),
            .I(N__59920));
    LocalMux I__7950 (
            .O(N__59920),
            .I(shift_srl_117Z0Z_1));
    InMux I__7949 (
            .O(N__59917),
            .I(N__59914));
    LocalMux I__7948 (
            .O(N__59914),
            .I(shift_srl_117Z0Z_2));
    InMux I__7947 (
            .O(N__59911),
            .I(N__59908));
    LocalMux I__7946 (
            .O(N__59908),
            .I(shift_srl_117Z0Z_3));
    InMux I__7945 (
            .O(N__59905),
            .I(N__59902));
    LocalMux I__7944 (
            .O(N__59902),
            .I(shift_srl_117Z0Z_4));
    InMux I__7943 (
            .O(N__59899),
            .I(N__59896));
    LocalMux I__7942 (
            .O(N__59896),
            .I(shift_srl_121Z0Z_3));
    InMux I__7941 (
            .O(N__59893),
            .I(N__59890));
    LocalMux I__7940 (
            .O(N__59890),
            .I(shift_srl_121Z0Z_4));
    InMux I__7939 (
            .O(N__59887),
            .I(N__59884));
    LocalMux I__7938 (
            .O(N__59884),
            .I(shift_srl_121Z0Z_5));
    InMux I__7937 (
            .O(N__59881),
            .I(N__59878));
    LocalMux I__7936 (
            .O(N__59878),
            .I(shift_srl_121Z0Z_6));
    InMux I__7935 (
            .O(N__59875),
            .I(N__59872));
    LocalMux I__7934 (
            .O(N__59872),
            .I(N__59869));
    Span4Mux_v I__7933 (
            .O(N__59869),
            .I(N__59866));
    Odrv4 I__7932 (
            .O(N__59866),
            .I(shift_srl_121Z0Z_7));
    CEMux I__7931 (
            .O(N__59863),
            .I(N__59859));
    CEMux I__7930 (
            .O(N__59862),
            .I(N__59856));
    LocalMux I__7929 (
            .O(N__59859),
            .I(N__59853));
    LocalMux I__7928 (
            .O(N__59856),
            .I(N__59850));
    Span4Mux_v I__7927 (
            .O(N__59853),
            .I(N__59847));
    Span4Mux_h I__7926 (
            .O(N__59850),
            .I(N__59844));
    Odrv4 I__7925 (
            .O(N__59847),
            .I(clk_en_121));
    Odrv4 I__7924 (
            .O(N__59844),
            .I(clk_en_121));
    InMux I__7923 (
            .O(N__59839),
            .I(N__59836));
    LocalMux I__7922 (
            .O(N__59836),
            .I(shift_srl_143Z0Z_10));
    InMux I__7921 (
            .O(N__59833),
            .I(N__59830));
    LocalMux I__7920 (
            .O(N__59830),
            .I(shift_srl_143Z0Z_11));
    InMux I__7919 (
            .O(N__59827),
            .I(N__59824));
    LocalMux I__7918 (
            .O(N__59824),
            .I(shift_srl_143Z0Z_12));
    InMux I__7917 (
            .O(N__59821),
            .I(N__59818));
    LocalMux I__7916 (
            .O(N__59818),
            .I(shift_srl_143Z0Z_13));
    InMux I__7915 (
            .O(N__59815),
            .I(N__59812));
    LocalMux I__7914 (
            .O(N__59812),
            .I(shift_srl_26Z0Z_2));
    InMux I__7913 (
            .O(N__59809),
            .I(N__59806));
    LocalMux I__7912 (
            .O(N__59806),
            .I(shift_srl_26Z0Z_3));
    InMux I__7911 (
            .O(N__59803),
            .I(N__59800));
    LocalMux I__7910 (
            .O(N__59800),
            .I(shift_srl_26Z0Z_4));
    InMux I__7909 (
            .O(N__59797),
            .I(N__59794));
    LocalMux I__7908 (
            .O(N__59794),
            .I(shift_srl_26Z0Z_5));
    InMux I__7907 (
            .O(N__59791),
            .I(N__59788));
    LocalMux I__7906 (
            .O(N__59788),
            .I(shift_srl_26Z0Z_6));
    InMux I__7905 (
            .O(N__59785),
            .I(N__59782));
    LocalMux I__7904 (
            .O(N__59782),
            .I(shift_srl_121Z0Z_0));
    InMux I__7903 (
            .O(N__59779),
            .I(N__59776));
    LocalMux I__7902 (
            .O(N__59776),
            .I(shift_srl_121Z0Z_1));
    InMux I__7901 (
            .O(N__59773),
            .I(N__59770));
    LocalMux I__7900 (
            .O(N__59770),
            .I(shift_srl_121Z0Z_2));
    InMux I__7899 (
            .O(N__59767),
            .I(N__59764));
    LocalMux I__7898 (
            .O(N__59764),
            .I(shift_srl_143Z0Z_0));
    InMux I__7897 (
            .O(N__59761),
            .I(N__59758));
    LocalMux I__7896 (
            .O(N__59758),
            .I(shift_srl_143Z0Z_1));
    InMux I__7895 (
            .O(N__59755),
            .I(N__59752));
    LocalMux I__7894 (
            .O(N__59752),
            .I(shift_srl_143Z0Z_2));
    InMux I__7893 (
            .O(N__59749),
            .I(N__59746));
    LocalMux I__7892 (
            .O(N__59746),
            .I(shift_srl_143Z0Z_3));
    InMux I__7891 (
            .O(N__59743),
            .I(N__59740));
    LocalMux I__7890 (
            .O(N__59740),
            .I(shift_srl_143Z0Z_4));
    InMux I__7889 (
            .O(N__59737),
            .I(N__59734));
    LocalMux I__7888 (
            .O(N__59734),
            .I(shift_srl_143Z0Z_5));
    InMux I__7887 (
            .O(N__59731),
            .I(N__59728));
    LocalMux I__7886 (
            .O(N__59728),
            .I(shift_srl_143Z0Z_6));
    InMux I__7885 (
            .O(N__59725),
            .I(N__59722));
    LocalMux I__7884 (
            .O(N__59722),
            .I(shift_srl_26Z0Z_0));
    InMux I__7883 (
            .O(N__59719),
            .I(N__59716));
    LocalMux I__7882 (
            .O(N__59716),
            .I(shift_srl_26Z0Z_1));
    InMux I__7881 (
            .O(N__59713),
            .I(N__59710));
    LocalMux I__7880 (
            .O(N__59710),
            .I(shift_srl_89Z0Z_13));
    InMux I__7879 (
            .O(N__59707),
            .I(N__59704));
    LocalMux I__7878 (
            .O(N__59704),
            .I(shift_srl_89Z0Z_9));
    InMux I__7877 (
            .O(N__59701),
            .I(N__59698));
    LocalMux I__7876 (
            .O(N__59698),
            .I(shift_srl_89Z0Z_7));
    InMux I__7875 (
            .O(N__59695),
            .I(N__59692));
    LocalMux I__7874 (
            .O(N__59692),
            .I(shift_srl_89Z0Z_8));
    InMux I__7873 (
            .O(N__59689),
            .I(N__59686));
    LocalMux I__7872 (
            .O(N__59686),
            .I(shift_srl_24Z0Z_0));
    InMux I__7871 (
            .O(N__59683),
            .I(N__59680));
    LocalMux I__7870 (
            .O(N__59680),
            .I(shift_srl_24Z0Z_1));
    InMux I__7869 (
            .O(N__59677),
            .I(N__59674));
    LocalMux I__7868 (
            .O(N__59674),
            .I(shift_srl_24Z0Z_2));
    InMux I__7867 (
            .O(N__59671),
            .I(N__59668));
    LocalMux I__7866 (
            .O(N__59668),
            .I(shift_srl_89Z0Z_2));
    InMux I__7865 (
            .O(N__59665),
            .I(N__59662));
    LocalMux I__7864 (
            .O(N__59662),
            .I(shift_srl_89Z0Z_3));
    InMux I__7863 (
            .O(N__59659),
            .I(N__59656));
    LocalMux I__7862 (
            .O(N__59656),
            .I(shift_srl_89Z0Z_4));
    InMux I__7861 (
            .O(N__59653),
            .I(N__59650));
    LocalMux I__7860 (
            .O(N__59650),
            .I(shift_srl_89Z0Z_5));
    InMux I__7859 (
            .O(N__59647),
            .I(N__59644));
    LocalMux I__7858 (
            .O(N__59644),
            .I(shift_srl_89Z0Z_6));
    InMux I__7857 (
            .O(N__59641),
            .I(N__59638));
    LocalMux I__7856 (
            .O(N__59638),
            .I(shift_srl_89Z0Z_10));
    InMux I__7855 (
            .O(N__59635),
            .I(N__59632));
    LocalMux I__7854 (
            .O(N__59632),
            .I(shift_srl_89Z0Z_11));
    InMux I__7853 (
            .O(N__59629),
            .I(N__59626));
    LocalMux I__7852 (
            .O(N__59626),
            .I(shift_srl_89Z0Z_12));
    InMux I__7851 (
            .O(N__59623),
            .I(N__59620));
    LocalMux I__7850 (
            .O(N__59620),
            .I(shift_srl_25Z0Z_11));
    InMux I__7849 (
            .O(N__59617),
            .I(N__59614));
    LocalMux I__7848 (
            .O(N__59614),
            .I(shift_srl_25Z0Z_12));
    InMux I__7847 (
            .O(N__59611),
            .I(N__59608));
    LocalMux I__7846 (
            .O(N__59608),
            .I(shift_srl_25Z0Z_13));
    InMux I__7845 (
            .O(N__59605),
            .I(N__59602));
    LocalMux I__7844 (
            .O(N__59602),
            .I(shift_srl_25Z0Z_14));
    InMux I__7843 (
            .O(N__59599),
            .I(N__59596));
    LocalMux I__7842 (
            .O(N__59596),
            .I(shift_srl_25Z0Z_9));
    InMux I__7841 (
            .O(N__59593),
            .I(N__59590));
    LocalMux I__7840 (
            .O(N__59590),
            .I(shift_srl_25Z0Z_7));
    InMux I__7839 (
            .O(N__59587),
            .I(N__59584));
    LocalMux I__7838 (
            .O(N__59584),
            .I(shift_srl_25Z0Z_8));
    CEMux I__7837 (
            .O(N__59581),
            .I(N__59578));
    LocalMux I__7836 (
            .O(N__59578),
            .I(N__59575));
    Span4Mux_v I__7835 (
            .O(N__59575),
            .I(N__59569));
    CEMux I__7834 (
            .O(N__59574),
            .I(N__59566));
    CEMux I__7833 (
            .O(N__59573),
            .I(N__59563));
    CEMux I__7832 (
            .O(N__59572),
            .I(N__59560));
    Sp12to4 I__7831 (
            .O(N__59569),
            .I(N__59555));
    LocalMux I__7830 (
            .O(N__59566),
            .I(N__59555));
    LocalMux I__7829 (
            .O(N__59563),
            .I(N__59552));
    LocalMux I__7828 (
            .O(N__59560),
            .I(N__59549));
    Odrv12 I__7827 (
            .O(N__59555),
            .I(clk_en_25));
    Odrv12 I__7826 (
            .O(N__59552),
            .I(clk_en_25));
    Odrv4 I__7825 (
            .O(N__59549),
            .I(clk_en_25));
    InMux I__7824 (
            .O(N__59542),
            .I(N__59539));
    LocalMux I__7823 (
            .O(N__59539),
            .I(shift_srl_89Z0Z_0));
    InMux I__7822 (
            .O(N__59536),
            .I(N__59533));
    LocalMux I__7821 (
            .O(N__59533),
            .I(shift_srl_89Z0Z_1));
    InMux I__7820 (
            .O(N__59530),
            .I(N__59527));
    LocalMux I__7819 (
            .O(N__59527),
            .I(shift_srl_91Z0Z_3));
    InMux I__7818 (
            .O(N__59524),
            .I(N__59521));
    LocalMux I__7817 (
            .O(N__59521),
            .I(shift_srl_91Z0Z_4));
    InMux I__7816 (
            .O(N__59518),
            .I(N__59515));
    LocalMux I__7815 (
            .O(N__59515),
            .I(shift_srl_91Z0Z_5));
    InMux I__7814 (
            .O(N__59512),
            .I(N__59509));
    LocalMux I__7813 (
            .O(N__59509),
            .I(shift_srl_91Z0Z_6));
    InMux I__7812 (
            .O(N__59506),
            .I(N__59503));
    LocalMux I__7811 (
            .O(N__59503),
            .I(shift_srl_91Z0Z_7));
    InMux I__7810 (
            .O(N__59500),
            .I(N__59497));
    LocalMux I__7809 (
            .O(N__59497),
            .I(shift_srl_25Z0Z_4));
    InMux I__7808 (
            .O(N__59494),
            .I(N__59491));
    LocalMux I__7807 (
            .O(N__59491),
            .I(shift_srl_25Z0Z_5));
    InMux I__7806 (
            .O(N__59488),
            .I(N__59485));
    LocalMux I__7805 (
            .O(N__59485),
            .I(shift_srl_25Z0Z_6));
    InMux I__7804 (
            .O(N__59482),
            .I(N__59479));
    LocalMux I__7803 (
            .O(N__59479),
            .I(shift_srl_25Z0Z_10));
    InMux I__7802 (
            .O(N__59476),
            .I(N__59473));
    LocalMux I__7801 (
            .O(N__59473),
            .I(shift_srl_91Z0Z_11));
    InMux I__7800 (
            .O(N__59470),
            .I(N__59467));
    LocalMux I__7799 (
            .O(N__59467),
            .I(shift_srl_91Z0Z_12));
    InMux I__7798 (
            .O(N__59464),
            .I(N__59461));
    LocalMux I__7797 (
            .O(N__59461),
            .I(shift_srl_91Z0Z_13));
    InMux I__7796 (
            .O(N__59458),
            .I(N__59455));
    LocalMux I__7795 (
            .O(N__59455),
            .I(shift_srl_91Z0Z_14));
    InMux I__7794 (
            .O(N__59452),
            .I(N__59449));
    LocalMux I__7793 (
            .O(N__59449),
            .I(shift_srl_91Z0Z_9));
    InMux I__7792 (
            .O(N__59446),
            .I(N__59443));
    LocalMux I__7791 (
            .O(N__59443),
            .I(shift_srl_91Z0Z_8));
    InMux I__7790 (
            .O(N__59440),
            .I(N__59437));
    LocalMux I__7789 (
            .O(N__59437),
            .I(shift_srl_91Z0Z_0));
    InMux I__7788 (
            .O(N__59434),
            .I(N__59431));
    LocalMux I__7787 (
            .O(N__59431),
            .I(shift_srl_91Z0Z_1));
    InMux I__7786 (
            .O(N__59428),
            .I(N__59425));
    LocalMux I__7785 (
            .O(N__59425),
            .I(shift_srl_91Z0Z_2));
    InMux I__7784 (
            .O(N__59422),
            .I(N__59419));
    LocalMux I__7783 (
            .O(N__59419),
            .I(N__59416));
    Odrv4 I__7782 (
            .O(N__59416),
            .I(shift_srl_103Z0Z_6));
    IoInMux I__7781 (
            .O(N__59413),
            .I(N__59410));
    LocalMux I__7780 (
            .O(N__59410),
            .I(N__59407));
    Span12Mux_s3_v I__7779 (
            .O(N__59407),
            .I(N__59404));
    Odrv12 I__7778 (
            .O(N__59404),
            .I(rco_c_165));
    InMux I__7777 (
            .O(N__59401),
            .I(N__59398));
    LocalMux I__7776 (
            .O(N__59398),
            .I(shift_srl_90Z0Z_9));
    InMux I__7775 (
            .O(N__59395),
            .I(N__59392));
    LocalMux I__7774 (
            .O(N__59392),
            .I(shift_srl_90Z0Z_8));
    InMux I__7773 (
            .O(N__59389),
            .I(N__59386));
    LocalMux I__7772 (
            .O(N__59386),
            .I(shift_srl_90Z0Z_6));
    InMux I__7771 (
            .O(N__59383),
            .I(N__59380));
    LocalMux I__7770 (
            .O(N__59380),
            .I(shift_srl_90Z0Z_7));
    InMux I__7769 (
            .O(N__59377),
            .I(N__59374));
    LocalMux I__7768 (
            .O(N__59374),
            .I(shift_srl_91Z0Z_10));
    InMux I__7767 (
            .O(N__59371),
            .I(N__59368));
    LocalMux I__7766 (
            .O(N__59368),
            .I(shift_srl_103Z0Z_1));
    InMux I__7765 (
            .O(N__59365),
            .I(N__59362));
    LocalMux I__7764 (
            .O(N__59362),
            .I(shift_srl_103Z0Z_2));
    InMux I__7763 (
            .O(N__59359),
            .I(N__59356));
    LocalMux I__7762 (
            .O(N__59356),
            .I(shift_srl_103Z0Z_3));
    InMux I__7761 (
            .O(N__59353),
            .I(N__59350));
    LocalMux I__7760 (
            .O(N__59350),
            .I(shift_srl_103Z0Z_4));
    InMux I__7759 (
            .O(N__59347),
            .I(N__59344));
    LocalMux I__7758 (
            .O(N__59344),
            .I(shift_srl_103Z0Z_5));
    InMux I__7757 (
            .O(N__59341),
            .I(N__59338));
    LocalMux I__7756 (
            .O(N__59338),
            .I(shift_srl_100Z0Z_9));
    InMux I__7755 (
            .O(N__59335),
            .I(N__59332));
    LocalMux I__7754 (
            .O(N__59332),
            .I(shift_srl_100Z0Z_8));
    InMux I__7753 (
            .O(N__59329),
            .I(N__59326));
    LocalMux I__7752 (
            .O(N__59326),
            .I(N__59323));
    Span4Mux_v I__7751 (
            .O(N__59323),
            .I(N__59320));
    Odrv4 I__7750 (
            .O(N__59320),
            .I(shift_srl_100Z0Z_6));
    InMux I__7749 (
            .O(N__59317),
            .I(N__59314));
    LocalMux I__7748 (
            .O(N__59314),
            .I(shift_srl_100Z0Z_7));
    CascadeMux I__7747 (
            .O(N__59311),
            .I(shift_srl_102_RNIN8GNZ0Z_15_cascade_));
    CEMux I__7746 (
            .O(N__59308),
            .I(N__59304));
    CEMux I__7745 (
            .O(N__59307),
            .I(N__59301));
    LocalMux I__7744 (
            .O(N__59304),
            .I(clk_en_104));
    LocalMux I__7743 (
            .O(N__59301),
            .I(clk_en_104));
    InMux I__7742 (
            .O(N__59296),
            .I(N__59293));
    LocalMux I__7741 (
            .O(N__59293),
            .I(shift_srl_101Z0Z_14));
    InMux I__7740 (
            .O(N__59290),
            .I(N__59285));
    InMux I__7739 (
            .O(N__59289),
            .I(N__59275));
    InMux I__7738 (
            .O(N__59288),
            .I(N__59275));
    LocalMux I__7737 (
            .O(N__59285),
            .I(N__59272));
    InMux I__7736 (
            .O(N__59284),
            .I(N__59263));
    InMux I__7735 (
            .O(N__59283),
            .I(N__59263));
    InMux I__7734 (
            .O(N__59282),
            .I(N__59263));
    InMux I__7733 (
            .O(N__59281),
            .I(N__59263));
    InMux I__7732 (
            .O(N__59280),
            .I(N__59260));
    LocalMux I__7731 (
            .O(N__59275),
            .I(shift_srl_105Z0Z_15));
    Odrv4 I__7730 (
            .O(N__59272),
            .I(shift_srl_105Z0Z_15));
    LocalMux I__7729 (
            .O(N__59263),
            .I(shift_srl_105Z0Z_15));
    LocalMux I__7728 (
            .O(N__59260),
            .I(shift_srl_105Z0Z_15));
    InMux I__7727 (
            .O(N__59251),
            .I(N__59247));
    CascadeMux I__7726 (
            .O(N__59250),
            .I(N__59243));
    LocalMux I__7725 (
            .O(N__59247),
            .I(N__59239));
    CascadeMux I__7724 (
            .O(N__59246),
            .I(N__59236));
    InMux I__7723 (
            .O(N__59243),
            .I(N__59231));
    InMux I__7722 (
            .O(N__59242),
            .I(N__59228));
    Span4Mux_h I__7721 (
            .O(N__59239),
            .I(N__59225));
    InMux I__7720 (
            .O(N__59236),
            .I(N__59218));
    InMux I__7719 (
            .O(N__59235),
            .I(N__59218));
    InMux I__7718 (
            .O(N__59234),
            .I(N__59218));
    LocalMux I__7717 (
            .O(N__59231),
            .I(N__59215));
    LocalMux I__7716 (
            .O(N__59228),
            .I(shift_srl_106Z0Z_15));
    Odrv4 I__7715 (
            .O(N__59225),
            .I(shift_srl_106Z0Z_15));
    LocalMux I__7714 (
            .O(N__59218),
            .I(shift_srl_106Z0Z_15));
    Odrv4 I__7713 (
            .O(N__59215),
            .I(shift_srl_106Z0Z_15));
    CEMux I__7712 (
            .O(N__59206),
            .I(N__59201));
    CEMux I__7711 (
            .O(N__59205),
            .I(N__59198));
    CEMux I__7710 (
            .O(N__59204),
            .I(N__59195));
    LocalMux I__7709 (
            .O(N__59201),
            .I(N__59189));
    LocalMux I__7708 (
            .O(N__59198),
            .I(N__59189));
    LocalMux I__7707 (
            .O(N__59195),
            .I(N__59186));
    CEMux I__7706 (
            .O(N__59194),
            .I(N__59183));
    Span4Mux_v I__7705 (
            .O(N__59189),
            .I(N__59180));
    Span4Mux_v I__7704 (
            .O(N__59186),
            .I(N__59175));
    LocalMux I__7703 (
            .O(N__59183),
            .I(N__59175));
    Odrv4 I__7702 (
            .O(N__59180),
            .I(clk_en_101));
    Odrv4 I__7701 (
            .O(N__59175),
            .I(clk_en_101));
    CascadeMux I__7700 (
            .O(N__59170),
            .I(clk_en_0_a3_0_a2_sx_103_cascade_));
    IoInMux I__7699 (
            .O(N__59167),
            .I(N__59164));
    LocalMux I__7698 (
            .O(N__59164),
            .I(N__59161));
    IoSpan4Mux I__7697 (
            .O(N__59161),
            .I(N__59158));
    Span4Mux_s1_h I__7696 (
            .O(N__59158),
            .I(N__59155));
    Sp12to4 I__7695 (
            .O(N__59155),
            .I(N__59152));
    Span12Mux_h I__7694 (
            .O(N__59152),
            .I(N__59148));
    InMux I__7693 (
            .O(N__59151),
            .I(N__59145));
    Odrv12 I__7692 (
            .O(N__59148),
            .I(rco_c_102));
    LocalMux I__7691 (
            .O(N__59145),
            .I(rco_c_102));
    IoInMux I__7690 (
            .O(N__59140),
            .I(N__59137));
    LocalMux I__7689 (
            .O(N__59137),
            .I(N__59134));
    IoSpan4Mux I__7688 (
            .O(N__59134),
            .I(N__59131));
    Span4Mux_s3_h I__7687 (
            .O(N__59131),
            .I(N__59128));
    Span4Mux_h I__7686 (
            .O(N__59128),
            .I(N__59125));
    Span4Mux_h I__7685 (
            .O(N__59125),
            .I(N__59122));
    Odrv4 I__7684 (
            .O(N__59122),
            .I(rco_c_103));
    InMux I__7683 (
            .O(N__59119),
            .I(N__59116));
    LocalMux I__7682 (
            .O(N__59116),
            .I(shift_srl_103Z0Z_0));
    InMux I__7681 (
            .O(N__59113),
            .I(N__59110));
    LocalMux I__7680 (
            .O(N__59110),
            .I(shift_srl_104Z0Z_10));
    InMux I__7679 (
            .O(N__59107),
            .I(N__59104));
    LocalMux I__7678 (
            .O(N__59104),
            .I(shift_srl_104Z0Z_11));
    InMux I__7677 (
            .O(N__59101),
            .I(N__59098));
    LocalMux I__7676 (
            .O(N__59098),
            .I(shift_srl_104Z0Z_12));
    InMux I__7675 (
            .O(N__59095),
            .I(N__59092));
    LocalMux I__7674 (
            .O(N__59092),
            .I(shift_srl_104Z0Z_13));
    InMux I__7673 (
            .O(N__59089),
            .I(N__59086));
    LocalMux I__7672 (
            .O(N__59086),
            .I(shift_srl_104Z0Z_14));
    InMux I__7671 (
            .O(N__59083),
            .I(N__59080));
    LocalMux I__7670 (
            .O(N__59080),
            .I(shift_srl_104Z0Z_9));
    InMux I__7669 (
            .O(N__59077),
            .I(N__59074));
    LocalMux I__7668 (
            .O(N__59074),
            .I(shift_srl_104Z0Z_7));
    InMux I__7667 (
            .O(N__59071),
            .I(N__59068));
    LocalMux I__7666 (
            .O(N__59068),
            .I(shift_srl_104Z0Z_8));
    InMux I__7665 (
            .O(N__59065),
            .I(N__59062));
    LocalMux I__7664 (
            .O(N__59062),
            .I(shift_srl_118Z0Z_5));
    InMux I__7663 (
            .O(N__59059),
            .I(N__59056));
    LocalMux I__7662 (
            .O(N__59056),
            .I(shift_srl_118Z0Z_6));
    InMux I__7661 (
            .O(N__59053),
            .I(N__59050));
    LocalMux I__7660 (
            .O(N__59050),
            .I(N__59047));
    Span4Mux_v I__7659 (
            .O(N__59047),
            .I(N__59044));
    Odrv4 I__7658 (
            .O(N__59044),
            .I(shift_srl_118Z0Z_7));
    InMux I__7657 (
            .O(N__59041),
            .I(N__59038));
    LocalMux I__7656 (
            .O(N__59038),
            .I(shift_srl_100Z0Z_0));
    InMux I__7655 (
            .O(N__59035),
            .I(N__59032));
    LocalMux I__7654 (
            .O(N__59032),
            .I(shift_srl_100Z0Z_1));
    InMux I__7653 (
            .O(N__59029),
            .I(N__59026));
    LocalMux I__7652 (
            .O(N__59026),
            .I(shift_srl_100Z0Z_2));
    InMux I__7651 (
            .O(N__59023),
            .I(N__59020));
    LocalMux I__7650 (
            .O(N__59020),
            .I(shift_srl_100Z0Z_3));
    InMux I__7649 (
            .O(N__59017),
            .I(N__59014));
    LocalMux I__7648 (
            .O(N__59014),
            .I(shift_srl_100Z0Z_4));
    InMux I__7647 (
            .O(N__59011),
            .I(N__59008));
    LocalMux I__7646 (
            .O(N__59008),
            .I(shift_srl_100Z0Z_5));
    InMux I__7645 (
            .O(N__59005),
            .I(N__59002));
    LocalMux I__7644 (
            .O(N__59002),
            .I(shift_srl_114Z0Z_4));
    InMux I__7643 (
            .O(N__58999),
            .I(N__58996));
    LocalMux I__7642 (
            .O(N__58996),
            .I(shift_srl_114Z0Z_5));
    InMux I__7641 (
            .O(N__58993),
            .I(N__58990));
    LocalMux I__7640 (
            .O(N__58990),
            .I(shift_srl_114Z0Z_6));
    InMux I__7639 (
            .O(N__58987),
            .I(N__58984));
    LocalMux I__7638 (
            .O(N__58984),
            .I(shift_srl_114Z0Z_7));
    InMux I__7637 (
            .O(N__58981),
            .I(N__58978));
    LocalMux I__7636 (
            .O(N__58978),
            .I(shift_srl_118Z0Z_0));
    InMux I__7635 (
            .O(N__58975),
            .I(N__58972));
    LocalMux I__7634 (
            .O(N__58972),
            .I(shift_srl_118Z0Z_1));
    InMux I__7633 (
            .O(N__58969),
            .I(N__58966));
    LocalMux I__7632 (
            .O(N__58966),
            .I(shift_srl_118Z0Z_2));
    InMux I__7631 (
            .O(N__58963),
            .I(N__58960));
    LocalMux I__7630 (
            .O(N__58960),
            .I(shift_srl_118Z0Z_3));
    InMux I__7629 (
            .O(N__58957),
            .I(N__58954));
    LocalMux I__7628 (
            .O(N__58954),
            .I(shift_srl_118Z0Z_4));
    InMux I__7627 (
            .O(N__58951),
            .I(N__58948));
    LocalMux I__7626 (
            .O(N__58948),
            .I(shift_srl_114Z0Z_13));
    InMux I__7625 (
            .O(N__58945),
            .I(N__58942));
    LocalMux I__7624 (
            .O(N__58942),
            .I(shift_srl_114Z0Z_14));
    InMux I__7623 (
            .O(N__58939),
            .I(N__58936));
    LocalMux I__7622 (
            .O(N__58936),
            .I(shift_srl_114Z0Z_9));
    InMux I__7621 (
            .O(N__58933),
            .I(N__58930));
    LocalMux I__7620 (
            .O(N__58930),
            .I(shift_srl_114Z0Z_8));
    InMux I__7619 (
            .O(N__58927),
            .I(N__58924));
    LocalMux I__7618 (
            .O(N__58924),
            .I(N__58921));
    Span4Mux_v I__7617 (
            .O(N__58921),
            .I(N__58913));
    InMux I__7616 (
            .O(N__58920),
            .I(N__58904));
    InMux I__7615 (
            .O(N__58919),
            .I(N__58904));
    InMux I__7614 (
            .O(N__58918),
            .I(N__58904));
    InMux I__7613 (
            .O(N__58917),
            .I(N__58904));
    InMux I__7612 (
            .O(N__58916),
            .I(N__58900));
    Span4Mux_h I__7611 (
            .O(N__58913),
            .I(N__58895));
    LocalMux I__7610 (
            .O(N__58904),
            .I(N__58895));
    InMux I__7609 (
            .O(N__58903),
            .I(N__58892));
    LocalMux I__7608 (
            .O(N__58900),
            .I(shift_srl_114Z0Z_15));
    Odrv4 I__7607 (
            .O(N__58895),
            .I(shift_srl_114Z0Z_15));
    LocalMux I__7606 (
            .O(N__58892),
            .I(shift_srl_114Z0Z_15));
    InMux I__7605 (
            .O(N__58885),
            .I(N__58882));
    LocalMux I__7604 (
            .O(N__58882),
            .I(shift_srl_114Z0Z_0));
    InMux I__7603 (
            .O(N__58879),
            .I(N__58876));
    LocalMux I__7602 (
            .O(N__58876),
            .I(shift_srl_114Z0Z_1));
    InMux I__7601 (
            .O(N__58873),
            .I(N__58870));
    LocalMux I__7600 (
            .O(N__58870),
            .I(shift_srl_114Z0Z_2));
    InMux I__7599 (
            .O(N__58867),
            .I(N__58864));
    LocalMux I__7598 (
            .O(N__58864),
            .I(shift_srl_114Z0Z_3));
    InMux I__7597 (
            .O(N__58861),
            .I(N__58858));
    LocalMux I__7596 (
            .O(N__58858),
            .I(shift_srl_117Z0Z_14));
    InMux I__7595 (
            .O(N__58855),
            .I(N__58852));
    LocalMux I__7594 (
            .O(N__58852),
            .I(shift_srl_117Z0Z_13));
    InMux I__7593 (
            .O(N__58849),
            .I(N__58846));
    LocalMux I__7592 (
            .O(N__58846),
            .I(shift_srl_117Z0Z_12));
    InMux I__7591 (
            .O(N__58843),
            .I(N__58840));
    LocalMux I__7590 (
            .O(N__58840),
            .I(shift_srl_117Z0Z_11));
    InMux I__7589 (
            .O(N__58837),
            .I(N__58834));
    LocalMux I__7588 (
            .O(N__58834),
            .I(shift_srl_117Z0Z_10));
    InMux I__7587 (
            .O(N__58831),
            .I(N__58828));
    LocalMux I__7586 (
            .O(N__58828),
            .I(shift_srl_114Z0Z_10));
    InMux I__7585 (
            .O(N__58825),
            .I(N__58822));
    LocalMux I__7584 (
            .O(N__58822),
            .I(shift_srl_114Z0Z_11));
    InMux I__7583 (
            .O(N__58819),
            .I(N__58816));
    LocalMux I__7582 (
            .O(N__58816),
            .I(shift_srl_114Z0Z_12));
    CascadeMux I__7581 (
            .O(N__58813),
            .I(N__58810));
    InMux I__7580 (
            .O(N__58810),
            .I(N__58804));
    InMux I__7579 (
            .O(N__58809),
            .I(N__58804));
    LocalMux I__7578 (
            .O(N__58804),
            .I(N__58797));
    CascadeMux I__7577 (
            .O(N__58803),
            .I(N__58794));
    InMux I__7576 (
            .O(N__58802),
            .I(N__58791));
    InMux I__7575 (
            .O(N__58801),
            .I(N__58788));
    InMux I__7574 (
            .O(N__58800),
            .I(N__58782));
    Span4Mux_v I__7573 (
            .O(N__58797),
            .I(N__58779));
    InMux I__7572 (
            .O(N__58794),
            .I(N__58776));
    LocalMux I__7571 (
            .O(N__58791),
            .I(N__58773));
    LocalMux I__7570 (
            .O(N__58788),
            .I(N__58770));
    InMux I__7569 (
            .O(N__58787),
            .I(N__58767));
    InMux I__7568 (
            .O(N__58786),
            .I(N__58762));
    InMux I__7567 (
            .O(N__58785),
            .I(N__58762));
    LocalMux I__7566 (
            .O(N__58782),
            .I(N__58755));
    Sp12to4 I__7565 (
            .O(N__58779),
            .I(N__58755));
    LocalMux I__7564 (
            .O(N__58776),
            .I(N__58755));
    Odrv4 I__7563 (
            .O(N__58773),
            .I(shift_srl_116Z0Z_15));
    Odrv4 I__7562 (
            .O(N__58770),
            .I(shift_srl_116Z0Z_15));
    LocalMux I__7561 (
            .O(N__58767),
            .I(shift_srl_116Z0Z_15));
    LocalMux I__7560 (
            .O(N__58762),
            .I(shift_srl_116Z0Z_15));
    Odrv12 I__7559 (
            .O(N__58755),
            .I(shift_srl_116Z0Z_15));
    CascadeMux I__7558 (
            .O(N__58744),
            .I(rco_int_0_a2_1_a2_1_118_cascade_));
    CascadeMux I__7557 (
            .O(N__58741),
            .I(rco_c_118_cascade_));
    InMux I__7556 (
            .O(N__58738),
            .I(N__58735));
    LocalMux I__7555 (
            .O(N__58735),
            .I(N__58732));
    Span4Mux_h I__7554 (
            .O(N__58732),
            .I(N__58729));
    Span4Mux_h I__7553 (
            .O(N__58729),
            .I(N__58726));
    Odrv4 I__7552 (
            .O(N__58726),
            .I(rco_int_0_a2_1_a2_1_123));
    CEMux I__7551 (
            .O(N__58723),
            .I(N__58719));
    CEMux I__7550 (
            .O(N__58722),
            .I(N__58715));
    LocalMux I__7549 (
            .O(N__58719),
            .I(N__58712));
    CEMux I__7548 (
            .O(N__58718),
            .I(N__58709));
    LocalMux I__7547 (
            .O(N__58715),
            .I(N__58706));
    Span4Mux_h I__7546 (
            .O(N__58712),
            .I(N__58703));
    LocalMux I__7545 (
            .O(N__58709),
            .I(N__58700));
    Span4Mux_h I__7544 (
            .O(N__58706),
            .I(N__58697));
    Odrv4 I__7543 (
            .O(N__58703),
            .I(clk_en_124));
    Odrv12 I__7542 (
            .O(N__58700),
            .I(clk_en_124));
    Odrv4 I__7541 (
            .O(N__58697),
            .I(clk_en_124));
    InMux I__7540 (
            .O(N__58690),
            .I(N__58687));
    LocalMux I__7539 (
            .O(N__58687),
            .I(shift_srl_144Z0Z_6));
    InMux I__7538 (
            .O(N__58684),
            .I(N__58681));
    LocalMux I__7537 (
            .O(N__58681),
            .I(shift_srl_144Z0Z_10));
    InMux I__7536 (
            .O(N__58678),
            .I(N__58675));
    LocalMux I__7535 (
            .O(N__58675),
            .I(shift_srl_144Z0Z_11));
    InMux I__7534 (
            .O(N__58672),
            .I(N__58669));
    LocalMux I__7533 (
            .O(N__58669),
            .I(shift_srl_144Z0Z_12));
    InMux I__7532 (
            .O(N__58666),
            .I(N__58663));
    LocalMux I__7531 (
            .O(N__58663),
            .I(shift_srl_144Z0Z_13));
    InMux I__7530 (
            .O(N__58660),
            .I(N__58657));
    LocalMux I__7529 (
            .O(N__58657),
            .I(shift_srl_144Z0Z_14));
    InMux I__7528 (
            .O(N__58654),
            .I(N__58651));
    LocalMux I__7527 (
            .O(N__58651),
            .I(shift_srl_144Z0Z_9));
    InMux I__7526 (
            .O(N__58648),
            .I(N__58645));
    LocalMux I__7525 (
            .O(N__58645),
            .I(shift_srl_144Z0Z_7));
    InMux I__7524 (
            .O(N__58642),
            .I(N__58639));
    LocalMux I__7523 (
            .O(N__58639),
            .I(shift_srl_144Z0Z_8));
    InMux I__7522 (
            .O(N__58636),
            .I(N__58633));
    LocalMux I__7521 (
            .O(N__58633),
            .I(shift_srl_124Z0Z_5));
    InMux I__7520 (
            .O(N__58630),
            .I(N__58627));
    LocalMux I__7519 (
            .O(N__58627),
            .I(shift_srl_124Z0Z_6));
    InMux I__7518 (
            .O(N__58624),
            .I(N__58621));
    LocalMux I__7517 (
            .O(N__58621),
            .I(shift_srl_124Z0Z_7));
    InMux I__7516 (
            .O(N__58618),
            .I(N__58615));
    LocalMux I__7515 (
            .O(N__58615),
            .I(shift_srl_144Z0Z_0));
    InMux I__7514 (
            .O(N__58612),
            .I(N__58609));
    LocalMux I__7513 (
            .O(N__58609),
            .I(shift_srl_144Z0Z_1));
    InMux I__7512 (
            .O(N__58606),
            .I(N__58603));
    LocalMux I__7511 (
            .O(N__58603),
            .I(shift_srl_144Z0Z_2));
    InMux I__7510 (
            .O(N__58600),
            .I(N__58597));
    LocalMux I__7509 (
            .O(N__58597),
            .I(shift_srl_144Z0Z_3));
    InMux I__7508 (
            .O(N__58594),
            .I(N__58591));
    LocalMux I__7507 (
            .O(N__58591),
            .I(shift_srl_144Z0Z_4));
    InMux I__7506 (
            .O(N__58588),
            .I(N__58585));
    LocalMux I__7505 (
            .O(N__58585),
            .I(shift_srl_144Z0Z_5));
    InMux I__7504 (
            .O(N__58582),
            .I(N__58579));
    LocalMux I__7503 (
            .O(N__58579),
            .I(shift_srl_155Z0Z_14));
    InMux I__7502 (
            .O(N__58576),
            .I(N__58573));
    LocalMux I__7501 (
            .O(N__58573),
            .I(shift_srl_155Z0Z_2));
    InMux I__7500 (
            .O(N__58570),
            .I(N__58567));
    LocalMux I__7499 (
            .O(N__58567),
            .I(shift_srl_155Z0Z_3));
    InMux I__7498 (
            .O(N__58564),
            .I(N__58561));
    LocalMux I__7497 (
            .O(N__58561),
            .I(shift_srl_155Z0Z_10));
    InMux I__7496 (
            .O(N__58558),
            .I(N__58555));
    LocalMux I__7495 (
            .O(N__58555),
            .I(shift_srl_155Z0Z_11));
    CEMux I__7494 (
            .O(N__58552),
            .I(N__58548));
    CEMux I__7493 (
            .O(N__58551),
            .I(N__58545));
    LocalMux I__7492 (
            .O(N__58548),
            .I(clk_en_155));
    LocalMux I__7491 (
            .O(N__58545),
            .I(clk_en_155));
    InMux I__7490 (
            .O(N__58540),
            .I(N__58537));
    LocalMux I__7489 (
            .O(N__58537),
            .I(shift_srl_124Z0Z_0));
    InMux I__7488 (
            .O(N__58534),
            .I(N__58531));
    LocalMux I__7487 (
            .O(N__58531),
            .I(shift_srl_124Z0Z_1));
    InMux I__7486 (
            .O(N__58528),
            .I(N__58525));
    LocalMux I__7485 (
            .O(N__58525),
            .I(shift_srl_124Z0Z_2));
    InMux I__7484 (
            .O(N__58522),
            .I(N__58519));
    LocalMux I__7483 (
            .O(N__58519),
            .I(shift_srl_124Z0Z_3));
    InMux I__7482 (
            .O(N__58516),
            .I(N__58513));
    LocalMux I__7481 (
            .O(N__58513),
            .I(shift_srl_124Z0Z_4));
    InMux I__7480 (
            .O(N__58510),
            .I(N__58507));
    LocalMux I__7479 (
            .O(N__58507),
            .I(shift_srl_155Z0Z_6));
    InMux I__7478 (
            .O(N__58504),
            .I(N__58501));
    LocalMux I__7477 (
            .O(N__58501),
            .I(shift_srl_155Z0Z_9));
    InMux I__7476 (
            .O(N__58498),
            .I(N__58495));
    LocalMux I__7475 (
            .O(N__58495),
            .I(shift_srl_155Z0Z_5));
    InMux I__7474 (
            .O(N__58492),
            .I(N__58489));
    LocalMux I__7473 (
            .O(N__58489),
            .I(shift_srl_155Z0Z_4));
    InMux I__7472 (
            .O(N__58486),
            .I(N__58483));
    LocalMux I__7471 (
            .O(N__58483),
            .I(shift_srl_155Z0Z_7));
    InMux I__7470 (
            .O(N__58480),
            .I(N__58477));
    LocalMux I__7469 (
            .O(N__58477),
            .I(shift_srl_155Z0Z_8));
    InMux I__7468 (
            .O(N__58474),
            .I(N__58471));
    LocalMux I__7467 (
            .O(N__58471),
            .I(shift_srl_155Z0Z_12));
    InMux I__7466 (
            .O(N__58468),
            .I(N__58465));
    LocalMux I__7465 (
            .O(N__58465),
            .I(shift_srl_155Z0Z_13));
    InMux I__7464 (
            .O(N__58462),
            .I(N__58459));
    LocalMux I__7463 (
            .O(N__58459),
            .I(shift_srl_157Z0Z_2));
    InMux I__7462 (
            .O(N__58456),
            .I(N__58453));
    LocalMux I__7461 (
            .O(N__58453),
            .I(shift_srl_157Z0Z_3));
    InMux I__7460 (
            .O(N__58450),
            .I(N__58447));
    LocalMux I__7459 (
            .O(N__58447),
            .I(shift_srl_157Z0Z_4));
    InMux I__7458 (
            .O(N__58444),
            .I(N__58441));
    LocalMux I__7457 (
            .O(N__58441),
            .I(shift_srl_157Z0Z_12));
    InMux I__7456 (
            .O(N__58438),
            .I(N__58435));
    LocalMux I__7455 (
            .O(N__58435),
            .I(shift_srl_157Z0Z_13));
    InMux I__7454 (
            .O(N__58432),
            .I(N__58429));
    LocalMux I__7453 (
            .O(N__58429),
            .I(shift_srl_157Z0Z_14));
    InMux I__7452 (
            .O(N__58426),
            .I(N__58423));
    LocalMux I__7451 (
            .O(N__58423),
            .I(shift_srl_157Z0Z_6));
    InMux I__7450 (
            .O(N__58420),
            .I(N__58417));
    LocalMux I__7449 (
            .O(N__58417),
            .I(shift_srl_157Z0Z_7));
    CEMux I__7448 (
            .O(N__58414),
            .I(N__58410));
    CEMux I__7447 (
            .O(N__58413),
            .I(N__58407));
    LocalMux I__7446 (
            .O(N__58410),
            .I(clk_en_157));
    LocalMux I__7445 (
            .O(N__58407),
            .I(clk_en_157));
    InMux I__7444 (
            .O(N__58402),
            .I(N__58399));
    LocalMux I__7443 (
            .O(N__58399),
            .I(shift_srl_155Z0Z_0));
    InMux I__7442 (
            .O(N__58396),
            .I(N__58393));
    LocalMux I__7441 (
            .O(N__58393),
            .I(shift_srl_155Z0Z_1));
    InMux I__7440 (
            .O(N__58390),
            .I(N__58387));
    LocalMux I__7439 (
            .O(N__58387),
            .I(shift_srl_25Z0Z_3));
    InMux I__7438 (
            .O(N__58384),
            .I(N__58381));
    LocalMux I__7437 (
            .O(N__58381),
            .I(shift_srl_25Z0Z_0));
    InMux I__7436 (
            .O(N__58378),
            .I(N__58375));
    LocalMux I__7435 (
            .O(N__58375),
            .I(shift_srl_25Z0Z_1));
    InMux I__7434 (
            .O(N__58372),
            .I(N__58369));
    LocalMux I__7433 (
            .O(N__58369),
            .I(shift_srl_25Z0Z_2));
    IoInMux I__7432 (
            .O(N__58366),
            .I(N__58363));
    LocalMux I__7431 (
            .O(N__58363),
            .I(N__58360));
    Span12Mux_s2_h I__7430 (
            .O(N__58360),
            .I(N__58356));
    InMux I__7429 (
            .O(N__58359),
            .I(N__58353));
    Odrv12 I__7428 (
            .O(N__58356),
            .I(rco_c_24));
    LocalMux I__7427 (
            .O(N__58353),
            .I(rco_c_24));
    InMux I__7426 (
            .O(N__58348),
            .I(N__58345));
    LocalMux I__7425 (
            .O(N__58345),
            .I(shift_srl_157Z0Z_0));
    InMux I__7424 (
            .O(N__58342),
            .I(N__58339));
    LocalMux I__7423 (
            .O(N__58339),
            .I(shift_srl_157Z0Z_1));
    InMux I__7422 (
            .O(N__58336),
            .I(N__58333));
    LocalMux I__7421 (
            .O(N__58333),
            .I(shift_srl_101Z0Z_3));
    InMux I__7420 (
            .O(N__58330),
            .I(N__58327));
    LocalMux I__7419 (
            .O(N__58327),
            .I(shift_srl_101Z0Z_4));
    InMux I__7418 (
            .O(N__58324),
            .I(N__58321));
    LocalMux I__7417 (
            .O(N__58321),
            .I(shift_srl_101Z0Z_5));
    InMux I__7416 (
            .O(N__58318),
            .I(N__58315));
    LocalMux I__7415 (
            .O(N__58315),
            .I(N__58312));
    Odrv4 I__7414 (
            .O(N__58312),
            .I(shift_srl_101Z0Z_6));
    InMux I__7413 (
            .O(N__58309),
            .I(N__58306));
    LocalMux I__7412 (
            .O(N__58306),
            .I(N__58303));
    Span4Mux_v I__7411 (
            .O(N__58303),
            .I(N__58300));
    Span4Mux_v I__7410 (
            .O(N__58300),
            .I(N__58297));
    Odrv4 I__7409 (
            .O(N__58297),
            .I(shift_srl_149_RNIU42SZ0Z_15));
    IoInMux I__7408 (
            .O(N__58294),
            .I(N__58291));
    LocalMux I__7407 (
            .O(N__58291),
            .I(N__58288));
    Span4Mux_s1_v I__7406 (
            .O(N__58288),
            .I(N__58285));
    Span4Mux_h I__7405 (
            .O(N__58285),
            .I(N__58282));
    Odrv4 I__7404 (
            .O(N__58282),
            .I(rco_c_149));
    InMux I__7403 (
            .O(N__58279),
            .I(N__58276));
    LocalMux I__7402 (
            .O(N__58276),
            .I(shift_srl_148Z0Z_6));
    InMux I__7401 (
            .O(N__58273),
            .I(N__58270));
    LocalMux I__7400 (
            .O(N__58270),
            .I(shift_srl_148Z0Z_7));
    InMux I__7399 (
            .O(N__58267),
            .I(N__58264));
    LocalMux I__7398 (
            .O(N__58264),
            .I(shift_srl_148Z0Z_2));
    InMux I__7397 (
            .O(N__58261),
            .I(N__58258));
    LocalMux I__7396 (
            .O(N__58258),
            .I(shift_srl_148Z0Z_3));
    InMux I__7395 (
            .O(N__58255),
            .I(N__58252));
    LocalMux I__7394 (
            .O(N__58252),
            .I(shift_srl_148Z0Z_4));
    InMux I__7393 (
            .O(N__58249),
            .I(N__58246));
    LocalMux I__7392 (
            .O(N__58246),
            .I(shift_srl_148Z0Z_5));
    CEMux I__7391 (
            .O(N__58243),
            .I(N__58240));
    LocalMux I__7390 (
            .O(N__58240),
            .I(N__58237));
    Span4Mux_v I__7389 (
            .O(N__58237),
            .I(N__58232));
    CEMux I__7388 (
            .O(N__58236),
            .I(N__58229));
    CEMux I__7387 (
            .O(N__58235),
            .I(N__58226));
    Span4Mux_h I__7386 (
            .O(N__58232),
            .I(N__58223));
    LocalMux I__7385 (
            .O(N__58229),
            .I(N__58220));
    LocalMux I__7384 (
            .O(N__58226),
            .I(N__58217));
    Odrv4 I__7383 (
            .O(N__58223),
            .I(clk_en_148));
    Odrv12 I__7382 (
            .O(N__58220),
            .I(clk_en_148));
    Odrv4 I__7381 (
            .O(N__58217),
            .I(clk_en_148));
    InMux I__7380 (
            .O(N__58210),
            .I(N__58207));
    LocalMux I__7379 (
            .O(N__58207),
            .I(shift_srl_101Z0Z_13));
    InMux I__7378 (
            .O(N__58204),
            .I(N__58201));
    LocalMux I__7377 (
            .O(N__58201),
            .I(shift_srl_101Z0Z_9));
    InMux I__7376 (
            .O(N__58198),
            .I(N__58195));
    LocalMux I__7375 (
            .O(N__58195),
            .I(shift_srl_101Z0Z_8));
    InMux I__7374 (
            .O(N__58192),
            .I(N__58189));
    LocalMux I__7373 (
            .O(N__58189),
            .I(shift_srl_101Z0Z_7));
    IoInMux I__7372 (
            .O(N__58186),
            .I(N__58183));
    LocalMux I__7371 (
            .O(N__58183),
            .I(N__58180));
    IoSpan4Mux I__7370 (
            .O(N__58180),
            .I(N__58177));
    Span4Mux_s3_v I__7369 (
            .O(N__58177),
            .I(N__58174));
    Odrv4 I__7368 (
            .O(N__58174),
            .I(rco_c_101));
    InMux I__7367 (
            .O(N__58171),
            .I(N__58168));
    LocalMux I__7366 (
            .O(N__58168),
            .I(shift_srl_101Z0Z_0));
    InMux I__7365 (
            .O(N__58165),
            .I(N__58162));
    LocalMux I__7364 (
            .O(N__58162),
            .I(shift_srl_101Z0Z_1));
    InMux I__7363 (
            .O(N__58159),
            .I(N__58156));
    LocalMux I__7362 (
            .O(N__58156),
            .I(shift_srl_101Z0Z_2));
    InMux I__7361 (
            .O(N__58153),
            .I(N__58150));
    LocalMux I__7360 (
            .O(N__58150),
            .I(shift_srl_104Z0Z_2));
    InMux I__7359 (
            .O(N__58147),
            .I(N__58144));
    LocalMux I__7358 (
            .O(N__58144),
            .I(shift_srl_104Z0Z_3));
    InMux I__7357 (
            .O(N__58141),
            .I(N__58138));
    LocalMux I__7356 (
            .O(N__58138),
            .I(shift_srl_104Z0Z_4));
    InMux I__7355 (
            .O(N__58135),
            .I(N__58132));
    LocalMux I__7354 (
            .O(N__58132),
            .I(shift_srl_104Z0Z_5));
    InMux I__7353 (
            .O(N__58129),
            .I(N__58126));
    LocalMux I__7352 (
            .O(N__58126),
            .I(shift_srl_104Z0Z_6));
    InMux I__7351 (
            .O(N__58123),
            .I(N__58120));
    LocalMux I__7350 (
            .O(N__58120),
            .I(shift_srl_101Z0Z_10));
    InMux I__7349 (
            .O(N__58117),
            .I(N__58114));
    LocalMux I__7348 (
            .O(N__58114),
            .I(shift_srl_101Z0Z_11));
    InMux I__7347 (
            .O(N__58111),
            .I(N__58108));
    LocalMux I__7346 (
            .O(N__58108),
            .I(shift_srl_101Z0Z_12));
    InMux I__7345 (
            .O(N__58105),
            .I(N__58102));
    LocalMux I__7344 (
            .O(N__58102),
            .I(shift_srl_105Z0Z_11));
    InMux I__7343 (
            .O(N__58099),
            .I(N__58096));
    LocalMux I__7342 (
            .O(N__58096),
            .I(shift_srl_105Z0Z_12));
    InMux I__7341 (
            .O(N__58093),
            .I(N__58090));
    LocalMux I__7340 (
            .O(N__58090),
            .I(shift_srl_105Z0Z_13));
    InMux I__7339 (
            .O(N__58087),
            .I(N__58084));
    LocalMux I__7338 (
            .O(N__58084),
            .I(shift_srl_105Z0Z_14));
    InMux I__7337 (
            .O(N__58081),
            .I(N__58078));
    LocalMux I__7336 (
            .O(N__58078),
            .I(shift_srl_105Z0Z_9));
    InMux I__7335 (
            .O(N__58075),
            .I(N__58072));
    LocalMux I__7334 (
            .O(N__58072),
            .I(N__58069));
    Odrv4 I__7333 (
            .O(N__58069),
            .I(shift_srl_105Z0Z_7));
    InMux I__7332 (
            .O(N__58066),
            .I(N__58063));
    LocalMux I__7331 (
            .O(N__58063),
            .I(shift_srl_105Z0Z_8));
    CEMux I__7330 (
            .O(N__58060),
            .I(N__58056));
    CEMux I__7329 (
            .O(N__58059),
            .I(N__58052));
    LocalMux I__7328 (
            .O(N__58056),
            .I(N__58049));
    CEMux I__7327 (
            .O(N__58055),
            .I(N__58046));
    LocalMux I__7326 (
            .O(N__58052),
            .I(N__58043));
    Span4Mux_v I__7325 (
            .O(N__58049),
            .I(N__58040));
    LocalMux I__7324 (
            .O(N__58046),
            .I(N__58037));
    Span4Mux_v I__7323 (
            .O(N__58043),
            .I(N__58034));
    Odrv4 I__7322 (
            .O(N__58040),
            .I(clk_en_105));
    Odrv12 I__7321 (
            .O(N__58037),
            .I(clk_en_105));
    Odrv4 I__7320 (
            .O(N__58034),
            .I(clk_en_105));
    InMux I__7319 (
            .O(N__58027),
            .I(N__58024));
    LocalMux I__7318 (
            .O(N__58024),
            .I(shift_srl_104Z0Z_0));
    InMux I__7317 (
            .O(N__58021),
            .I(N__58018));
    LocalMux I__7316 (
            .O(N__58018),
            .I(shift_srl_104Z0Z_1));
    InMux I__7315 (
            .O(N__58015),
            .I(N__58012));
    LocalMux I__7314 (
            .O(N__58012),
            .I(shift_srl_109Z0Z_6));
    InMux I__7313 (
            .O(N__58009),
            .I(N__58006));
    LocalMux I__7312 (
            .O(N__58006),
            .I(shift_srl_109Z0Z_7));
    CEMux I__7311 (
            .O(N__58003),
            .I(N__58000));
    LocalMux I__7310 (
            .O(N__58000),
            .I(N__57996));
    CEMux I__7309 (
            .O(N__57999),
            .I(N__57993));
    Span4Mux_h I__7308 (
            .O(N__57996),
            .I(N__57990));
    LocalMux I__7307 (
            .O(N__57993),
            .I(N__57987));
    Odrv4 I__7306 (
            .O(N__57990),
            .I(clk_en_109));
    Odrv12 I__7305 (
            .O(N__57987),
            .I(clk_en_109));
    IoInMux I__7304 (
            .O(N__57982),
            .I(N__57979));
    LocalMux I__7303 (
            .O(N__57979),
            .I(N__57976));
    Span4Mux_s3_v I__7302 (
            .O(N__57976),
            .I(N__57973));
    Span4Mux_v I__7301 (
            .O(N__57973),
            .I(N__57970));
    Odrv4 I__7300 (
            .O(N__57970),
            .I(rco_c_105));
    InMux I__7299 (
            .O(N__57967),
            .I(N__57964));
    LocalMux I__7298 (
            .O(N__57964),
            .I(shift_srl_105Z0Z_0));
    InMux I__7297 (
            .O(N__57961),
            .I(N__57958));
    LocalMux I__7296 (
            .O(N__57958),
            .I(shift_srl_105Z0Z_1));
    InMux I__7295 (
            .O(N__57955),
            .I(N__57952));
    LocalMux I__7294 (
            .O(N__57952),
            .I(shift_srl_105Z0Z_2));
    InMux I__7293 (
            .O(N__57949),
            .I(N__57946));
    LocalMux I__7292 (
            .O(N__57946),
            .I(shift_srl_105Z0Z_3));
    InMux I__7291 (
            .O(N__57943),
            .I(N__57940));
    LocalMux I__7290 (
            .O(N__57940),
            .I(N__57937));
    Span4Mux_v I__7289 (
            .O(N__57937),
            .I(N__57934));
    Odrv4 I__7288 (
            .O(N__57934),
            .I(shift_srl_105Z0Z_4));
    InMux I__7287 (
            .O(N__57931),
            .I(N__57928));
    LocalMux I__7286 (
            .O(N__57928),
            .I(shift_srl_105Z0Z_10));
    InMux I__7285 (
            .O(N__57925),
            .I(N__57922));
    LocalMux I__7284 (
            .O(N__57922),
            .I(shift_srl_109Z0Z_14));
    InMux I__7283 (
            .O(N__57919),
            .I(N__57916));
    LocalMux I__7282 (
            .O(N__57916),
            .I(shift_srl_109Z0Z_9));
    InMux I__7281 (
            .O(N__57913),
            .I(N__57910));
    LocalMux I__7280 (
            .O(N__57910),
            .I(shift_srl_109Z0Z_8));
    InMux I__7279 (
            .O(N__57907),
            .I(N__57904));
    LocalMux I__7278 (
            .O(N__57904),
            .I(shift_srl_109Z0Z_0));
    InMux I__7277 (
            .O(N__57901),
            .I(N__57898));
    LocalMux I__7276 (
            .O(N__57898),
            .I(shift_srl_109Z0Z_1));
    InMux I__7275 (
            .O(N__57895),
            .I(N__57892));
    LocalMux I__7274 (
            .O(N__57892),
            .I(shift_srl_109Z0Z_2));
    InMux I__7273 (
            .O(N__57889),
            .I(N__57886));
    LocalMux I__7272 (
            .O(N__57886),
            .I(shift_srl_109Z0Z_3));
    InMux I__7271 (
            .O(N__57883),
            .I(N__57880));
    LocalMux I__7270 (
            .O(N__57880),
            .I(shift_srl_109Z0Z_4));
    InMux I__7269 (
            .O(N__57877),
            .I(N__57874));
    LocalMux I__7268 (
            .O(N__57874),
            .I(shift_srl_109Z0Z_5));
    InMux I__7267 (
            .O(N__57871),
            .I(N__57868));
    LocalMux I__7266 (
            .O(N__57868),
            .I(shift_srl_112Z0Z_12));
    InMux I__7265 (
            .O(N__57865),
            .I(N__57862));
    LocalMux I__7264 (
            .O(N__57862),
            .I(shift_srl_112Z0Z_13));
    InMux I__7263 (
            .O(N__57859),
            .I(N__57856));
    LocalMux I__7262 (
            .O(N__57856),
            .I(shift_srl_112Z0Z_14));
    InMux I__7261 (
            .O(N__57853),
            .I(N__57850));
    LocalMux I__7260 (
            .O(N__57850),
            .I(shift_srl_112Z0Z_9));
    InMux I__7259 (
            .O(N__57847),
            .I(N__57844));
    LocalMux I__7258 (
            .O(N__57844),
            .I(N__57841));
    Odrv12 I__7257 (
            .O(N__57841),
            .I(shift_srl_112Z0Z_7));
    InMux I__7256 (
            .O(N__57838),
            .I(N__57835));
    LocalMux I__7255 (
            .O(N__57835),
            .I(shift_srl_112Z0Z_8));
    InMux I__7254 (
            .O(N__57832),
            .I(N__57829));
    LocalMux I__7253 (
            .O(N__57829),
            .I(shift_srl_109Z0Z_10));
    InMux I__7252 (
            .O(N__57826),
            .I(N__57823));
    LocalMux I__7251 (
            .O(N__57823),
            .I(shift_srl_109Z0Z_11));
    InMux I__7250 (
            .O(N__57820),
            .I(N__57817));
    LocalMux I__7249 (
            .O(N__57817),
            .I(shift_srl_109Z0Z_12));
    InMux I__7248 (
            .O(N__57814),
            .I(N__57811));
    LocalMux I__7247 (
            .O(N__57811),
            .I(shift_srl_109Z0Z_13));
    InMux I__7246 (
            .O(N__57808),
            .I(N__57805));
    LocalMux I__7245 (
            .O(N__57805),
            .I(shift_srl_113Z0Z_14));
    InMux I__7244 (
            .O(N__57802),
            .I(N__57799));
    LocalMux I__7243 (
            .O(N__57799),
            .I(shift_srl_113Z0Z_13));
    InMux I__7242 (
            .O(N__57796),
            .I(N__57793));
    LocalMux I__7241 (
            .O(N__57793),
            .I(shift_srl_113Z0Z_12));
    InMux I__7240 (
            .O(N__57790),
            .I(N__57787));
    LocalMux I__7239 (
            .O(N__57787),
            .I(shift_srl_113Z0Z_11));
    InMux I__7238 (
            .O(N__57784),
            .I(N__57781));
    LocalMux I__7237 (
            .O(N__57781),
            .I(shift_srl_113Z0Z_10));
    InMux I__7236 (
            .O(N__57778),
            .I(N__57775));
    LocalMux I__7235 (
            .O(N__57775),
            .I(N__57772));
    Span4Mux_v I__7234 (
            .O(N__57772),
            .I(N__57769));
    Odrv4 I__7233 (
            .O(N__57769),
            .I(shift_srl_113Z0Z_8));
    InMux I__7232 (
            .O(N__57766),
            .I(N__57763));
    LocalMux I__7231 (
            .O(N__57763),
            .I(shift_srl_113Z0Z_9));
    CEMux I__7230 (
            .O(N__57760),
            .I(N__57756));
    CEMux I__7229 (
            .O(N__57759),
            .I(N__57753));
    LocalMux I__7228 (
            .O(N__57756),
            .I(N__57749));
    LocalMux I__7227 (
            .O(N__57753),
            .I(N__57746));
    CEMux I__7226 (
            .O(N__57752),
            .I(N__57743));
    Span4Mux_h I__7225 (
            .O(N__57749),
            .I(N__57738));
    Span4Mux_v I__7224 (
            .O(N__57746),
            .I(N__57738));
    LocalMux I__7223 (
            .O(N__57743),
            .I(N__57735));
    Span4Mux_h I__7222 (
            .O(N__57738),
            .I(N__57732));
    Span4Mux_v I__7221 (
            .O(N__57735),
            .I(N__57729));
    Odrv4 I__7220 (
            .O(N__57732),
            .I(clk_en_113));
    Odrv4 I__7219 (
            .O(N__57729),
            .I(clk_en_113));
    InMux I__7218 (
            .O(N__57724),
            .I(N__57721));
    LocalMux I__7217 (
            .O(N__57721),
            .I(shift_srl_112Z0Z_10));
    InMux I__7216 (
            .O(N__57718),
            .I(N__57715));
    LocalMux I__7215 (
            .O(N__57715),
            .I(shift_srl_112Z0Z_11));
    InMux I__7214 (
            .O(N__57712),
            .I(N__57709));
    LocalMux I__7213 (
            .O(N__57709),
            .I(shift_srl_122Z0Z_10));
    InMux I__7212 (
            .O(N__57706),
            .I(N__57703));
    LocalMux I__7211 (
            .O(N__57703),
            .I(shift_srl_122Z0Z_11));
    InMux I__7210 (
            .O(N__57700),
            .I(N__57697));
    LocalMux I__7209 (
            .O(N__57697),
            .I(shift_srl_122Z0Z_12));
    InMux I__7208 (
            .O(N__57694),
            .I(N__57691));
    LocalMux I__7207 (
            .O(N__57691),
            .I(shift_srl_122Z0Z_13));
    InMux I__7206 (
            .O(N__57688),
            .I(N__57685));
    LocalMux I__7205 (
            .O(N__57685),
            .I(shift_srl_122Z0Z_14));
    InMux I__7204 (
            .O(N__57682),
            .I(N__57679));
    LocalMux I__7203 (
            .O(N__57679),
            .I(shift_srl_122Z0Z_9));
    InMux I__7202 (
            .O(N__57676),
            .I(N__57673));
    LocalMux I__7201 (
            .O(N__57673),
            .I(shift_srl_122Z0Z_8));
    InMux I__7200 (
            .O(N__57670),
            .I(N__57667));
    LocalMux I__7199 (
            .O(N__57667),
            .I(shift_srl_126Z0Z_5));
    InMux I__7198 (
            .O(N__57664),
            .I(N__57661));
    LocalMux I__7197 (
            .O(N__57661),
            .I(shift_srl_126Z0Z_6));
    InMux I__7196 (
            .O(N__57658),
            .I(N__57655));
    LocalMux I__7195 (
            .O(N__57655),
            .I(shift_srl_126Z0Z_13));
    InMux I__7194 (
            .O(N__57652),
            .I(N__57649));
    LocalMux I__7193 (
            .O(N__57649),
            .I(shift_srl_126Z0Z_14));
    IoInMux I__7192 (
            .O(N__57646),
            .I(N__57643));
    LocalMux I__7191 (
            .O(N__57643),
            .I(N__57640));
    IoSpan4Mux I__7190 (
            .O(N__57640),
            .I(N__57637));
    Span4Mux_s1_h I__7189 (
            .O(N__57637),
            .I(N__57634));
    Sp12to4 I__7188 (
            .O(N__57634),
            .I(N__57631));
    Span12Mux_s10_h I__7187 (
            .O(N__57631),
            .I(N__57628));
    Odrv12 I__7186 (
            .O(N__57628),
            .I(rco_c_126));
    IoInMux I__7185 (
            .O(N__57625),
            .I(N__57621));
    InMux I__7184 (
            .O(N__57624),
            .I(N__57618));
    LocalMux I__7183 (
            .O(N__57621),
            .I(N__57613));
    LocalMux I__7182 (
            .O(N__57618),
            .I(N__57609));
    InMux I__7181 (
            .O(N__57617),
            .I(N__57606));
    InMux I__7180 (
            .O(N__57616),
            .I(N__57602));
    Span4Mux_s3_h I__7179 (
            .O(N__57613),
            .I(N__57597));
    InMux I__7178 (
            .O(N__57612),
            .I(N__57594));
    Sp12to4 I__7177 (
            .O(N__57609),
            .I(N__57589));
    LocalMux I__7176 (
            .O(N__57606),
            .I(N__57589));
    InMux I__7175 (
            .O(N__57605),
            .I(N__57586));
    LocalMux I__7174 (
            .O(N__57602),
            .I(N__57583));
    InMux I__7173 (
            .O(N__57601),
            .I(N__57578));
    InMux I__7172 (
            .O(N__57600),
            .I(N__57578));
    Sp12to4 I__7171 (
            .O(N__57597),
            .I(N__57573));
    LocalMux I__7170 (
            .O(N__57594),
            .I(N__57570));
    Span12Mux_v I__7169 (
            .O(N__57589),
            .I(N__57561));
    LocalMux I__7168 (
            .O(N__57586),
            .I(N__57561));
    Span12Mux_s3_h I__7167 (
            .O(N__57583),
            .I(N__57561));
    LocalMux I__7166 (
            .O(N__57578),
            .I(N__57561));
    InMux I__7165 (
            .O(N__57577),
            .I(N__57556));
    InMux I__7164 (
            .O(N__57576),
            .I(N__57556));
    Odrv12 I__7163 (
            .O(N__57573),
            .I(rco_c_123));
    Odrv4 I__7162 (
            .O(N__57570),
            .I(rco_c_123));
    Odrv12 I__7161 (
            .O(N__57561),
            .I(rco_c_123));
    LocalMux I__7160 (
            .O(N__57556),
            .I(rco_c_123));
    CEMux I__7159 (
            .O(N__57547),
            .I(N__57543));
    CEMux I__7158 (
            .O(N__57546),
            .I(N__57540));
    LocalMux I__7157 (
            .O(N__57543),
            .I(clk_en_126));
    LocalMux I__7156 (
            .O(N__57540),
            .I(clk_en_126));
    InMux I__7155 (
            .O(N__57535),
            .I(N__57532));
    LocalMux I__7154 (
            .O(N__57532),
            .I(N__57529));
    Odrv4 I__7153 (
            .O(N__57529),
            .I(shift_srl_124Z0Z_14));
    CascadeMux I__7152 (
            .O(N__57526),
            .I(rco_int_0_a2_1_a2_0_127_cascade_));
    InMux I__7151 (
            .O(N__57523),
            .I(N__57520));
    LocalMux I__7150 (
            .O(N__57520),
            .I(N__57517));
    Odrv12 I__7149 (
            .O(N__57517),
            .I(rco_int_0_a2_0_a2_1_sx_sx_145));
    CascadeMux I__7148 (
            .O(N__57514),
            .I(rco_int_0_a2_0_a2_1_sx_145_cascade_));
    InMux I__7147 (
            .O(N__57511),
            .I(N__57508));
    LocalMux I__7146 (
            .O(N__57508),
            .I(shift_srl_124Z0Z_13));
    InMux I__7145 (
            .O(N__57505),
            .I(N__57502));
    LocalMux I__7144 (
            .O(N__57502),
            .I(shift_srl_124Z0Z_9));
    InMux I__7143 (
            .O(N__57499),
            .I(N__57496));
    LocalMux I__7142 (
            .O(N__57496),
            .I(shift_srl_124Z0Z_8));
    InMux I__7141 (
            .O(N__57493),
            .I(N__57490));
    LocalMux I__7140 (
            .O(N__57490),
            .I(shift_srl_126Z0Z_12));
    InMux I__7139 (
            .O(N__57487),
            .I(N__57484));
    LocalMux I__7138 (
            .O(N__57484),
            .I(shift_srl_126Z0Z_0));
    InMux I__7137 (
            .O(N__57481),
            .I(N__57478));
    LocalMux I__7136 (
            .O(N__57478),
            .I(shift_srl_126Z0Z_1));
    InMux I__7135 (
            .O(N__57475),
            .I(N__57472));
    LocalMux I__7134 (
            .O(N__57472),
            .I(shift_srl_126Z0Z_2));
    InMux I__7133 (
            .O(N__57469),
            .I(N__57466));
    LocalMux I__7132 (
            .O(N__57466),
            .I(shift_srl_126Z0Z_3));
    InMux I__7131 (
            .O(N__57463),
            .I(N__57460));
    LocalMux I__7130 (
            .O(N__57460),
            .I(shift_srl_126Z0Z_4));
    InMux I__7129 (
            .O(N__57457),
            .I(N__57454));
    LocalMux I__7128 (
            .O(N__57454),
            .I(shift_srl_161Z0Z_2));
    InMux I__7127 (
            .O(N__57451),
            .I(N__57448));
    LocalMux I__7126 (
            .O(N__57448),
            .I(shift_srl_161Z0Z_3));
    InMux I__7125 (
            .O(N__57445),
            .I(N__57442));
    LocalMux I__7124 (
            .O(N__57442),
            .I(shift_srl_161Z0Z_4));
    InMux I__7123 (
            .O(N__57439),
            .I(N__57436));
    LocalMux I__7122 (
            .O(N__57436),
            .I(shift_srl_161Z0Z_5));
    InMux I__7121 (
            .O(N__57433),
            .I(N__57430));
    LocalMux I__7120 (
            .O(N__57430),
            .I(shift_srl_161Z0Z_6));
    InMux I__7119 (
            .O(N__57427),
            .I(N__57424));
    LocalMux I__7118 (
            .O(N__57424),
            .I(shift_srl_161Z0Z_7));
    CEMux I__7117 (
            .O(N__57421),
            .I(N__57417));
    CEMux I__7116 (
            .O(N__57420),
            .I(N__57414));
    LocalMux I__7115 (
            .O(N__57417),
            .I(N__57411));
    LocalMux I__7114 (
            .O(N__57414),
            .I(N__57408));
    Span4Mux_h I__7113 (
            .O(N__57411),
            .I(N__57403));
    Span4Mux_h I__7112 (
            .O(N__57408),
            .I(N__57403));
    Odrv4 I__7111 (
            .O(N__57403),
            .I(clk_en_161));
    InMux I__7110 (
            .O(N__57400),
            .I(N__57397));
    LocalMux I__7109 (
            .O(N__57397),
            .I(shift_srl_124Z0Z_10));
    InMux I__7108 (
            .O(N__57394),
            .I(N__57391));
    LocalMux I__7107 (
            .O(N__57391),
            .I(shift_srl_124Z0Z_11));
    InMux I__7106 (
            .O(N__57388),
            .I(N__57385));
    LocalMux I__7105 (
            .O(N__57385),
            .I(shift_srl_124Z0Z_12));
    InMux I__7104 (
            .O(N__57382),
            .I(N__57379));
    LocalMux I__7103 (
            .O(N__57379),
            .I(shift_srl_154Z0Z_14));
    InMux I__7102 (
            .O(N__57376),
            .I(N__57373));
    LocalMux I__7101 (
            .O(N__57373),
            .I(shift_srl_154Z0Z_13));
    InMux I__7100 (
            .O(N__57370),
            .I(N__57367));
    LocalMux I__7099 (
            .O(N__57367),
            .I(N__57364));
    Odrv4 I__7098 (
            .O(N__57364),
            .I(shift_srl_154Z0Z_11));
    InMux I__7097 (
            .O(N__57361),
            .I(N__57358));
    LocalMux I__7096 (
            .O(N__57358),
            .I(shift_srl_154Z0Z_12));
    CEMux I__7095 (
            .O(N__57355),
            .I(N__57352));
    LocalMux I__7094 (
            .O(N__57352),
            .I(N__57349));
    Span4Mux_v I__7093 (
            .O(N__57349),
            .I(N__57345));
    CEMux I__7092 (
            .O(N__57348),
            .I(N__57342));
    Span4Mux_h I__7091 (
            .O(N__57345),
            .I(N__57335));
    LocalMux I__7090 (
            .O(N__57342),
            .I(N__57335));
    CEMux I__7089 (
            .O(N__57341),
            .I(N__57332));
    CEMux I__7088 (
            .O(N__57340),
            .I(N__57329));
    Span4Mux_h I__7087 (
            .O(N__57335),
            .I(N__57326));
    LocalMux I__7086 (
            .O(N__57332),
            .I(N__57321));
    LocalMux I__7085 (
            .O(N__57329),
            .I(N__57321));
    Odrv4 I__7084 (
            .O(N__57326),
            .I(clk_en_154));
    Odrv12 I__7083 (
            .O(N__57321),
            .I(clk_en_154));
    InMux I__7082 (
            .O(N__57316),
            .I(N__57313));
    LocalMux I__7081 (
            .O(N__57313),
            .I(shift_srl_161Z0Z_0));
    InMux I__7080 (
            .O(N__57310),
            .I(N__57307));
    LocalMux I__7079 (
            .O(N__57307),
            .I(shift_srl_161Z0Z_1));
    InMux I__7078 (
            .O(N__57304),
            .I(N__57301));
    LocalMux I__7077 (
            .O(N__57301),
            .I(shift_srl_157Z0Z_10));
    InMux I__7076 (
            .O(N__57298),
            .I(N__57295));
    LocalMux I__7075 (
            .O(N__57295),
            .I(shift_srl_157Z0Z_11));
    InMux I__7074 (
            .O(N__57292),
            .I(N__57289));
    LocalMux I__7073 (
            .O(N__57289),
            .I(shift_srl_157Z0Z_5));
    InMux I__7072 (
            .O(N__57286),
            .I(N__57283));
    LocalMux I__7071 (
            .O(N__57283),
            .I(shift_srl_157Z0Z_9));
    InMux I__7070 (
            .O(N__57280),
            .I(N__57277));
    LocalMux I__7069 (
            .O(N__57277),
            .I(shift_srl_157Z0Z_8));
    CEMux I__7068 (
            .O(N__57274),
            .I(N__57271));
    LocalMux I__7067 (
            .O(N__57271),
            .I(N__57267));
    CEMux I__7066 (
            .O(N__57270),
            .I(N__57264));
    Span4Mux_v I__7065 (
            .O(N__57267),
            .I(N__57261));
    LocalMux I__7064 (
            .O(N__57264),
            .I(N__57258));
    Span4Mux_h I__7063 (
            .O(N__57261),
            .I(N__57253));
    Span4Mux_v I__7062 (
            .O(N__57258),
            .I(N__57253));
    Odrv4 I__7061 (
            .O(N__57253),
            .I(clk_en_160));
    InMux I__7060 (
            .O(N__57250),
            .I(N__57247));
    LocalMux I__7059 (
            .O(N__57247),
            .I(N__57242));
    CEMux I__7058 (
            .O(N__57246),
            .I(N__57239));
    CEMux I__7057 (
            .O(N__57245),
            .I(N__57236));
    Span4Mux_v I__7056 (
            .O(N__57242),
            .I(N__57227));
    LocalMux I__7055 (
            .O(N__57239),
            .I(N__57227));
    LocalMux I__7054 (
            .O(N__57236),
            .I(N__57227));
    CEMux I__7053 (
            .O(N__57235),
            .I(N__57224));
    InMux I__7052 (
            .O(N__57234),
            .I(N__57221));
    Span4Mux_v I__7051 (
            .O(N__57227),
            .I(N__57213));
    LocalMux I__7050 (
            .O(N__57224),
            .I(N__57213));
    LocalMux I__7049 (
            .O(N__57221),
            .I(N__57210));
    InMux I__7048 (
            .O(N__57220),
            .I(N__57207));
    InMux I__7047 (
            .O(N__57219),
            .I(N__57202));
    InMux I__7046 (
            .O(N__57218),
            .I(N__57202));
    Span4Mux_v I__7045 (
            .O(N__57213),
            .I(N__57199));
    Span4Mux_h I__7044 (
            .O(N__57210),
            .I(N__57194));
    LocalMux I__7043 (
            .O(N__57207),
            .I(N__57194));
    LocalMux I__7042 (
            .O(N__57202),
            .I(N__57191));
    Sp12to4 I__7041 (
            .O(N__57199),
            .I(N__57188));
    Span4Mux_h I__7040 (
            .O(N__57194),
            .I(N__57185));
    Span12Mux_h I__7039 (
            .O(N__57191),
            .I(N__57182));
    Span12Mux_h I__7038 (
            .O(N__57188),
            .I(N__57179));
    Span4Mux_v I__7037 (
            .O(N__57185),
            .I(N__57176));
    Odrv12 I__7036 (
            .O(N__57182),
            .I(en_in_c));
    Odrv12 I__7035 (
            .O(N__57179),
            .I(en_in_c));
    Odrv4 I__7034 (
            .O(N__57176),
            .I(en_in_c));
    InMux I__7033 (
            .O(N__57169),
            .I(N__57166));
    LocalMux I__7032 (
            .O(N__57166),
            .I(N__57162));
    InMux I__7031 (
            .O(N__57165),
            .I(N__57159));
    Span4Mux_v I__7030 (
            .O(N__57162),
            .I(N__57154));
    LocalMux I__7029 (
            .O(N__57159),
            .I(N__57154));
    Span4Mux_h I__7028 (
            .O(N__57154),
            .I(N__57148));
    InMux I__7027 (
            .O(N__57153),
            .I(N__57145));
    InMux I__7026 (
            .O(N__57152),
            .I(N__57140));
    InMux I__7025 (
            .O(N__57151),
            .I(N__57140));
    Odrv4 I__7024 (
            .O(N__57148),
            .I(shift_srl_1Z0Z_15));
    LocalMux I__7023 (
            .O(N__57145),
            .I(shift_srl_1Z0Z_15));
    LocalMux I__7022 (
            .O(N__57140),
            .I(shift_srl_1Z0Z_15));
    IoInMux I__7021 (
            .O(N__57133),
            .I(N__57130));
    LocalMux I__7020 (
            .O(N__57130),
            .I(N__57127));
    IoSpan4Mux I__7019 (
            .O(N__57127),
            .I(N__57124));
    Span4Mux_s0_v I__7018 (
            .O(N__57124),
            .I(N__57121));
    Sp12to4 I__7017 (
            .O(N__57121),
            .I(N__57118));
    Span12Mux_s11_v I__7016 (
            .O(N__57118),
            .I(N__57115));
    Odrv12 I__7015 (
            .O(N__57115),
            .I(N_452_i));
    InMux I__7014 (
            .O(N__57112),
            .I(N__57109));
    LocalMux I__7013 (
            .O(N__57109),
            .I(shift_srl_154Z0Z_10));
    InMux I__7012 (
            .O(N__57106),
            .I(N__57103));
    LocalMux I__7011 (
            .O(N__57103),
            .I(shift_srl_154Z0Z_9));
    InMux I__7010 (
            .O(N__57100),
            .I(N__57097));
    LocalMux I__7009 (
            .O(N__57097),
            .I(shift_srl_154Z0Z_8));
    InMux I__7008 (
            .O(N__57094),
            .I(N__57091));
    LocalMux I__7007 (
            .O(N__57091),
            .I(shift_srl_154Z0Z_7));
    InMux I__7006 (
            .O(N__57088),
            .I(N__57085));
    LocalMux I__7005 (
            .O(N__57085),
            .I(shift_srl_154Z0Z_6));
    InMux I__7004 (
            .O(N__57082),
            .I(N__57079));
    LocalMux I__7003 (
            .O(N__57079),
            .I(shift_srl_154Z0Z_5));
    InMux I__7002 (
            .O(N__57076),
            .I(N__57073));
    LocalMux I__7001 (
            .O(N__57073),
            .I(N__57070));
    Span4Mux_v I__7000 (
            .O(N__57070),
            .I(N__57067));
    Odrv4 I__6999 (
            .O(N__57067),
            .I(shift_srl_154Z0Z_3));
    InMux I__6998 (
            .O(N__57064),
            .I(N__57061));
    LocalMux I__6997 (
            .O(N__57061),
            .I(shift_srl_154Z0Z_4));
    InMux I__6996 (
            .O(N__57058),
            .I(N__57055));
    LocalMux I__6995 (
            .O(N__57055),
            .I(shift_srl_148Z0Z_12));
    InMux I__6994 (
            .O(N__57052),
            .I(N__57049));
    LocalMux I__6993 (
            .O(N__57049),
            .I(shift_srl_148Z0Z_13));
    InMux I__6992 (
            .O(N__57046),
            .I(N__57043));
    LocalMux I__6991 (
            .O(N__57043),
            .I(shift_srl_148Z0Z_14));
    InMux I__6990 (
            .O(N__57040),
            .I(N__57037));
    LocalMux I__6989 (
            .O(N__57037),
            .I(shift_srl_148Z0Z_9));
    InMux I__6988 (
            .O(N__57034),
            .I(N__57031));
    LocalMux I__6987 (
            .O(N__57031),
            .I(shift_srl_148Z0Z_8));
    InMux I__6986 (
            .O(N__57028),
            .I(N__57020));
    InMux I__6985 (
            .O(N__57027),
            .I(N__57010));
    InMux I__6984 (
            .O(N__57026),
            .I(N__57010));
    InMux I__6983 (
            .O(N__57025),
            .I(N__57010));
    InMux I__6982 (
            .O(N__57024),
            .I(N__57010));
    InMux I__6981 (
            .O(N__57023),
            .I(N__57007));
    LocalMux I__6980 (
            .O(N__57020),
            .I(N__57004));
    InMux I__6979 (
            .O(N__57019),
            .I(N__57001));
    LocalMux I__6978 (
            .O(N__57010),
            .I(N__56998));
    LocalMux I__6977 (
            .O(N__57007),
            .I(shift_srl_147Z0Z_15));
    Odrv4 I__6976 (
            .O(N__57004),
            .I(shift_srl_147Z0Z_15));
    LocalMux I__6975 (
            .O(N__57001),
            .I(shift_srl_147Z0Z_15));
    Odrv12 I__6974 (
            .O(N__56998),
            .I(shift_srl_147Z0Z_15));
    CascadeMux I__6973 (
            .O(N__56989),
            .I(N__56986));
    InMux I__6972 (
            .O(N__56986),
            .I(N__56983));
    LocalMux I__6971 (
            .O(N__56983),
            .I(N__56977));
    InMux I__6970 (
            .O(N__56982),
            .I(N__56974));
    InMux I__6969 (
            .O(N__56981),
            .I(N__56969));
    InMux I__6968 (
            .O(N__56980),
            .I(N__56969));
    Sp12to4 I__6967 (
            .O(N__56977),
            .I(N__56961));
    LocalMux I__6966 (
            .O(N__56974),
            .I(N__56961));
    LocalMux I__6965 (
            .O(N__56969),
            .I(N__56961));
    InMux I__6964 (
            .O(N__56968),
            .I(N__56958));
    Span12Mux_v I__6963 (
            .O(N__56961),
            .I(N__56955));
    LocalMux I__6962 (
            .O(N__56958),
            .I(shift_srl_148Z0Z_15));
    Odrv12 I__6961 (
            .O(N__56955),
            .I(shift_srl_148Z0Z_15));
    InMux I__6960 (
            .O(N__56950),
            .I(N__56947));
    LocalMux I__6959 (
            .O(N__56947),
            .I(shift_srl_148Z0Z_0));
    InMux I__6958 (
            .O(N__56944),
            .I(N__56941));
    LocalMux I__6957 (
            .O(N__56941),
            .I(shift_srl_148Z0Z_1));
    InMux I__6956 (
            .O(N__56938),
            .I(N__56935));
    LocalMux I__6955 (
            .O(N__56935),
            .I(shift_srl_108Z0Z_7));
    InMux I__6954 (
            .O(N__56932),
            .I(N__56929));
    LocalMux I__6953 (
            .O(N__56929),
            .I(shift_srl_108Z0Z_8));
    CEMux I__6952 (
            .O(N__56926),
            .I(N__56922));
    CEMux I__6951 (
            .O(N__56925),
            .I(N__56918));
    LocalMux I__6950 (
            .O(N__56922),
            .I(N__56915));
    CEMux I__6949 (
            .O(N__56921),
            .I(N__56912));
    LocalMux I__6948 (
            .O(N__56918),
            .I(N__56909));
    Span4Mux_v I__6947 (
            .O(N__56915),
            .I(N__56906));
    LocalMux I__6946 (
            .O(N__56912),
            .I(N__56903));
    Span4Mux_h I__6945 (
            .O(N__56909),
            .I(N__56898));
    Span4Mux_h I__6944 (
            .O(N__56906),
            .I(N__56898));
    Span4Mux_h I__6943 (
            .O(N__56903),
            .I(N__56895));
    Odrv4 I__6942 (
            .O(N__56898),
            .I(clk_en_108));
    Odrv4 I__6941 (
            .O(N__56895),
            .I(clk_en_108));
    InMux I__6940 (
            .O(N__56890),
            .I(N__56887));
    LocalMux I__6939 (
            .O(N__56887),
            .I(shift_srl_0Z0Z_10));
    InMux I__6938 (
            .O(N__56884),
            .I(N__56881));
    LocalMux I__6937 (
            .O(N__56881),
            .I(shift_srl_0Z0Z_11));
    InMux I__6936 (
            .O(N__56878),
            .I(N__56875));
    LocalMux I__6935 (
            .O(N__56875),
            .I(shift_srl_0Z0Z_12));
    InMux I__6934 (
            .O(N__56872),
            .I(N__56869));
    LocalMux I__6933 (
            .O(N__56869),
            .I(shift_srl_0Z0Z_13));
    InMux I__6932 (
            .O(N__56866),
            .I(N__56863));
    LocalMux I__6931 (
            .O(N__56863),
            .I(shift_srl_0Z0Z_14));
    InMux I__6930 (
            .O(N__56860),
            .I(N__56857));
    LocalMux I__6929 (
            .O(N__56857),
            .I(shift_srl_148Z0Z_10));
    InMux I__6928 (
            .O(N__56854),
            .I(N__56851));
    LocalMux I__6927 (
            .O(N__56851),
            .I(shift_srl_148Z0Z_11));
    InMux I__6926 (
            .O(N__56848),
            .I(N__56845));
    LocalMux I__6925 (
            .O(N__56845),
            .I(shift_srl_108Z0Z_0));
    InMux I__6924 (
            .O(N__56842),
            .I(N__56839));
    LocalMux I__6923 (
            .O(N__56839),
            .I(shift_srl_108Z0Z_1));
    InMux I__6922 (
            .O(N__56836),
            .I(N__56833));
    LocalMux I__6921 (
            .O(N__56833),
            .I(shift_srl_108Z0Z_2));
    InMux I__6920 (
            .O(N__56830),
            .I(N__56827));
    LocalMux I__6919 (
            .O(N__56827),
            .I(shift_srl_108Z0Z_3));
    InMux I__6918 (
            .O(N__56824),
            .I(N__56821));
    LocalMux I__6917 (
            .O(N__56821),
            .I(shift_srl_108Z0Z_4));
    InMux I__6916 (
            .O(N__56818),
            .I(N__56815));
    LocalMux I__6915 (
            .O(N__56815),
            .I(shift_srl_108Z0Z_5));
    InMux I__6914 (
            .O(N__56812),
            .I(N__56809));
    LocalMux I__6913 (
            .O(N__56809),
            .I(shift_srl_108Z0Z_6));
    InMux I__6912 (
            .O(N__56806),
            .I(N__56803));
    LocalMux I__6911 (
            .O(N__56803),
            .I(shift_srl_108Z0Z_10));
    InMux I__6910 (
            .O(N__56800),
            .I(N__56797));
    LocalMux I__6909 (
            .O(N__56797),
            .I(N__56794));
    Span4Mux_v I__6908 (
            .O(N__56794),
            .I(N__56791));
    Odrv4 I__6907 (
            .O(N__56791),
            .I(shift_srl_108Z0Z_11));
    InMux I__6906 (
            .O(N__56788),
            .I(N__56785));
    LocalMux I__6905 (
            .O(N__56785),
            .I(shift_srl_108Z0Z_9));
    InMux I__6904 (
            .O(N__56782),
            .I(N__56779));
    LocalMux I__6903 (
            .O(N__56779),
            .I(shift_srl_106Z0Z_10));
    InMux I__6902 (
            .O(N__56776),
            .I(N__56773));
    LocalMux I__6901 (
            .O(N__56773),
            .I(shift_srl_106Z0Z_11));
    InMux I__6900 (
            .O(N__56770),
            .I(N__56767));
    LocalMux I__6899 (
            .O(N__56767),
            .I(shift_srl_106Z0Z_12));
    InMux I__6898 (
            .O(N__56764),
            .I(N__56761));
    LocalMux I__6897 (
            .O(N__56761),
            .I(shift_srl_106Z0Z_13));
    InMux I__6896 (
            .O(N__56758),
            .I(N__56755));
    LocalMux I__6895 (
            .O(N__56755),
            .I(shift_srl_106Z0Z_14));
    InMux I__6894 (
            .O(N__56752),
            .I(N__56749));
    LocalMux I__6893 (
            .O(N__56749),
            .I(shift_srl_106Z0Z_8));
    InMux I__6892 (
            .O(N__56746),
            .I(N__56743));
    LocalMux I__6891 (
            .O(N__56743),
            .I(shift_srl_106Z0Z_9));
    InMux I__6890 (
            .O(N__56740),
            .I(N__56737));
    LocalMux I__6889 (
            .O(N__56737),
            .I(shift_srl_106Z0Z_0));
    InMux I__6888 (
            .O(N__56734),
            .I(N__56731));
    LocalMux I__6887 (
            .O(N__56731),
            .I(shift_srl_106Z0Z_1));
    CEMux I__6886 (
            .O(N__56728),
            .I(N__56725));
    LocalMux I__6885 (
            .O(N__56725),
            .I(N__56721));
    CEMux I__6884 (
            .O(N__56724),
            .I(N__56718));
    Span4Mux_h I__6883 (
            .O(N__56721),
            .I(N__56713));
    LocalMux I__6882 (
            .O(N__56718),
            .I(N__56713));
    Span4Mux_h I__6881 (
            .O(N__56713),
            .I(N__56710));
    Odrv4 I__6880 (
            .O(N__56710),
            .I(clk_en_106));
    InMux I__6879 (
            .O(N__56707),
            .I(N__56704));
    LocalMux I__6878 (
            .O(N__56704),
            .I(N__56701));
    Odrv4 I__6877 (
            .O(N__56701),
            .I(shift_srl_107Z0Z_7));
    InMux I__6876 (
            .O(N__56698),
            .I(N__56695));
    LocalMux I__6875 (
            .O(N__56695),
            .I(shift_srl_107Z0Z_8));
    CEMux I__6874 (
            .O(N__56692),
            .I(N__56688));
    CEMux I__6873 (
            .O(N__56691),
            .I(N__56684));
    LocalMux I__6872 (
            .O(N__56688),
            .I(N__56680));
    CEMux I__6871 (
            .O(N__56687),
            .I(N__56677));
    LocalMux I__6870 (
            .O(N__56684),
            .I(N__56674));
    CEMux I__6869 (
            .O(N__56683),
            .I(N__56671));
    Span4Mux_v I__6868 (
            .O(N__56680),
            .I(N__56668));
    LocalMux I__6867 (
            .O(N__56677),
            .I(N__56665));
    Span4Mux_h I__6866 (
            .O(N__56674),
            .I(N__56660));
    LocalMux I__6865 (
            .O(N__56671),
            .I(N__56660));
    Span4Mux_h I__6864 (
            .O(N__56668),
            .I(N__56657));
    Span4Mux_h I__6863 (
            .O(N__56665),
            .I(N__56652));
    Span4Mux_v I__6862 (
            .O(N__56660),
            .I(N__56652));
    Odrv4 I__6861 (
            .O(N__56657),
            .I(clk_en_107));
    Odrv4 I__6860 (
            .O(N__56652),
            .I(clk_en_107));
    IoInMux I__6859 (
            .O(N__56647),
            .I(N__56644));
    LocalMux I__6858 (
            .O(N__56644),
            .I(N__56641));
    Span4Mux_s0_v I__6857 (
            .O(N__56641),
            .I(N__56638));
    Span4Mux_v I__6856 (
            .O(N__56638),
            .I(N__56635));
    Sp12to4 I__6855 (
            .O(N__56635),
            .I(N__56630));
    InMux I__6854 (
            .O(N__56634),
            .I(N__56625));
    InMux I__6853 (
            .O(N__56633),
            .I(N__56625));
    Span12Mux_s10_h I__6852 (
            .O(N__56630),
            .I(N__56622));
    LocalMux I__6851 (
            .O(N__56625),
            .I(N__56619));
    Span12Mux_h I__6850 (
            .O(N__56622),
            .I(N__56616));
    Span4Mux_s3_v I__6849 (
            .O(N__56619),
            .I(N__56613));
    Odrv12 I__6848 (
            .O(N__56616),
            .I(rco_c_106));
    Odrv4 I__6847 (
            .O(N__56613),
            .I(rco_c_106));
    InMux I__6846 (
            .O(N__56608),
            .I(N__56605));
    LocalMux I__6845 (
            .O(N__56605),
            .I(shift_srl_106_RNIPC6S1Z0Z_15));
    CascadeMux I__6844 (
            .O(N__56602),
            .I(shift_srl_106_RNIPC6S1Z0Z_15_cascade_));
    CascadeMux I__6843 (
            .O(N__56599),
            .I(rco_int_0_a3_0_a2_out_0_cascade_));
    CascadeMux I__6842 (
            .O(N__56596),
            .I(N__56593));
    InMux I__6841 (
            .O(N__56593),
            .I(N__56590));
    LocalMux I__6840 (
            .O(N__56590),
            .I(N__56587));
    Odrv12 I__6839 (
            .O(N__56587),
            .I(clk_en_0_a3_0_a2_sx_109));
    InMux I__6838 (
            .O(N__56584),
            .I(N__56581));
    LocalMux I__6837 (
            .O(N__56581),
            .I(shift_srl_110Z0Z_8));
    InMux I__6836 (
            .O(N__56578),
            .I(N__56575));
    LocalMux I__6835 (
            .O(N__56575),
            .I(shift_srl_110Z0Z_6));
    InMux I__6834 (
            .O(N__56572),
            .I(N__56569));
    LocalMux I__6833 (
            .O(N__56569),
            .I(shift_srl_110Z0Z_7));
    InMux I__6832 (
            .O(N__56566),
            .I(N__56563));
    LocalMux I__6831 (
            .O(N__56563),
            .I(shift_srl_107Z0Z_10));
    InMux I__6830 (
            .O(N__56560),
            .I(N__56557));
    LocalMux I__6829 (
            .O(N__56557),
            .I(shift_srl_107Z0Z_11));
    InMux I__6828 (
            .O(N__56554),
            .I(N__56551));
    LocalMux I__6827 (
            .O(N__56551),
            .I(shift_srl_107Z0Z_12));
    InMux I__6826 (
            .O(N__56548),
            .I(N__56545));
    LocalMux I__6825 (
            .O(N__56545),
            .I(shift_srl_107Z0Z_13));
    InMux I__6824 (
            .O(N__56542),
            .I(N__56539));
    LocalMux I__6823 (
            .O(N__56539),
            .I(shift_srl_107Z0Z_14));
    InMux I__6822 (
            .O(N__56536),
            .I(N__56533));
    LocalMux I__6821 (
            .O(N__56533),
            .I(shift_srl_107Z0Z_9));
    InMux I__6820 (
            .O(N__56530),
            .I(N__56527));
    LocalMux I__6819 (
            .O(N__56527),
            .I(shift_srl_108Z0Z_14));
    InMux I__6818 (
            .O(N__56524),
            .I(N__56521));
    LocalMux I__6817 (
            .O(N__56521),
            .I(shift_srl_108Z0Z_13));
    InMux I__6816 (
            .O(N__56518),
            .I(N__56515));
    LocalMux I__6815 (
            .O(N__56515),
            .I(shift_srl_108Z0Z_12));
    InMux I__6814 (
            .O(N__56512),
            .I(N__56509));
    LocalMux I__6813 (
            .O(N__56509),
            .I(shift_srl_110Z0Z_0));
    InMux I__6812 (
            .O(N__56506),
            .I(N__56503));
    LocalMux I__6811 (
            .O(N__56503),
            .I(shift_srl_110Z0Z_1));
    InMux I__6810 (
            .O(N__56500),
            .I(N__56497));
    LocalMux I__6809 (
            .O(N__56497),
            .I(shift_srl_110Z0Z_2));
    InMux I__6808 (
            .O(N__56494),
            .I(N__56491));
    LocalMux I__6807 (
            .O(N__56491),
            .I(shift_srl_110Z0Z_3));
    InMux I__6806 (
            .O(N__56488),
            .I(N__56485));
    LocalMux I__6805 (
            .O(N__56485),
            .I(shift_srl_110Z0Z_4));
    InMux I__6804 (
            .O(N__56482),
            .I(N__56479));
    LocalMux I__6803 (
            .O(N__56479),
            .I(shift_srl_110Z0Z_5));
    CascadeMux I__6802 (
            .O(N__56476),
            .I(g0_9_1_cascade_));
    InMux I__6801 (
            .O(N__56473),
            .I(N__56470));
    LocalMux I__6800 (
            .O(N__56470),
            .I(N__56467));
    Span4Mux_h I__6799 (
            .O(N__56467),
            .I(N__56464));
    Span4Mux_h I__6798 (
            .O(N__56464),
            .I(N__56461));
    Odrv4 I__6797 (
            .O(N__56461),
            .I(g0_14));
    InMux I__6796 (
            .O(N__56458),
            .I(N__56455));
    LocalMux I__6795 (
            .O(N__56455),
            .I(N__56452));
    Span4Mux_v I__6794 (
            .O(N__56452),
            .I(N__56449));
    Sp12to4 I__6793 (
            .O(N__56449),
            .I(N__56446));
    Odrv12 I__6792 (
            .O(N__56446),
            .I(g0_9_0));
    InMux I__6791 (
            .O(N__56443),
            .I(N__56440));
    LocalMux I__6790 (
            .O(N__56440),
            .I(N__56437));
    Span4Mux_h I__6789 (
            .O(N__56437),
            .I(N__56434));
    Odrv4 I__6788 (
            .O(N__56434),
            .I(g0_8_2));
    CascadeMux I__6787 (
            .O(N__56431),
            .I(clk_en_0_a3_0_a2_sx_110_cascade_));
    InMux I__6786 (
            .O(N__56428),
            .I(N__56425));
    LocalMux I__6785 (
            .O(N__56425),
            .I(clk_en_0_a3_0_a2_1_110));
    InMux I__6784 (
            .O(N__56422),
            .I(N__56419));
    LocalMux I__6783 (
            .O(N__56419),
            .I(shift_srl_125Z0Z_10));
    InMux I__6782 (
            .O(N__56416),
            .I(N__56413));
    LocalMux I__6781 (
            .O(N__56413),
            .I(shift_srl_125Z0Z_11));
    InMux I__6780 (
            .O(N__56410),
            .I(N__56407));
    LocalMux I__6779 (
            .O(N__56407),
            .I(shift_srl_125Z0Z_12));
    InMux I__6778 (
            .O(N__56404),
            .I(N__56401));
    LocalMux I__6777 (
            .O(N__56401),
            .I(shift_srl_125Z0Z_13));
    InMux I__6776 (
            .O(N__56398),
            .I(N__56395));
    LocalMux I__6775 (
            .O(N__56395),
            .I(shift_srl_125Z0Z_14));
    InMux I__6774 (
            .O(N__56392),
            .I(N__56389));
    LocalMux I__6773 (
            .O(N__56389),
            .I(shift_srl_125Z0Z_9));
    InMux I__6772 (
            .O(N__56386),
            .I(N__56383));
    LocalMux I__6771 (
            .O(N__56383),
            .I(shift_srl_125Z0Z_7));
    InMux I__6770 (
            .O(N__56380),
            .I(N__56377));
    LocalMux I__6769 (
            .O(N__56377),
            .I(shift_srl_125Z0Z_8));
    CEMux I__6768 (
            .O(N__56374),
            .I(N__56370));
    CEMux I__6767 (
            .O(N__56373),
            .I(N__56367));
    LocalMux I__6766 (
            .O(N__56370),
            .I(N__56364));
    LocalMux I__6765 (
            .O(N__56367),
            .I(N__56361));
    Span4Mux_v I__6764 (
            .O(N__56364),
            .I(N__56358));
    Span4Mux_v I__6763 (
            .O(N__56361),
            .I(N__56355));
    Span4Mux_h I__6762 (
            .O(N__56358),
            .I(N__56352));
    Span4Mux_h I__6761 (
            .O(N__56355),
            .I(N__56349));
    Odrv4 I__6760 (
            .O(N__56352),
            .I(clk_en_125));
    Odrv4 I__6759 (
            .O(N__56349),
            .I(clk_en_125));
    InMux I__6758 (
            .O(N__56344),
            .I(N__56341));
    LocalMux I__6757 (
            .O(N__56341),
            .I(shift_srl_121Z0Z_10));
    InMux I__6756 (
            .O(N__56338),
            .I(N__56335));
    LocalMux I__6755 (
            .O(N__56335),
            .I(shift_srl_121Z0Z_11));
    InMux I__6754 (
            .O(N__56332),
            .I(N__56329));
    LocalMux I__6753 (
            .O(N__56329),
            .I(shift_srl_121Z0Z_12));
    InMux I__6752 (
            .O(N__56326),
            .I(N__56323));
    LocalMux I__6751 (
            .O(N__56323),
            .I(shift_srl_121Z0Z_13));
    InMux I__6750 (
            .O(N__56320),
            .I(N__56317));
    LocalMux I__6749 (
            .O(N__56317),
            .I(shift_srl_121Z0Z_14));
    InMux I__6748 (
            .O(N__56314),
            .I(N__56311));
    LocalMux I__6747 (
            .O(N__56311),
            .I(shift_srl_121Z0Z_9));
    InMux I__6746 (
            .O(N__56308),
            .I(N__56305));
    LocalMux I__6745 (
            .O(N__56305),
            .I(shift_srl_121Z0Z_8));
    InMux I__6744 (
            .O(N__56302),
            .I(N__56299));
    LocalMux I__6743 (
            .O(N__56299),
            .I(shift_srl_126Z0Z_9));
    InMux I__6742 (
            .O(N__56296),
            .I(N__56293));
    LocalMux I__6741 (
            .O(N__56293),
            .I(shift_srl_126Z0Z_7));
    InMux I__6740 (
            .O(N__56290),
            .I(N__56287));
    LocalMux I__6739 (
            .O(N__56287),
            .I(shift_srl_126Z0Z_8));
    CascadeMux I__6738 (
            .O(N__56284),
            .I(clk_en_0_a2_0_a2_sx_128_cascade_));
    CEMux I__6737 (
            .O(N__56281),
            .I(N__56276));
    CEMux I__6736 (
            .O(N__56280),
            .I(N__56273));
    CEMux I__6735 (
            .O(N__56279),
            .I(N__56270));
    LocalMux I__6734 (
            .O(N__56276),
            .I(N__56267));
    LocalMux I__6733 (
            .O(N__56273),
            .I(N__56264));
    LocalMux I__6732 (
            .O(N__56270),
            .I(N__56261));
    Span4Mux_h I__6731 (
            .O(N__56267),
            .I(N__56258));
    Span4Mux_v I__6730 (
            .O(N__56264),
            .I(N__56253));
    Span4Mux_h I__6729 (
            .O(N__56261),
            .I(N__56253));
    Odrv4 I__6728 (
            .O(N__56258),
            .I(clk_en_128));
    Odrv4 I__6727 (
            .O(N__56253),
            .I(clk_en_128));
    InMux I__6726 (
            .O(N__56248),
            .I(N__56245));
    LocalMux I__6725 (
            .O(N__56245),
            .I(N__56242));
    Odrv4 I__6724 (
            .O(N__56242),
            .I(shift_srl_123Z0Z_14));
    InMux I__6723 (
            .O(N__56239),
            .I(N__56233));
    InMux I__6722 (
            .O(N__56238),
            .I(N__56233));
    LocalMux I__6721 (
            .O(N__56233),
            .I(shift_srl_123Z0Z_15));
    InMux I__6720 (
            .O(N__56230),
            .I(N__56227));
    LocalMux I__6719 (
            .O(N__56227),
            .I(shift_srl_123Z0Z_0));
    InMux I__6718 (
            .O(N__56224),
            .I(N__56221));
    LocalMux I__6717 (
            .O(N__56221),
            .I(shift_srl_123Z0Z_1));
    InMux I__6716 (
            .O(N__56218),
            .I(N__56215));
    LocalMux I__6715 (
            .O(N__56215),
            .I(N__56212));
    Span4Mux_v I__6714 (
            .O(N__56212),
            .I(N__56209));
    Odrv4 I__6713 (
            .O(N__56209),
            .I(shift_srl_123Z0Z_2));
    CEMux I__6712 (
            .O(N__56206),
            .I(N__56202));
    CEMux I__6711 (
            .O(N__56205),
            .I(N__56199));
    LocalMux I__6710 (
            .O(N__56202),
            .I(N__56195));
    LocalMux I__6709 (
            .O(N__56199),
            .I(N__56192));
    CEMux I__6708 (
            .O(N__56198),
            .I(N__56189));
    Span4Mux_v I__6707 (
            .O(N__56195),
            .I(N__56186));
    Span4Mux_v I__6706 (
            .O(N__56192),
            .I(N__56183));
    LocalMux I__6705 (
            .O(N__56189),
            .I(N__56180));
    Span4Mux_h I__6704 (
            .O(N__56186),
            .I(N__56175));
    Span4Mux_h I__6703 (
            .O(N__56183),
            .I(N__56175));
    Span4Mux_v I__6702 (
            .O(N__56180),
            .I(N__56172));
    Odrv4 I__6701 (
            .O(N__56175),
            .I(clk_en_123));
    Odrv4 I__6700 (
            .O(N__56172),
            .I(clk_en_123));
    InMux I__6699 (
            .O(N__56167),
            .I(N__56164));
    LocalMux I__6698 (
            .O(N__56164),
            .I(N__56161));
    Odrv4 I__6697 (
            .O(N__56161),
            .I(shift_srl_146Z0Z_14));
    CEMux I__6696 (
            .O(N__56158),
            .I(N__56154));
    CEMux I__6695 (
            .O(N__56157),
            .I(N__56150));
    LocalMux I__6694 (
            .O(N__56154),
            .I(N__56147));
    CEMux I__6693 (
            .O(N__56153),
            .I(N__56144));
    LocalMux I__6692 (
            .O(N__56150),
            .I(N__56141));
    Span4Mux_h I__6691 (
            .O(N__56147),
            .I(N__56135));
    LocalMux I__6690 (
            .O(N__56144),
            .I(N__56135));
    Span4Mux_h I__6689 (
            .O(N__56141),
            .I(N__56132));
    CEMux I__6688 (
            .O(N__56140),
            .I(N__56129));
    Span4Mux_v I__6687 (
            .O(N__56135),
            .I(N__56122));
    Span4Mux_h I__6686 (
            .O(N__56132),
            .I(N__56122));
    LocalMux I__6685 (
            .O(N__56129),
            .I(N__56122));
    Odrv4 I__6684 (
            .O(N__56122),
            .I(clk_en_146));
    InMux I__6683 (
            .O(N__56119),
            .I(N__56116));
    LocalMux I__6682 (
            .O(N__56116),
            .I(N__56112));
    InMux I__6681 (
            .O(N__56115),
            .I(N__56108));
    Span4Mux_v I__6680 (
            .O(N__56112),
            .I(N__56105));
    InMux I__6679 (
            .O(N__56111),
            .I(N__56102));
    LocalMux I__6678 (
            .O(N__56108),
            .I(shift_srl_149Z0Z_15));
    Odrv4 I__6677 (
            .O(N__56105),
            .I(shift_srl_149Z0Z_15));
    LocalMux I__6676 (
            .O(N__56102),
            .I(shift_srl_149Z0Z_15));
    CascadeMux I__6675 (
            .O(N__56095),
            .I(N__56092));
    InMux I__6674 (
            .O(N__56092),
            .I(N__56089));
    LocalMux I__6673 (
            .O(N__56089),
            .I(N__56085));
    InMux I__6672 (
            .O(N__56088),
            .I(N__56082));
    Span4Mux_v I__6671 (
            .O(N__56085),
            .I(N__56079));
    LocalMux I__6670 (
            .O(N__56082),
            .I(shift_srl_150Z0Z_15));
    Odrv4 I__6669 (
            .O(N__56079),
            .I(shift_srl_150Z0Z_15));
    CascadeMux I__6668 (
            .O(N__56074),
            .I(shift_srl_150_RNIPH7TZ0Z_15_cascade_));
    CascadeMux I__6667 (
            .O(N__56071),
            .I(shift_srl_146_RNIVSUTZ0Z_15_cascade_));
    InMux I__6666 (
            .O(N__56068),
            .I(N__56065));
    LocalMux I__6665 (
            .O(N__56065),
            .I(shift_srl_126Z0Z_10));
    InMux I__6664 (
            .O(N__56062),
            .I(N__56059));
    LocalMux I__6663 (
            .O(N__56059),
            .I(shift_srl_126Z0Z_11));
    InMux I__6662 (
            .O(N__56056),
            .I(N__56053));
    LocalMux I__6661 (
            .O(N__56053),
            .I(shift_srl_161Z0Z_12));
    InMux I__6660 (
            .O(N__56050),
            .I(N__56047));
    LocalMux I__6659 (
            .O(N__56047),
            .I(shift_srl_161Z0Z_13));
    InMux I__6658 (
            .O(N__56044),
            .I(N__56041));
    LocalMux I__6657 (
            .O(N__56041),
            .I(shift_srl_161Z0Z_14));
    InMux I__6656 (
            .O(N__56038),
            .I(N__56035));
    LocalMux I__6655 (
            .O(N__56035),
            .I(shift_srl_161Z0Z_9));
    InMux I__6654 (
            .O(N__56032),
            .I(N__56029));
    LocalMux I__6653 (
            .O(N__56029),
            .I(shift_srl_161Z0Z_8));
    IoInMux I__6652 (
            .O(N__56026),
            .I(N__56023));
    LocalMux I__6651 (
            .O(N__56023),
            .I(N__56020));
    IoSpan4Mux I__6650 (
            .O(N__56020),
            .I(N__56017));
    Span4Mux_s1_h I__6649 (
            .O(N__56017),
            .I(N__56014));
    Span4Mux_h I__6648 (
            .O(N__56014),
            .I(N__56011));
    Sp12to4 I__6647 (
            .O(N__56011),
            .I(N__56008));
    Span12Mux_v I__6646 (
            .O(N__56008),
            .I(N__56005));
    Odrv12 I__6645 (
            .O(N__56005),
            .I(rco_c_148));
    IoInMux I__6644 (
            .O(N__56002),
            .I(N__55999));
    LocalMux I__6643 (
            .O(N__55999),
            .I(N__55996));
    Span4Mux_s0_h I__6642 (
            .O(N__55996),
            .I(N__55993));
    Span4Mux_h I__6641 (
            .O(N__55993),
            .I(N__55990));
    Sp12to4 I__6640 (
            .O(N__55990),
            .I(N__55987));
    Span12Mux_v I__6639 (
            .O(N__55987),
            .I(N__55984));
    Odrv12 I__6638 (
            .O(N__55984),
            .I(rco_c_147));
    CascadeMux I__6637 (
            .O(N__55981),
            .I(clk_en_0_a3_0_a2_sx_149_cascade_));
    CEMux I__6636 (
            .O(N__55978),
            .I(N__55974));
    CEMux I__6635 (
            .O(N__55977),
            .I(N__55971));
    LocalMux I__6634 (
            .O(N__55974),
            .I(clk_en_149));
    LocalMux I__6633 (
            .O(N__55971),
            .I(clk_en_149));
    InMux I__6632 (
            .O(N__55966),
            .I(N__55963));
    LocalMux I__6631 (
            .O(N__55963),
            .I(shift_srl_160Z0Z_7));
    InMux I__6630 (
            .O(N__55960),
            .I(N__55957));
    LocalMux I__6629 (
            .O(N__55957),
            .I(shift_srl_160Z0Z_0));
    InMux I__6628 (
            .O(N__55954),
            .I(N__55951));
    LocalMux I__6627 (
            .O(N__55951),
            .I(shift_srl_160Z0Z_11));
    InMux I__6626 (
            .O(N__55948),
            .I(N__55945));
    LocalMux I__6625 (
            .O(N__55945),
            .I(shift_srl_160Z0Z_4));
    InMux I__6624 (
            .O(N__55942),
            .I(N__55939));
    LocalMux I__6623 (
            .O(N__55939),
            .I(shift_srl_160Z0Z_5));
    InMux I__6622 (
            .O(N__55936),
            .I(N__55933));
    LocalMux I__6621 (
            .O(N__55933),
            .I(shift_srl_160Z0Z_6));
    InMux I__6620 (
            .O(N__55930),
            .I(N__55927));
    LocalMux I__6619 (
            .O(N__55927),
            .I(shift_srl_160Z0Z_12));
    InMux I__6618 (
            .O(N__55924),
            .I(N__55921));
    LocalMux I__6617 (
            .O(N__55921),
            .I(shift_srl_160Z0Z_13));
    InMux I__6616 (
            .O(N__55918),
            .I(N__55915));
    LocalMux I__6615 (
            .O(N__55915),
            .I(shift_srl_161Z0Z_10));
    InMux I__6614 (
            .O(N__55912),
            .I(N__55909));
    LocalMux I__6613 (
            .O(N__55909),
            .I(shift_srl_161Z0Z_11));
    InMux I__6612 (
            .O(N__55906),
            .I(N__55903));
    LocalMux I__6611 (
            .O(N__55903),
            .I(shift_srl_160Z0Z_10));
    InMux I__6610 (
            .O(N__55900),
            .I(N__55897));
    LocalMux I__6609 (
            .O(N__55897),
            .I(shift_srl_160Z0Z_3));
    InMux I__6608 (
            .O(N__55894),
            .I(N__55891));
    LocalMux I__6607 (
            .O(N__55891),
            .I(shift_srl_160Z0Z_1));
    InMux I__6606 (
            .O(N__55888),
            .I(N__55885));
    LocalMux I__6605 (
            .O(N__55885),
            .I(shift_srl_160Z0Z_2));
    InMux I__6604 (
            .O(N__55882),
            .I(N__55879));
    LocalMux I__6603 (
            .O(N__55879),
            .I(shift_srl_160Z0Z_9));
    InMux I__6602 (
            .O(N__55876),
            .I(N__55873));
    LocalMux I__6601 (
            .O(N__55873),
            .I(shift_srl_160Z0Z_8));
    InMux I__6600 (
            .O(N__55870),
            .I(N__55867));
    LocalMux I__6599 (
            .O(N__55867),
            .I(shift_srl_160Z0Z_14));
    InMux I__6598 (
            .O(N__55864),
            .I(N__55861));
    LocalMux I__6597 (
            .O(N__55861),
            .I(shift_srl_147Z0Z_4));
    InMux I__6596 (
            .O(N__55858),
            .I(N__55855));
    LocalMux I__6595 (
            .O(N__55855),
            .I(shift_srl_147Z0Z_9));
    InMux I__6594 (
            .O(N__55852),
            .I(N__55849));
    LocalMux I__6593 (
            .O(N__55849),
            .I(shift_srl_147Z0Z_7));
    InMux I__6592 (
            .O(N__55846),
            .I(N__55843));
    LocalMux I__6591 (
            .O(N__55843),
            .I(shift_srl_147Z0Z_8));
    CEMux I__6590 (
            .O(N__55840),
            .I(N__55837));
    LocalMux I__6589 (
            .O(N__55837),
            .I(N__55833));
    CEMux I__6588 (
            .O(N__55836),
            .I(N__55829));
    Sp12to4 I__6587 (
            .O(N__55833),
            .I(N__55826));
    CEMux I__6586 (
            .O(N__55832),
            .I(N__55823));
    LocalMux I__6585 (
            .O(N__55829),
            .I(clk_en_147));
    Odrv12 I__6584 (
            .O(N__55826),
            .I(clk_en_147));
    LocalMux I__6583 (
            .O(N__55823),
            .I(clk_en_147));
    InMux I__6582 (
            .O(N__55816),
            .I(N__55813));
    LocalMux I__6581 (
            .O(N__55813),
            .I(shift_srl_146Z0Z_0));
    InMux I__6580 (
            .O(N__55810),
            .I(N__55807));
    LocalMux I__6579 (
            .O(N__55807),
            .I(shift_srl_146Z0Z_1));
    InMux I__6578 (
            .O(N__55804),
            .I(N__55801));
    LocalMux I__6577 (
            .O(N__55801),
            .I(shift_srl_146Z0Z_2));
    InMux I__6576 (
            .O(N__55798),
            .I(N__55795));
    LocalMux I__6575 (
            .O(N__55795),
            .I(shift_srl_147Z0Z_14));
    InMux I__6574 (
            .O(N__55792),
            .I(N__55789));
    LocalMux I__6573 (
            .O(N__55789),
            .I(shift_srl_147Z0Z_13));
    InMux I__6572 (
            .O(N__55786),
            .I(N__55783));
    LocalMux I__6571 (
            .O(N__55783),
            .I(shift_srl_147Z0Z_12));
    InMux I__6570 (
            .O(N__55780),
            .I(N__55777));
    LocalMux I__6569 (
            .O(N__55777),
            .I(shift_srl_147Z0Z_11));
    InMux I__6568 (
            .O(N__55774),
            .I(N__55771));
    LocalMux I__6567 (
            .O(N__55771),
            .I(shift_srl_147Z0Z_10));
    InMux I__6566 (
            .O(N__55768),
            .I(N__55765));
    LocalMux I__6565 (
            .O(N__55765),
            .I(shift_srl_147Z0Z_0));
    InMux I__6564 (
            .O(N__55762),
            .I(N__55759));
    LocalMux I__6563 (
            .O(N__55759),
            .I(shift_srl_147Z0Z_1));
    InMux I__6562 (
            .O(N__55756),
            .I(N__55753));
    LocalMux I__6561 (
            .O(N__55753),
            .I(shift_srl_147Z0Z_2));
    InMux I__6560 (
            .O(N__55750),
            .I(N__55747));
    LocalMux I__6559 (
            .O(N__55747),
            .I(shift_srl_147Z0Z_3));
    InMux I__6558 (
            .O(N__55744),
            .I(N__55741));
    LocalMux I__6557 (
            .O(N__55741),
            .I(shift_srl_10Z0Z_5));
    InMux I__6556 (
            .O(N__55738),
            .I(N__55735));
    LocalMux I__6555 (
            .O(N__55735),
            .I(shift_srl_10Z0Z_6));
    InMux I__6554 (
            .O(N__55732),
            .I(N__55725));
    InMux I__6553 (
            .O(N__55731),
            .I(N__55725));
    CascadeMux I__6552 (
            .O(N__55730),
            .I(N__55721));
    LocalMux I__6551 (
            .O(N__55725),
            .I(N__55716));
    InMux I__6550 (
            .O(N__55724),
            .I(N__55711));
    InMux I__6549 (
            .O(N__55721),
            .I(N__55711));
    InMux I__6548 (
            .O(N__55720),
            .I(N__55704));
    InMux I__6547 (
            .O(N__55719),
            .I(N__55704));
    Span4Mux_v I__6546 (
            .O(N__55716),
            .I(N__55701));
    LocalMux I__6545 (
            .O(N__55711),
            .I(N__55698));
    InMux I__6544 (
            .O(N__55710),
            .I(N__55695));
    InMux I__6543 (
            .O(N__55709),
            .I(N__55692));
    LocalMux I__6542 (
            .O(N__55704),
            .I(N__55689));
    Span4Mux_h I__6541 (
            .O(N__55701),
            .I(N__55686));
    Span12Mux_s8_h I__6540 (
            .O(N__55698),
            .I(N__55683));
    LocalMux I__6539 (
            .O(N__55695),
            .I(N__55680));
    LocalMux I__6538 (
            .O(N__55692),
            .I(shift_srl_10Z0Z_15));
    Odrv4 I__6537 (
            .O(N__55689),
            .I(shift_srl_10Z0Z_15));
    Odrv4 I__6536 (
            .O(N__55686),
            .I(shift_srl_10Z0Z_15));
    Odrv12 I__6535 (
            .O(N__55683),
            .I(shift_srl_10Z0Z_15));
    Odrv4 I__6534 (
            .O(N__55680),
            .I(shift_srl_10Z0Z_15));
    InMux I__6533 (
            .O(N__55669),
            .I(N__55666));
    LocalMux I__6532 (
            .O(N__55666),
            .I(shift_srl_10Z0Z_0));
    InMux I__6531 (
            .O(N__55663),
            .I(N__55660));
    LocalMux I__6530 (
            .O(N__55660),
            .I(shift_srl_10Z0Z_1));
    InMux I__6529 (
            .O(N__55657),
            .I(N__55654));
    LocalMux I__6528 (
            .O(N__55654),
            .I(shift_srl_10Z0Z_2));
    InMux I__6527 (
            .O(N__55651),
            .I(N__55648));
    LocalMux I__6526 (
            .O(N__55648),
            .I(shift_srl_10Z0Z_3));
    CEMux I__6525 (
            .O(N__55645),
            .I(N__55642));
    LocalMux I__6524 (
            .O(N__55642),
            .I(N__55637));
    CEMux I__6523 (
            .O(N__55641),
            .I(N__55634));
    CEMux I__6522 (
            .O(N__55640),
            .I(N__55631));
    Sp12to4 I__6521 (
            .O(N__55637),
            .I(N__55626));
    LocalMux I__6520 (
            .O(N__55634),
            .I(N__55626));
    LocalMux I__6519 (
            .O(N__55631),
            .I(N__55623));
    Odrv12 I__6518 (
            .O(N__55626),
            .I(clk_en_10));
    Odrv4 I__6517 (
            .O(N__55623),
            .I(clk_en_10));
    CascadeMux I__6516 (
            .O(N__55618),
            .I(shift_srl_149_RNIU42SZ0Z_15_cascade_));
    CEMux I__6515 (
            .O(N__55615),
            .I(N__55611));
    CEMux I__6514 (
            .O(N__55614),
            .I(N__55608));
    LocalMux I__6513 (
            .O(N__55611),
            .I(clk_en_150));
    LocalMux I__6512 (
            .O(N__55608),
            .I(clk_en_150));
    InMux I__6511 (
            .O(N__55603),
            .I(N__55600));
    LocalMux I__6510 (
            .O(N__55600),
            .I(shift_srl_0Z0Z_7));
    InMux I__6509 (
            .O(N__55597),
            .I(N__55594));
    LocalMux I__6508 (
            .O(N__55594),
            .I(shift_srl_0Z0Z_5));
    InMux I__6507 (
            .O(N__55591),
            .I(N__55588));
    LocalMux I__6506 (
            .O(N__55588),
            .I(shift_srl_0Z0Z_6));
    InMux I__6505 (
            .O(N__55585),
            .I(N__55582));
    LocalMux I__6504 (
            .O(N__55582),
            .I(shift_srl_0Z0Z_8));
    InMux I__6503 (
            .O(N__55579),
            .I(N__55576));
    LocalMux I__6502 (
            .O(N__55576),
            .I(shift_srl_0Z0Z_9));
    IoInMux I__6501 (
            .O(N__55573),
            .I(N__55570));
    LocalMux I__6500 (
            .O(N__55570),
            .I(N__55567));
    IoSpan4Mux I__6499 (
            .O(N__55567),
            .I(N__55564));
    Span4Mux_s3_v I__6498 (
            .O(N__55564),
            .I(N__55561));
    Odrv4 I__6497 (
            .O(N__55561),
            .I(rco_c_152));
    InMux I__6496 (
            .O(N__55558),
            .I(N__55555));
    LocalMux I__6495 (
            .O(N__55555),
            .I(shift_srl_10Z0Z_4));
    InMux I__6494 (
            .O(N__55552),
            .I(N__55549));
    LocalMux I__6493 (
            .O(N__55549),
            .I(shift_srl_10Z0Z_7));
    IoInMux I__6492 (
            .O(N__55546),
            .I(N__55543));
    LocalMux I__6491 (
            .O(N__55543),
            .I(N__55540));
    IoSpan4Mux I__6490 (
            .O(N__55540),
            .I(N__55537));
    Odrv4 I__6489 (
            .O(N__55537),
            .I(rco_c_108));
    CascadeMux I__6488 (
            .O(N__55534),
            .I(rco_c_108_cascade_));
    IoInMux I__6487 (
            .O(N__55531),
            .I(N__55528));
    LocalMux I__6486 (
            .O(N__55528),
            .I(N__55525));
    IoSpan4Mux I__6485 (
            .O(N__55525),
            .I(N__55522));
    Odrv4 I__6484 (
            .O(N__55522),
            .I(rco_c_109));
    IoInMux I__6483 (
            .O(N__55519),
            .I(N__55516));
    LocalMux I__6482 (
            .O(N__55516),
            .I(N__55513));
    Span4Mux_s0_v I__6481 (
            .O(N__55513),
            .I(N__55510));
    Span4Mux_h I__6480 (
            .O(N__55510),
            .I(N__55507));
    Odrv4 I__6479 (
            .O(N__55507),
            .I(rco_c_107));
    InMux I__6478 (
            .O(N__55504),
            .I(N__55501));
    LocalMux I__6477 (
            .O(N__55501),
            .I(shift_srl_0Z0Z_0));
    InMux I__6476 (
            .O(N__55498),
            .I(N__55495));
    LocalMux I__6475 (
            .O(N__55495),
            .I(shift_srl_0Z0Z_1));
    InMux I__6474 (
            .O(N__55492),
            .I(N__55489));
    LocalMux I__6473 (
            .O(N__55489),
            .I(shift_srl_0Z0Z_2));
    InMux I__6472 (
            .O(N__55486),
            .I(N__55483));
    LocalMux I__6471 (
            .O(N__55483),
            .I(shift_srl_0Z0Z_3));
    InMux I__6470 (
            .O(N__55480),
            .I(N__55477));
    LocalMux I__6469 (
            .O(N__55477),
            .I(shift_srl_0Z0Z_4));
    InMux I__6468 (
            .O(N__55474),
            .I(N__55471));
    LocalMux I__6467 (
            .O(N__55471),
            .I(shift_srl_106Z0Z_2));
    InMux I__6466 (
            .O(N__55468),
            .I(N__55465));
    LocalMux I__6465 (
            .O(N__55465),
            .I(shift_srl_106Z0Z_3));
    InMux I__6464 (
            .O(N__55462),
            .I(N__55459));
    LocalMux I__6463 (
            .O(N__55459),
            .I(shift_srl_106Z0Z_4));
    InMux I__6462 (
            .O(N__55456),
            .I(N__55453));
    LocalMux I__6461 (
            .O(N__55453),
            .I(shift_srl_106Z0Z_5));
    InMux I__6460 (
            .O(N__55450),
            .I(N__55447));
    LocalMux I__6459 (
            .O(N__55447),
            .I(shift_srl_106Z0Z_6));
    InMux I__6458 (
            .O(N__55444),
            .I(N__55441));
    LocalMux I__6457 (
            .O(N__55441),
            .I(shift_srl_106Z0Z_7));
    InMux I__6456 (
            .O(N__55438),
            .I(N__55435));
    LocalMux I__6455 (
            .O(N__55435),
            .I(shift_srl_118Z0Z_10));
    InMux I__6454 (
            .O(N__55432),
            .I(N__55429));
    LocalMux I__6453 (
            .O(N__55429),
            .I(N__55426));
    Odrv12 I__6452 (
            .O(N__55426),
            .I(shift_srl_118Z0Z_11));
    InMux I__6451 (
            .O(N__55423),
            .I(N__55420));
    LocalMux I__6450 (
            .O(N__55420),
            .I(shift_srl_118Z0Z_9));
    InMux I__6449 (
            .O(N__55417),
            .I(N__55414));
    LocalMux I__6448 (
            .O(N__55414),
            .I(shift_srl_118Z0Z_8));
    InMux I__6447 (
            .O(N__55411),
            .I(N__55408));
    LocalMux I__6446 (
            .O(N__55408),
            .I(shift_srl_133Z0Z_0));
    InMux I__6445 (
            .O(N__55405),
            .I(N__55402));
    LocalMux I__6444 (
            .O(N__55402),
            .I(shift_srl_133Z0Z_1));
    InMux I__6443 (
            .O(N__55399),
            .I(N__55396));
    LocalMux I__6442 (
            .O(N__55396),
            .I(shift_srl_133Z0Z_2));
    InMux I__6441 (
            .O(N__55393),
            .I(N__55390));
    LocalMux I__6440 (
            .O(N__55390),
            .I(N__55387));
    Sp12to4 I__6439 (
            .O(N__55387),
            .I(N__55384));
    Span12Mux_v I__6438 (
            .O(N__55384),
            .I(N__55381));
    Odrv12 I__6437 (
            .O(N__55381),
            .I(shift_srl_133Z0Z_3));
    CEMux I__6436 (
            .O(N__55378),
            .I(N__55366));
    CEMux I__6435 (
            .O(N__55377),
            .I(N__55366));
    CEMux I__6434 (
            .O(N__55376),
            .I(N__55366));
    CEMux I__6433 (
            .O(N__55375),
            .I(N__55366));
    GlobalMux I__6432 (
            .O(N__55366),
            .I(N__55363));
    gio2CtrlBuf I__6431 (
            .O(N__55363),
            .I(clk_en_g_133));
    InMux I__6430 (
            .O(N__55360),
            .I(N__55357));
    LocalMux I__6429 (
            .O(N__55357),
            .I(shift_srl_105Z0Z_6));
    InMux I__6428 (
            .O(N__55354),
            .I(N__55351));
    LocalMux I__6427 (
            .O(N__55351),
            .I(shift_srl_105Z0Z_5));
    InMux I__6426 (
            .O(N__55348),
            .I(N__55345));
    LocalMux I__6425 (
            .O(N__55345),
            .I(shift_srl_110Z0Z_10));
    InMux I__6424 (
            .O(N__55342),
            .I(N__55339));
    LocalMux I__6423 (
            .O(N__55339),
            .I(shift_srl_110Z0Z_11));
    InMux I__6422 (
            .O(N__55336),
            .I(N__55333));
    LocalMux I__6421 (
            .O(N__55333),
            .I(shift_srl_110Z0Z_12));
    InMux I__6420 (
            .O(N__55330),
            .I(N__55327));
    LocalMux I__6419 (
            .O(N__55327),
            .I(shift_srl_110Z0Z_13));
    InMux I__6418 (
            .O(N__55324),
            .I(N__55321));
    LocalMux I__6417 (
            .O(N__55321),
            .I(shift_srl_110Z0Z_9));
    IoInMux I__6416 (
            .O(N__55318),
            .I(N__55315));
    LocalMux I__6415 (
            .O(N__55315),
            .I(N__55312));
    Span4Mux_s3_v I__6414 (
            .O(N__55312),
            .I(N__55309));
    Span4Mux_v I__6413 (
            .O(N__55309),
            .I(N__55306));
    Sp12to4 I__6412 (
            .O(N__55306),
            .I(N__55303));
    Span12Mux_h I__6411 (
            .O(N__55303),
            .I(N__55300));
    Odrv12 I__6410 (
            .O(N__55300),
            .I(rco_c_122));
    InMux I__6409 (
            .O(N__55297),
            .I(N__55294));
    LocalMux I__6408 (
            .O(N__55294),
            .I(shift_srl_113Z0Z_7));
    InMux I__6407 (
            .O(N__55291),
            .I(N__55288));
    LocalMux I__6406 (
            .O(N__55288),
            .I(shift_srl_113Z0Z_6));
    InMux I__6405 (
            .O(N__55285),
            .I(N__55282));
    LocalMux I__6404 (
            .O(N__55282),
            .I(shift_srl_113Z0Z_0));
    InMux I__6403 (
            .O(N__55279),
            .I(N__55276));
    LocalMux I__6402 (
            .O(N__55276),
            .I(shift_srl_113Z0Z_1));
    InMux I__6401 (
            .O(N__55273),
            .I(N__55270));
    LocalMux I__6400 (
            .O(N__55270),
            .I(shift_srl_113Z0Z_2));
    InMux I__6399 (
            .O(N__55267),
            .I(N__55264));
    LocalMux I__6398 (
            .O(N__55264),
            .I(shift_srl_113Z0Z_3));
    InMux I__6397 (
            .O(N__55261),
            .I(N__55258));
    LocalMux I__6396 (
            .O(N__55258),
            .I(shift_srl_113Z0Z_4));
    InMux I__6395 (
            .O(N__55255),
            .I(N__55252));
    LocalMux I__6394 (
            .O(N__55252),
            .I(shift_srl_113Z0Z_5));
    InMux I__6393 (
            .O(N__55249),
            .I(N__55246));
    LocalMux I__6392 (
            .O(N__55246),
            .I(shift_srl_118Z0Z_13));
    InMux I__6391 (
            .O(N__55243),
            .I(N__55240));
    LocalMux I__6390 (
            .O(N__55240),
            .I(shift_srl_118Z0Z_12));
    InMux I__6389 (
            .O(N__55237),
            .I(N__55234));
    LocalMux I__6388 (
            .O(N__55234),
            .I(shift_srl_125Z0Z_0));
    InMux I__6387 (
            .O(N__55231),
            .I(N__55228));
    LocalMux I__6386 (
            .O(N__55228),
            .I(shift_srl_125Z0Z_1));
    InMux I__6385 (
            .O(N__55225),
            .I(N__55222));
    LocalMux I__6384 (
            .O(N__55222),
            .I(shift_srl_125Z0Z_2));
    InMux I__6383 (
            .O(N__55219),
            .I(N__55216));
    LocalMux I__6382 (
            .O(N__55216),
            .I(shift_srl_125Z0Z_3));
    InMux I__6381 (
            .O(N__55213),
            .I(N__55210));
    LocalMux I__6380 (
            .O(N__55210),
            .I(shift_srl_125Z0Z_4));
    InMux I__6379 (
            .O(N__55207),
            .I(N__55204));
    LocalMux I__6378 (
            .O(N__55204),
            .I(shift_srl_125Z0Z_5));
    InMux I__6377 (
            .O(N__55201),
            .I(N__55198));
    LocalMux I__6376 (
            .O(N__55198),
            .I(shift_srl_125Z0Z_6));
    InMux I__6375 (
            .O(N__55195),
            .I(N__55192));
    LocalMux I__6374 (
            .O(N__55192),
            .I(shift_srl_123Z0Z_9));
    InMux I__6373 (
            .O(N__55189),
            .I(N__55186));
    LocalMux I__6372 (
            .O(N__55186),
            .I(shift_srl_123Z0Z_8));
    InMux I__6371 (
            .O(N__55183),
            .I(N__55180));
    LocalMux I__6370 (
            .O(N__55180),
            .I(N__55177));
    Span4Mux_h I__6369 (
            .O(N__55177),
            .I(N__55174));
    Odrv4 I__6368 (
            .O(N__55174),
            .I(shift_srl_123Z0Z_6));
    InMux I__6367 (
            .O(N__55171),
            .I(N__55168));
    LocalMux I__6366 (
            .O(N__55168),
            .I(shift_srl_123Z0Z_7));
    CascadeMux I__6365 (
            .O(N__55165),
            .I(clk_en_0_a3_0_a2_sx_123_cascade_));
    CascadeMux I__6364 (
            .O(N__55162),
            .I(clk_en_0_a3_0_a2_sx_125_cascade_));
    InMux I__6363 (
            .O(N__55159),
            .I(N__55156));
    LocalMux I__6362 (
            .O(N__55156),
            .I(shift_srl_118Z0Z_14));
    InMux I__6361 (
            .O(N__55153),
            .I(N__55150));
    LocalMux I__6360 (
            .O(N__55150),
            .I(shift_srl_149Z0Z_3));
    InMux I__6359 (
            .O(N__55147),
            .I(N__55144));
    LocalMux I__6358 (
            .O(N__55144),
            .I(shift_srl_149Z0Z_4));
    InMux I__6357 (
            .O(N__55141),
            .I(N__55138));
    LocalMux I__6356 (
            .O(N__55138),
            .I(shift_srl_149Z0Z_5));
    InMux I__6355 (
            .O(N__55135),
            .I(N__55132));
    LocalMux I__6354 (
            .O(N__55132),
            .I(shift_srl_149Z0Z_6));
    InMux I__6353 (
            .O(N__55129),
            .I(N__55126));
    LocalMux I__6352 (
            .O(N__55126),
            .I(shift_srl_149Z0Z_7));
    InMux I__6351 (
            .O(N__55123),
            .I(N__55120));
    LocalMux I__6350 (
            .O(N__55120),
            .I(shift_srl_123Z0Z_10));
    InMux I__6349 (
            .O(N__55117),
            .I(N__55114));
    LocalMux I__6348 (
            .O(N__55114),
            .I(shift_srl_123Z0Z_11));
    InMux I__6347 (
            .O(N__55111),
            .I(N__55108));
    LocalMux I__6346 (
            .O(N__55108),
            .I(shift_srl_123Z0Z_12));
    InMux I__6345 (
            .O(N__55105),
            .I(N__55102));
    LocalMux I__6344 (
            .O(N__55102),
            .I(shift_srl_123Z0Z_13));
    InMux I__6343 (
            .O(N__55099),
            .I(N__55096));
    LocalMux I__6342 (
            .O(N__55096),
            .I(shift_srl_149Z0Z_12));
    InMux I__6341 (
            .O(N__55093),
            .I(N__55090));
    LocalMux I__6340 (
            .O(N__55090),
            .I(shift_srl_149Z0Z_13));
    InMux I__6339 (
            .O(N__55087),
            .I(N__55084));
    LocalMux I__6338 (
            .O(N__55084),
            .I(shift_srl_149Z0Z_14));
    InMux I__6337 (
            .O(N__55081),
            .I(N__55078));
    LocalMux I__6336 (
            .O(N__55078),
            .I(shift_srl_149Z0Z_9));
    InMux I__6335 (
            .O(N__55075),
            .I(N__55072));
    LocalMux I__6334 (
            .O(N__55072),
            .I(shift_srl_149Z0Z_8));
    InMux I__6333 (
            .O(N__55069),
            .I(N__55066));
    LocalMux I__6332 (
            .O(N__55066),
            .I(shift_srl_149Z0Z_0));
    InMux I__6331 (
            .O(N__55063),
            .I(N__55060));
    LocalMux I__6330 (
            .O(N__55060),
            .I(shift_srl_149Z0Z_1));
    InMux I__6329 (
            .O(N__55057),
            .I(N__55054));
    LocalMux I__6328 (
            .O(N__55054),
            .I(shift_srl_149Z0Z_2));
    InMux I__6327 (
            .O(N__55051),
            .I(N__55048));
    LocalMux I__6326 (
            .O(N__55048),
            .I(shift_srl_27Z0Z_11));
    InMux I__6325 (
            .O(N__55045),
            .I(N__55042));
    LocalMux I__6324 (
            .O(N__55042),
            .I(shift_srl_27Z0Z_12));
    InMux I__6323 (
            .O(N__55039),
            .I(N__55036));
    LocalMux I__6322 (
            .O(N__55036),
            .I(shift_srl_27Z0Z_7));
    InMux I__6321 (
            .O(N__55033),
            .I(N__55030));
    LocalMux I__6320 (
            .O(N__55030),
            .I(shift_srl_27Z0Z_13));
    InMux I__6319 (
            .O(N__55027),
            .I(N__55024));
    LocalMux I__6318 (
            .O(N__55024),
            .I(shift_srl_27Z0Z_14));
    InMux I__6317 (
            .O(N__55021),
            .I(N__55018));
    LocalMux I__6316 (
            .O(N__55018),
            .I(shift_srl_27Z0Z_8));
    InMux I__6315 (
            .O(N__55015),
            .I(N__55012));
    LocalMux I__6314 (
            .O(N__55012),
            .I(shift_srl_27Z0Z_9));
    CEMux I__6313 (
            .O(N__55009),
            .I(N__55006));
    LocalMux I__6312 (
            .O(N__55006),
            .I(N__55002));
    CEMux I__6311 (
            .O(N__55005),
            .I(N__54999));
    Span4Mux_v I__6310 (
            .O(N__55002),
            .I(N__54994));
    LocalMux I__6309 (
            .O(N__54999),
            .I(N__54994));
    Span4Mux_v I__6308 (
            .O(N__54994),
            .I(N__54991));
    Odrv4 I__6307 (
            .O(N__54991),
            .I(clk_en_27));
    InMux I__6306 (
            .O(N__54988),
            .I(N__54985));
    LocalMux I__6305 (
            .O(N__54985),
            .I(shift_srl_149Z0Z_10));
    InMux I__6304 (
            .O(N__54982),
            .I(N__54979));
    LocalMux I__6303 (
            .O(N__54979),
            .I(shift_srl_149Z0Z_11));
    InMux I__6302 (
            .O(N__54976),
            .I(N__54973));
    LocalMux I__6301 (
            .O(N__54973),
            .I(shift_srl_27Z0Z_0));
    InMux I__6300 (
            .O(N__54970),
            .I(N__54967));
    LocalMux I__6299 (
            .O(N__54967),
            .I(shift_srl_27Z0Z_1));
    InMux I__6298 (
            .O(N__54964),
            .I(N__54961));
    LocalMux I__6297 (
            .O(N__54961),
            .I(shift_srl_27Z0Z_2));
    InMux I__6296 (
            .O(N__54958),
            .I(N__54955));
    LocalMux I__6295 (
            .O(N__54955),
            .I(shift_srl_27Z0Z_3));
    InMux I__6294 (
            .O(N__54952),
            .I(N__54949));
    LocalMux I__6293 (
            .O(N__54949),
            .I(shift_srl_27Z0Z_4));
    InMux I__6292 (
            .O(N__54946),
            .I(N__54943));
    LocalMux I__6291 (
            .O(N__54943),
            .I(shift_srl_27Z0Z_5));
    InMux I__6290 (
            .O(N__54940),
            .I(N__54937));
    LocalMux I__6289 (
            .O(N__54937),
            .I(shift_srl_27Z0Z_6));
    InMux I__6288 (
            .O(N__54934),
            .I(N__54931));
    LocalMux I__6287 (
            .O(N__54931),
            .I(shift_srl_27Z0Z_10));
    InMux I__6286 (
            .O(N__54928),
            .I(N__54925));
    LocalMux I__6285 (
            .O(N__54925),
            .I(shift_srl_146Z0Z_3));
    InMux I__6284 (
            .O(N__54922),
            .I(N__54919));
    LocalMux I__6283 (
            .O(N__54919),
            .I(shift_srl_146Z0Z_4));
    InMux I__6282 (
            .O(N__54916),
            .I(N__54913));
    LocalMux I__6281 (
            .O(N__54913),
            .I(shift_srl_146Z0Z_10));
    InMux I__6280 (
            .O(N__54910),
            .I(N__54907));
    LocalMux I__6279 (
            .O(N__54907),
            .I(shift_srl_146Z0Z_11));
    InMux I__6278 (
            .O(N__54904),
            .I(N__54901));
    LocalMux I__6277 (
            .O(N__54901),
            .I(shift_srl_146Z0Z_12));
    InMux I__6276 (
            .O(N__54898),
            .I(N__54895));
    LocalMux I__6275 (
            .O(N__54895),
            .I(shift_srl_146Z0Z_13));
    InMux I__6274 (
            .O(N__54892),
            .I(N__54889));
    LocalMux I__6273 (
            .O(N__54889),
            .I(shift_srl_146Z0Z_9));
    InMux I__6272 (
            .O(N__54886),
            .I(N__54883));
    LocalMux I__6271 (
            .O(N__54883),
            .I(shift_srl_146Z0Z_8));
    InMux I__6270 (
            .O(N__54880),
            .I(N__54877));
    LocalMux I__6269 (
            .O(N__54877),
            .I(shift_srl_146Z0Z_6));
    InMux I__6268 (
            .O(N__54874),
            .I(N__54871));
    LocalMux I__6267 (
            .O(N__54871),
            .I(shift_srl_146Z0Z_7));
    InMux I__6266 (
            .O(N__54868),
            .I(N__54865));
    LocalMux I__6265 (
            .O(N__54865),
            .I(shift_srl_150Z0Z_14));
    InMux I__6264 (
            .O(N__54862),
            .I(N__54859));
    LocalMux I__6263 (
            .O(N__54859),
            .I(shift_srl_150Z0Z_9));
    InMux I__6262 (
            .O(N__54856),
            .I(N__54853));
    LocalMux I__6261 (
            .O(N__54853),
            .I(shift_srl_150Z0Z_7));
    InMux I__6260 (
            .O(N__54850),
            .I(N__54847));
    LocalMux I__6259 (
            .O(N__54847),
            .I(shift_srl_150Z0Z_8));
    InMux I__6258 (
            .O(N__54844),
            .I(N__54841));
    LocalMux I__6257 (
            .O(N__54841),
            .I(shift_srl_147Z0Z_5));
    InMux I__6256 (
            .O(N__54838),
            .I(N__54835));
    LocalMux I__6255 (
            .O(N__54835),
            .I(shift_srl_147Z0Z_6));
    InMux I__6254 (
            .O(N__54832),
            .I(N__54829));
    LocalMux I__6253 (
            .O(N__54829),
            .I(shift_srl_146Z0Z_5));
    InMux I__6252 (
            .O(N__54826),
            .I(N__54823));
    LocalMux I__6251 (
            .O(N__54823),
            .I(shift_srl_150Z0Z_3));
    InMux I__6250 (
            .O(N__54820),
            .I(N__54817));
    LocalMux I__6249 (
            .O(N__54817),
            .I(shift_srl_150Z0Z_4));
    InMux I__6248 (
            .O(N__54814),
            .I(N__54811));
    LocalMux I__6247 (
            .O(N__54811),
            .I(shift_srl_150Z0Z_5));
    InMux I__6246 (
            .O(N__54808),
            .I(N__54805));
    LocalMux I__6245 (
            .O(N__54805),
            .I(shift_srl_150Z0Z_6));
    InMux I__6244 (
            .O(N__54802),
            .I(N__54799));
    LocalMux I__6243 (
            .O(N__54799),
            .I(shift_srl_150Z0Z_10));
    InMux I__6242 (
            .O(N__54796),
            .I(N__54793));
    LocalMux I__6241 (
            .O(N__54793),
            .I(shift_srl_150Z0Z_11));
    InMux I__6240 (
            .O(N__54790),
            .I(N__54787));
    LocalMux I__6239 (
            .O(N__54787),
            .I(shift_srl_150Z0Z_12));
    InMux I__6238 (
            .O(N__54784),
            .I(N__54781));
    LocalMux I__6237 (
            .O(N__54781),
            .I(shift_srl_150Z0Z_13));
    InMux I__6236 (
            .O(N__54778),
            .I(N__54775));
    LocalMux I__6235 (
            .O(N__54775),
            .I(shift_srl_10Z0Z_11));
    InMux I__6234 (
            .O(N__54772),
            .I(N__54769));
    LocalMux I__6233 (
            .O(N__54769),
            .I(shift_srl_10Z0Z_12));
    InMux I__6232 (
            .O(N__54766),
            .I(N__54763));
    LocalMux I__6231 (
            .O(N__54763),
            .I(shift_srl_10Z0Z_13));
    InMux I__6230 (
            .O(N__54760),
            .I(N__54757));
    LocalMux I__6229 (
            .O(N__54757),
            .I(shift_srl_10Z0Z_14));
    InMux I__6228 (
            .O(N__54754),
            .I(N__54751));
    LocalMux I__6227 (
            .O(N__54751),
            .I(shift_srl_10Z0Z_9));
    InMux I__6226 (
            .O(N__54748),
            .I(N__54745));
    LocalMux I__6225 (
            .O(N__54745),
            .I(shift_srl_10Z0Z_8));
    InMux I__6224 (
            .O(N__54742),
            .I(N__54739));
    LocalMux I__6223 (
            .O(N__54739),
            .I(shift_srl_150Z0Z_0));
    InMux I__6222 (
            .O(N__54736),
            .I(N__54733));
    LocalMux I__6221 (
            .O(N__54733),
            .I(shift_srl_150Z0Z_1));
    InMux I__6220 (
            .O(N__54730),
            .I(N__54727));
    LocalMux I__6219 (
            .O(N__54727),
            .I(shift_srl_150Z0Z_2));
    InMux I__6218 (
            .O(N__54724),
            .I(N__54721));
    LocalMux I__6217 (
            .O(N__54721),
            .I(shift_srl_107Z0Z_1));
    InMux I__6216 (
            .O(N__54718),
            .I(N__54715));
    LocalMux I__6215 (
            .O(N__54715),
            .I(shift_srl_107Z0Z_2));
    IoInMux I__6214 (
            .O(N__54712),
            .I(N__54709));
    LocalMux I__6213 (
            .O(N__54709),
            .I(N__54706));
    Odrv12 I__6212 (
            .O(N__54706),
            .I(rco_c_151));
    InMux I__6211 (
            .O(N__54703),
            .I(N__54700));
    LocalMux I__6210 (
            .O(N__54700),
            .I(shift_srl_1Z0Z_0));
    InMux I__6209 (
            .O(N__54697),
            .I(N__54694));
    LocalMux I__6208 (
            .O(N__54694),
            .I(shift_srl_1Z0Z_1));
    InMux I__6207 (
            .O(N__54691),
            .I(N__54688));
    LocalMux I__6206 (
            .O(N__54688),
            .I(shift_srl_1Z0Z_2));
    InMux I__6205 (
            .O(N__54685),
            .I(N__54682));
    LocalMux I__6204 (
            .O(N__54682),
            .I(N__54679));
    Span4Mux_h I__6203 (
            .O(N__54679),
            .I(N__54676));
    Odrv4 I__6202 (
            .O(N__54676),
            .I(shift_srl_1Z0Z_3));
    CEMux I__6201 (
            .O(N__54673),
            .I(N__54670));
    LocalMux I__6200 (
            .O(N__54670),
            .I(N__54666));
    CEMux I__6199 (
            .O(N__54669),
            .I(N__54663));
    Span4Mux_v I__6198 (
            .O(N__54666),
            .I(N__54658));
    LocalMux I__6197 (
            .O(N__54663),
            .I(N__54658));
    Span4Mux_v I__6196 (
            .O(N__54658),
            .I(N__54654));
    CEMux I__6195 (
            .O(N__54657),
            .I(N__54651));
    Span4Mux_s2_v I__6194 (
            .O(N__54654),
            .I(N__54647));
    LocalMux I__6193 (
            .O(N__54651),
            .I(N__54644));
    CEMux I__6192 (
            .O(N__54650),
            .I(N__54641));
    Span4Mux_v I__6191 (
            .O(N__54647),
            .I(N__54638));
    Span4Mux_h I__6190 (
            .O(N__54644),
            .I(N__54635));
    LocalMux I__6189 (
            .O(N__54641),
            .I(N__54632));
    Odrv4 I__6188 (
            .O(N__54638),
            .I(N_10_i));
    Odrv4 I__6187 (
            .O(N__54635),
            .I(N_10_i));
    Odrv4 I__6186 (
            .O(N__54632),
            .I(N_10_i));
    InMux I__6185 (
            .O(N__54625),
            .I(N__54622));
    LocalMux I__6184 (
            .O(N__54622),
            .I(shift_srl_10Z0Z_10));
    InMux I__6183 (
            .O(N__54619),
            .I(N__54616));
    LocalMux I__6182 (
            .O(N__54616),
            .I(shift_srl_123Z0Z_4));
    InMux I__6181 (
            .O(N__54613),
            .I(N__54610));
    LocalMux I__6180 (
            .O(N__54610),
            .I(shift_srl_123Z0Z_5));
    InMux I__6179 (
            .O(N__54607),
            .I(N__54604));
    LocalMux I__6178 (
            .O(N__54604),
            .I(shift_srl_123Z0Z_3));
    InMux I__6177 (
            .O(N__54601),
            .I(N__54598));
    LocalMux I__6176 (
            .O(N__54598),
            .I(shift_srl_107Z0Z_3));
    InMux I__6175 (
            .O(N__54595),
            .I(N__54592));
    LocalMux I__6174 (
            .O(N__54592),
            .I(shift_srl_107Z0Z_4));
    InMux I__6173 (
            .O(N__54589),
            .I(N__54586));
    LocalMux I__6172 (
            .O(N__54586),
            .I(shift_srl_107Z0Z_5));
    InMux I__6171 (
            .O(N__54583),
            .I(N__54580));
    LocalMux I__6170 (
            .O(N__54580),
            .I(shift_srl_107Z0Z_6));
    CEMux I__6169 (
            .O(N__54577),
            .I(N__54573));
    CEMux I__6168 (
            .O(N__54576),
            .I(N__54570));
    LocalMux I__6167 (
            .O(N__54573),
            .I(N__54566));
    LocalMux I__6166 (
            .O(N__54570),
            .I(N__54563));
    CEMux I__6165 (
            .O(N__54569),
            .I(N__54560));
    Span4Mux_v I__6164 (
            .O(N__54566),
            .I(N__54557));
    Span4Mux_h I__6163 (
            .O(N__54563),
            .I(N__54554));
    LocalMux I__6162 (
            .O(N__54560),
            .I(N__54551));
    Odrv4 I__6161 (
            .O(N__54557),
            .I(clk_en_116));
    Odrv4 I__6160 (
            .O(N__54554),
            .I(clk_en_116));
    Odrv12 I__6159 (
            .O(N__54551),
            .I(clk_en_116));
    InMux I__6158 (
            .O(N__54544),
            .I(N__54541));
    LocalMux I__6157 (
            .O(N__54541),
            .I(shift_srl_112Z0Z_0));
    InMux I__6156 (
            .O(N__54538),
            .I(N__54535));
    LocalMux I__6155 (
            .O(N__54535),
            .I(shift_srl_112Z0Z_1));
    InMux I__6154 (
            .O(N__54532),
            .I(N__54529));
    LocalMux I__6153 (
            .O(N__54529),
            .I(shift_srl_112Z0Z_2));
    InMux I__6152 (
            .O(N__54526),
            .I(N__54523));
    LocalMux I__6151 (
            .O(N__54523),
            .I(shift_srl_112Z0Z_3));
    InMux I__6150 (
            .O(N__54520),
            .I(N__54517));
    LocalMux I__6149 (
            .O(N__54517),
            .I(shift_srl_112Z0Z_4));
    InMux I__6148 (
            .O(N__54514),
            .I(N__54511));
    LocalMux I__6147 (
            .O(N__54511),
            .I(shift_srl_112Z0Z_5));
    InMux I__6146 (
            .O(N__54508),
            .I(N__54505));
    LocalMux I__6145 (
            .O(N__54505),
            .I(shift_srl_112Z0Z_6));
    InMux I__6144 (
            .O(N__54502),
            .I(N__54499));
    LocalMux I__6143 (
            .O(N__54499),
            .I(N__54496));
    Span4Mux_h I__6142 (
            .O(N__54496),
            .I(N__54493));
    Odrv4 I__6141 (
            .O(N__54493),
            .I(g0_9_3));
    CascadeMux I__6140 (
            .O(N__54490),
            .I(N__54487));
    InMux I__6139 (
            .O(N__54487),
            .I(N__54484));
    LocalMux I__6138 (
            .O(N__54484),
            .I(rco_int_0_a2_0_a2_1_1_sx_145));
    CascadeMux I__6137 (
            .O(N__54481),
            .I(N__54478));
    InMux I__6136 (
            .O(N__54478),
            .I(N__54475));
    LocalMux I__6135 (
            .O(N__54475),
            .I(N__54469));
    InMux I__6134 (
            .O(N__54474),
            .I(N__54461));
    InMux I__6133 (
            .O(N__54473),
            .I(N__54461));
    InMux I__6132 (
            .O(N__54472),
            .I(N__54461));
    Span4Mux_h I__6131 (
            .O(N__54469),
            .I(N__54457));
    InMux I__6130 (
            .O(N__54468),
            .I(N__54454));
    LocalMux I__6129 (
            .O(N__54461),
            .I(N__54451));
    InMux I__6128 (
            .O(N__54460),
            .I(N__54448));
    Span4Mux_h I__6127 (
            .O(N__54457),
            .I(N__54445));
    LocalMux I__6126 (
            .O(N__54454),
            .I(N__54440));
    Span4Mux_v I__6125 (
            .O(N__54451),
            .I(N__54440));
    LocalMux I__6124 (
            .O(N__54448),
            .I(shift_srl_136Z0Z_15));
    Odrv4 I__6123 (
            .O(N__54445),
            .I(shift_srl_136Z0Z_15));
    Odrv4 I__6122 (
            .O(N__54440),
            .I(shift_srl_136Z0Z_15));
    InMux I__6121 (
            .O(N__54433),
            .I(N__54430));
    LocalMux I__6120 (
            .O(N__54430),
            .I(N__54427));
    Span4Mux_s2_h I__6119 (
            .O(N__54427),
            .I(N__54424));
    Span4Mux_h I__6118 (
            .O(N__54424),
            .I(N__54421));
    Odrv4 I__6117 (
            .O(N__54421),
            .I(g0_10));
    InMux I__6116 (
            .O(N__54418),
            .I(N__54415));
    LocalMux I__6115 (
            .O(N__54415),
            .I(shift_srl_116Z0Z_14));
    InMux I__6114 (
            .O(N__54412),
            .I(N__54409));
    LocalMux I__6113 (
            .O(N__54409),
            .I(shift_srl_116Z0Z_13));
    InMux I__6112 (
            .O(N__54406),
            .I(N__54403));
    LocalMux I__6111 (
            .O(N__54403),
            .I(shift_srl_116Z0Z_12));
    InMux I__6110 (
            .O(N__54400),
            .I(N__54397));
    LocalMux I__6109 (
            .O(N__54397),
            .I(shift_srl_116Z0Z_11));
    InMux I__6108 (
            .O(N__54394),
            .I(N__54391));
    LocalMux I__6107 (
            .O(N__54391),
            .I(shift_srl_116Z0Z_10));
    InMux I__6106 (
            .O(N__54388),
            .I(N__54385));
    LocalMux I__6105 (
            .O(N__54385),
            .I(N__54382));
    Span4Mux_h I__6104 (
            .O(N__54382),
            .I(N__54379));
    Odrv4 I__6103 (
            .O(N__54379),
            .I(shift_srl_116Z0Z_8));
    InMux I__6102 (
            .O(N__54376),
            .I(N__54373));
    LocalMux I__6101 (
            .O(N__54373),
            .I(shift_srl_116Z0Z_9));
    CascadeMux I__6100 (
            .O(N__54370),
            .I(N__54366));
    InMux I__6099 (
            .O(N__54369),
            .I(N__54362));
    InMux I__6098 (
            .O(N__54366),
            .I(N__54356));
    InMux I__6097 (
            .O(N__54365),
            .I(N__54356));
    LocalMux I__6096 (
            .O(N__54362),
            .I(N__54351));
    InMux I__6095 (
            .O(N__54361),
            .I(N__54348));
    LocalMux I__6094 (
            .O(N__54356),
            .I(N__54345));
    InMux I__6093 (
            .O(N__54355),
            .I(N__54342));
    InMux I__6092 (
            .O(N__54354),
            .I(N__54337));
    Span4Mux_s3_h I__6091 (
            .O(N__54351),
            .I(N__54334));
    LocalMux I__6090 (
            .O(N__54348),
            .I(N__54327));
    Span4Mux_h I__6089 (
            .O(N__54345),
            .I(N__54327));
    LocalMux I__6088 (
            .O(N__54342),
            .I(N__54327));
    InMux I__6087 (
            .O(N__54341),
            .I(N__54324));
    InMux I__6086 (
            .O(N__54340),
            .I(N__54321));
    LocalMux I__6085 (
            .O(N__54337),
            .I(shift_srl_132Z0Z_15));
    Odrv4 I__6084 (
            .O(N__54334),
            .I(shift_srl_132Z0Z_15));
    Odrv4 I__6083 (
            .O(N__54327),
            .I(shift_srl_132Z0Z_15));
    LocalMux I__6082 (
            .O(N__54324),
            .I(shift_srl_132Z0Z_15));
    LocalMux I__6081 (
            .O(N__54321),
            .I(shift_srl_132Z0Z_15));
    InMux I__6080 (
            .O(N__54310),
            .I(N__54301));
    InMux I__6079 (
            .O(N__54309),
            .I(N__54301));
    InMux I__6078 (
            .O(N__54308),
            .I(N__54293));
    InMux I__6077 (
            .O(N__54307),
            .I(N__54290));
    InMux I__6076 (
            .O(N__54306),
            .I(N__54287));
    LocalMux I__6075 (
            .O(N__54301),
            .I(N__54284));
    InMux I__6074 (
            .O(N__54300),
            .I(N__54281));
    CascadeMux I__6073 (
            .O(N__54299),
            .I(N__54278));
    InMux I__6072 (
            .O(N__54298),
            .I(N__54275));
    InMux I__6071 (
            .O(N__54297),
            .I(N__54272));
    InMux I__6070 (
            .O(N__54296),
            .I(N__54269));
    LocalMux I__6069 (
            .O(N__54293),
            .I(N__54266));
    LocalMux I__6068 (
            .O(N__54290),
            .I(N__54263));
    LocalMux I__6067 (
            .O(N__54287),
            .I(N__54258));
    Span4Mux_h I__6066 (
            .O(N__54284),
            .I(N__54258));
    LocalMux I__6065 (
            .O(N__54281),
            .I(N__54255));
    InMux I__6064 (
            .O(N__54278),
            .I(N__54252));
    LocalMux I__6063 (
            .O(N__54275),
            .I(shift_srl_131Z0Z_15));
    LocalMux I__6062 (
            .O(N__54272),
            .I(shift_srl_131Z0Z_15));
    LocalMux I__6061 (
            .O(N__54269),
            .I(shift_srl_131Z0Z_15));
    Odrv4 I__6060 (
            .O(N__54266),
            .I(shift_srl_131Z0Z_15));
    Odrv4 I__6059 (
            .O(N__54263),
            .I(shift_srl_131Z0Z_15));
    Odrv4 I__6058 (
            .O(N__54258),
            .I(shift_srl_131Z0Z_15));
    Odrv4 I__6057 (
            .O(N__54255),
            .I(shift_srl_131Z0Z_15));
    LocalMux I__6056 (
            .O(N__54252),
            .I(shift_srl_131Z0Z_15));
    InMux I__6055 (
            .O(N__54235),
            .I(N__54225));
    InMux I__6054 (
            .O(N__54234),
            .I(N__54222));
    CascadeMux I__6053 (
            .O(N__54233),
            .I(N__54219));
    CascadeMux I__6052 (
            .O(N__54232),
            .I(N__54216));
    InMux I__6051 (
            .O(N__54231),
            .I(N__54213));
    InMux I__6050 (
            .O(N__54230),
            .I(N__54206));
    InMux I__6049 (
            .O(N__54229),
            .I(N__54206));
    InMux I__6048 (
            .O(N__54228),
            .I(N__54206));
    LocalMux I__6047 (
            .O(N__54225),
            .I(N__54200));
    LocalMux I__6046 (
            .O(N__54222),
            .I(N__54200));
    InMux I__6045 (
            .O(N__54219),
            .I(N__54195));
    InMux I__6044 (
            .O(N__54216),
            .I(N__54195));
    LocalMux I__6043 (
            .O(N__54213),
            .I(N__54190));
    LocalMux I__6042 (
            .O(N__54206),
            .I(N__54190));
    InMux I__6041 (
            .O(N__54205),
            .I(N__54187));
    Span4Mux_v I__6040 (
            .O(N__54200),
            .I(N__54181));
    LocalMux I__6039 (
            .O(N__54195),
            .I(N__54181));
    Span4Mux_v I__6038 (
            .O(N__54190),
            .I(N__54176));
    LocalMux I__6037 (
            .O(N__54187),
            .I(N__54173));
    InMux I__6036 (
            .O(N__54186),
            .I(N__54170));
    Span4Mux_h I__6035 (
            .O(N__54181),
            .I(N__54167));
    InMux I__6034 (
            .O(N__54180),
            .I(N__54162));
    InMux I__6033 (
            .O(N__54179),
            .I(N__54162));
    Odrv4 I__6032 (
            .O(N__54176),
            .I(shift_srl_129Z0Z_15));
    Odrv4 I__6031 (
            .O(N__54173),
            .I(shift_srl_129Z0Z_15));
    LocalMux I__6030 (
            .O(N__54170),
            .I(shift_srl_129Z0Z_15));
    Odrv4 I__6029 (
            .O(N__54167),
            .I(shift_srl_129Z0Z_15));
    LocalMux I__6028 (
            .O(N__54162),
            .I(shift_srl_129Z0Z_15));
    InMux I__6027 (
            .O(N__54151),
            .I(N__54148));
    LocalMux I__6026 (
            .O(N__54148),
            .I(N__54145));
    Span4Mux_h I__6025 (
            .O(N__54145),
            .I(N__54142));
    Odrv4 I__6024 (
            .O(N__54142),
            .I(g0_3));
    InMux I__6023 (
            .O(N__54139),
            .I(N__54136));
    LocalMux I__6022 (
            .O(N__54136),
            .I(shift_srl_128Z0Z_14));
    InMux I__6021 (
            .O(N__54133),
            .I(N__54130));
    LocalMux I__6020 (
            .O(N__54130),
            .I(shift_srl_128Z0Z_13));
    InMux I__6019 (
            .O(N__54127),
            .I(N__54124));
    LocalMux I__6018 (
            .O(N__54124),
            .I(shift_srl_128Z0Z_12));
    InMux I__6017 (
            .O(N__54121),
            .I(N__54118));
    LocalMux I__6016 (
            .O(N__54118),
            .I(shift_srl_128Z0Z_11));
    InMux I__6015 (
            .O(N__54115),
            .I(N__54112));
    LocalMux I__6014 (
            .O(N__54112),
            .I(shift_srl_128Z0Z_10));
    InMux I__6013 (
            .O(N__54109),
            .I(N__54106));
    LocalMux I__6012 (
            .O(N__54106),
            .I(N__54103));
    Odrv4 I__6011 (
            .O(N__54103),
            .I(shift_srl_128Z0Z_8));
    InMux I__6010 (
            .O(N__54100),
            .I(N__54097));
    LocalMux I__6009 (
            .O(N__54097),
            .I(shift_srl_128Z0Z_9));
    InMux I__6008 (
            .O(N__54094),
            .I(N__54091));
    LocalMux I__6007 (
            .O(N__54091),
            .I(shift_srl_9Z0Z_6));
    InMux I__6006 (
            .O(N__54088),
            .I(N__54085));
    LocalMux I__6005 (
            .O(N__54085),
            .I(shift_srl_9Z0Z_7));
    CEMux I__6004 (
            .O(N__54082),
            .I(N__54078));
    CEMux I__6003 (
            .O(N__54081),
            .I(N__54075));
    LocalMux I__6002 (
            .O(N__54078),
            .I(N__54072));
    LocalMux I__6001 (
            .O(N__54075),
            .I(N__54068));
    Span4Mux_v I__6000 (
            .O(N__54072),
            .I(N__54065));
    CEMux I__5999 (
            .O(N__54071),
            .I(N__54062));
    Span4Mux_h I__5998 (
            .O(N__54068),
            .I(N__54059));
    Span4Mux_h I__5997 (
            .O(N__54065),
            .I(N__54054));
    LocalMux I__5996 (
            .O(N__54062),
            .I(N__54054));
    Odrv4 I__5995 (
            .O(N__54059),
            .I(clk_en_9));
    Odrv4 I__5994 (
            .O(N__54054),
            .I(clk_en_9));
    InMux I__5993 (
            .O(N__54049),
            .I(N__54046));
    LocalMux I__5992 (
            .O(N__54046),
            .I(shift_srl_128Z0Z_0));
    InMux I__5991 (
            .O(N__54043),
            .I(N__54040));
    LocalMux I__5990 (
            .O(N__54040),
            .I(shift_srl_128Z0Z_1));
    InMux I__5989 (
            .O(N__54037),
            .I(N__54034));
    LocalMux I__5988 (
            .O(N__54034),
            .I(shift_srl_128Z0Z_2));
    InMux I__5987 (
            .O(N__54031),
            .I(N__54028));
    LocalMux I__5986 (
            .O(N__54028),
            .I(shift_srl_128Z0Z_3));
    InMux I__5985 (
            .O(N__54025),
            .I(N__54022));
    LocalMux I__5984 (
            .O(N__54022),
            .I(shift_srl_128Z0Z_4));
    InMux I__5983 (
            .O(N__54019),
            .I(N__54016));
    LocalMux I__5982 (
            .O(N__54016),
            .I(shift_srl_128Z0Z_5));
    InMux I__5981 (
            .O(N__54013),
            .I(N__54010));
    LocalMux I__5980 (
            .O(N__54010),
            .I(shift_srl_128Z0Z_6));
    InMux I__5979 (
            .O(N__54007),
            .I(N__54004));
    LocalMux I__5978 (
            .O(N__54004),
            .I(N__54001));
    Span4Mux_v I__5977 (
            .O(N__54001),
            .I(N__53998));
    Odrv4 I__5976 (
            .O(N__53998),
            .I(shift_srl_129Z0Z_14));
    CEMux I__5975 (
            .O(N__53995),
            .I(N__53991));
    CEMux I__5974 (
            .O(N__53994),
            .I(N__53988));
    LocalMux I__5973 (
            .O(N__53991),
            .I(N__53983));
    LocalMux I__5972 (
            .O(N__53988),
            .I(N__53980));
    CEMux I__5971 (
            .O(N__53987),
            .I(N__53977));
    CEMux I__5970 (
            .O(N__53986),
            .I(N__53974));
    Span4Mux_h I__5969 (
            .O(N__53983),
            .I(N__53971));
    Span4Mux_h I__5968 (
            .O(N__53980),
            .I(N__53968));
    LocalMux I__5967 (
            .O(N__53977),
            .I(N__53965));
    LocalMux I__5966 (
            .O(N__53974),
            .I(N__53962));
    Odrv4 I__5965 (
            .O(N__53971),
            .I(clk_en_129));
    Odrv4 I__5964 (
            .O(N__53968),
            .I(clk_en_129));
    Odrv4 I__5963 (
            .O(N__53965),
            .I(clk_en_129));
    Odrv4 I__5962 (
            .O(N__53962),
            .I(clk_en_129));
    CascadeMux I__5961 (
            .O(N__53953),
            .I(N_4016_i_cascade_));
    IoInMux I__5960 (
            .O(N__53950),
            .I(N__53947));
    LocalMux I__5959 (
            .O(N__53947),
            .I(N__53944));
    Span4Mux_s1_h I__5958 (
            .O(N__53944),
            .I(N__53941));
    Span4Mux_h I__5957 (
            .O(N__53941),
            .I(N__53938));
    Sp12to4 I__5956 (
            .O(N__53938),
            .I(N__53935));
    Span12Mux_v I__5955 (
            .O(N__53935),
            .I(N__53930));
    InMux I__5954 (
            .O(N__53934),
            .I(N__53925));
    InMux I__5953 (
            .O(N__53933),
            .I(N__53925));
    Odrv12 I__5952 (
            .O(N__53930),
            .I(rco_c_25));
    LocalMux I__5951 (
            .O(N__53925),
            .I(rco_c_25));
    InMux I__5950 (
            .O(N__53920),
            .I(N__53916));
    InMux I__5949 (
            .O(N__53919),
            .I(N__53913));
    LocalMux I__5948 (
            .O(N__53916),
            .I(shift_srl_9Z0Z_15));
    LocalMux I__5947 (
            .O(N__53913),
            .I(shift_srl_9Z0Z_15));
    InMux I__5946 (
            .O(N__53908),
            .I(N__53905));
    LocalMux I__5945 (
            .O(N__53905),
            .I(shift_srl_9Z0Z_10));
    InMux I__5944 (
            .O(N__53902),
            .I(N__53899));
    LocalMux I__5943 (
            .O(N__53899),
            .I(shift_srl_9Z0Z_11));
    InMux I__5942 (
            .O(N__53896),
            .I(N__53893));
    LocalMux I__5941 (
            .O(N__53893),
            .I(shift_srl_9Z0Z_12));
    InMux I__5940 (
            .O(N__53890),
            .I(N__53887));
    LocalMux I__5939 (
            .O(N__53887),
            .I(shift_srl_9Z0Z_13));
    InMux I__5938 (
            .O(N__53884),
            .I(N__53881));
    LocalMux I__5937 (
            .O(N__53881),
            .I(shift_srl_9Z0Z_14));
    InMux I__5936 (
            .O(N__53878),
            .I(N__53875));
    LocalMux I__5935 (
            .O(N__53875),
            .I(shift_srl_9Z0Z_9));
    InMux I__5934 (
            .O(N__53872),
            .I(N__53869));
    LocalMux I__5933 (
            .O(N__53869),
            .I(shift_srl_9Z0Z_8));
    InMux I__5932 (
            .O(N__53866),
            .I(N__53863));
    LocalMux I__5931 (
            .O(N__53863),
            .I(shift_srl_154Z0Z_0));
    InMux I__5930 (
            .O(N__53860),
            .I(N__53857));
    LocalMux I__5929 (
            .O(N__53857),
            .I(shift_srl_154Z0Z_1));
    InMux I__5928 (
            .O(N__53854),
            .I(N__53851));
    LocalMux I__5927 (
            .O(N__53851),
            .I(shift_srl_154Z0Z_2));
    IoInMux I__5926 (
            .O(N__53848),
            .I(N__53845));
    LocalMux I__5925 (
            .O(N__53845),
            .I(N__53842));
    IoSpan4Mux I__5924 (
            .O(N__53842),
            .I(N__53839));
    Sp12to4 I__5923 (
            .O(N__53839),
            .I(N__53836));
    Span12Mux_s6_h I__5922 (
            .O(N__53836),
            .I(N__53833));
    Odrv12 I__5921 (
            .O(N__53833),
            .I(rco_c_26));
    InMux I__5920 (
            .O(N__53830),
            .I(N__53827));
    LocalMux I__5919 (
            .O(N__53827),
            .I(N__53823));
    InMux I__5918 (
            .O(N__53826),
            .I(N__53819));
    Span4Mux_h I__5917 (
            .O(N__53823),
            .I(N__53816));
    InMux I__5916 (
            .O(N__53822),
            .I(N__53813));
    LocalMux I__5915 (
            .O(N__53819),
            .I(shift_srl_8Z0Z_15));
    Odrv4 I__5914 (
            .O(N__53816),
            .I(shift_srl_8Z0Z_15));
    LocalMux I__5913 (
            .O(N__53813),
            .I(shift_srl_8Z0Z_15));
    InMux I__5912 (
            .O(N__53806),
            .I(N__53797));
    InMux I__5911 (
            .O(N__53805),
            .I(N__53797));
    InMux I__5910 (
            .O(N__53804),
            .I(N__53794));
    InMux I__5909 (
            .O(N__53803),
            .I(N__53789));
    InMux I__5908 (
            .O(N__53802),
            .I(N__53789));
    LocalMux I__5907 (
            .O(N__53797),
            .I(N__53786));
    LocalMux I__5906 (
            .O(N__53794),
            .I(N__53781));
    LocalMux I__5905 (
            .O(N__53789),
            .I(N__53781));
    Span4Mux_v I__5904 (
            .O(N__53786),
            .I(N__53778));
    Span4Mux_v I__5903 (
            .O(N__53781),
            .I(N__53775));
    Odrv4 I__5902 (
            .O(N__53778),
            .I(rco_int_0_a2_0_9));
    Odrv4 I__5901 (
            .O(N__53775),
            .I(rco_int_0_a2_0_9));
    InMux I__5900 (
            .O(N__53770),
            .I(N__53767));
    LocalMux I__5899 (
            .O(N__53767),
            .I(N__53763));
    CascadeMux I__5898 (
            .O(N__53766),
            .I(N__53757));
    Span4Mux_v I__5897 (
            .O(N__53763),
            .I(N__53753));
    InMux I__5896 (
            .O(N__53762),
            .I(N__53750));
    InMux I__5895 (
            .O(N__53761),
            .I(N__53747));
    InMux I__5894 (
            .O(N__53760),
            .I(N__53740));
    InMux I__5893 (
            .O(N__53757),
            .I(N__53740));
    InMux I__5892 (
            .O(N__53756),
            .I(N__53740));
    Span4Mux_h I__5891 (
            .O(N__53753),
            .I(N__53737));
    LocalMux I__5890 (
            .O(N__53750),
            .I(shift_srl_7Z0Z_15));
    LocalMux I__5889 (
            .O(N__53747),
            .I(shift_srl_7Z0Z_15));
    LocalMux I__5888 (
            .O(N__53740),
            .I(shift_srl_7Z0Z_15));
    Odrv4 I__5887 (
            .O(N__53737),
            .I(shift_srl_7Z0Z_15));
    InMux I__5886 (
            .O(N__53728),
            .I(N__53717));
    InMux I__5885 (
            .O(N__53727),
            .I(N__53717));
    InMux I__5884 (
            .O(N__53726),
            .I(N__53714));
    InMux I__5883 (
            .O(N__53725),
            .I(N__53709));
    InMux I__5882 (
            .O(N__53724),
            .I(N__53709));
    InMux I__5881 (
            .O(N__53723),
            .I(N__53704));
    InMux I__5880 (
            .O(N__53722),
            .I(N__53704));
    LocalMux I__5879 (
            .O(N__53717),
            .I(N__53696));
    LocalMux I__5878 (
            .O(N__53714),
            .I(N__53696));
    LocalMux I__5877 (
            .O(N__53709),
            .I(N__53693));
    LocalMux I__5876 (
            .O(N__53704),
            .I(N__53690));
    InMux I__5875 (
            .O(N__53703),
            .I(N__53685));
    InMux I__5874 (
            .O(N__53702),
            .I(N__53685));
    InMux I__5873 (
            .O(N__53701),
            .I(N__53682));
    Span4Mux_v I__5872 (
            .O(N__53696),
            .I(N__53677));
    Span4Mux_s1_h I__5871 (
            .O(N__53693),
            .I(N__53677));
    Span4Mux_v I__5870 (
            .O(N__53690),
            .I(N__53671));
    LocalMux I__5869 (
            .O(N__53685),
            .I(N__53671));
    LocalMux I__5868 (
            .O(N__53682),
            .I(N__53668));
    Span4Mux_h I__5867 (
            .O(N__53677),
            .I(N__53665));
    InMux I__5866 (
            .O(N__53676),
            .I(N__53662));
    Span4Mux_v I__5865 (
            .O(N__53671),
            .I(N__53659));
    Span4Mux_v I__5864 (
            .O(N__53668),
            .I(N__53656));
    Odrv4 I__5863 (
            .O(N__53665),
            .I(N_453));
    LocalMux I__5862 (
            .O(N__53662),
            .I(N_453));
    Odrv4 I__5861 (
            .O(N__53659),
            .I(N_453));
    Odrv4 I__5860 (
            .O(N__53656),
            .I(N_453));
    CascadeMux I__5859 (
            .O(N__53647),
            .I(rco_int_0_a2_0_9_cascade_));
    CascadeMux I__5858 (
            .O(N__53644),
            .I(N__53640));
    InMux I__5857 (
            .O(N__53643),
            .I(N__53636));
    InMux I__5856 (
            .O(N__53640),
            .I(N__53633));
    InMux I__5855 (
            .O(N__53639),
            .I(N__53630));
    LocalMux I__5854 (
            .O(N__53636),
            .I(N__53627));
    LocalMux I__5853 (
            .O(N__53633),
            .I(N__53624));
    LocalMux I__5852 (
            .O(N__53630),
            .I(N__53619));
    Span4Mux_h I__5851 (
            .O(N__53627),
            .I(N__53619));
    Span4Mux_h I__5850 (
            .O(N__53624),
            .I(N__53616));
    Span4Mux_h I__5849 (
            .O(N__53619),
            .I(N__53613));
    Odrv4 I__5848 (
            .O(N__53616),
            .I(rco_int_0_a2_out_1));
    Odrv4 I__5847 (
            .O(N__53613),
            .I(rco_int_0_a2_out_1));
    CascadeMux I__5846 (
            .O(N__53608),
            .I(rco_c_9_cascade_));
    InMux I__5845 (
            .O(N__53605),
            .I(N__53602));
    LocalMux I__5844 (
            .O(N__53602),
            .I(shift_srl_23Z0Z_3));
    InMux I__5843 (
            .O(N__53599),
            .I(N__53596));
    LocalMux I__5842 (
            .O(N__53596),
            .I(shift_srl_23Z0Z_4));
    InMux I__5841 (
            .O(N__53593),
            .I(N__53590));
    LocalMux I__5840 (
            .O(N__53590),
            .I(shift_srl_23Z0Z_5));
    InMux I__5839 (
            .O(N__53587),
            .I(N__53584));
    LocalMux I__5838 (
            .O(N__53584),
            .I(shift_srl_23Z0Z_6));
    CEMux I__5837 (
            .O(N__53581),
            .I(N__53576));
    CEMux I__5836 (
            .O(N__53580),
            .I(N__53573));
    CEMux I__5835 (
            .O(N__53579),
            .I(N__53570));
    LocalMux I__5834 (
            .O(N__53576),
            .I(N_702));
    LocalMux I__5833 (
            .O(N__53573),
            .I(N_702));
    LocalMux I__5832 (
            .O(N__53570),
            .I(N_702));
    IoInMux I__5831 (
            .O(N__53563),
            .I(N__53560));
    LocalMux I__5830 (
            .O(N__53560),
            .I(N__53557));
    Span4Mux_s3_h I__5829 (
            .O(N__53557),
            .I(N__53554));
    Span4Mux_v I__5828 (
            .O(N__53554),
            .I(N__53551));
    Span4Mux_h I__5827 (
            .O(N__53551),
            .I(N__53548));
    Odrv4 I__5826 (
            .O(N__53548),
            .I(rco_c_155));
    IoInMux I__5825 (
            .O(N__53545),
            .I(N__53542));
    LocalMux I__5824 (
            .O(N__53542),
            .I(N__53539));
    Span4Mux_s2_h I__5823 (
            .O(N__53539),
            .I(N__53536));
    Span4Mux_v I__5822 (
            .O(N__53536),
            .I(N__53533));
    Span4Mux_h I__5821 (
            .O(N__53533),
            .I(N__53530));
    Odrv4 I__5820 (
            .O(N__53530),
            .I(rco_c_154));
    IoInMux I__5819 (
            .O(N__53527),
            .I(N__53524));
    LocalMux I__5818 (
            .O(N__53524),
            .I(N__53521));
    IoSpan4Mux I__5817 (
            .O(N__53521),
            .I(N__53518));
    Span4Mux_s2_h I__5816 (
            .O(N__53518),
            .I(N__53515));
    Span4Mux_h I__5815 (
            .O(N__53515),
            .I(N__53512));
    Odrv4 I__5814 (
            .O(N__53512),
            .I(rco_c_156));
    IoInMux I__5813 (
            .O(N__53509),
            .I(N__53506));
    LocalMux I__5812 (
            .O(N__53506),
            .I(N__53503));
    Span4Mux_s2_h I__5811 (
            .O(N__53503),
            .I(N__53500));
    Span4Mux_v I__5810 (
            .O(N__53500),
            .I(N__53497));
    Span4Mux_h I__5809 (
            .O(N__53497),
            .I(N__53494));
    Odrv4 I__5808 (
            .O(N__53494),
            .I(rco_c_159));
    IoInMux I__5807 (
            .O(N__53491),
            .I(N__53488));
    LocalMux I__5806 (
            .O(N__53488),
            .I(N__53485));
    Span4Mux_s2_h I__5805 (
            .O(N__53485),
            .I(N__53482));
    Span4Mux_v I__5804 (
            .O(N__53482),
            .I(N__53479));
    Span4Mux_h I__5803 (
            .O(N__53479),
            .I(N__53476));
    Odrv4 I__5802 (
            .O(N__53476),
            .I(rco_c_160));
    IoInMux I__5801 (
            .O(N__53473),
            .I(N__53470));
    LocalMux I__5800 (
            .O(N__53470),
            .I(N__53467));
    Span4Mux_s3_h I__5799 (
            .O(N__53467),
            .I(N__53464));
    Span4Mux_h I__5798 (
            .O(N__53464),
            .I(N__53461));
    Odrv4 I__5797 (
            .O(N__53461),
            .I(rco_c_161));
    InMux I__5796 (
            .O(N__53458),
            .I(N__53455));
    LocalMux I__5795 (
            .O(N__53455),
            .I(shift_srl_1Z0Z_10));
    InMux I__5794 (
            .O(N__53452),
            .I(N__53449));
    LocalMux I__5793 (
            .O(N__53449),
            .I(shift_srl_1Z0Z_8));
    InMux I__5792 (
            .O(N__53446),
            .I(N__53443));
    LocalMux I__5791 (
            .O(N__53443),
            .I(shift_srl_1Z0Z_9));
    InMux I__5790 (
            .O(N__53440),
            .I(N__53437));
    LocalMux I__5789 (
            .O(N__53437),
            .I(shift_srl_1Z0Z_14));
    InMux I__5788 (
            .O(N__53434),
            .I(N__53430));
    InMux I__5787 (
            .O(N__53433),
            .I(N__53427));
    LocalMux I__5786 (
            .O(N__53430),
            .I(N__53423));
    LocalMux I__5785 (
            .O(N__53427),
            .I(N__53420));
    InMux I__5784 (
            .O(N__53426),
            .I(N__53416));
    Span4Mux_h I__5783 (
            .O(N__53423),
            .I(N__53413));
    Span4Mux_v I__5782 (
            .O(N__53420),
            .I(N__53410));
    InMux I__5781 (
            .O(N__53419),
            .I(N__53407));
    LocalMux I__5780 (
            .O(N__53416),
            .I(N__53404));
    Odrv4 I__5779 (
            .O(N__53413),
            .I(shift_srl_22Z0Z_15));
    Odrv4 I__5778 (
            .O(N__53410),
            .I(shift_srl_22Z0Z_15));
    LocalMux I__5777 (
            .O(N__53407),
            .I(shift_srl_22Z0Z_15));
    Odrv4 I__5776 (
            .O(N__53404),
            .I(shift_srl_22Z0Z_15));
    InMux I__5775 (
            .O(N__53395),
            .I(N__53392));
    LocalMux I__5774 (
            .O(N__53392),
            .I(shift_srl_23Z0Z_14));
    InMux I__5773 (
            .O(N__53389),
            .I(N__53383));
    InMux I__5772 (
            .O(N__53388),
            .I(N__53383));
    LocalMux I__5771 (
            .O(N__53383),
            .I(shift_srl_23Z0Z_15));
    InMux I__5770 (
            .O(N__53380),
            .I(N__53377));
    LocalMux I__5769 (
            .O(N__53377),
            .I(shift_srl_23Z0Z_0));
    InMux I__5768 (
            .O(N__53374),
            .I(N__53371));
    LocalMux I__5767 (
            .O(N__53371),
            .I(shift_srl_23Z0Z_1));
    InMux I__5766 (
            .O(N__53368),
            .I(N__53365));
    LocalMux I__5765 (
            .O(N__53365),
            .I(shift_srl_23Z0Z_2));
    InMux I__5764 (
            .O(N__53362),
            .I(N__53359));
    LocalMux I__5763 (
            .O(N__53359),
            .I(shift_srl_1Z0Z_7));
    InMux I__5762 (
            .O(N__53356),
            .I(N__53353));
    LocalMux I__5761 (
            .O(N__53353),
            .I(shift_srl_1Z0Z_6));
    InMux I__5760 (
            .O(N__53350),
            .I(N__53347));
    LocalMux I__5759 (
            .O(N__53347),
            .I(shift_srl_1Z0Z_5));
    InMux I__5758 (
            .O(N__53344),
            .I(N__53341));
    LocalMux I__5757 (
            .O(N__53341),
            .I(shift_srl_1Z0Z_4));
    CEMux I__5756 (
            .O(N__53338),
            .I(N__53334));
    CEMux I__5755 (
            .O(N__53337),
            .I(N__53330));
    LocalMux I__5754 (
            .O(N__53334),
            .I(N__53327));
    CEMux I__5753 (
            .O(N__53333),
            .I(N__53324));
    LocalMux I__5752 (
            .O(N__53330),
            .I(N__53321));
    Span4Mux_v I__5751 (
            .O(N__53327),
            .I(N__53316));
    LocalMux I__5750 (
            .O(N__53324),
            .I(N__53316));
    Span4Mux_v I__5749 (
            .O(N__53321),
            .I(N__53311));
    Span4Mux_v I__5748 (
            .O(N__53316),
            .I(N__53311));
    Odrv4 I__5747 (
            .O(N__53311),
            .I(N_12_i));
    InMux I__5746 (
            .O(N__53308),
            .I(N__53305));
    LocalMux I__5745 (
            .O(N__53305),
            .I(shift_srl_1Z0Z_13));
    InMux I__5744 (
            .O(N__53302),
            .I(N__53299));
    LocalMux I__5743 (
            .O(N__53299),
            .I(shift_srl_1Z0Z_12));
    InMux I__5742 (
            .O(N__53296),
            .I(N__53293));
    LocalMux I__5741 (
            .O(N__53293),
            .I(shift_srl_1Z0Z_11));
    InMux I__5740 (
            .O(N__53290),
            .I(N__53287));
    LocalMux I__5739 (
            .O(N__53287),
            .I(shift_srl_116Z0Z_3));
    InMux I__5738 (
            .O(N__53284),
            .I(N__53281));
    LocalMux I__5737 (
            .O(N__53281),
            .I(shift_srl_116Z0Z_4));
    InMux I__5736 (
            .O(N__53278),
            .I(N__53275));
    LocalMux I__5735 (
            .O(N__53275),
            .I(shift_srl_116Z0Z_5));
    InMux I__5734 (
            .O(N__53272),
            .I(N__53269));
    LocalMux I__5733 (
            .O(N__53269),
            .I(shift_srl_116Z0Z_6));
    InMux I__5732 (
            .O(N__53266),
            .I(N__53263));
    LocalMux I__5731 (
            .O(N__53263),
            .I(shift_srl_116Z0Z_7));
    IoInMux I__5730 (
            .O(N__53260),
            .I(N__53257));
    LocalMux I__5729 (
            .O(N__53257),
            .I(N__53254));
    Span4Mux_s0_v I__5728 (
            .O(N__53254),
            .I(N__53251));
    Span4Mux_v I__5727 (
            .O(N__53251),
            .I(N__53248));
    Span4Mux_v I__5726 (
            .O(N__53248),
            .I(N__53245));
    Odrv4 I__5725 (
            .O(N__53245),
            .I(rco_c_113));
    InMux I__5724 (
            .O(N__53242),
            .I(N__53239));
    LocalMux I__5723 (
            .O(N__53239),
            .I(shift_srl_107Z0Z_0));
    IoInMux I__5722 (
            .O(N__53236),
            .I(N__53233));
    LocalMux I__5721 (
            .O(N__53233),
            .I(N__53230));
    Span12Mux_s1_v I__5720 (
            .O(N__53230),
            .I(N__53227));
    Odrv12 I__5719 (
            .O(N__53227),
            .I(rco_c_164));
    InMux I__5718 (
            .O(N__53224),
            .I(N__53221));
    LocalMux I__5717 (
            .O(N__53221),
            .I(shift_srl_135Z0Z_2));
    InMux I__5716 (
            .O(N__53218),
            .I(N__53215));
    LocalMux I__5715 (
            .O(N__53215),
            .I(shift_srl_135Z0Z_3));
    InMux I__5714 (
            .O(N__53212),
            .I(N__53209));
    LocalMux I__5713 (
            .O(N__53209),
            .I(shift_srl_135Z0Z_4));
    InMux I__5712 (
            .O(N__53206),
            .I(N__53203));
    LocalMux I__5711 (
            .O(N__53203),
            .I(shift_srl_135Z0Z_0));
    InMux I__5710 (
            .O(N__53200),
            .I(N__53197));
    LocalMux I__5709 (
            .O(N__53197),
            .I(shift_srl_135Z0Z_1));
    InMux I__5708 (
            .O(N__53194),
            .I(N__53191));
    LocalMux I__5707 (
            .O(N__53191),
            .I(shift_srl_135Z0Z_5));
    InMux I__5706 (
            .O(N__53188),
            .I(N__53185));
    LocalMux I__5705 (
            .O(N__53185),
            .I(shift_srl_135Z0Z_6));
    InMux I__5704 (
            .O(N__53182),
            .I(N__53179));
    LocalMux I__5703 (
            .O(N__53179),
            .I(shift_srl_135Z0Z_7));
    CEMux I__5702 (
            .O(N__53176),
            .I(N__53172));
    CEMux I__5701 (
            .O(N__53175),
            .I(N__53169));
    LocalMux I__5700 (
            .O(N__53172),
            .I(N__53166));
    LocalMux I__5699 (
            .O(N__53169),
            .I(N__53163));
    Odrv4 I__5698 (
            .O(N__53166),
            .I(clk_en_135));
    Odrv4 I__5697 (
            .O(N__53163),
            .I(clk_en_135));
    InMux I__5696 (
            .O(N__53158),
            .I(N__53155));
    LocalMux I__5695 (
            .O(N__53155),
            .I(shift_srl_116Z0Z_0));
    InMux I__5694 (
            .O(N__53152),
            .I(N__53149));
    LocalMux I__5693 (
            .O(N__53149),
            .I(shift_srl_116Z0Z_1));
    InMux I__5692 (
            .O(N__53146),
            .I(N__53143));
    LocalMux I__5691 (
            .O(N__53143),
            .I(shift_srl_116Z0Z_2));
    InMux I__5690 (
            .O(N__53140),
            .I(N__53137));
    LocalMux I__5689 (
            .O(N__53137),
            .I(g0_10_0));
    CascadeMux I__5688 (
            .O(N__53134),
            .I(g0_9_2_cascade_));
    InMux I__5687 (
            .O(N__53131),
            .I(N__53128));
    LocalMux I__5686 (
            .O(N__53128),
            .I(N__53125));
    Span4Mux_v I__5685 (
            .O(N__53125),
            .I(N__53122));
    Odrv4 I__5684 (
            .O(N__53122),
            .I(g0_11_1));
    CascadeMux I__5683 (
            .O(N__53119),
            .I(g0_12_0_cascade_));
    InMux I__5682 (
            .O(N__53116),
            .I(N__53113));
    LocalMux I__5681 (
            .O(N__53113),
            .I(g0_16_2));
    InMux I__5680 (
            .O(N__53110),
            .I(N__53107));
    LocalMux I__5679 (
            .O(N__53107),
            .I(shift_srl_135Z0Z_8));
    InMux I__5678 (
            .O(N__53104),
            .I(N__53100));
    InMux I__5677 (
            .O(N__53103),
            .I(N__53096));
    LocalMux I__5676 (
            .O(N__53100),
            .I(N__53092));
    CascadeMux I__5675 (
            .O(N__53099),
            .I(N__53089));
    LocalMux I__5674 (
            .O(N__53096),
            .I(N__53086));
    InMux I__5673 (
            .O(N__53095),
            .I(N__53082));
    Span4Mux_h I__5672 (
            .O(N__53092),
            .I(N__53079));
    InMux I__5671 (
            .O(N__53089),
            .I(N__53076));
    Span4Mux_v I__5670 (
            .O(N__53086),
            .I(N__53073));
    InMux I__5669 (
            .O(N__53085),
            .I(N__53070));
    LocalMux I__5668 (
            .O(N__53082),
            .I(shift_srl_135Z0Z_15));
    Odrv4 I__5667 (
            .O(N__53079),
            .I(shift_srl_135Z0Z_15));
    LocalMux I__5666 (
            .O(N__53076),
            .I(shift_srl_135Z0Z_15));
    Odrv4 I__5665 (
            .O(N__53073),
            .I(shift_srl_135Z0Z_15));
    LocalMux I__5664 (
            .O(N__53070),
            .I(shift_srl_135Z0Z_15));
    InMux I__5663 (
            .O(N__53059),
            .I(N__53056));
    LocalMux I__5662 (
            .O(N__53056),
            .I(shift_srl_134Z0Z_0));
    InMux I__5661 (
            .O(N__53053),
            .I(N__53050));
    LocalMux I__5660 (
            .O(N__53050),
            .I(shift_srl_134Z0Z_1));
    InMux I__5659 (
            .O(N__53047),
            .I(N__53044));
    LocalMux I__5658 (
            .O(N__53044),
            .I(shift_srl_134Z0Z_2));
    InMux I__5657 (
            .O(N__53041),
            .I(N__53038));
    LocalMux I__5656 (
            .O(N__53038),
            .I(shift_srl_134Z0Z_3));
    InMux I__5655 (
            .O(N__53035),
            .I(N__53032));
    LocalMux I__5654 (
            .O(N__53032),
            .I(shift_srl_134Z0Z_4));
    InMux I__5653 (
            .O(N__53029),
            .I(N__53026));
    LocalMux I__5652 (
            .O(N__53026),
            .I(shift_srl_134Z0Z_5));
    InMux I__5651 (
            .O(N__53023),
            .I(N__53020));
    LocalMux I__5650 (
            .O(N__53020),
            .I(shift_srl_134Z0Z_6));
    InMux I__5649 (
            .O(N__53017),
            .I(N__53014));
    LocalMux I__5648 (
            .O(N__53014),
            .I(N__53011));
    Span4Mux_h I__5647 (
            .O(N__53011),
            .I(N__53008));
    Odrv4 I__5646 (
            .O(N__53008),
            .I(shift_srl_134Z0Z_7));
    CEMux I__5645 (
            .O(N__53005),
            .I(N__53000));
    CEMux I__5644 (
            .O(N__53004),
            .I(N__52997));
    CEMux I__5643 (
            .O(N__53003),
            .I(N__52994));
    LocalMux I__5642 (
            .O(N__53000),
            .I(clk_en_134));
    LocalMux I__5641 (
            .O(N__52997),
            .I(clk_en_134));
    LocalMux I__5640 (
            .O(N__52994),
            .I(clk_en_134));
    InMux I__5639 (
            .O(N__52987),
            .I(N__52984));
    LocalMux I__5638 (
            .O(N__52984),
            .I(shift_srl_132Z0Z_4));
    InMux I__5637 (
            .O(N__52981),
            .I(N__52978));
    LocalMux I__5636 (
            .O(N__52978),
            .I(shift_srl_132Z0Z_5));
    InMux I__5635 (
            .O(N__52975),
            .I(N__52972));
    LocalMux I__5634 (
            .O(N__52972),
            .I(shift_srl_132Z0Z_6));
    InMux I__5633 (
            .O(N__52969),
            .I(N__52966));
    LocalMux I__5632 (
            .O(N__52966),
            .I(shift_srl_132Z0Z_7));
    InMux I__5631 (
            .O(N__52963),
            .I(N__52960));
    LocalMux I__5630 (
            .O(N__52960),
            .I(shift_srl_132Z0Z_14));
    CascadeMux I__5629 (
            .O(N__52957),
            .I(g0_43_1_cascade_));
    CEMux I__5628 (
            .O(N__52954),
            .I(N__52949));
    CEMux I__5627 (
            .O(N__52953),
            .I(N__52946));
    CEMux I__5626 (
            .O(N__52952),
            .I(N__52943));
    LocalMux I__5625 (
            .O(N__52949),
            .I(clk_en_132));
    LocalMux I__5624 (
            .O(N__52946),
            .I(clk_en_132));
    LocalMux I__5623 (
            .O(N__52943),
            .I(clk_en_132));
    InMux I__5622 (
            .O(N__52936),
            .I(N__52933));
    LocalMux I__5621 (
            .O(N__52933),
            .I(N__52924));
    CascadeMux I__5620 (
            .O(N__52932),
            .I(N__52921));
    CascadeMux I__5619 (
            .O(N__52931),
            .I(N__52918));
    InMux I__5618 (
            .O(N__52930),
            .I(N__52914));
    InMux I__5617 (
            .O(N__52929),
            .I(N__52905));
    InMux I__5616 (
            .O(N__52928),
            .I(N__52905));
    InMux I__5615 (
            .O(N__52927),
            .I(N__52902));
    Span4Mux_h I__5614 (
            .O(N__52924),
            .I(N__52899));
    InMux I__5613 (
            .O(N__52921),
            .I(N__52892));
    InMux I__5612 (
            .O(N__52918),
            .I(N__52892));
    InMux I__5611 (
            .O(N__52917),
            .I(N__52892));
    LocalMux I__5610 (
            .O(N__52914),
            .I(N__52889));
    InMux I__5609 (
            .O(N__52913),
            .I(N__52884));
    InMux I__5608 (
            .O(N__52912),
            .I(N__52884));
    InMux I__5607 (
            .O(N__52911),
            .I(N__52879));
    InMux I__5606 (
            .O(N__52910),
            .I(N__52879));
    LocalMux I__5605 (
            .O(N__52905),
            .I(N__52876));
    LocalMux I__5604 (
            .O(N__52902),
            .I(shift_srl_130Z0Z_15));
    Odrv4 I__5603 (
            .O(N__52899),
            .I(shift_srl_130Z0Z_15));
    LocalMux I__5602 (
            .O(N__52892),
            .I(shift_srl_130Z0Z_15));
    Odrv4 I__5601 (
            .O(N__52889),
            .I(shift_srl_130Z0Z_15));
    LocalMux I__5600 (
            .O(N__52884),
            .I(shift_srl_130Z0Z_15));
    LocalMux I__5599 (
            .O(N__52879),
            .I(shift_srl_130Z0Z_15));
    Odrv4 I__5598 (
            .O(N__52876),
            .I(shift_srl_130Z0Z_15));
    CascadeMux I__5597 (
            .O(N__52861),
            .I(shift_srl_132_RNI731TZ0Z_15_cascade_));
    CascadeMux I__5596 (
            .O(N__52858),
            .I(rco_int_0_a3_0_a2_0_132_cascade_));
    InMux I__5595 (
            .O(N__52855),
            .I(N__52852));
    LocalMux I__5594 (
            .O(N__52852),
            .I(shift_srl_8Z0Z_14));
    InMux I__5593 (
            .O(N__52849),
            .I(N__52846));
    LocalMux I__5592 (
            .O(N__52846),
            .I(shift_srl_8Z0Z_8));
    InMux I__5591 (
            .O(N__52843),
            .I(N__52840));
    LocalMux I__5590 (
            .O(N__52840),
            .I(shift_srl_8Z0Z_9));
    CEMux I__5589 (
            .O(N__52837),
            .I(N__52833));
    CEMux I__5588 (
            .O(N__52836),
            .I(N__52830));
    LocalMux I__5587 (
            .O(N__52833),
            .I(N__52826));
    LocalMux I__5586 (
            .O(N__52830),
            .I(N__52823));
    CEMux I__5585 (
            .O(N__52829),
            .I(N__52820));
    Span4Mux_h I__5584 (
            .O(N__52826),
            .I(N__52817));
    Span4Mux_h I__5583 (
            .O(N__52823),
            .I(N__52814));
    LocalMux I__5582 (
            .O(N__52820),
            .I(N__52811));
    Odrv4 I__5581 (
            .O(N__52817),
            .I(clk_en_8));
    Odrv4 I__5580 (
            .O(N__52814),
            .I(clk_en_8));
    Odrv4 I__5579 (
            .O(N__52811),
            .I(clk_en_8));
    InMux I__5578 (
            .O(N__52804),
            .I(N__52801));
    LocalMux I__5577 (
            .O(N__52801),
            .I(shift_srl_128Z0Z_7));
    InMux I__5576 (
            .O(N__52798),
            .I(N__52795));
    LocalMux I__5575 (
            .O(N__52795),
            .I(shift_srl_132Z0Z_0));
    InMux I__5574 (
            .O(N__52792),
            .I(N__52789));
    LocalMux I__5573 (
            .O(N__52789),
            .I(shift_srl_132Z0Z_1));
    InMux I__5572 (
            .O(N__52786),
            .I(N__52783));
    LocalMux I__5571 (
            .O(N__52783),
            .I(shift_srl_132Z0Z_2));
    InMux I__5570 (
            .O(N__52780),
            .I(N__52777));
    LocalMux I__5569 (
            .O(N__52777),
            .I(shift_srl_132Z0Z_3));
    InMux I__5568 (
            .O(N__52774),
            .I(N__52771));
    LocalMux I__5567 (
            .O(N__52771),
            .I(shift_srl_9Z0Z_2));
    InMux I__5566 (
            .O(N__52768),
            .I(N__52765));
    LocalMux I__5565 (
            .O(N__52765),
            .I(shift_srl_9Z0Z_3));
    InMux I__5564 (
            .O(N__52762),
            .I(N__52759));
    LocalMux I__5563 (
            .O(N__52759),
            .I(shift_srl_9Z0Z_4));
    InMux I__5562 (
            .O(N__52756),
            .I(N__52753));
    LocalMux I__5561 (
            .O(N__52753),
            .I(shift_srl_9Z0Z_5));
    InMux I__5560 (
            .O(N__52750),
            .I(N__52747));
    LocalMux I__5559 (
            .O(N__52747),
            .I(shift_srl_8Z0Z_10));
    InMux I__5558 (
            .O(N__52744),
            .I(N__52741));
    LocalMux I__5557 (
            .O(N__52741),
            .I(shift_srl_8Z0Z_11));
    InMux I__5556 (
            .O(N__52738),
            .I(N__52735));
    LocalMux I__5555 (
            .O(N__52735),
            .I(shift_srl_8Z0Z_12));
    InMux I__5554 (
            .O(N__52732),
            .I(N__52729));
    LocalMux I__5553 (
            .O(N__52729),
            .I(shift_srl_8Z0Z_13));
    InMux I__5552 (
            .O(N__52726),
            .I(N__52723));
    LocalMux I__5551 (
            .O(N__52723),
            .I(shift_srl_17Z0Z_11));
    InMux I__5550 (
            .O(N__52720),
            .I(N__52717));
    LocalMux I__5549 (
            .O(N__52717),
            .I(shift_srl_17Z0Z_12));
    InMux I__5548 (
            .O(N__52714),
            .I(N__52711));
    LocalMux I__5547 (
            .O(N__52711),
            .I(shift_srl_17Z0Z_13));
    InMux I__5546 (
            .O(N__52708),
            .I(N__52705));
    LocalMux I__5545 (
            .O(N__52705),
            .I(N__52702));
    Span4Mux_v I__5544 (
            .O(N__52702),
            .I(N__52699));
    Odrv4 I__5543 (
            .O(N__52699),
            .I(shift_srl_17Z0Z_14));
    InMux I__5542 (
            .O(N__52696),
            .I(N__52693));
    LocalMux I__5541 (
            .O(N__52693),
            .I(shift_srl_17Z0Z_9));
    InMux I__5540 (
            .O(N__52690),
            .I(N__52687));
    LocalMux I__5539 (
            .O(N__52687),
            .I(shift_srl_17Z0Z_7));
    InMux I__5538 (
            .O(N__52684),
            .I(N__52681));
    LocalMux I__5537 (
            .O(N__52681),
            .I(shift_srl_17Z0Z_8));
    CEMux I__5536 (
            .O(N__52678),
            .I(N__52673));
    CEMux I__5535 (
            .O(N__52677),
            .I(N__52670));
    CEMux I__5534 (
            .O(N__52676),
            .I(N__52667));
    LocalMux I__5533 (
            .O(N__52673),
            .I(N__52664));
    LocalMux I__5532 (
            .O(N__52670),
            .I(N__52659));
    LocalMux I__5531 (
            .O(N__52667),
            .I(N__52659));
    Span4Mux_v I__5530 (
            .O(N__52664),
            .I(N__52656));
    Span4Mux_h I__5529 (
            .O(N__52659),
            .I(N__52653));
    Span4Mux_h I__5528 (
            .O(N__52656),
            .I(N__52650));
    Span4Mux_s3_h I__5527 (
            .O(N__52653),
            .I(N__52647));
    Odrv4 I__5526 (
            .O(N__52650),
            .I(clk_en_17));
    Odrv4 I__5525 (
            .O(N__52647),
            .I(clk_en_17));
    InMux I__5524 (
            .O(N__52642),
            .I(N__52638));
    IoInMux I__5523 (
            .O(N__52641),
            .I(N__52635));
    LocalMux I__5522 (
            .O(N__52638),
            .I(N__52632));
    LocalMux I__5521 (
            .O(N__52635),
            .I(N__52629));
    Span4Mux_h I__5520 (
            .O(N__52632),
            .I(N__52626));
    Odrv4 I__5519 (
            .O(N__52629),
            .I(rco_c_8));
    Odrv4 I__5518 (
            .O(N__52626),
            .I(rco_c_8));
    InMux I__5517 (
            .O(N__52621),
            .I(N__52618));
    LocalMux I__5516 (
            .O(N__52618),
            .I(shift_srl_9Z0Z_0));
    InMux I__5515 (
            .O(N__52615),
            .I(N__52612));
    LocalMux I__5514 (
            .O(N__52612),
            .I(shift_srl_9Z0Z_1));
    InMux I__5513 (
            .O(N__52609),
            .I(N__52606));
    LocalMux I__5512 (
            .O(N__52606),
            .I(shift_srl_17Z0Z_0));
    InMux I__5511 (
            .O(N__52603),
            .I(N__52600));
    LocalMux I__5510 (
            .O(N__52600),
            .I(shift_srl_17Z0Z_1));
    InMux I__5509 (
            .O(N__52597),
            .I(N__52594));
    LocalMux I__5508 (
            .O(N__52594),
            .I(shift_srl_17Z0Z_2));
    InMux I__5507 (
            .O(N__52591),
            .I(N__52588));
    LocalMux I__5506 (
            .O(N__52588),
            .I(shift_srl_17Z0Z_3));
    InMux I__5505 (
            .O(N__52585),
            .I(N__52582));
    LocalMux I__5504 (
            .O(N__52582),
            .I(shift_srl_17Z0Z_4));
    InMux I__5503 (
            .O(N__52579),
            .I(N__52576));
    LocalMux I__5502 (
            .O(N__52576),
            .I(shift_srl_17Z0Z_5));
    InMux I__5501 (
            .O(N__52573),
            .I(N__52570));
    LocalMux I__5500 (
            .O(N__52570),
            .I(shift_srl_17Z0Z_6));
    InMux I__5499 (
            .O(N__52567),
            .I(N__52564));
    LocalMux I__5498 (
            .O(N__52564),
            .I(shift_srl_17Z0Z_10));
    InMux I__5497 (
            .O(N__52561),
            .I(N__52554));
    InMux I__5496 (
            .O(N__52560),
            .I(N__52551));
    InMux I__5495 (
            .O(N__52559),
            .I(N__52544));
    InMux I__5494 (
            .O(N__52558),
            .I(N__52544));
    InMux I__5493 (
            .O(N__52557),
            .I(N__52544));
    LocalMux I__5492 (
            .O(N__52554),
            .I(N__52540));
    LocalMux I__5491 (
            .O(N__52551),
            .I(N__52535));
    LocalMux I__5490 (
            .O(N__52544),
            .I(N__52535));
    InMux I__5489 (
            .O(N__52543),
            .I(N__52532));
    Span4Mux_h I__5488 (
            .O(N__52540),
            .I(N__52529));
    Span4Mux_h I__5487 (
            .O(N__52535),
            .I(N__52526));
    LocalMux I__5486 (
            .O(N__52532),
            .I(shift_srl_19Z0Z_15));
    Odrv4 I__5485 (
            .O(N__52529),
            .I(shift_srl_19Z0Z_15));
    Odrv4 I__5484 (
            .O(N__52526),
            .I(shift_srl_19Z0Z_15));
    InMux I__5483 (
            .O(N__52519),
            .I(N__52516));
    LocalMux I__5482 (
            .O(N__52516),
            .I(shift_srl_19Z0Z_0));
    InMux I__5481 (
            .O(N__52513),
            .I(N__52510));
    LocalMux I__5480 (
            .O(N__52510),
            .I(shift_srl_19Z0Z_1));
    InMux I__5479 (
            .O(N__52507),
            .I(N__52504));
    LocalMux I__5478 (
            .O(N__52504),
            .I(shift_srl_19Z0Z_2));
    InMux I__5477 (
            .O(N__52501),
            .I(N__52498));
    LocalMux I__5476 (
            .O(N__52498),
            .I(shift_srl_19Z0Z_3));
    InMux I__5475 (
            .O(N__52495),
            .I(N__52492));
    LocalMux I__5474 (
            .O(N__52492),
            .I(shift_srl_19Z0Z_4));
    InMux I__5473 (
            .O(N__52489),
            .I(N__52486));
    LocalMux I__5472 (
            .O(N__52486),
            .I(shift_srl_19Z0Z_5));
    InMux I__5471 (
            .O(N__52483),
            .I(N__52480));
    LocalMux I__5470 (
            .O(N__52480),
            .I(shift_srl_19Z0Z_11));
    InMux I__5469 (
            .O(N__52477),
            .I(N__52474));
    LocalMux I__5468 (
            .O(N__52474),
            .I(shift_srl_19Z0Z_12));
    InMux I__5467 (
            .O(N__52471),
            .I(N__52468));
    LocalMux I__5466 (
            .O(N__52468),
            .I(shift_srl_19Z0Z_13));
    CEMux I__5465 (
            .O(N__52465),
            .I(N__52461));
    CEMux I__5464 (
            .O(N__52464),
            .I(N__52458));
    LocalMux I__5463 (
            .O(N__52461),
            .I(N__52455));
    LocalMux I__5462 (
            .O(N__52458),
            .I(N__52452));
    Span4Mux_h I__5461 (
            .O(N__52455),
            .I(N__52449));
    Span4Mux_h I__5460 (
            .O(N__52452),
            .I(N__52446));
    Odrv4 I__5459 (
            .O(N__52449),
            .I(clk_en_19));
    Odrv4 I__5458 (
            .O(N__52446),
            .I(clk_en_19));
    InMux I__5457 (
            .O(N__52441),
            .I(N__52435));
    InMux I__5456 (
            .O(N__52440),
            .I(N__52432));
    CascadeMux I__5455 (
            .O(N__52439),
            .I(N__52426));
    InMux I__5454 (
            .O(N__52438),
            .I(N__52423));
    LocalMux I__5453 (
            .O(N__52435),
            .I(N__52418));
    LocalMux I__5452 (
            .O(N__52432),
            .I(N__52418));
    InMux I__5451 (
            .O(N__52431),
            .I(N__52415));
    InMux I__5450 (
            .O(N__52430),
            .I(N__52410));
    InMux I__5449 (
            .O(N__52429),
            .I(N__52410));
    InMux I__5448 (
            .O(N__52426),
            .I(N__52407));
    LocalMux I__5447 (
            .O(N__52423),
            .I(shift_srl_17Z0Z_15));
    Odrv12 I__5446 (
            .O(N__52418),
            .I(shift_srl_17Z0Z_15));
    LocalMux I__5445 (
            .O(N__52415),
            .I(shift_srl_17Z0Z_15));
    LocalMux I__5444 (
            .O(N__52410),
            .I(shift_srl_17Z0Z_15));
    LocalMux I__5443 (
            .O(N__52407),
            .I(shift_srl_17Z0Z_15));
    InMux I__5442 (
            .O(N__52396),
            .I(N__52393));
    LocalMux I__5441 (
            .O(N__52393),
            .I(shift_srl_23Z0Z_8));
    InMux I__5440 (
            .O(N__52390),
            .I(N__52387));
    LocalMux I__5439 (
            .O(N__52387),
            .I(shift_srl_23Z0Z_7));
    InMux I__5438 (
            .O(N__52384),
            .I(N__52381));
    LocalMux I__5437 (
            .O(N__52381),
            .I(shift_srl_19Z0Z_10));
    InMux I__5436 (
            .O(N__52378),
            .I(N__52375));
    LocalMux I__5435 (
            .O(N__52375),
            .I(shift_srl_19Z0Z_6));
    InMux I__5434 (
            .O(N__52372),
            .I(N__52369));
    LocalMux I__5433 (
            .O(N__52369),
            .I(shift_srl_19Z0Z_14));
    InMux I__5432 (
            .O(N__52366),
            .I(N__52363));
    LocalMux I__5431 (
            .O(N__52363),
            .I(shift_srl_19Z0Z_9));
    InMux I__5430 (
            .O(N__52360),
            .I(N__52357));
    LocalMux I__5429 (
            .O(N__52357),
            .I(shift_srl_19Z0Z_7));
    InMux I__5428 (
            .O(N__52354),
            .I(N__52351));
    LocalMux I__5427 (
            .O(N__52351),
            .I(shift_srl_19Z0Z_8));
    InMux I__5426 (
            .O(N__52348),
            .I(N__52344));
    InMux I__5425 (
            .O(N__52347),
            .I(N__52341));
    LocalMux I__5424 (
            .O(N__52344),
            .I(N__52336));
    LocalMux I__5423 (
            .O(N__52341),
            .I(N__52336));
    Span4Mux_h I__5422 (
            .O(N__52336),
            .I(N__52333));
    Odrv4 I__5421 (
            .O(N__52333),
            .I(shift_srl_7_RNI00TC1Z0Z_15));
    CascadeMux I__5420 (
            .O(N__52330),
            .I(N_453_cascade_));
    IoInMux I__5419 (
            .O(N__52327),
            .I(N__52324));
    LocalMux I__5418 (
            .O(N__52324),
            .I(N__52321));
    IoSpan4Mux I__5417 (
            .O(N__52321),
            .I(N__52318));
    IoSpan4Mux I__5416 (
            .O(N__52318),
            .I(N__52315));
    IoSpan4Mux I__5415 (
            .O(N__52315),
            .I(N__52312));
    Span4Mux_s3_h I__5414 (
            .O(N__52312),
            .I(N__52308));
    InMux I__5413 (
            .O(N__52311),
            .I(N__52305));
    Odrv4 I__5412 (
            .O(N__52308),
            .I(rco_c_10));
    LocalMux I__5411 (
            .O(N__52305),
            .I(rco_c_10));
    InMux I__5410 (
            .O(N__52300),
            .I(N__52295));
    InMux I__5409 (
            .O(N__52299),
            .I(N__52290));
    InMux I__5408 (
            .O(N__52298),
            .I(N__52290));
    LocalMux I__5407 (
            .O(N__52295),
            .I(shift_srl_2Z0Z_15));
    LocalMux I__5406 (
            .O(N__52290),
            .I(shift_srl_2Z0Z_15));
    IoInMux I__5405 (
            .O(N__52285),
            .I(N__52282));
    LocalMux I__5404 (
            .O(N__52282),
            .I(N__52279));
    Span4Mux_s2_h I__5403 (
            .O(N__52279),
            .I(N__52276));
    Sp12to4 I__5402 (
            .O(N__52276),
            .I(N__52273));
    Span12Mux_v I__5401 (
            .O(N__52273),
            .I(N__52270));
    Odrv12 I__5400 (
            .O(N__52270),
            .I(N_453_i));
    InMux I__5399 (
            .O(N__52267),
            .I(N__52264));
    LocalMux I__5398 (
            .O(N__52264),
            .I(shift_srl_23Z0Z_10));
    InMux I__5397 (
            .O(N__52261),
            .I(N__52258));
    LocalMux I__5396 (
            .O(N__52258),
            .I(shift_srl_23Z0Z_11));
    InMux I__5395 (
            .O(N__52255),
            .I(N__52252));
    LocalMux I__5394 (
            .O(N__52252),
            .I(shift_srl_23Z0Z_12));
    InMux I__5393 (
            .O(N__52249),
            .I(N__52246));
    LocalMux I__5392 (
            .O(N__52246),
            .I(shift_srl_23Z0Z_13));
    InMux I__5391 (
            .O(N__52243),
            .I(N__52240));
    LocalMux I__5390 (
            .O(N__52240),
            .I(shift_srl_23Z0Z_9));
    InMux I__5389 (
            .O(N__52237),
            .I(N__52234));
    LocalMux I__5388 (
            .O(N__52234),
            .I(shift_srl_2Z0Z_3));
    InMux I__5387 (
            .O(N__52231),
            .I(N__52228));
    LocalMux I__5386 (
            .O(N__52228),
            .I(shift_srl_2Z0Z_4));
    InMux I__5385 (
            .O(N__52225),
            .I(N__52222));
    LocalMux I__5384 (
            .O(N__52222),
            .I(shift_srl_2Z0Z_5));
    InMux I__5383 (
            .O(N__52219),
            .I(N__52216));
    LocalMux I__5382 (
            .O(N__52216),
            .I(shift_srl_2Z0Z_6));
    InMux I__5381 (
            .O(N__52213),
            .I(N__52210));
    LocalMux I__5380 (
            .O(N__52210),
            .I(shift_srl_2Z0Z_7));
    CEMux I__5379 (
            .O(N__52207),
            .I(N__52203));
    CEMux I__5378 (
            .O(N__52206),
            .I(N__52198));
    LocalMux I__5377 (
            .O(N__52203),
            .I(N__52194));
    CEMux I__5376 (
            .O(N__52202),
            .I(N__52191));
    CEMux I__5375 (
            .O(N__52201),
            .I(N__52188));
    LocalMux I__5374 (
            .O(N__52198),
            .I(N__52185));
    CEMux I__5373 (
            .O(N__52197),
            .I(N__52182));
    Span4Mux_s2_h I__5372 (
            .O(N__52194),
            .I(N__52177));
    LocalMux I__5371 (
            .O(N__52191),
            .I(N__52177));
    LocalMux I__5370 (
            .O(N__52188),
            .I(N__52174));
    Span4Mux_v I__5369 (
            .O(N__52185),
            .I(N__52171));
    LocalMux I__5368 (
            .O(N__52182),
            .I(N__52168));
    Span4Mux_h I__5367 (
            .O(N__52177),
            .I(N__52165));
    Span12Mux_s8_v I__5366 (
            .O(N__52174),
            .I(N__52162));
    Span4Mux_h I__5365 (
            .O(N__52171),
            .I(N__52157));
    Span4Mux_v I__5364 (
            .O(N__52168),
            .I(N__52157));
    Odrv4 I__5363 (
            .O(N__52165),
            .I(N_701));
    Odrv12 I__5362 (
            .O(N__52162),
            .I(N_701));
    Odrv4 I__5361 (
            .O(N__52157),
            .I(N_701));
    CascadeMux I__5360 (
            .O(N__52150),
            .I(shift_srl_10_RNIQHCJ1Z0Z_15_cascade_));
    IoInMux I__5359 (
            .O(N__52147),
            .I(N__52144));
    LocalMux I__5358 (
            .O(N__52144),
            .I(N__52140));
    InMux I__5357 (
            .O(N__52143),
            .I(N__52137));
    Span12Mux_s11_h I__5356 (
            .O(N__52140),
            .I(N__52134));
    LocalMux I__5355 (
            .O(N__52137),
            .I(N__52131));
    Span12Mux_v I__5354 (
            .O(N__52134),
            .I(N__52127));
    Span12Mux_s5_h I__5353 (
            .O(N__52131),
            .I(N__52124));
    InMux I__5352 (
            .O(N__52130),
            .I(N__52121));
    Odrv12 I__5351 (
            .O(N__52127),
            .I(rco_c_21));
    Odrv12 I__5350 (
            .O(N__52124),
            .I(rco_c_21));
    LocalMux I__5349 (
            .O(N__52121),
            .I(rco_c_21));
    CascadeMux I__5348 (
            .O(N__52114),
            .I(rco_c_21_cascade_));
    InMux I__5347 (
            .O(N__52111),
            .I(N__52108));
    LocalMux I__5346 (
            .O(N__52108),
            .I(shift_srl_2Z0Z_14));
    InMux I__5345 (
            .O(N__52105),
            .I(N__52102));
    LocalMux I__5344 (
            .O(N__52102),
            .I(shift_srl_2Z0Z_11));
    InMux I__5343 (
            .O(N__52099),
            .I(N__52096));
    LocalMux I__5342 (
            .O(N__52096),
            .I(shift_srl_2Z0Z_12));
    InMux I__5341 (
            .O(N__52093),
            .I(N__52090));
    LocalMux I__5340 (
            .O(N__52090),
            .I(shift_srl_2Z0Z_8));
    InMux I__5339 (
            .O(N__52087),
            .I(N__52084));
    LocalMux I__5338 (
            .O(N__52084),
            .I(shift_srl_2Z0Z_9));
    InMux I__5337 (
            .O(N__52081),
            .I(N__52078));
    LocalMux I__5336 (
            .O(N__52078),
            .I(shift_srl_2Z0Z_2));
    InMux I__5335 (
            .O(N__52075),
            .I(N__52072));
    LocalMux I__5334 (
            .O(N__52072),
            .I(shift_srl_2Z0Z_0));
    InMux I__5333 (
            .O(N__52069),
            .I(N__52066));
    LocalMux I__5332 (
            .O(N__52066),
            .I(shift_srl_2Z0Z_1));
    InMux I__5331 (
            .O(N__52063),
            .I(N__52060));
    LocalMux I__5330 (
            .O(N__52060),
            .I(shift_srl_2Z0Z_13));
    InMux I__5329 (
            .O(N__52057),
            .I(N__52054));
    LocalMux I__5328 (
            .O(N__52054),
            .I(shift_srl_135Z0Z_12));
    InMux I__5327 (
            .O(N__52051),
            .I(N__52048));
    LocalMux I__5326 (
            .O(N__52048),
            .I(shift_srl_135Z0Z_13));
    InMux I__5325 (
            .O(N__52045),
            .I(N__52042));
    LocalMux I__5324 (
            .O(N__52042),
            .I(shift_srl_135Z0Z_14));
    InMux I__5323 (
            .O(N__52039),
            .I(N__52036));
    LocalMux I__5322 (
            .O(N__52036),
            .I(shift_srl_135Z0Z_9));
    InMux I__5321 (
            .O(N__52033),
            .I(N__52030));
    LocalMux I__5320 (
            .O(N__52030),
            .I(shift_srl_135Z0Z_10));
    InMux I__5319 (
            .O(N__52027),
            .I(N__52024));
    LocalMux I__5318 (
            .O(N__52024),
            .I(shift_srl_2Z0Z_10));
    InMux I__5317 (
            .O(N__52021),
            .I(N__52017));
    InMux I__5316 (
            .O(N__52020),
            .I(N__52012));
    LocalMux I__5315 (
            .O(N__52017),
            .I(N__52009));
    InMux I__5314 (
            .O(N__52016),
            .I(N__52003));
    InMux I__5313 (
            .O(N__52015),
            .I(N__52000));
    LocalMux I__5312 (
            .O(N__52012),
            .I(N__51997));
    Span4Mux_s3_h I__5311 (
            .O(N__52009),
            .I(N__51994));
    InMux I__5310 (
            .O(N__52008),
            .I(N__51987));
    InMux I__5309 (
            .O(N__52007),
            .I(N__51987));
    InMux I__5308 (
            .O(N__52006),
            .I(N__51987));
    LocalMux I__5307 (
            .O(N__52003),
            .I(shift_srl_134Z0Z_15));
    LocalMux I__5306 (
            .O(N__52000),
            .I(shift_srl_134Z0Z_15));
    Odrv12 I__5305 (
            .O(N__51997),
            .I(shift_srl_134Z0Z_15));
    Odrv4 I__5304 (
            .O(N__51994),
            .I(shift_srl_134Z0Z_15));
    LocalMux I__5303 (
            .O(N__51987),
            .I(shift_srl_134Z0Z_15));
    CascadeMux I__5302 (
            .O(N__51976),
            .I(g0_2_cascade_));
    CascadeMux I__5301 (
            .O(N__51973),
            .I(g0_13_0_cascade_));
    CascadeMux I__5300 (
            .O(N__51970),
            .I(g0_10_1_cascade_));
    InMux I__5299 (
            .O(N__51967),
            .I(N__51964));
    LocalMux I__5298 (
            .O(N__51964),
            .I(g0_14_0));
    InMux I__5297 (
            .O(N__51961),
            .I(N__51958));
    LocalMux I__5296 (
            .O(N__51958),
            .I(g0_12_1));
    InMux I__5295 (
            .O(N__51955),
            .I(N__51952));
    LocalMux I__5294 (
            .O(N__51952),
            .I(shift_srl_135Z0Z_11));
    InMux I__5293 (
            .O(N__51949),
            .I(N__51946));
    LocalMux I__5292 (
            .O(N__51946),
            .I(shift_srl_132Z0Z_8));
    InMux I__5291 (
            .O(N__51943),
            .I(N__51940));
    LocalMux I__5290 (
            .O(N__51940),
            .I(shift_srl_131Z0Z_10));
    InMux I__5289 (
            .O(N__51937),
            .I(N__51934));
    LocalMux I__5288 (
            .O(N__51934),
            .I(shift_srl_131Z0Z_11));
    InMux I__5287 (
            .O(N__51931),
            .I(N__51928));
    LocalMux I__5286 (
            .O(N__51928),
            .I(shift_srl_131Z0Z_12));
    InMux I__5285 (
            .O(N__51925),
            .I(N__51922));
    LocalMux I__5284 (
            .O(N__51922),
            .I(shift_srl_131Z0Z_13));
    InMux I__5283 (
            .O(N__51919),
            .I(N__51916));
    LocalMux I__5282 (
            .O(N__51916),
            .I(shift_srl_131Z0Z_14));
    InMux I__5281 (
            .O(N__51913),
            .I(N__51910));
    LocalMux I__5280 (
            .O(N__51910),
            .I(shift_srl_131Z0Z_8));
    InMux I__5279 (
            .O(N__51907),
            .I(N__51904));
    LocalMux I__5278 (
            .O(N__51904),
            .I(shift_srl_131Z0Z_9));
    InMux I__5277 (
            .O(N__51901),
            .I(N__51898));
    LocalMux I__5276 (
            .O(N__51898),
            .I(shift_srl_131Z0Z_0));
    InMux I__5275 (
            .O(N__51895),
            .I(N__51892));
    LocalMux I__5274 (
            .O(N__51892),
            .I(shift_srl_131Z0Z_1));
    CEMux I__5273 (
            .O(N__51889),
            .I(N__51885));
    CEMux I__5272 (
            .O(N__51888),
            .I(N__51882));
    LocalMux I__5271 (
            .O(N__51885),
            .I(N__51879));
    LocalMux I__5270 (
            .O(N__51882),
            .I(N__51876));
    Span4Mux_v I__5269 (
            .O(N__51879),
            .I(N__51873));
    Span4Mux_h I__5268 (
            .O(N__51876),
            .I(N__51870));
    Odrv4 I__5267 (
            .O(N__51873),
            .I(clk_en_131));
    Odrv4 I__5266 (
            .O(N__51870),
            .I(clk_en_131));
    InMux I__5265 (
            .O(N__51865),
            .I(N__51862));
    LocalMux I__5264 (
            .O(N__51862),
            .I(shift_srl_133Z0Z_7));
    InMux I__5263 (
            .O(N__51859),
            .I(N__51856));
    LocalMux I__5262 (
            .O(N__51856),
            .I(shift_srl_133Z0Z_10));
    InMux I__5261 (
            .O(N__51853),
            .I(N__51850));
    LocalMux I__5260 (
            .O(N__51850),
            .I(shift_srl_133Z0Z_8));
    InMux I__5259 (
            .O(N__51847),
            .I(N__51844));
    LocalMux I__5258 (
            .O(N__51844),
            .I(shift_srl_133Z0Z_9));
    InMux I__5257 (
            .O(N__51841),
            .I(N__51838));
    LocalMux I__5256 (
            .O(N__51838),
            .I(shift_srl_132Z0Z_10));
    InMux I__5255 (
            .O(N__51835),
            .I(N__51832));
    LocalMux I__5254 (
            .O(N__51832),
            .I(shift_srl_132Z0Z_11));
    InMux I__5253 (
            .O(N__51829),
            .I(N__51826));
    LocalMux I__5252 (
            .O(N__51826),
            .I(shift_srl_132Z0Z_12));
    InMux I__5251 (
            .O(N__51823),
            .I(N__51820));
    LocalMux I__5250 (
            .O(N__51820),
            .I(shift_srl_132Z0Z_13));
    InMux I__5249 (
            .O(N__51817),
            .I(N__51814));
    LocalMux I__5248 (
            .O(N__51814),
            .I(shift_srl_132Z0Z_9));
    InMux I__5247 (
            .O(N__51811),
            .I(N__51808));
    LocalMux I__5246 (
            .O(N__51808),
            .I(shift_srl_8Z0Z_3));
    InMux I__5245 (
            .O(N__51805),
            .I(N__51802));
    LocalMux I__5244 (
            .O(N__51802),
            .I(shift_srl_8Z0Z_6));
    InMux I__5243 (
            .O(N__51799),
            .I(N__51796));
    LocalMux I__5242 (
            .O(N__51796),
            .I(shift_srl_8Z0Z_4));
    InMux I__5241 (
            .O(N__51793),
            .I(N__51790));
    LocalMux I__5240 (
            .O(N__51790),
            .I(shift_srl_8Z0Z_5));
    InMux I__5239 (
            .O(N__51787),
            .I(N__51784));
    LocalMux I__5238 (
            .O(N__51784),
            .I(shift_srl_8Z0Z_7));
    InMux I__5237 (
            .O(N__51781),
            .I(N__51778));
    LocalMux I__5236 (
            .O(N__51778),
            .I(shift_srl_133Z0Z_4));
    InMux I__5235 (
            .O(N__51775),
            .I(N__51772));
    LocalMux I__5234 (
            .O(N__51772),
            .I(shift_srl_133Z0Z_5));
    InMux I__5233 (
            .O(N__51769),
            .I(N__51766));
    LocalMux I__5232 (
            .O(N__51766),
            .I(shift_srl_133Z0Z_6));
    InMux I__5231 (
            .O(N__51763),
            .I(N__51760));
    LocalMux I__5230 (
            .O(N__51760),
            .I(shift_srl_20Z0Z_13));
    InMux I__5229 (
            .O(N__51757),
            .I(N__51754));
    LocalMux I__5228 (
            .O(N__51754),
            .I(shift_srl_20Z0Z_14));
    InMux I__5227 (
            .O(N__51751),
            .I(N__51747));
    InMux I__5226 (
            .O(N__51750),
            .I(N__51742));
    LocalMux I__5225 (
            .O(N__51747),
            .I(N__51739));
    InMux I__5224 (
            .O(N__51746),
            .I(N__51734));
    InMux I__5223 (
            .O(N__51745),
            .I(N__51734));
    LocalMux I__5222 (
            .O(N__51742),
            .I(shift_srl_20Z0Z_15));
    Odrv4 I__5221 (
            .O(N__51739),
            .I(shift_srl_20Z0Z_15));
    LocalMux I__5220 (
            .O(N__51734),
            .I(shift_srl_20Z0Z_15));
    InMux I__5219 (
            .O(N__51727),
            .I(N__51724));
    LocalMux I__5218 (
            .O(N__51724),
            .I(shift_srl_20Z0Z_11));
    InMux I__5217 (
            .O(N__51721),
            .I(N__51718));
    LocalMux I__5216 (
            .O(N__51718),
            .I(shift_srl_20Z0Z_12));
    InMux I__5215 (
            .O(N__51715),
            .I(N__51712));
    LocalMux I__5214 (
            .O(N__51712),
            .I(shift_srl_20Z0Z_7));
    InMux I__5213 (
            .O(N__51709),
            .I(N__51706));
    LocalMux I__5212 (
            .O(N__51706),
            .I(shift_srl_20Z0Z_8));
    CEMux I__5211 (
            .O(N__51703),
            .I(N__51699));
    CEMux I__5210 (
            .O(N__51702),
            .I(N__51696));
    LocalMux I__5209 (
            .O(N__51699),
            .I(clk_en_20));
    LocalMux I__5208 (
            .O(N__51696),
            .I(clk_en_20));
    InMux I__5207 (
            .O(N__51691),
            .I(N__51687));
    IoInMux I__5206 (
            .O(N__51690),
            .I(N__51684));
    LocalMux I__5205 (
            .O(N__51687),
            .I(N__51681));
    LocalMux I__5204 (
            .O(N__51684),
            .I(N__51678));
    Span4Mux_h I__5203 (
            .O(N__51681),
            .I(N__51675));
    Odrv4 I__5202 (
            .O(N__51678),
            .I(rco_c_7));
    Odrv4 I__5201 (
            .O(N__51675),
            .I(rco_c_7));
    InMux I__5200 (
            .O(N__51670),
            .I(N__51667));
    LocalMux I__5199 (
            .O(N__51667),
            .I(shift_srl_8Z0Z_0));
    InMux I__5198 (
            .O(N__51664),
            .I(N__51661));
    LocalMux I__5197 (
            .O(N__51661),
            .I(shift_srl_8Z0Z_1));
    InMux I__5196 (
            .O(N__51658),
            .I(N__51655));
    LocalMux I__5195 (
            .O(N__51655),
            .I(shift_srl_8Z0Z_2));
    InMux I__5194 (
            .O(N__51652),
            .I(N__51649));
    LocalMux I__5193 (
            .O(N__51649),
            .I(shift_srl_20Z0Z_2));
    InMux I__5192 (
            .O(N__51646),
            .I(N__51643));
    LocalMux I__5191 (
            .O(N__51643),
            .I(shift_srl_20Z0Z_0));
    InMux I__5190 (
            .O(N__51640),
            .I(N__51637));
    LocalMux I__5189 (
            .O(N__51637),
            .I(shift_srl_20Z0Z_3));
    InMux I__5188 (
            .O(N__51634),
            .I(N__51631));
    LocalMux I__5187 (
            .O(N__51631),
            .I(shift_srl_20Z0Z_4));
    InMux I__5186 (
            .O(N__51628),
            .I(N__51625));
    LocalMux I__5185 (
            .O(N__51625),
            .I(shift_srl_20Z0Z_5));
    InMux I__5184 (
            .O(N__51622),
            .I(N__51619));
    LocalMux I__5183 (
            .O(N__51619),
            .I(shift_srl_20Z0Z_6));
    InMux I__5182 (
            .O(N__51616),
            .I(N__51613));
    LocalMux I__5181 (
            .O(N__51613),
            .I(shift_srl_20Z0Z_10));
    InMux I__5180 (
            .O(N__51610),
            .I(N__51607));
    LocalMux I__5179 (
            .O(N__51607),
            .I(shift_srl_20Z0Z_9));
    InMux I__5178 (
            .O(N__51604),
            .I(N__51601));
    LocalMux I__5177 (
            .O(N__51601),
            .I(shift_srl_16Z0Z_1));
    InMux I__5176 (
            .O(N__51598),
            .I(N__51595));
    LocalMux I__5175 (
            .O(N__51595),
            .I(shift_srl_16Z0Z_7));
    InMux I__5174 (
            .O(N__51592),
            .I(N__51589));
    LocalMux I__5173 (
            .O(N__51589),
            .I(shift_srl_16Z0Z_2));
    InMux I__5172 (
            .O(N__51586),
            .I(N__51583));
    LocalMux I__5171 (
            .O(N__51583),
            .I(shift_srl_16Z0Z_3));
    InMux I__5170 (
            .O(N__51580),
            .I(N__51577));
    LocalMux I__5169 (
            .O(N__51577),
            .I(shift_srl_16Z0Z_4));
    InMux I__5168 (
            .O(N__51574),
            .I(N__51571));
    LocalMux I__5167 (
            .O(N__51571),
            .I(shift_srl_16Z0Z_5));
    InMux I__5166 (
            .O(N__51568),
            .I(N__51565));
    LocalMux I__5165 (
            .O(N__51565),
            .I(shift_srl_16Z0Z_6));
    InMux I__5164 (
            .O(N__51562),
            .I(N__51559));
    LocalMux I__5163 (
            .O(N__51559),
            .I(shift_srl_16Z0Z_8));
    InMux I__5162 (
            .O(N__51556),
            .I(N__51553));
    LocalMux I__5161 (
            .O(N__51553),
            .I(shift_srl_16Z0Z_9));
    CEMux I__5160 (
            .O(N__51550),
            .I(N__51546));
    CEMux I__5159 (
            .O(N__51549),
            .I(N__51543));
    LocalMux I__5158 (
            .O(N__51546),
            .I(N__51540));
    LocalMux I__5157 (
            .O(N__51543),
            .I(N__51537));
    Span4Mux_v I__5156 (
            .O(N__51540),
            .I(N__51534));
    Span4Mux_v I__5155 (
            .O(N__51537),
            .I(N__51531));
    Span4Mux_h I__5154 (
            .O(N__51534),
            .I(N__51528));
    Span4Mux_s3_h I__5153 (
            .O(N__51531),
            .I(N__51525));
    Odrv4 I__5152 (
            .O(N__51528),
            .I(clk_en_16));
    Odrv4 I__5151 (
            .O(N__51525),
            .I(clk_en_16));
    InMux I__5150 (
            .O(N__51520),
            .I(N__51517));
    LocalMux I__5149 (
            .O(N__51517),
            .I(shift_srl_20Z0Z_1));
    InMux I__5148 (
            .O(N__51514),
            .I(N__51511));
    LocalMux I__5147 (
            .O(N__51511),
            .I(shift_srl_11Z0Z_0));
    InMux I__5146 (
            .O(N__51508),
            .I(N__51505));
    LocalMux I__5145 (
            .O(N__51505),
            .I(shift_srl_11Z0Z_1));
    InMux I__5144 (
            .O(N__51502),
            .I(N__51499));
    LocalMux I__5143 (
            .O(N__51499),
            .I(shift_srl_11Z0Z_2));
    InMux I__5142 (
            .O(N__51496),
            .I(N__51493));
    LocalMux I__5141 (
            .O(N__51493),
            .I(shift_srl_11Z0Z_3));
    InMux I__5140 (
            .O(N__51490),
            .I(N__51487));
    LocalMux I__5139 (
            .O(N__51487),
            .I(shift_srl_11Z0Z_4));
    InMux I__5138 (
            .O(N__51484),
            .I(N__51481));
    LocalMux I__5137 (
            .O(N__51481),
            .I(shift_srl_11Z0Z_7));
    InMux I__5136 (
            .O(N__51478),
            .I(N__51475));
    LocalMux I__5135 (
            .O(N__51475),
            .I(shift_srl_11Z0Z_8));
    InMux I__5134 (
            .O(N__51472),
            .I(N__51469));
    LocalMux I__5133 (
            .O(N__51469),
            .I(shift_srl_11Z0Z_5));
    InMux I__5132 (
            .O(N__51466),
            .I(N__51463));
    LocalMux I__5131 (
            .O(N__51463),
            .I(shift_srl_11Z0Z_6));
    CEMux I__5130 (
            .O(N__51460),
            .I(N__51457));
    LocalMux I__5129 (
            .O(N__51457),
            .I(N__51453));
    CEMux I__5128 (
            .O(N__51456),
            .I(N__51450));
    Span4Mux_h I__5127 (
            .O(N__51453),
            .I(N__51444));
    LocalMux I__5126 (
            .O(N__51450),
            .I(N__51444));
    CEMux I__5125 (
            .O(N__51449),
            .I(N__51441));
    Span4Mux_h I__5124 (
            .O(N__51444),
            .I(N__51438));
    LocalMux I__5123 (
            .O(N__51441),
            .I(N__51435));
    Odrv4 I__5122 (
            .O(N__51438),
            .I(clk_en_11));
    Odrv4 I__5121 (
            .O(N__51435),
            .I(clk_en_11));
    InMux I__5120 (
            .O(N__51430),
            .I(N__51427));
    LocalMux I__5119 (
            .O(N__51427),
            .I(shift_srl_16Z0Z_0));
    InMux I__5118 (
            .O(N__51424),
            .I(N__51421));
    LocalMux I__5117 (
            .O(N__51421),
            .I(shift_srl_22Z0Z_10));
    InMux I__5116 (
            .O(N__51418),
            .I(N__51415));
    LocalMux I__5115 (
            .O(N__51415),
            .I(shift_srl_22Z0Z_11));
    InMux I__5114 (
            .O(N__51412),
            .I(N__51409));
    LocalMux I__5113 (
            .O(N__51409),
            .I(shift_srl_22Z0Z_12));
    InMux I__5112 (
            .O(N__51406),
            .I(N__51403));
    LocalMux I__5111 (
            .O(N__51403),
            .I(shift_srl_22Z0Z_13));
    InMux I__5110 (
            .O(N__51400),
            .I(N__51397));
    LocalMux I__5109 (
            .O(N__51397),
            .I(N__51394));
    Odrv4 I__5108 (
            .O(N__51394),
            .I(shift_srl_22Z0Z_7));
    InMux I__5107 (
            .O(N__51391),
            .I(N__51388));
    LocalMux I__5106 (
            .O(N__51388),
            .I(shift_srl_22Z0Z_14));
    InMux I__5105 (
            .O(N__51385),
            .I(N__51382));
    LocalMux I__5104 (
            .O(N__51382),
            .I(shift_srl_22Z0Z_8));
    InMux I__5103 (
            .O(N__51379),
            .I(N__51376));
    LocalMux I__5102 (
            .O(N__51376),
            .I(shift_srl_22Z0Z_9));
    CascadeMux I__5101 (
            .O(N__51373),
            .I(N__51367));
    CascadeMux I__5100 (
            .O(N__51372),
            .I(N__51364));
    InMux I__5099 (
            .O(N__51371),
            .I(N__51359));
    InMux I__5098 (
            .O(N__51370),
            .I(N__51359));
    InMux I__5097 (
            .O(N__51367),
            .I(N__51355));
    InMux I__5096 (
            .O(N__51364),
            .I(N__51352));
    LocalMux I__5095 (
            .O(N__51359),
            .I(N__51349));
    InMux I__5094 (
            .O(N__51358),
            .I(N__51345));
    LocalMux I__5093 (
            .O(N__51355),
            .I(N__51340));
    LocalMux I__5092 (
            .O(N__51352),
            .I(N__51340));
    Span4Mux_v I__5091 (
            .O(N__51349),
            .I(N__51337));
    InMux I__5090 (
            .O(N__51348),
            .I(N__51334));
    LocalMux I__5089 (
            .O(N__51345),
            .I(shift_srl_11Z0Z_15));
    Odrv12 I__5088 (
            .O(N__51340),
            .I(shift_srl_11Z0Z_15));
    Odrv4 I__5087 (
            .O(N__51337),
            .I(shift_srl_11Z0Z_15));
    LocalMux I__5086 (
            .O(N__51334),
            .I(shift_srl_11Z0Z_15));
    InMux I__5085 (
            .O(N__51325),
            .I(N__51321));
    InMux I__5084 (
            .O(N__51324),
            .I(N__51318));
    LocalMux I__5083 (
            .O(N__51321),
            .I(N__51315));
    LocalMux I__5082 (
            .O(N__51318),
            .I(shift_srl_138Z0Z_15));
    Odrv4 I__5081 (
            .O(N__51315),
            .I(shift_srl_138Z0Z_15));
    CascadeMux I__5080 (
            .O(N__51310),
            .I(shift_srl_133_fast_RNIML0IZ0Z_15_cascade_));
    IoInMux I__5079 (
            .O(N__51307),
            .I(N__51304));
    LocalMux I__5078 (
            .O(N__51304),
            .I(N__51301));
    IoSpan4Mux I__5077 (
            .O(N__51301),
            .I(N__51298));
    Span4Mux_s3_v I__5076 (
            .O(N__51298),
            .I(N__51295));
    Span4Mux_v I__5075 (
            .O(N__51295),
            .I(N__51292));
    Odrv4 I__5074 (
            .O(N__51292),
            .I(rco_c_136));
    InMux I__5073 (
            .O(N__51289),
            .I(N__51286));
    LocalMux I__5072 (
            .O(N__51286),
            .I(N__51282));
    InMux I__5071 (
            .O(N__51285),
            .I(N__51279));
    Odrv12 I__5070 (
            .O(N__51282),
            .I(shift_srl_133Z0Z_14));
    LocalMux I__5069 (
            .O(N__51279),
            .I(shift_srl_133Z0Z_14));
    InMux I__5068 (
            .O(N__51274),
            .I(N__51271));
    LocalMux I__5067 (
            .O(N__51271),
            .I(shift_srl_133_fastZ0Z_15));
    InMux I__5066 (
            .O(N__51268),
            .I(N__51265));
    LocalMux I__5065 (
            .O(N__51265),
            .I(N__51259));
    InMux I__5064 (
            .O(N__51264),
            .I(N__51252));
    InMux I__5063 (
            .O(N__51263),
            .I(N__51252));
    InMux I__5062 (
            .O(N__51262),
            .I(N__51252));
    Span4Mux_s3_h I__5061 (
            .O(N__51259),
            .I(N__51247));
    LocalMux I__5060 (
            .O(N__51252),
            .I(N__51247));
    Odrv4 I__5059 (
            .O(N__51247),
            .I(shift_srl_137Z0Z_15));
    InMux I__5058 (
            .O(N__51244),
            .I(N__51241));
    LocalMux I__5057 (
            .O(N__51241),
            .I(N__51238));
    Odrv4 I__5056 (
            .O(N__51238),
            .I(g0_7));
    IoInMux I__5055 (
            .O(N__51235),
            .I(N__51232));
    LocalMux I__5054 (
            .O(N__51232),
            .I(N__51229));
    IoSpan4Mux I__5053 (
            .O(N__51229),
            .I(N__51226));
    Span4Mux_s3_v I__5052 (
            .O(N__51226),
            .I(N__51223));
    Span4Mux_v I__5051 (
            .O(N__51223),
            .I(N__51220));
    Odrv4 I__5050 (
            .O(N__51220),
            .I(rco_c_134));
    CascadeMux I__5049 (
            .O(N__51217),
            .I(N__51213));
    InMux I__5048 (
            .O(N__51216),
            .I(N__51209));
    InMux I__5047 (
            .O(N__51213),
            .I(N__51204));
    InMux I__5046 (
            .O(N__51212),
            .I(N__51204));
    LocalMux I__5045 (
            .O(N__51209),
            .I(shift_srl_133_fast_RNIML0IZ0Z_15));
    LocalMux I__5044 (
            .O(N__51204),
            .I(shift_srl_133_fast_RNIML0IZ0Z_15));
    IoInMux I__5043 (
            .O(N__51199),
            .I(N__51196));
    LocalMux I__5042 (
            .O(N__51196),
            .I(N__51193));
    Span4Mux_s1_v I__5041 (
            .O(N__51193),
            .I(N__51190));
    Span4Mux_v I__5040 (
            .O(N__51190),
            .I(N__51187));
    Span4Mux_v I__5039 (
            .O(N__51187),
            .I(N__51184));
    Odrv4 I__5038 (
            .O(N__51184),
            .I(rco_c_135));
    IoInMux I__5037 (
            .O(N__51181),
            .I(N__51178));
    LocalMux I__5036 (
            .O(N__51178),
            .I(N__51175));
    IoSpan4Mux I__5035 (
            .O(N__51175),
            .I(N__51172));
    Span4Mux_s3_h I__5034 (
            .O(N__51172),
            .I(N__51169));
    Odrv4 I__5033 (
            .O(N__51169),
            .I(rco_c_125));
    InMux I__5032 (
            .O(N__51166),
            .I(N__51163));
    LocalMux I__5031 (
            .O(N__51163),
            .I(shift_srl_134Z0Z_10));
    InMux I__5030 (
            .O(N__51160),
            .I(N__51157));
    LocalMux I__5029 (
            .O(N__51157),
            .I(shift_srl_134Z0Z_11));
    InMux I__5028 (
            .O(N__51154),
            .I(N__51151));
    LocalMux I__5027 (
            .O(N__51151),
            .I(shift_srl_134Z0Z_12));
    InMux I__5026 (
            .O(N__51148),
            .I(N__51145));
    LocalMux I__5025 (
            .O(N__51145),
            .I(shift_srl_134Z0Z_13));
    InMux I__5024 (
            .O(N__51142),
            .I(N__51139));
    LocalMux I__5023 (
            .O(N__51139),
            .I(shift_srl_134Z0Z_14));
    InMux I__5022 (
            .O(N__51136),
            .I(N__51133));
    LocalMux I__5021 (
            .O(N__51133),
            .I(shift_srl_134Z0Z_9));
    InMux I__5020 (
            .O(N__51130),
            .I(N__51127));
    LocalMux I__5019 (
            .O(N__51127),
            .I(shift_srl_134Z0Z_8));
    IoInMux I__5018 (
            .O(N__51124),
            .I(N__51121));
    LocalMux I__5017 (
            .O(N__51121),
            .I(N__51118));
    Span4Mux_s2_v I__5016 (
            .O(N__51118),
            .I(N__51115));
    Span4Mux_v I__5015 (
            .O(N__51115),
            .I(N__51112));
    Span4Mux_v I__5014 (
            .O(N__51112),
            .I(N__51109));
    Odrv4 I__5013 (
            .O(N__51109),
            .I(rco_c_137));
    InMux I__5012 (
            .O(N__51106),
            .I(N__51103));
    LocalMux I__5011 (
            .O(N__51103),
            .I(g0_2_1));
    InMux I__5010 (
            .O(N__51100),
            .I(N__51097));
    LocalMux I__5009 (
            .O(N__51097),
            .I(g0_11_0));
    InMux I__5008 (
            .O(N__51094),
            .I(N__51091));
    LocalMux I__5007 (
            .O(N__51091),
            .I(g0_6));
    InMux I__5006 (
            .O(N__51088),
            .I(N__51085));
    LocalMux I__5005 (
            .O(N__51085),
            .I(shift_srl_129Z0Z_13));
    InMux I__5004 (
            .O(N__51082),
            .I(N__51079));
    LocalMux I__5003 (
            .O(N__51079),
            .I(shift_srl_129Z0Z_12));
    InMux I__5002 (
            .O(N__51076),
            .I(N__51073));
    LocalMux I__5001 (
            .O(N__51073),
            .I(shift_srl_129Z0Z_11));
    InMux I__5000 (
            .O(N__51070),
            .I(N__51067));
    LocalMux I__4999 (
            .O(N__51067),
            .I(N__51064));
    Span4Mux_v I__4998 (
            .O(N__51064),
            .I(N__51061));
    Odrv4 I__4997 (
            .O(N__51061),
            .I(shift_srl_129Z0Z_9));
    InMux I__4996 (
            .O(N__51058),
            .I(N__51055));
    LocalMux I__4995 (
            .O(N__51055),
            .I(shift_srl_129Z0Z_10));
    InMux I__4994 (
            .O(N__51052),
            .I(N__51049));
    LocalMux I__4993 (
            .O(N__51049),
            .I(shift_srl_131Z0Z_4));
    InMux I__4992 (
            .O(N__51046),
            .I(N__51043));
    LocalMux I__4991 (
            .O(N__51043),
            .I(shift_srl_131Z0Z_5));
    InMux I__4990 (
            .O(N__51040),
            .I(N__51037));
    LocalMux I__4989 (
            .O(N__51037),
            .I(shift_srl_131Z0Z_6));
    InMux I__4988 (
            .O(N__51034),
            .I(N__51031));
    LocalMux I__4987 (
            .O(N__51031),
            .I(shift_srl_131Z0Z_7));
    CascadeMux I__4986 (
            .O(N__51028),
            .I(rco_obuf_RNO_0Z0Z_131_cascade_));
    IoInMux I__4985 (
            .O(N__51025),
            .I(N__51022));
    LocalMux I__4984 (
            .O(N__51022),
            .I(N__51019));
    IoSpan4Mux I__4983 (
            .O(N__51019),
            .I(N__51016));
    Span4Mux_s3_h I__4982 (
            .O(N__51016),
            .I(N__51013));
    Span4Mux_v I__4981 (
            .O(N__51013),
            .I(N__51010));
    Odrv4 I__4980 (
            .O(N__51010),
            .I(rco_c_131));
    IoInMux I__4979 (
            .O(N__51007),
            .I(N__51004));
    LocalMux I__4978 (
            .O(N__51004),
            .I(N__51001));
    Span4Mux_s3_h I__4977 (
            .O(N__51001),
            .I(N__50998));
    Span4Mux_v I__4976 (
            .O(N__50998),
            .I(N__50995));
    Span4Mux_v I__4975 (
            .O(N__50995),
            .I(N__50992));
    Odrv4 I__4974 (
            .O(N__50992),
            .I(rco_c_130));
    InMux I__4973 (
            .O(N__50989),
            .I(N__50986));
    LocalMux I__4972 (
            .O(N__50986),
            .I(g0_2_0));
    CascadeMux I__4971 (
            .O(N__50983),
            .I(rco_c_123_cascade_));
    IoInMux I__4970 (
            .O(N__50980),
            .I(N__50977));
    LocalMux I__4969 (
            .O(N__50977),
            .I(N__50974));
    Span4Mux_s3_h I__4968 (
            .O(N__50974),
            .I(N__50971));
    Odrv4 I__4967 (
            .O(N__50971),
            .I(clk_en_133));
    InMux I__4966 (
            .O(N__50968),
            .I(N__50965));
    LocalMux I__4965 (
            .O(N__50965),
            .I(shift_srl_133Z0Z_13));
    InMux I__4964 (
            .O(N__50962),
            .I(N__50959));
    LocalMux I__4963 (
            .O(N__50959),
            .I(shift_srl_133Z0Z_12));
    InMux I__4962 (
            .O(N__50956),
            .I(N__50953));
    LocalMux I__4961 (
            .O(N__50953),
            .I(shift_srl_133Z0Z_11));
    InMux I__4960 (
            .O(N__50950),
            .I(N__50947));
    LocalMux I__4959 (
            .O(N__50947),
            .I(shift_srl_131Z0Z_2));
    InMux I__4958 (
            .O(N__50944),
            .I(N__50941));
    LocalMux I__4957 (
            .O(N__50941),
            .I(shift_srl_131Z0Z_3));
    InMux I__4956 (
            .O(N__50938),
            .I(N__50935));
    LocalMux I__4955 (
            .O(N__50935),
            .I(shift_srl_21Z0Z_5));
    InMux I__4954 (
            .O(N__50932),
            .I(N__50929));
    LocalMux I__4953 (
            .O(N__50929),
            .I(shift_srl_21Z0Z_6));
    InMux I__4952 (
            .O(N__50926),
            .I(N__50923));
    LocalMux I__4951 (
            .O(N__50923),
            .I(shift_srl_21Z0Z_7));
    CEMux I__4950 (
            .O(N__50920),
            .I(N__50916));
    CEMux I__4949 (
            .O(N__50919),
            .I(N__50913));
    LocalMux I__4948 (
            .O(N__50916),
            .I(N__50910));
    LocalMux I__4947 (
            .O(N__50913),
            .I(N__50907));
    Span4Mux_h I__4946 (
            .O(N__50910),
            .I(N__50902));
    Span4Mux_h I__4945 (
            .O(N__50907),
            .I(N__50902));
    Odrv4 I__4944 (
            .O(N__50902),
            .I(clk_en_21));
    InMux I__4943 (
            .O(N__50899),
            .I(N__50896));
    LocalMux I__4942 (
            .O(N__50896),
            .I(N__50893));
    Odrv4 I__4941 (
            .O(N__50893),
            .I(shift_srl_18Z0Z_1));
    InMux I__4940 (
            .O(N__50890),
            .I(N__50887));
    LocalMux I__4939 (
            .O(N__50887),
            .I(shift_srl_18Z0Z_2));
    InMux I__4938 (
            .O(N__50884),
            .I(N__50881));
    LocalMux I__4937 (
            .O(N__50881),
            .I(shift_srl_18Z0Z_3));
    InMux I__4936 (
            .O(N__50878),
            .I(N__50875));
    LocalMux I__4935 (
            .O(N__50875),
            .I(shift_srl_18Z0Z_4));
    InMux I__4934 (
            .O(N__50872),
            .I(N__50869));
    LocalMux I__4933 (
            .O(N__50869),
            .I(shift_srl_18Z0Z_5));
    InMux I__4932 (
            .O(N__50866),
            .I(N__50863));
    LocalMux I__4931 (
            .O(N__50863),
            .I(shift_srl_18Z0Z_6));
    InMux I__4930 (
            .O(N__50860),
            .I(N__50857));
    LocalMux I__4929 (
            .O(N__50857),
            .I(shift_srl_18Z0Z_7));
    CEMux I__4928 (
            .O(N__50854),
            .I(N__50849));
    CEMux I__4927 (
            .O(N__50853),
            .I(N__50846));
    CEMux I__4926 (
            .O(N__50852),
            .I(N__50843));
    LocalMux I__4925 (
            .O(N__50849),
            .I(N__50840));
    LocalMux I__4924 (
            .O(N__50846),
            .I(N__50835));
    LocalMux I__4923 (
            .O(N__50843),
            .I(N__50835));
    Span4Mux_v I__4922 (
            .O(N__50840),
            .I(N__50832));
    Span4Mux_v I__4921 (
            .O(N__50835),
            .I(N__50829));
    Span4Mux_s3_h I__4920 (
            .O(N__50832),
            .I(N__50826));
    Span4Mux_s3_h I__4919 (
            .O(N__50829),
            .I(N__50823));
    Odrv4 I__4918 (
            .O(N__50826),
            .I(clk_en_18));
    Odrv4 I__4917 (
            .O(N__50823),
            .I(clk_en_18));
    InMux I__4916 (
            .O(N__50818),
            .I(N__50811));
    InMux I__4915 (
            .O(N__50817),
            .I(N__50806));
    InMux I__4914 (
            .O(N__50816),
            .I(N__50806));
    InMux I__4913 (
            .O(N__50815),
            .I(N__50801));
    InMux I__4912 (
            .O(N__50814),
            .I(N__50798));
    LocalMux I__4911 (
            .O(N__50811),
            .I(N__50793));
    LocalMux I__4910 (
            .O(N__50806),
            .I(N__50793));
    InMux I__4909 (
            .O(N__50805),
            .I(N__50788));
    InMux I__4908 (
            .O(N__50804),
            .I(N__50788));
    LocalMux I__4907 (
            .O(N__50801),
            .I(shift_srl_12Z0Z_15));
    LocalMux I__4906 (
            .O(N__50798),
            .I(shift_srl_12Z0Z_15));
    Odrv4 I__4905 (
            .O(N__50793),
            .I(shift_srl_12Z0Z_15));
    LocalMux I__4904 (
            .O(N__50788),
            .I(shift_srl_12Z0Z_15));
    CascadeMux I__4903 (
            .O(N__50779),
            .I(N__50772));
    InMux I__4902 (
            .O(N__50778),
            .I(N__50768));
    InMux I__4901 (
            .O(N__50777),
            .I(N__50764));
    InMux I__4900 (
            .O(N__50776),
            .I(N__50761));
    InMux I__4899 (
            .O(N__50775),
            .I(N__50758));
    InMux I__4898 (
            .O(N__50772),
            .I(N__50753));
    InMux I__4897 (
            .O(N__50771),
            .I(N__50753));
    LocalMux I__4896 (
            .O(N__50768),
            .I(N__50750));
    InMux I__4895 (
            .O(N__50767),
            .I(N__50747));
    LocalMux I__4894 (
            .O(N__50764),
            .I(N__50738));
    LocalMux I__4893 (
            .O(N__50761),
            .I(N__50738));
    LocalMux I__4892 (
            .O(N__50758),
            .I(N__50738));
    LocalMux I__4891 (
            .O(N__50753),
            .I(N__50738));
    Odrv4 I__4890 (
            .O(N__50750),
            .I(shift_srl_13Z0Z_15));
    LocalMux I__4889 (
            .O(N__50747),
            .I(shift_srl_13Z0Z_15));
    Odrv4 I__4888 (
            .O(N__50738),
            .I(shift_srl_13Z0Z_15));
    InMux I__4887 (
            .O(N__50731),
            .I(N__50728));
    LocalMux I__4886 (
            .O(N__50728),
            .I(N__50725));
    Span4Mux_h I__4885 (
            .O(N__50725),
            .I(N__50722));
    Odrv4 I__4884 (
            .O(N__50722),
            .I(rco_int_0_a2_sx_13));
    CascadeMux I__4883 (
            .O(N__50719),
            .I(N__50714));
    CascadeMux I__4882 (
            .O(N__50718),
            .I(N__50711));
    InMux I__4881 (
            .O(N__50717),
            .I(N__50707));
    InMux I__4880 (
            .O(N__50714),
            .I(N__50704));
    InMux I__4879 (
            .O(N__50711),
            .I(N__50699));
    CascadeMux I__4878 (
            .O(N__50710),
            .I(N__50696));
    LocalMux I__4877 (
            .O(N__50707),
            .I(N__50692));
    LocalMux I__4876 (
            .O(N__50704),
            .I(N__50689));
    InMux I__4875 (
            .O(N__50703),
            .I(N__50684));
    InMux I__4874 (
            .O(N__50702),
            .I(N__50684));
    LocalMux I__4873 (
            .O(N__50699),
            .I(N__50681));
    InMux I__4872 (
            .O(N__50696),
            .I(N__50676));
    InMux I__4871 (
            .O(N__50695),
            .I(N__50676));
    Span4Mux_h I__4870 (
            .O(N__50692),
            .I(N__50669));
    Span4Mux_h I__4869 (
            .O(N__50689),
            .I(N__50669));
    LocalMux I__4868 (
            .O(N__50684),
            .I(N__50669));
    Span4Mux_h I__4867 (
            .O(N__50681),
            .I(N__50666));
    LocalMux I__4866 (
            .O(N__50676),
            .I(N__50663));
    Span4Mux_v I__4865 (
            .O(N__50669),
            .I(N__50660));
    Span4Mux_v I__4864 (
            .O(N__50666),
            .I(N__50657));
    Odrv12 I__4863 (
            .O(N__50663),
            .I(shift_srl_18Z0Z_15));
    Odrv4 I__4862 (
            .O(N__50660),
            .I(shift_srl_18Z0Z_15));
    Odrv4 I__4861 (
            .O(N__50657),
            .I(shift_srl_18Z0Z_15));
    InMux I__4860 (
            .O(N__50650),
            .I(N__50647));
    LocalMux I__4859 (
            .O(N__50647),
            .I(shift_srl_18Z0Z_0));
    InMux I__4858 (
            .O(N__50644),
            .I(N__50640));
    InMux I__4857 (
            .O(N__50643),
            .I(N__50637));
    LocalMux I__4856 (
            .O(N__50640),
            .I(N__50634));
    LocalMux I__4855 (
            .O(N__50637),
            .I(shift_srl_21Z0Z_15));
    Odrv4 I__4854 (
            .O(N__50634),
            .I(shift_srl_21Z0Z_15));
    InMux I__4853 (
            .O(N__50629),
            .I(N__50626));
    LocalMux I__4852 (
            .O(N__50626),
            .I(shift_srl_21Z0Z_0));
    InMux I__4851 (
            .O(N__50623),
            .I(N__50620));
    LocalMux I__4850 (
            .O(N__50620),
            .I(shift_srl_21Z0Z_1));
    InMux I__4849 (
            .O(N__50617),
            .I(N__50614));
    LocalMux I__4848 (
            .O(N__50614),
            .I(shift_srl_21Z0Z_2));
    InMux I__4847 (
            .O(N__50611),
            .I(N__50608));
    LocalMux I__4846 (
            .O(N__50608),
            .I(shift_srl_21Z0Z_3));
    InMux I__4845 (
            .O(N__50605),
            .I(N__50602));
    LocalMux I__4844 (
            .O(N__50602),
            .I(shift_srl_21Z0Z_4));
    IoInMux I__4843 (
            .O(N__50599),
            .I(N__50596));
    LocalMux I__4842 (
            .O(N__50596),
            .I(N__50593));
    Span12Mux_s3_h I__4841 (
            .O(N__50593),
            .I(N__50589));
    InMux I__4840 (
            .O(N__50592),
            .I(N__50586));
    Odrv12 I__4839 (
            .O(N__50589),
            .I(rco_c_14));
    LocalMux I__4838 (
            .O(N__50586),
            .I(rco_c_14));
    CascadeMux I__4837 (
            .O(N__50581),
            .I(rco_int_0_a2_21_m6_0_a2_s_6_cascade_));
    IoInMux I__4836 (
            .O(N__50578),
            .I(N__50575));
    LocalMux I__4835 (
            .O(N__50575),
            .I(N__50572));
    IoSpan4Mux I__4834 (
            .O(N__50572),
            .I(N__50569));
    Span4Mux_s3_h I__4833 (
            .O(N__50569),
            .I(N__50566));
    Span4Mux_v I__4832 (
            .O(N__50566),
            .I(N__50563));
    Odrv4 I__4831 (
            .O(N__50563),
            .I(rco_c_18));
    CascadeMux I__4830 (
            .O(N__50560),
            .I(rco_c_18_cascade_));
    InMux I__4829 (
            .O(N__50557),
            .I(N__50551));
    InMux I__4828 (
            .O(N__50556),
            .I(N__50551));
    LocalMux I__4827 (
            .O(N__50551),
            .I(N__50543));
    InMux I__4826 (
            .O(N__50550),
            .I(N__50538));
    InMux I__4825 (
            .O(N__50549),
            .I(N__50538));
    InMux I__4824 (
            .O(N__50548),
            .I(N__50535));
    InMux I__4823 (
            .O(N__50547),
            .I(N__50532));
    InMux I__4822 (
            .O(N__50546),
            .I(N__50529));
    Sp12to4 I__4821 (
            .O(N__50543),
            .I(N__50522));
    LocalMux I__4820 (
            .O(N__50538),
            .I(N__50522));
    LocalMux I__4819 (
            .O(N__50535),
            .I(N__50522));
    LocalMux I__4818 (
            .O(N__50532),
            .I(N__50519));
    LocalMux I__4817 (
            .O(N__50529),
            .I(shift_srl_15Z0Z_15));
    Odrv12 I__4816 (
            .O(N__50522),
            .I(shift_srl_15Z0Z_15));
    Odrv4 I__4815 (
            .O(N__50519),
            .I(shift_srl_15Z0Z_15));
    CascadeMux I__4814 (
            .O(N__50512),
            .I(rco_int_0_a2_sx_15_cascade_));
    InMux I__4813 (
            .O(N__50509),
            .I(N__50504));
    InMux I__4812 (
            .O(N__50508),
            .I(N__50496));
    InMux I__4811 (
            .O(N__50507),
            .I(N__50496));
    LocalMux I__4810 (
            .O(N__50504),
            .I(N__50493));
    InMux I__4809 (
            .O(N__50503),
            .I(N__50490));
    InMux I__4808 (
            .O(N__50502),
            .I(N__50487));
    InMux I__4807 (
            .O(N__50501),
            .I(N__50483));
    LocalMux I__4806 (
            .O(N__50496),
            .I(N__50480));
    Sp12to4 I__4805 (
            .O(N__50493),
            .I(N__50473));
    LocalMux I__4804 (
            .O(N__50490),
            .I(N__50473));
    LocalMux I__4803 (
            .O(N__50487),
            .I(N__50473));
    InMux I__4802 (
            .O(N__50486),
            .I(N__50470));
    LocalMux I__4801 (
            .O(N__50483),
            .I(shift_srl_14Z0Z_15));
    Odrv4 I__4800 (
            .O(N__50480),
            .I(shift_srl_14Z0Z_15));
    Odrv12 I__4799 (
            .O(N__50473),
            .I(shift_srl_14Z0Z_15));
    LocalMux I__4798 (
            .O(N__50470),
            .I(shift_srl_14Z0Z_15));
    IoInMux I__4797 (
            .O(N__50461),
            .I(N__50458));
    LocalMux I__4796 (
            .O(N__50458),
            .I(N__50455));
    IoSpan4Mux I__4795 (
            .O(N__50455),
            .I(N__50452));
    Span4Mux_s3_h I__4794 (
            .O(N__50452),
            .I(N__50448));
    CascadeMux I__4793 (
            .O(N__50451),
            .I(N__50445));
    Sp12to4 I__4792 (
            .O(N__50448),
            .I(N__50442));
    InMux I__4791 (
            .O(N__50445),
            .I(N__50439));
    Odrv12 I__4790 (
            .O(N__50442),
            .I(rco_c_15));
    LocalMux I__4789 (
            .O(N__50439),
            .I(rco_c_15));
    CascadeMux I__4788 (
            .O(N__50434),
            .I(rco_c_15_cascade_));
    InMux I__4787 (
            .O(N__50431),
            .I(N__50423));
    InMux I__4786 (
            .O(N__50430),
            .I(N__50423));
    InMux I__4785 (
            .O(N__50429),
            .I(N__50417));
    InMux I__4784 (
            .O(N__50428),
            .I(N__50414));
    LocalMux I__4783 (
            .O(N__50423),
            .I(N__50411));
    InMux I__4782 (
            .O(N__50422),
            .I(N__50404));
    InMux I__4781 (
            .O(N__50421),
            .I(N__50404));
    InMux I__4780 (
            .O(N__50420),
            .I(N__50404));
    LocalMux I__4779 (
            .O(N__50417),
            .I(shift_srl_16Z0Z_15));
    LocalMux I__4778 (
            .O(N__50414),
            .I(shift_srl_16Z0Z_15));
    Odrv4 I__4777 (
            .O(N__50411),
            .I(shift_srl_16Z0Z_15));
    LocalMux I__4776 (
            .O(N__50404),
            .I(shift_srl_16Z0Z_15));
    InMux I__4775 (
            .O(N__50395),
            .I(N__50392));
    LocalMux I__4774 (
            .O(N__50392),
            .I(shift_srl_16Z0Z_12));
    InMux I__4773 (
            .O(N__50389),
            .I(N__50386));
    LocalMux I__4772 (
            .O(N__50386),
            .I(shift_srl_16Z0Z_13));
    InMux I__4771 (
            .O(N__50383),
            .I(N__50380));
    LocalMux I__4770 (
            .O(N__50380),
            .I(shift_srl_16Z0Z_14));
    IoInMux I__4769 (
            .O(N__50377),
            .I(N__50374));
    LocalMux I__4768 (
            .O(N__50374),
            .I(N__50370));
    InMux I__4767 (
            .O(N__50373),
            .I(N__50367));
    Span4Mux_s2_h I__4766 (
            .O(N__50370),
            .I(N__50362));
    LocalMux I__4765 (
            .O(N__50367),
            .I(N__50359));
    InMux I__4764 (
            .O(N__50366),
            .I(N__50356));
    InMux I__4763 (
            .O(N__50365),
            .I(N__50353));
    Odrv4 I__4762 (
            .O(N__50362),
            .I(rco_c_11));
    Odrv4 I__4761 (
            .O(N__50359),
            .I(rco_c_11));
    LocalMux I__4760 (
            .O(N__50356),
            .I(rco_c_11));
    LocalMux I__4759 (
            .O(N__50353),
            .I(rco_c_11));
    CascadeMux I__4758 (
            .O(N__50344),
            .I(rco_c_14_cascade_));
    CascadeMux I__4757 (
            .O(N__50341),
            .I(rco_c_17_cascade_));
    IoInMux I__4756 (
            .O(N__50338),
            .I(N__50335));
    LocalMux I__4755 (
            .O(N__50335),
            .I(N__50332));
    IoSpan4Mux I__4754 (
            .O(N__50332),
            .I(N__50329));
    Span4Mux_s2_h I__4753 (
            .O(N__50329),
            .I(N__50326));
    Span4Mux_v I__4752 (
            .O(N__50326),
            .I(N__50323));
    Span4Mux_v I__4751 (
            .O(N__50323),
            .I(N__50320));
    Odrv4 I__4750 (
            .O(N__50320),
            .I(rco_c_20));
    IoInMux I__4749 (
            .O(N__50317),
            .I(N__50314));
    LocalMux I__4748 (
            .O(N__50314),
            .I(N__50311));
    Span12Mux_s3_h I__4747 (
            .O(N__50311),
            .I(N__50307));
    InMux I__4746 (
            .O(N__50310),
            .I(N__50304));
    Odrv12 I__4745 (
            .O(N__50307),
            .I(rco_c_17));
    LocalMux I__4744 (
            .O(N__50304),
            .I(rco_c_17));
    InMux I__4743 (
            .O(N__50299),
            .I(N__50296));
    LocalMux I__4742 (
            .O(N__50296),
            .I(shift_srl_11Z0Z_14));
    InMux I__4741 (
            .O(N__50293),
            .I(N__50290));
    LocalMux I__4740 (
            .O(N__50290),
            .I(shift_srl_11Z0Z_13));
    InMux I__4739 (
            .O(N__50287),
            .I(N__50284));
    LocalMux I__4738 (
            .O(N__50284),
            .I(shift_srl_11Z0Z_12));
    InMux I__4737 (
            .O(N__50281),
            .I(N__50278));
    LocalMux I__4736 (
            .O(N__50278),
            .I(shift_srl_11Z0Z_11));
    InMux I__4735 (
            .O(N__50275),
            .I(N__50272));
    LocalMux I__4734 (
            .O(N__50272),
            .I(shift_srl_11Z0Z_10));
    InMux I__4733 (
            .O(N__50269),
            .I(N__50266));
    LocalMux I__4732 (
            .O(N__50266),
            .I(shift_srl_11Z0Z_9));
    InMux I__4731 (
            .O(N__50263),
            .I(N__50260));
    LocalMux I__4730 (
            .O(N__50260),
            .I(shift_srl_16Z0Z_10));
    InMux I__4729 (
            .O(N__50257),
            .I(N__50254));
    LocalMux I__4728 (
            .O(N__50254),
            .I(shift_srl_16Z0Z_11));
    InMux I__4727 (
            .O(N__50251),
            .I(N__50248));
    LocalMux I__4726 (
            .O(N__50248),
            .I(shift_srl_14Z0Z_0));
    InMux I__4725 (
            .O(N__50245),
            .I(N__50242));
    LocalMux I__4724 (
            .O(N__50242),
            .I(shift_srl_14Z0Z_1));
    InMux I__4723 (
            .O(N__50239),
            .I(N__50236));
    LocalMux I__4722 (
            .O(N__50236),
            .I(shift_srl_14Z0Z_2));
    InMux I__4721 (
            .O(N__50233),
            .I(N__50230));
    LocalMux I__4720 (
            .O(N__50230),
            .I(shift_srl_14Z0Z_3));
    InMux I__4719 (
            .O(N__50227),
            .I(N__50224));
    LocalMux I__4718 (
            .O(N__50224),
            .I(shift_srl_14Z0Z_4));
    InMux I__4717 (
            .O(N__50221),
            .I(N__50218));
    LocalMux I__4716 (
            .O(N__50218),
            .I(shift_srl_14Z0Z_12));
    InMux I__4715 (
            .O(N__50215),
            .I(N__50212));
    LocalMux I__4714 (
            .O(N__50212),
            .I(shift_srl_14Z0Z_13));
    InMux I__4713 (
            .O(N__50209),
            .I(N__50206));
    LocalMux I__4712 (
            .O(N__50206),
            .I(shift_srl_14Z0Z_14));
    CEMux I__4711 (
            .O(N__50203),
            .I(N__50199));
    CEMux I__4710 (
            .O(N__50202),
            .I(N__50196));
    LocalMux I__4709 (
            .O(N__50199),
            .I(N__50193));
    LocalMux I__4708 (
            .O(N__50196),
            .I(N__50190));
    Span4Mux_h I__4707 (
            .O(N__50193),
            .I(N__50187));
    Span4Mux_v I__4706 (
            .O(N__50190),
            .I(N__50184));
    Odrv4 I__4705 (
            .O(N__50187),
            .I(clk_en_14));
    Odrv4 I__4704 (
            .O(N__50184),
            .I(clk_en_14));
    IoInMux I__4703 (
            .O(N__50179),
            .I(N__50176));
    LocalMux I__4702 (
            .O(N__50176),
            .I(N__50173));
    Span4Mux_s2_h I__4701 (
            .O(N__50173),
            .I(N__50170));
    Odrv4 I__4700 (
            .O(N__50170),
            .I(rco_c_124));
    InMux I__4699 (
            .O(N__50167),
            .I(N__50164));
    LocalMux I__4698 (
            .O(N__50164),
            .I(shift_srl_15Z0Z_10));
    InMux I__4697 (
            .O(N__50161),
            .I(N__50158));
    LocalMux I__4696 (
            .O(N__50158),
            .I(shift_srl_15Z0Z_11));
    InMux I__4695 (
            .O(N__50155),
            .I(N__50152));
    LocalMux I__4694 (
            .O(N__50152),
            .I(shift_srl_15Z0Z_12));
    InMux I__4693 (
            .O(N__50149),
            .I(N__50146));
    LocalMux I__4692 (
            .O(N__50146),
            .I(shift_srl_15Z0Z_13));
    InMux I__4691 (
            .O(N__50143),
            .I(N__50140));
    LocalMux I__4690 (
            .O(N__50140),
            .I(shift_srl_15Z0Z_14));
    InMux I__4689 (
            .O(N__50137),
            .I(N__50134));
    LocalMux I__4688 (
            .O(N__50134),
            .I(shift_srl_15Z0Z_9));
    InMux I__4687 (
            .O(N__50131),
            .I(N__50128));
    LocalMux I__4686 (
            .O(N__50128),
            .I(shift_srl_15Z0Z_7));
    InMux I__4685 (
            .O(N__50125),
            .I(N__50122));
    LocalMux I__4684 (
            .O(N__50122),
            .I(shift_srl_15Z0Z_8));
    CEMux I__4683 (
            .O(N__50119),
            .I(N__50115));
    CEMux I__4682 (
            .O(N__50118),
            .I(N__50112));
    LocalMux I__4681 (
            .O(N__50115),
            .I(N__50109));
    LocalMux I__4680 (
            .O(N__50112),
            .I(N__50106));
    Span4Mux_v I__4679 (
            .O(N__50109),
            .I(N__50103));
    Span4Mux_v I__4678 (
            .O(N__50106),
            .I(N__50100));
    Odrv4 I__4677 (
            .O(N__50103),
            .I(clk_en_15));
    Odrv4 I__4676 (
            .O(N__50100),
            .I(clk_en_15));
    CascadeMux I__4675 (
            .O(N__50095),
            .I(g0_8_0_cascade_));
    InMux I__4674 (
            .O(N__50092),
            .I(N__50089));
    LocalMux I__4673 (
            .O(N__50089),
            .I(shift_srl_138Z0Z_9));
    InMux I__4672 (
            .O(N__50086),
            .I(N__50083));
    LocalMux I__4671 (
            .O(N__50083),
            .I(shift_srl_138Z0Z_11));
    InMux I__4670 (
            .O(N__50080),
            .I(N__50077));
    LocalMux I__4669 (
            .O(N__50077),
            .I(shift_srl_138Z0Z_12));
    InMux I__4668 (
            .O(N__50074),
            .I(N__50071));
    LocalMux I__4667 (
            .O(N__50071),
            .I(shift_srl_138Z0Z_13));
    InMux I__4666 (
            .O(N__50068),
            .I(N__50065));
    LocalMux I__4665 (
            .O(N__50065),
            .I(shift_srl_138Z0Z_14));
    InMux I__4664 (
            .O(N__50062),
            .I(N__50059));
    LocalMux I__4663 (
            .O(N__50059),
            .I(shift_srl_138Z0Z_5));
    InMux I__4662 (
            .O(N__50056),
            .I(N__50053));
    LocalMux I__4661 (
            .O(N__50053),
            .I(shift_srl_138Z0Z_6));
    InMux I__4660 (
            .O(N__50050),
            .I(N__50047));
    LocalMux I__4659 (
            .O(N__50047),
            .I(shift_srl_138Z0Z_7));
    InMux I__4658 (
            .O(N__50044),
            .I(N__50041));
    LocalMux I__4657 (
            .O(N__50041),
            .I(shift_srl_138Z0Z_8));
    CEMux I__4656 (
            .O(N__50038),
            .I(N__50034));
    CEMux I__4655 (
            .O(N__50037),
            .I(N__50031));
    LocalMux I__4654 (
            .O(N__50034),
            .I(N__50028));
    LocalMux I__4653 (
            .O(N__50031),
            .I(N__50025));
    Odrv4 I__4652 (
            .O(N__50028),
            .I(clk_en_138));
    Odrv12 I__4651 (
            .O(N__50025),
            .I(clk_en_138));
    InMux I__4650 (
            .O(N__50020),
            .I(N__50017));
    LocalMux I__4649 (
            .O(N__50017),
            .I(shift_srl_137Z0Z_14));
    InMux I__4648 (
            .O(N__50014),
            .I(N__50011));
    LocalMux I__4647 (
            .O(N__50011),
            .I(shift_srl_137Z0Z_9));
    InMux I__4646 (
            .O(N__50008),
            .I(N__50005));
    LocalMux I__4645 (
            .O(N__50005),
            .I(N__50002));
    Span4Mux_h I__4644 (
            .O(N__50002),
            .I(N__49999));
    Odrv4 I__4643 (
            .O(N__49999),
            .I(shift_srl_137Z0Z_7));
    InMux I__4642 (
            .O(N__49996),
            .I(N__49993));
    LocalMux I__4641 (
            .O(N__49993),
            .I(shift_srl_137Z0Z_8));
    CEMux I__4640 (
            .O(N__49990),
            .I(N__49987));
    LocalMux I__4639 (
            .O(N__49987),
            .I(N__49983));
    CEMux I__4638 (
            .O(N__49986),
            .I(N__49980));
    Span4Mux_v I__4637 (
            .O(N__49983),
            .I(N__49977));
    LocalMux I__4636 (
            .O(N__49980),
            .I(N__49974));
    Odrv4 I__4635 (
            .O(N__49977),
            .I(clk_en_137));
    Odrv4 I__4634 (
            .O(N__49974),
            .I(clk_en_137));
    CascadeMux I__4633 (
            .O(N__49969),
            .I(g0_4_0_cascade_));
    CascadeMux I__4632 (
            .O(N__49966),
            .I(g0_13_cascade_));
    InMux I__4631 (
            .O(N__49963),
            .I(N__49960));
    LocalMux I__4630 (
            .O(N__49960),
            .I(g0_15_0));
    CascadeMux I__4629 (
            .O(N__49957),
            .I(g0_16_1_cascade_));
    CEMux I__4628 (
            .O(N__49954),
            .I(N__49949));
    CEMux I__4627 (
            .O(N__49953),
            .I(N__49946));
    CEMux I__4626 (
            .O(N__49952),
            .I(N__49943));
    LocalMux I__4625 (
            .O(N__49949),
            .I(N__49940));
    LocalMux I__4624 (
            .O(N__49946),
            .I(N__49937));
    LocalMux I__4623 (
            .O(N__49943),
            .I(N__49934));
    Span4Mux_s2_h I__4622 (
            .O(N__49940),
            .I(N__49931));
    Span4Mux_s3_h I__4621 (
            .O(N__49937),
            .I(N__49928));
    Span4Mux_s3_h I__4620 (
            .O(N__49934),
            .I(N__49925));
    Odrv4 I__4619 (
            .O(N__49931),
            .I(clk_en_136));
    Odrv4 I__4618 (
            .O(N__49928),
            .I(clk_en_136));
    Odrv4 I__4617 (
            .O(N__49925),
            .I(clk_en_136));
    InMux I__4616 (
            .O(N__49918),
            .I(N__49915));
    LocalMux I__4615 (
            .O(N__49915),
            .I(shift_srl_130Z0Z_13));
    InMux I__4614 (
            .O(N__49912),
            .I(N__49909));
    LocalMux I__4613 (
            .O(N__49909),
            .I(shift_srl_130Z0Z_12));
    InMux I__4612 (
            .O(N__49906),
            .I(N__49903));
    LocalMux I__4611 (
            .O(N__49903),
            .I(shift_srl_130Z0Z_11));
    InMux I__4610 (
            .O(N__49900),
            .I(N__49897));
    LocalMux I__4609 (
            .O(N__49897),
            .I(N__49894));
    Span4Mux_h I__4608 (
            .O(N__49894),
            .I(N__49891));
    Odrv4 I__4607 (
            .O(N__49891),
            .I(shift_srl_130Z0Z_9));
    InMux I__4606 (
            .O(N__49888),
            .I(N__49885));
    LocalMux I__4605 (
            .O(N__49885),
            .I(shift_srl_130Z0Z_10));
    CEMux I__4604 (
            .O(N__49882),
            .I(N__49878));
    CEMux I__4603 (
            .O(N__49881),
            .I(N__49874));
    LocalMux I__4602 (
            .O(N__49878),
            .I(N__49871));
    CEMux I__4601 (
            .O(N__49877),
            .I(N__49868));
    LocalMux I__4600 (
            .O(N__49874),
            .I(N__49865));
    Sp12to4 I__4599 (
            .O(N__49871),
            .I(N__49860));
    LocalMux I__4598 (
            .O(N__49868),
            .I(N__49860));
    Odrv12 I__4597 (
            .O(N__49865),
            .I(clk_en_130));
    Odrv12 I__4596 (
            .O(N__49860),
            .I(clk_en_130));
    InMux I__4595 (
            .O(N__49855),
            .I(N__49852));
    LocalMux I__4594 (
            .O(N__49852),
            .I(shift_srl_137Z0Z_10));
    InMux I__4593 (
            .O(N__49849),
            .I(N__49846));
    LocalMux I__4592 (
            .O(N__49846),
            .I(shift_srl_137Z0Z_11));
    InMux I__4591 (
            .O(N__49843),
            .I(N__49840));
    LocalMux I__4590 (
            .O(N__49840),
            .I(shift_srl_137Z0Z_12));
    InMux I__4589 (
            .O(N__49837),
            .I(N__49834));
    LocalMux I__4588 (
            .O(N__49834),
            .I(shift_srl_137Z0Z_13));
    InMux I__4587 (
            .O(N__49831),
            .I(N__49828));
    LocalMux I__4586 (
            .O(N__49828),
            .I(shift_srl_129Z0Z_2));
    InMux I__4585 (
            .O(N__49825),
            .I(N__49822));
    LocalMux I__4584 (
            .O(N__49822),
            .I(shift_srl_129Z0Z_3));
    InMux I__4583 (
            .O(N__49819),
            .I(N__49816));
    LocalMux I__4582 (
            .O(N__49816),
            .I(shift_srl_129Z0Z_4));
    InMux I__4581 (
            .O(N__49813),
            .I(N__49810));
    LocalMux I__4580 (
            .O(N__49810),
            .I(shift_srl_129Z0Z_5));
    InMux I__4579 (
            .O(N__49807),
            .I(N__49804));
    LocalMux I__4578 (
            .O(N__49804),
            .I(shift_srl_129Z0Z_6));
    InMux I__4577 (
            .O(N__49801),
            .I(N__49798));
    LocalMux I__4576 (
            .O(N__49798),
            .I(shift_srl_129Z0Z_7));
    InMux I__4575 (
            .O(N__49795),
            .I(N__49792));
    LocalMux I__4574 (
            .O(N__49792),
            .I(g0_8_1));
    InMux I__4573 (
            .O(N__49789),
            .I(N__49786));
    LocalMux I__4572 (
            .O(N__49786),
            .I(shift_srl_130Z0Z_14));
    InMux I__4571 (
            .O(N__49783),
            .I(N__49780));
    LocalMux I__4570 (
            .O(N__49780),
            .I(shift_srl_18Z0Z_11));
    InMux I__4569 (
            .O(N__49777),
            .I(N__49774));
    LocalMux I__4568 (
            .O(N__49774),
            .I(shift_srl_18Z0Z_12));
    InMux I__4567 (
            .O(N__49771),
            .I(N__49768));
    LocalMux I__4566 (
            .O(N__49768),
            .I(shift_srl_18Z0Z_13));
    InMux I__4565 (
            .O(N__49765),
            .I(N__49762));
    LocalMux I__4564 (
            .O(N__49762),
            .I(shift_srl_18Z0Z_14));
    InMux I__4563 (
            .O(N__49759),
            .I(N__49756));
    LocalMux I__4562 (
            .O(N__49756),
            .I(shift_srl_18Z0Z_9));
    InMux I__4561 (
            .O(N__49753),
            .I(N__49750));
    LocalMux I__4560 (
            .O(N__49750),
            .I(shift_srl_18Z0Z_8));
    InMux I__4559 (
            .O(N__49747),
            .I(N__49744));
    LocalMux I__4558 (
            .O(N__49744),
            .I(shift_srl_129Z0Z_0));
    InMux I__4557 (
            .O(N__49741),
            .I(N__49738));
    LocalMux I__4556 (
            .O(N__49738),
            .I(shift_srl_129Z0Z_1));
    InMux I__4555 (
            .O(N__49735),
            .I(N__49732));
    LocalMux I__4554 (
            .O(N__49732),
            .I(shift_srl_7Z0Z_10));
    InMux I__4553 (
            .O(N__49729),
            .I(N__49726));
    LocalMux I__4552 (
            .O(N__49726),
            .I(shift_srl_7Z0Z_11));
    InMux I__4551 (
            .O(N__49723),
            .I(N__49720));
    LocalMux I__4550 (
            .O(N__49720),
            .I(shift_srl_7Z0Z_12));
    InMux I__4549 (
            .O(N__49717),
            .I(N__49714));
    LocalMux I__4548 (
            .O(N__49714),
            .I(shift_srl_7Z0Z_13));
    InMux I__4547 (
            .O(N__49711),
            .I(N__49708));
    LocalMux I__4546 (
            .O(N__49708),
            .I(N__49705));
    Odrv4 I__4545 (
            .O(N__49705),
            .I(shift_srl_7Z0Z_14));
    InMux I__4544 (
            .O(N__49702),
            .I(N__49699));
    LocalMux I__4543 (
            .O(N__49699),
            .I(shift_srl_7Z0Z_9));
    InMux I__4542 (
            .O(N__49696),
            .I(N__49693));
    LocalMux I__4541 (
            .O(N__49693),
            .I(shift_srl_7Z0Z_8));
    InMux I__4540 (
            .O(N__49690),
            .I(N__49687));
    LocalMux I__4539 (
            .O(N__49687),
            .I(shift_srl_7Z0Z_6));
    InMux I__4538 (
            .O(N__49684),
            .I(N__49681));
    LocalMux I__4537 (
            .O(N__49681),
            .I(shift_srl_7Z0Z_7));
    CEMux I__4536 (
            .O(N__49678),
            .I(N__49672));
    CEMux I__4535 (
            .O(N__49677),
            .I(N__49669));
    CEMux I__4534 (
            .O(N__49676),
            .I(N__49666));
    CEMux I__4533 (
            .O(N__49675),
            .I(N__49663));
    LocalMux I__4532 (
            .O(N__49672),
            .I(clk_en_7));
    LocalMux I__4531 (
            .O(N__49669),
            .I(clk_en_7));
    LocalMux I__4530 (
            .O(N__49666),
            .I(clk_en_7));
    LocalMux I__4529 (
            .O(N__49663),
            .I(clk_en_7));
    InMux I__4528 (
            .O(N__49654),
            .I(N__49651));
    LocalMux I__4527 (
            .O(N__49651),
            .I(shift_srl_18Z0Z_10));
    CascadeMux I__4526 (
            .O(N__49648),
            .I(rco_c_7_cascade_));
    InMux I__4525 (
            .O(N__49645),
            .I(N__49642));
    LocalMux I__4524 (
            .O(N__49642),
            .I(shift_srl_21Z0Z_10));
    InMux I__4523 (
            .O(N__49639),
            .I(N__49636));
    LocalMux I__4522 (
            .O(N__49636),
            .I(shift_srl_21Z0Z_11));
    InMux I__4521 (
            .O(N__49633),
            .I(N__49630));
    LocalMux I__4520 (
            .O(N__49630),
            .I(shift_srl_21Z0Z_12));
    InMux I__4519 (
            .O(N__49627),
            .I(N__49624));
    LocalMux I__4518 (
            .O(N__49624),
            .I(shift_srl_21Z0Z_13));
    InMux I__4517 (
            .O(N__49621),
            .I(N__49618));
    LocalMux I__4516 (
            .O(N__49618),
            .I(shift_srl_21Z0Z_14));
    InMux I__4515 (
            .O(N__49615),
            .I(N__49612));
    LocalMux I__4514 (
            .O(N__49612),
            .I(shift_srl_21Z0Z_9));
    InMux I__4513 (
            .O(N__49609),
            .I(N__49606));
    LocalMux I__4512 (
            .O(N__49606),
            .I(shift_srl_21Z0Z_8));
    IoInMux I__4511 (
            .O(N__49603),
            .I(N__49600));
    LocalMux I__4510 (
            .O(N__49600),
            .I(N__49597));
    Span4Mux_s2_h I__4509 (
            .O(N__49597),
            .I(N__49593));
    InMux I__4508 (
            .O(N__49596),
            .I(N__49590));
    Odrv4 I__4507 (
            .O(N__49593),
            .I(rco_c_16));
    LocalMux I__4506 (
            .O(N__49590),
            .I(rco_c_16));
    IoInMux I__4505 (
            .O(N__49585),
            .I(N__49582));
    LocalMux I__4504 (
            .O(N__49582),
            .I(N__49579));
    Odrv12 I__4503 (
            .O(N__49579),
            .I(rco_c_19));
    CascadeMux I__4502 (
            .O(N__49576),
            .I(rco_c_12_cascade_));
    CEMux I__4501 (
            .O(N__49573),
            .I(N__49570));
    LocalMux I__4500 (
            .O(N__49570),
            .I(N__49565));
    CEMux I__4499 (
            .O(N__49569),
            .I(N__49562));
    CEMux I__4498 (
            .O(N__49568),
            .I(N__49559));
    Span4Mux_v I__4497 (
            .O(N__49565),
            .I(N__49556));
    LocalMux I__4496 (
            .O(N__49562),
            .I(N__49553));
    LocalMux I__4495 (
            .O(N__49559),
            .I(N__49550));
    Span4Mux_v I__4494 (
            .O(N__49556),
            .I(N__49547));
    Span4Mux_v I__4493 (
            .O(N__49553),
            .I(N__49544));
    Span4Mux_v I__4492 (
            .O(N__49550),
            .I(N__49541));
    Odrv4 I__4491 (
            .O(N__49547),
            .I(clk_en_13));
    Odrv4 I__4490 (
            .O(N__49544),
            .I(clk_en_13));
    Odrv4 I__4489 (
            .O(N__49541),
            .I(clk_en_13));
    InMux I__4488 (
            .O(N__49534),
            .I(N__49531));
    LocalMux I__4487 (
            .O(N__49531),
            .I(rco_int_0_a2_sx_12));
    IoInMux I__4486 (
            .O(N__49528),
            .I(N__49525));
    LocalMux I__4485 (
            .O(N__49525),
            .I(N__49522));
    IoSpan4Mux I__4484 (
            .O(N__49522),
            .I(N__49518));
    CascadeMux I__4483 (
            .O(N__49521),
            .I(N__49515));
    Span4Mux_s1_h I__4482 (
            .O(N__49518),
            .I(N__49512));
    InMux I__4481 (
            .O(N__49515),
            .I(N__49509));
    Odrv4 I__4480 (
            .O(N__49512),
            .I(rco_c_12));
    LocalMux I__4479 (
            .O(N__49509),
            .I(rco_c_12));
    CascadeMux I__4478 (
            .O(N__49504),
            .I(N__49501));
    InMux I__4477 (
            .O(N__49501),
            .I(N__49498));
    LocalMux I__4476 (
            .O(N__49498),
            .I(N__49495));
    Odrv12 I__4475 (
            .O(N__49495),
            .I(rco_int_0_a2_sx_11));
    CascadeMux I__4474 (
            .O(N__49492),
            .I(N__49489));
    InMux I__4473 (
            .O(N__49489),
            .I(N__49485));
    InMux I__4472 (
            .O(N__49488),
            .I(N__49482));
    LocalMux I__4471 (
            .O(N__49485),
            .I(shift_srl_6_RNI00BHZ0Z_15));
    LocalMux I__4470 (
            .O(N__49482),
            .I(shift_srl_6_RNI00BHZ0Z_15));
    InMux I__4469 (
            .O(N__49477),
            .I(N__49470));
    InMux I__4468 (
            .O(N__49476),
            .I(N__49465));
    InMux I__4467 (
            .O(N__49475),
            .I(N__49465));
    InMux I__4466 (
            .O(N__49474),
            .I(N__49459));
    InMux I__4465 (
            .O(N__49473),
            .I(N__49459));
    LocalMux I__4464 (
            .O(N__49470),
            .I(N__49452));
    LocalMux I__4463 (
            .O(N__49465),
            .I(N__49452));
    InMux I__4462 (
            .O(N__49464),
            .I(N__49449));
    LocalMux I__4461 (
            .O(N__49459),
            .I(N__49446));
    InMux I__4460 (
            .O(N__49458),
            .I(N__49441));
    InMux I__4459 (
            .O(N__49457),
            .I(N__49441));
    Span4Mux_v I__4458 (
            .O(N__49452),
            .I(N__49438));
    LocalMux I__4457 (
            .O(N__49449),
            .I(N__49435));
    Odrv12 I__4456 (
            .O(N__49446),
            .I(shift_srl_3Z0Z_15));
    LocalMux I__4455 (
            .O(N__49441),
            .I(shift_srl_3Z0Z_15));
    Odrv4 I__4454 (
            .O(N__49438),
            .I(shift_srl_3Z0Z_15));
    Odrv4 I__4453 (
            .O(N__49435),
            .I(shift_srl_3Z0Z_15));
    InMux I__4452 (
            .O(N__49426),
            .I(N__49423));
    LocalMux I__4451 (
            .O(N__49423),
            .I(shift_srl_12Z0Z_11));
    InMux I__4450 (
            .O(N__49420),
            .I(N__49417));
    LocalMux I__4449 (
            .O(N__49417),
            .I(shift_srl_12Z0Z_10));
    InMux I__4448 (
            .O(N__49414),
            .I(N__49411));
    LocalMux I__4447 (
            .O(N__49411),
            .I(N__49408));
    Odrv4 I__4446 (
            .O(N__49408),
            .I(shift_srl_12Z0Z_8));
    InMux I__4445 (
            .O(N__49405),
            .I(N__49402));
    LocalMux I__4444 (
            .O(N__49402),
            .I(shift_srl_12Z0Z_9));
    CEMux I__4443 (
            .O(N__49399),
            .I(N__49396));
    LocalMux I__4442 (
            .O(N__49396),
            .I(N__49391));
    CEMux I__4441 (
            .O(N__49395),
            .I(N__49388));
    CEMux I__4440 (
            .O(N__49394),
            .I(N__49385));
    Span4Mux_h I__4439 (
            .O(N__49391),
            .I(N__49382));
    LocalMux I__4438 (
            .O(N__49388),
            .I(N__49379));
    LocalMux I__4437 (
            .O(N__49385),
            .I(N__49376));
    Odrv4 I__4436 (
            .O(N__49382),
            .I(clk_en_12));
    Odrv12 I__4435 (
            .O(N__49379),
            .I(clk_en_12));
    Odrv4 I__4434 (
            .O(N__49376),
            .I(clk_en_12));
    InMux I__4433 (
            .O(N__49369),
            .I(N__49364));
    CascadeMux I__4432 (
            .O(N__49368),
            .I(N__49361));
    InMux I__4431 (
            .O(N__49367),
            .I(N__49358));
    LocalMux I__4430 (
            .O(N__49364),
            .I(N__49355));
    InMux I__4429 (
            .O(N__49361),
            .I(N__49352));
    LocalMux I__4428 (
            .O(N__49358),
            .I(shift_srl_6Z0Z_15));
    Odrv4 I__4427 (
            .O(N__49355),
            .I(shift_srl_6Z0Z_15));
    LocalMux I__4426 (
            .O(N__49352),
            .I(shift_srl_6Z0Z_15));
    InMux I__4425 (
            .O(N__49345),
            .I(N__49342));
    LocalMux I__4424 (
            .O(N__49342),
            .I(N__49337));
    InMux I__4423 (
            .O(N__49341),
            .I(N__49331));
    InMux I__4422 (
            .O(N__49340),
            .I(N__49331));
    Span4Mux_h I__4421 (
            .O(N__49337),
            .I(N__49328));
    InMux I__4420 (
            .O(N__49336),
            .I(N__49325));
    LocalMux I__4419 (
            .O(N__49331),
            .I(shift_srl_5Z0Z_15));
    Odrv4 I__4418 (
            .O(N__49328),
            .I(shift_srl_5Z0Z_15));
    LocalMux I__4417 (
            .O(N__49325),
            .I(shift_srl_5Z0Z_15));
    CascadeMux I__4416 (
            .O(N__49318),
            .I(N__49314));
    CascadeMux I__4415 (
            .O(N__49317),
            .I(N__49311));
    InMux I__4414 (
            .O(N__49314),
            .I(N__49305));
    InMux I__4413 (
            .O(N__49311),
            .I(N__49305));
    InMux I__4412 (
            .O(N__49310),
            .I(N__49300));
    LocalMux I__4411 (
            .O(N__49305),
            .I(N__49297));
    InMux I__4410 (
            .O(N__49304),
            .I(N__49294));
    InMux I__4409 (
            .O(N__49303),
            .I(N__49291));
    LocalMux I__4408 (
            .O(N__49300),
            .I(shift_srl_4Z0Z_15));
    Odrv4 I__4407 (
            .O(N__49297),
            .I(shift_srl_4Z0Z_15));
    LocalMux I__4406 (
            .O(N__49294),
            .I(shift_srl_4Z0Z_15));
    LocalMux I__4405 (
            .O(N__49291),
            .I(shift_srl_4Z0Z_15));
    CascadeMux I__4404 (
            .O(N__49282),
            .I(shift_srl_6_RNI00BHZ0Z_15_cascade_));
    CascadeMux I__4403 (
            .O(N__49279),
            .I(shift_srl_7_RNI00TC1Z0Z_15_cascade_));
    IoInMux I__4402 (
            .O(N__49276),
            .I(N__49273));
    LocalMux I__4401 (
            .O(N__49273),
            .I(N__49269));
    CascadeMux I__4400 (
            .O(N__49272),
            .I(N__49266));
    Span4Mux_s2_h I__4399 (
            .O(N__49269),
            .I(N__49263));
    InMux I__4398 (
            .O(N__49266),
            .I(N__49260));
    Odrv4 I__4397 (
            .O(N__49263),
            .I(rco_c_13));
    LocalMux I__4396 (
            .O(N__49260),
            .I(rco_c_13));
    CascadeMux I__4395 (
            .O(N__49255),
            .I(rco_c_13_cascade_));
    CascadeMux I__4394 (
            .O(N__49252),
            .I(rco_c_16_cascade_));
    InMux I__4393 (
            .O(N__49249),
            .I(N__49246));
    LocalMux I__4392 (
            .O(N__49246),
            .I(shift_srl_13Z0Z_13));
    InMux I__4391 (
            .O(N__49243),
            .I(N__49240));
    LocalMux I__4390 (
            .O(N__49240),
            .I(shift_srl_13Z0Z_14));
    InMux I__4389 (
            .O(N__49237),
            .I(N__49234));
    LocalMux I__4388 (
            .O(N__49234),
            .I(shift_srl_13Z0Z_9));
    InMux I__4387 (
            .O(N__49231),
            .I(N__49228));
    LocalMux I__4386 (
            .O(N__49228),
            .I(N__49225));
    Odrv4 I__4385 (
            .O(N__49225),
            .I(shift_srl_13Z0Z_7));
    InMux I__4384 (
            .O(N__49222),
            .I(N__49219));
    LocalMux I__4383 (
            .O(N__49219),
            .I(shift_srl_13Z0Z_8));
    InMux I__4382 (
            .O(N__49216),
            .I(N__49213));
    LocalMux I__4381 (
            .O(N__49213),
            .I(shift_srl_12Z0Z_14));
    InMux I__4380 (
            .O(N__49210),
            .I(N__49207));
    LocalMux I__4379 (
            .O(N__49207),
            .I(shift_srl_12Z0Z_13));
    InMux I__4378 (
            .O(N__49204),
            .I(N__49201));
    LocalMux I__4377 (
            .O(N__49201),
            .I(shift_srl_12Z0Z_12));
    InMux I__4376 (
            .O(N__49198),
            .I(N__49195));
    LocalMux I__4375 (
            .O(N__49195),
            .I(shift_srl_14Z0Z_5));
    InMux I__4374 (
            .O(N__49192),
            .I(N__49189));
    LocalMux I__4373 (
            .O(N__49189),
            .I(shift_srl_14Z0Z_6));
    InMux I__4372 (
            .O(N__49186),
            .I(N__49183));
    LocalMux I__4371 (
            .O(N__49183),
            .I(shift_srl_14Z0Z_9));
    InMux I__4370 (
            .O(N__49180),
            .I(N__49177));
    LocalMux I__4369 (
            .O(N__49177),
            .I(shift_srl_14Z0Z_7));
    InMux I__4368 (
            .O(N__49174),
            .I(N__49171));
    LocalMux I__4367 (
            .O(N__49171),
            .I(shift_srl_14Z0Z_8));
    InMux I__4366 (
            .O(N__49168),
            .I(N__49165));
    LocalMux I__4365 (
            .O(N__49165),
            .I(shift_srl_13Z0Z_10));
    InMux I__4364 (
            .O(N__49162),
            .I(N__49159));
    LocalMux I__4363 (
            .O(N__49159),
            .I(shift_srl_13Z0Z_11));
    InMux I__4362 (
            .O(N__49156),
            .I(N__49153));
    LocalMux I__4361 (
            .O(N__49153),
            .I(shift_srl_13Z0Z_12));
    InMux I__4360 (
            .O(N__49150),
            .I(N__49147));
    LocalMux I__4359 (
            .O(N__49147),
            .I(shift_srl_15Z0Z_1));
    InMux I__4358 (
            .O(N__49144),
            .I(N__49141));
    LocalMux I__4357 (
            .O(N__49141),
            .I(shift_srl_15Z0Z_2));
    InMux I__4356 (
            .O(N__49138),
            .I(N__49135));
    LocalMux I__4355 (
            .O(N__49135),
            .I(shift_srl_15Z0Z_3));
    InMux I__4354 (
            .O(N__49132),
            .I(N__49129));
    LocalMux I__4353 (
            .O(N__49129),
            .I(shift_srl_15Z0Z_4));
    InMux I__4352 (
            .O(N__49126),
            .I(N__49123));
    LocalMux I__4351 (
            .O(N__49123),
            .I(shift_srl_15Z0Z_5));
    InMux I__4350 (
            .O(N__49120),
            .I(N__49117));
    LocalMux I__4349 (
            .O(N__49117),
            .I(shift_srl_15Z0Z_6));
    InMux I__4348 (
            .O(N__49114),
            .I(N__49111));
    LocalMux I__4347 (
            .O(N__49111),
            .I(shift_srl_14Z0Z_10));
    InMux I__4346 (
            .O(N__49108),
            .I(N__49105));
    LocalMux I__4345 (
            .O(N__49105),
            .I(shift_srl_14Z0Z_11));
    InMux I__4344 (
            .O(N__49102),
            .I(N__49099));
    LocalMux I__4343 (
            .O(N__49099),
            .I(shift_srl_138Z0Z_1));
    InMux I__4342 (
            .O(N__49096),
            .I(N__49093));
    LocalMux I__4341 (
            .O(N__49093),
            .I(shift_srl_138Z0Z_2));
    InMux I__4340 (
            .O(N__49090),
            .I(N__49087));
    LocalMux I__4339 (
            .O(N__49087),
            .I(shift_srl_138Z0Z_3));
    InMux I__4338 (
            .O(N__49084),
            .I(N__49081));
    LocalMux I__4337 (
            .O(N__49081),
            .I(shift_srl_138Z0Z_4));
    InMux I__4336 (
            .O(N__49078),
            .I(N__49075));
    LocalMux I__4335 (
            .O(N__49075),
            .I(shift_srl_138Z0Z_0));
    InMux I__4334 (
            .O(N__49072),
            .I(N__49069));
    LocalMux I__4333 (
            .O(N__49069),
            .I(shift_srl_138Z0Z_10));
    InMux I__4332 (
            .O(N__49066),
            .I(N__49063));
    LocalMux I__4331 (
            .O(N__49063),
            .I(shift_srl_22Z0Z_1));
    InMux I__4330 (
            .O(N__49060),
            .I(N__49057));
    LocalMux I__4329 (
            .O(N__49057),
            .I(shift_srl_22Z0Z_2));
    InMux I__4328 (
            .O(N__49054),
            .I(N__49051));
    LocalMux I__4327 (
            .O(N__49051),
            .I(shift_srl_15Z0Z_0));
    InMux I__4326 (
            .O(N__49048),
            .I(N__49045));
    LocalMux I__4325 (
            .O(N__49045),
            .I(shift_srl_136Z0Z_0));
    InMux I__4324 (
            .O(N__49042),
            .I(N__49039));
    LocalMux I__4323 (
            .O(N__49039),
            .I(shift_srl_136Z0Z_1));
    InMux I__4322 (
            .O(N__49036),
            .I(N__49033));
    LocalMux I__4321 (
            .O(N__49033),
            .I(shift_srl_136Z0Z_2));
    InMux I__4320 (
            .O(N__49030),
            .I(N__49027));
    LocalMux I__4319 (
            .O(N__49027),
            .I(shift_srl_136Z0Z_3));
    InMux I__4318 (
            .O(N__49024),
            .I(N__49021));
    LocalMux I__4317 (
            .O(N__49021),
            .I(shift_srl_136Z0Z_4));
    InMux I__4316 (
            .O(N__49018),
            .I(N__49015));
    LocalMux I__4315 (
            .O(N__49015),
            .I(shift_srl_136Z0Z_5));
    InMux I__4314 (
            .O(N__49012),
            .I(N__49009));
    LocalMux I__4313 (
            .O(N__49009),
            .I(shift_srl_136Z0Z_6));
    InMux I__4312 (
            .O(N__49006),
            .I(N__49003));
    LocalMux I__4311 (
            .O(N__49003),
            .I(shift_srl_136Z0Z_7));
    CascadeMux I__4310 (
            .O(N__49000),
            .I(g0_11_cascade_));
    InMux I__4309 (
            .O(N__48997),
            .I(N__48994));
    LocalMux I__4308 (
            .O(N__48994),
            .I(g0_16_0));
    CascadeMux I__4307 (
            .O(N__48991),
            .I(g0_17_cascade_));
    InMux I__4306 (
            .O(N__48988),
            .I(N__48985));
    LocalMux I__4305 (
            .O(N__48985),
            .I(shift_srl_136Z0Z_10));
    InMux I__4304 (
            .O(N__48982),
            .I(N__48979));
    LocalMux I__4303 (
            .O(N__48979),
            .I(shift_srl_136Z0Z_11));
    InMux I__4302 (
            .O(N__48976),
            .I(N__48973));
    LocalMux I__4301 (
            .O(N__48973),
            .I(shift_srl_136Z0Z_12));
    InMux I__4300 (
            .O(N__48970),
            .I(N__48967));
    LocalMux I__4299 (
            .O(N__48967),
            .I(shift_srl_136Z0Z_13));
    InMux I__4298 (
            .O(N__48964),
            .I(N__48961));
    LocalMux I__4297 (
            .O(N__48961),
            .I(shift_srl_136Z0Z_14));
    InMux I__4296 (
            .O(N__48958),
            .I(N__48955));
    LocalMux I__4295 (
            .O(N__48955),
            .I(shift_srl_136Z0Z_9));
    InMux I__4294 (
            .O(N__48952),
            .I(N__48949));
    LocalMux I__4293 (
            .O(N__48949),
            .I(shift_srl_136Z0Z_8));
    InMux I__4292 (
            .O(N__48946),
            .I(N__48943));
    LocalMux I__4291 (
            .O(N__48943),
            .I(shift_srl_130Z0Z_0));
    InMux I__4290 (
            .O(N__48940),
            .I(N__48937));
    LocalMux I__4289 (
            .O(N__48937),
            .I(shift_srl_130Z0Z_1));
    InMux I__4288 (
            .O(N__48934),
            .I(N__48931));
    LocalMux I__4287 (
            .O(N__48931),
            .I(shift_srl_130Z0Z_2));
    InMux I__4286 (
            .O(N__48928),
            .I(N__48925));
    LocalMux I__4285 (
            .O(N__48925),
            .I(shift_srl_130Z0Z_3));
    InMux I__4284 (
            .O(N__48922),
            .I(N__48919));
    LocalMux I__4283 (
            .O(N__48919),
            .I(shift_srl_130Z0Z_4));
    InMux I__4282 (
            .O(N__48916),
            .I(N__48913));
    LocalMux I__4281 (
            .O(N__48913),
            .I(shift_srl_130Z0Z_5));
    CascadeMux I__4280 (
            .O(N__48910),
            .I(shift_srl_129_RNIDM4DZ0Z_15_cascade_));
    CascadeMux I__4279 (
            .O(N__48907),
            .I(rco_c_6_cascade_));
    InMux I__4278 (
            .O(N__48904),
            .I(N__48901));
    LocalMux I__4277 (
            .O(N__48901),
            .I(shift_srl_7Z0Z_0));
    InMux I__4276 (
            .O(N__48898),
            .I(N__48895));
    LocalMux I__4275 (
            .O(N__48895),
            .I(shift_srl_7Z0Z_1));
    InMux I__4274 (
            .O(N__48892),
            .I(N__48889));
    LocalMux I__4273 (
            .O(N__48889),
            .I(shift_srl_7Z0Z_2));
    InMux I__4272 (
            .O(N__48886),
            .I(N__48883));
    LocalMux I__4271 (
            .O(N__48883),
            .I(shift_srl_7Z0Z_3));
    InMux I__4270 (
            .O(N__48880),
            .I(N__48877));
    LocalMux I__4269 (
            .O(N__48877),
            .I(shift_srl_7Z0Z_4));
    InMux I__4268 (
            .O(N__48874),
            .I(N__48871));
    LocalMux I__4267 (
            .O(N__48871),
            .I(shift_srl_7Z0Z_5));
    InMux I__4266 (
            .O(N__48868),
            .I(N__48865));
    LocalMux I__4265 (
            .O(N__48865),
            .I(shift_srl_129Z0Z_8));
    InMux I__4264 (
            .O(N__48862),
            .I(N__48859));
    LocalMux I__4263 (
            .O(N__48859),
            .I(shift_srl_6Z0Z_0));
    InMux I__4262 (
            .O(N__48856),
            .I(N__48853));
    LocalMux I__4261 (
            .O(N__48853),
            .I(shift_srl_6Z0Z_1));
    InMux I__4260 (
            .O(N__48850),
            .I(N__48847));
    LocalMux I__4259 (
            .O(N__48847),
            .I(shift_srl_6Z0Z_2));
    InMux I__4258 (
            .O(N__48844),
            .I(N__48841));
    LocalMux I__4257 (
            .O(N__48841),
            .I(shift_srl_6Z0Z_3));
    InMux I__4256 (
            .O(N__48838),
            .I(N__48835));
    LocalMux I__4255 (
            .O(N__48835),
            .I(shift_srl_6Z0Z_4));
    InMux I__4254 (
            .O(N__48832),
            .I(N__48829));
    LocalMux I__4253 (
            .O(N__48829),
            .I(shift_srl_6Z0Z_5));
    InMux I__4252 (
            .O(N__48826),
            .I(N__48823));
    LocalMux I__4251 (
            .O(N__48823),
            .I(shift_srl_6Z0Z_6));
    CEMux I__4250 (
            .O(N__48820),
            .I(N__48817));
    LocalMux I__4249 (
            .O(N__48817),
            .I(N__48813));
    CEMux I__4248 (
            .O(N__48816),
            .I(N__48809));
    Span4Mux_v I__4247 (
            .O(N__48813),
            .I(N__48806));
    CEMux I__4246 (
            .O(N__48812),
            .I(N__48803));
    LocalMux I__4245 (
            .O(N__48809),
            .I(N__48798));
    Span4Mux_s1_h I__4244 (
            .O(N__48806),
            .I(N__48798));
    LocalMux I__4243 (
            .O(N__48803),
            .I(N__48795));
    Odrv4 I__4242 (
            .O(N__48798),
            .I(clk_en_6));
    Odrv4 I__4241 (
            .O(N__48795),
            .I(clk_en_6));
    IoInMux I__4240 (
            .O(N__48790),
            .I(N__48787));
    LocalMux I__4239 (
            .O(N__48787),
            .I(N__48784));
    Span4Mux_s0_h I__4238 (
            .O(N__48784),
            .I(N__48781));
    Span4Mux_v I__4237 (
            .O(N__48781),
            .I(N__48778));
    Odrv4 I__4236 (
            .O(N__48778),
            .I(rco_c_6));
    InMux I__4235 (
            .O(N__48775),
            .I(N__48772));
    LocalMux I__4234 (
            .O(N__48772),
            .I(shift_srl_4Z0Z_10));
    InMux I__4233 (
            .O(N__48769),
            .I(N__48766));
    LocalMux I__4232 (
            .O(N__48766),
            .I(shift_srl_4Z0Z_11));
    InMux I__4231 (
            .O(N__48763),
            .I(N__48760));
    LocalMux I__4230 (
            .O(N__48760),
            .I(shift_srl_4Z0Z_12));
    InMux I__4229 (
            .O(N__48757),
            .I(N__48754));
    LocalMux I__4228 (
            .O(N__48754),
            .I(shift_srl_4Z0Z_13));
    InMux I__4227 (
            .O(N__48751),
            .I(N__48748));
    LocalMux I__4226 (
            .O(N__48748),
            .I(shift_srl_4Z0Z_14));
    InMux I__4225 (
            .O(N__48745),
            .I(N__48742));
    LocalMux I__4224 (
            .O(N__48742),
            .I(shift_srl_4Z0Z_9));
    InMux I__4223 (
            .O(N__48739),
            .I(N__48736));
    LocalMux I__4222 (
            .O(N__48736),
            .I(shift_srl_4Z0Z_7));
    InMux I__4221 (
            .O(N__48733),
            .I(N__48730));
    LocalMux I__4220 (
            .O(N__48730),
            .I(shift_srl_4Z0Z_8));
    CEMux I__4219 (
            .O(N__48727),
            .I(N__48723));
    CEMux I__4218 (
            .O(N__48726),
            .I(N__48720));
    LocalMux I__4217 (
            .O(N__48723),
            .I(clk_en_4));
    LocalMux I__4216 (
            .O(N__48720),
            .I(clk_en_4));
    InMux I__4215 (
            .O(N__48715),
            .I(N__48712));
    LocalMux I__4214 (
            .O(N__48712),
            .I(shift_srl_6Z0Z_8));
    InMux I__4213 (
            .O(N__48709),
            .I(N__48706));
    LocalMux I__4212 (
            .O(N__48706),
            .I(shift_srl_6Z0Z_7));
    InMux I__4211 (
            .O(N__48703),
            .I(N__48700));
    LocalMux I__4210 (
            .O(N__48700),
            .I(shift_srl_12Z0Z_6));
    InMux I__4209 (
            .O(N__48697),
            .I(N__48694));
    LocalMux I__4208 (
            .O(N__48694),
            .I(shift_srl_12Z0Z_0));
    InMux I__4207 (
            .O(N__48691),
            .I(N__48688));
    LocalMux I__4206 (
            .O(N__48688),
            .I(shift_srl_12Z0Z_1));
    InMux I__4205 (
            .O(N__48685),
            .I(N__48682));
    LocalMux I__4204 (
            .O(N__48682),
            .I(shift_srl_12Z0Z_2));
    InMux I__4203 (
            .O(N__48679),
            .I(N__48676));
    LocalMux I__4202 (
            .O(N__48676),
            .I(shift_srl_12Z0Z_3));
    InMux I__4201 (
            .O(N__48673),
            .I(N__48670));
    LocalMux I__4200 (
            .O(N__48670),
            .I(shift_srl_12Z0Z_4));
    InMux I__4199 (
            .O(N__48667),
            .I(N__48664));
    LocalMux I__4198 (
            .O(N__48664),
            .I(shift_srl_12Z0Z_5));
    InMux I__4197 (
            .O(N__48661),
            .I(N__48658));
    LocalMux I__4196 (
            .O(N__48658),
            .I(shift_srl_13Z0Z_2));
    InMux I__4195 (
            .O(N__48655),
            .I(N__48652));
    LocalMux I__4194 (
            .O(N__48652),
            .I(shift_srl_13Z0Z_3));
    InMux I__4193 (
            .O(N__48649),
            .I(N__48646));
    LocalMux I__4192 (
            .O(N__48646),
            .I(shift_srl_13Z0Z_0));
    InMux I__4191 (
            .O(N__48643),
            .I(N__48640));
    LocalMux I__4190 (
            .O(N__48640),
            .I(shift_srl_13Z0Z_1));
    InMux I__4189 (
            .O(N__48637),
            .I(N__48634));
    LocalMux I__4188 (
            .O(N__48634),
            .I(shift_srl_13Z0Z_4));
    InMux I__4187 (
            .O(N__48631),
            .I(N__48628));
    LocalMux I__4186 (
            .O(N__48628),
            .I(shift_srl_13Z0Z_5));
    InMux I__4185 (
            .O(N__48625),
            .I(N__48622));
    LocalMux I__4184 (
            .O(N__48622),
            .I(shift_srl_13Z0Z_6));
    InMux I__4183 (
            .O(N__48619),
            .I(N__48616));
    LocalMux I__4182 (
            .O(N__48616),
            .I(shift_srl_12Z0Z_7));
    InMux I__4181 (
            .O(N__48613),
            .I(N__48610));
    LocalMux I__4180 (
            .O(N__48610),
            .I(shift_srl_137Z0Z_5));
    InMux I__4179 (
            .O(N__48607),
            .I(N__48604));
    LocalMux I__4178 (
            .O(N__48604),
            .I(shift_srl_137Z0Z_6));
    InMux I__4177 (
            .O(N__48601),
            .I(N__48598));
    LocalMux I__4176 (
            .O(N__48598),
            .I(shift_srl_22Z0Z_3));
    InMux I__4175 (
            .O(N__48595),
            .I(N__48592));
    LocalMux I__4174 (
            .O(N__48592),
            .I(shift_srl_22Z0Z_4));
    InMux I__4173 (
            .O(N__48589),
            .I(N__48586));
    LocalMux I__4172 (
            .O(N__48586),
            .I(shift_srl_22Z0Z_5));
    InMux I__4171 (
            .O(N__48583),
            .I(N__48580));
    LocalMux I__4170 (
            .O(N__48580),
            .I(shift_srl_22Z0Z_6));
    InMux I__4169 (
            .O(N__48577),
            .I(N__48574));
    LocalMux I__4168 (
            .O(N__48574),
            .I(shift_srl_22Z0Z_0));
    InMux I__4167 (
            .O(N__48571),
            .I(N__48568));
    LocalMux I__4166 (
            .O(N__48568),
            .I(shift_srl_130Z0Z_8));
    InMux I__4165 (
            .O(N__48565),
            .I(N__48562));
    LocalMux I__4164 (
            .O(N__48562),
            .I(shift_srl_130Z0Z_6));
    InMux I__4163 (
            .O(N__48559),
            .I(N__48556));
    LocalMux I__4162 (
            .O(N__48556),
            .I(shift_srl_130Z0Z_7));
    InMux I__4161 (
            .O(N__48553),
            .I(N__48550));
    LocalMux I__4160 (
            .O(N__48550),
            .I(shift_srl_137Z0Z_0));
    InMux I__4159 (
            .O(N__48547),
            .I(N__48544));
    LocalMux I__4158 (
            .O(N__48544),
            .I(shift_srl_137Z0Z_1));
    InMux I__4157 (
            .O(N__48541),
            .I(N__48538));
    LocalMux I__4156 (
            .O(N__48538),
            .I(shift_srl_137Z0Z_2));
    InMux I__4155 (
            .O(N__48535),
            .I(N__48532));
    LocalMux I__4154 (
            .O(N__48532),
            .I(shift_srl_137Z0Z_3));
    InMux I__4153 (
            .O(N__48529),
            .I(N__48526));
    LocalMux I__4152 (
            .O(N__48526),
            .I(shift_srl_137Z0Z_4));
    InMux I__4151 (
            .O(N__48523),
            .I(N__48520));
    LocalMux I__4150 (
            .O(N__48520),
            .I(shift_srl_5Z0Z_4));
    InMux I__4149 (
            .O(N__48517),
            .I(N__48514));
    LocalMux I__4148 (
            .O(N__48514),
            .I(shift_srl_5Z0Z_5));
    InMux I__4147 (
            .O(N__48511),
            .I(N__48508));
    LocalMux I__4146 (
            .O(N__48508),
            .I(shift_srl_5Z0Z_6));
    InMux I__4145 (
            .O(N__48505),
            .I(N__48502));
    LocalMux I__4144 (
            .O(N__48502),
            .I(N__48499));
    Odrv4 I__4143 (
            .O(N__48499),
            .I(shift_srl_5Z0Z_7));
    InMux I__4142 (
            .O(N__48496),
            .I(N__48493));
    LocalMux I__4141 (
            .O(N__48493),
            .I(shift_srl_5Z0Z_3));
    InMux I__4140 (
            .O(N__48490),
            .I(N__48487));
    LocalMux I__4139 (
            .O(N__48487),
            .I(shift_srl_5Z0Z_0));
    InMux I__4138 (
            .O(N__48484),
            .I(N__48481));
    LocalMux I__4137 (
            .O(N__48481),
            .I(shift_srl_5Z0Z_1));
    InMux I__4136 (
            .O(N__48478),
            .I(N__48475));
    LocalMux I__4135 (
            .O(N__48475),
            .I(shift_srl_5Z0Z_2));
    CEMux I__4134 (
            .O(N__48472),
            .I(N__48467));
    CEMux I__4133 (
            .O(N__48471),
            .I(N__48464));
    CEMux I__4132 (
            .O(N__48470),
            .I(N__48461));
    LocalMux I__4131 (
            .O(N__48467),
            .I(clk_en_5));
    LocalMux I__4130 (
            .O(N__48464),
            .I(clk_en_5));
    LocalMux I__4129 (
            .O(N__48461),
            .I(clk_en_5));
    InMux I__4128 (
            .O(N__48454),
            .I(N__48451));
    LocalMux I__4127 (
            .O(N__48451),
            .I(shift_srl_5Z0Z_12));
    InMux I__4126 (
            .O(N__48448),
            .I(N__48445));
    LocalMux I__4125 (
            .O(N__48445),
            .I(shift_srl_5Z0Z_13));
    InMux I__4124 (
            .O(N__48442),
            .I(N__48439));
    LocalMux I__4123 (
            .O(N__48439),
            .I(shift_srl_5Z0Z_14));
    InMux I__4122 (
            .O(N__48436),
            .I(N__48433));
    LocalMux I__4121 (
            .O(N__48433),
            .I(shift_srl_5Z0Z_9));
    InMux I__4120 (
            .O(N__48430),
            .I(N__48427));
    LocalMux I__4119 (
            .O(N__48427),
            .I(shift_srl_5Z0Z_8));
    IoInMux I__4118 (
            .O(N__48424),
            .I(N__48421));
    LocalMux I__4117 (
            .O(N__48421),
            .I(N__48418));
    Span4Mux_s2_h I__4116 (
            .O(N__48418),
            .I(N__48415));
    Span4Mux_v I__4115 (
            .O(N__48415),
            .I(N__48412));
    Odrv4 I__4114 (
            .O(N__48412),
            .I(rco_c_5));
    CascadeMux I__4113 (
            .O(N__48409),
            .I(rco_c_5_cascade_));
    IoInMux I__4112 (
            .O(N__48406),
            .I(N__48403));
    LocalMux I__4111 (
            .O(N__48403),
            .I(N__48400));
    IoSpan4Mux I__4110 (
            .O(N__48400),
            .I(N__48397));
    Odrv4 I__4109 (
            .O(N__48397),
            .I(rco_c_4));
    CascadeMux I__4108 (
            .O(N__48394),
            .I(rco_c_4_cascade_));
    InMux I__4107 (
            .O(N__48391),
            .I(N__48388));
    LocalMux I__4106 (
            .O(N__48388),
            .I(shift_srl_6Z0Z_14));
    InMux I__4105 (
            .O(N__48385),
            .I(N__48382));
    LocalMux I__4104 (
            .O(N__48382),
            .I(shift_srl_6Z0Z_13));
    InMux I__4103 (
            .O(N__48379),
            .I(N__48376));
    LocalMux I__4102 (
            .O(N__48376),
            .I(shift_srl_6Z0Z_12));
    InMux I__4101 (
            .O(N__48373),
            .I(N__48370));
    LocalMux I__4100 (
            .O(N__48370),
            .I(shift_srl_6Z0Z_11));
    InMux I__4099 (
            .O(N__48367),
            .I(N__48364));
    LocalMux I__4098 (
            .O(N__48364),
            .I(shift_srl_6Z0Z_10));
    InMux I__4097 (
            .O(N__48361),
            .I(N__48358));
    LocalMux I__4096 (
            .O(N__48358),
            .I(shift_srl_6Z0Z_9));
    InMux I__4095 (
            .O(N__48355),
            .I(N__48352));
    LocalMux I__4094 (
            .O(N__48352),
            .I(shift_srl_5Z0Z_10));
    InMux I__4093 (
            .O(N__48349),
            .I(N__48346));
    LocalMux I__4092 (
            .O(N__48346),
            .I(shift_srl_5Z0Z_11));
    InMux I__4091 (
            .O(N__48343),
            .I(N__48340));
    LocalMux I__4090 (
            .O(N__48340),
            .I(shift_srl_4Z0Z_0));
    InMux I__4089 (
            .O(N__48337),
            .I(N__48334));
    LocalMux I__4088 (
            .O(N__48334),
            .I(shift_srl_4Z0Z_1));
    InMux I__4087 (
            .O(N__48331),
            .I(N__48328));
    LocalMux I__4086 (
            .O(N__48328),
            .I(shift_srl_4Z0Z_2));
    InMux I__4085 (
            .O(N__48325),
            .I(N__48322));
    LocalMux I__4084 (
            .O(N__48322),
            .I(shift_srl_4Z0Z_3));
    InMux I__4083 (
            .O(N__48319),
            .I(N__48316));
    LocalMux I__4082 (
            .O(N__48316),
            .I(shift_srl_4Z0Z_4));
    InMux I__4081 (
            .O(N__48313),
            .I(N__48310));
    LocalMux I__4080 (
            .O(N__48310),
            .I(shift_srl_4Z0Z_5));
    InMux I__4079 (
            .O(N__48307),
            .I(N__48304));
    LocalMux I__4078 (
            .O(N__48304),
            .I(shift_srl_4Z0Z_6));
    InMux I__4077 (
            .O(N__48301),
            .I(N__48298));
    LocalMux I__4076 (
            .O(N__48298),
            .I(N__48295));
    Odrv4 I__4075 (
            .O(N__48295),
            .I(shift_srl_3Z0Z_13));
    InMux I__4074 (
            .O(N__48292),
            .I(N__48289));
    LocalMux I__4073 (
            .O(N__48289),
            .I(shift_srl_3Z0Z_14));
    InMux I__4072 (
            .O(N__48286),
            .I(N__48283));
    LocalMux I__4071 (
            .O(N__48283),
            .I(shift_srl_3Z0Z_3));
    InMux I__4070 (
            .O(N__48280),
            .I(N__48277));
    LocalMux I__4069 (
            .O(N__48277),
            .I(shift_srl_3Z0Z_4));
    IoInMux I__4068 (
            .O(N__48274),
            .I(N__48271));
    LocalMux I__4067 (
            .O(N__48271),
            .I(N__48268));
    IoSpan4Mux I__4066 (
            .O(N__48268),
            .I(N__48265));
    IoSpan4Mux I__4065 (
            .O(N__48265),
            .I(N__48262));
    Odrv4 I__4064 (
            .O(N__48262),
            .I(rco_c_3));
    CascadeMux I__4063 (
            .O(N__48259),
            .I(rco_c_3_cascade_));
    InMux I__4062 (
            .O(N__48256),
            .I(N__48253));
    LocalMux I__4061 (
            .O(N__48253),
            .I(shift_srl_3Z0Z_0));
    InMux I__4060 (
            .O(N__48250),
            .I(N__48247));
    LocalMux I__4059 (
            .O(N__48247),
            .I(shift_srl_3Z0Z_1));
    InMux I__4058 (
            .O(N__48244),
            .I(N__48241));
    LocalMux I__4057 (
            .O(N__48241),
            .I(shift_srl_3Z0Z_2));
    CEMux I__4056 (
            .O(N__48238),
            .I(N__48235));
    LocalMux I__4055 (
            .O(N__48235),
            .I(N__48230));
    CEMux I__4054 (
            .O(N__48234),
            .I(N__48227));
    CEMux I__4053 (
            .O(N__48233),
            .I(N__48224));
    Span4Mux_h I__4052 (
            .O(N__48230),
            .I(N__48221));
    LocalMux I__4051 (
            .O(N__48227),
            .I(N__48218));
    LocalMux I__4050 (
            .O(N__48224),
            .I(N__48215));
    Odrv4 I__4049 (
            .O(N__48221),
            .I(clk_en_3));
    Odrv12 I__4048 (
            .O(N__48218),
            .I(clk_en_3));
    Odrv4 I__4047 (
            .O(N__48215),
            .I(clk_en_3));
    InMux I__4046 (
            .O(N__48208),
            .I(N__48205));
    LocalMux I__4045 (
            .O(N__48205),
            .I(shift_srl_3Z0Z_10));
    InMux I__4044 (
            .O(N__48202),
            .I(N__48199));
    LocalMux I__4043 (
            .O(N__48199),
            .I(shift_srl_3Z0Z_11));
    InMux I__4042 (
            .O(N__48196),
            .I(N__48193));
    LocalMux I__4041 (
            .O(N__48193),
            .I(shift_srl_3Z0Z_12));
    InMux I__4040 (
            .O(N__48190),
            .I(N__48187));
    LocalMux I__4039 (
            .O(N__48187),
            .I(shift_srl_3Z0Z_8));
    InMux I__4038 (
            .O(N__48184),
            .I(N__48181));
    LocalMux I__4037 (
            .O(N__48181),
            .I(shift_srl_3Z0Z_9));
    InMux I__4036 (
            .O(N__48178),
            .I(N__48175));
    LocalMux I__4035 (
            .O(N__48175),
            .I(shift_srl_3Z0Z_5));
    InMux I__4034 (
            .O(N__48172),
            .I(N__48169));
    LocalMux I__4033 (
            .O(N__48169),
            .I(shift_srl_3Z0Z_6));
    InMux I__4032 (
            .O(N__48166),
            .I(N__48163));
    LocalMux I__4031 (
            .O(N__48163),
            .I(N__48160));
    Odrv4 I__4030 (
            .O(N__48160),
            .I(shift_srl_3Z0Z_7));
    IoInMux I__4029 (
            .O(N__48157),
            .I(N__48154));
    LocalMux I__4028 (
            .O(N__48154),
            .I(N__48151));
    Span4Mux_s1_h I__4027 (
            .O(N__48151),
            .I(N__48148));
    Span4Mux_v I__4026 (
            .O(N__48148),
            .I(N__48145));
    Odrv4 I__4025 (
            .O(N__48145),
            .I(N_4015_i));
    ICE_GB shift_srl_132_RNIOHTB11_0_15 (
            .USERSIGNALTOGLOBALBUFFER(N__50980),
            .GLOBALBUFFEROUTPUT(clk_en_g_133));
    ICE_GB shift_srl_0_RNIMIE4A_0_15 (
            .USERSIGNALTOGLOBALBUFFER(N__67267),
            .GLOBALBUFFEROUTPUT(clk_en_g_40));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam rco_obuf_RNO_22_LC_1_7_7.C_ON=1'b0;
    defparam rco_obuf_RNO_22_LC_1_7_7.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_22_LC_1_7_7.LUT_INIT=16'b1100110000000000;
    LogicCell40 rco_obuf_RNO_22_LC_1_7_7 (
            .in0(_gnd_net_),
            .in1(N__52143),
            .in2(_gnd_net_),
            .in3(N__53434),
            .lcout(N_4015_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_3_10_LC_1_8_0.C_ON=1'b0;
    defparam shift_srl_3_10_LC_1_8_0.SEQ_MODE=4'b1000;
    defparam shift_srl_3_10_LC_1_8_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_3_10_LC_1_8_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48184),
            .lcout(shift_srl_3Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92972),
            .ce(N__48238),
            .sr(_gnd_net_));
    defparam shift_srl_3_11_LC_1_8_1.C_ON=1'b0;
    defparam shift_srl_3_11_LC_1_8_1.SEQ_MODE=4'b1000;
    defparam shift_srl_3_11_LC_1_8_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_3_11_LC_1_8_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48208),
            .lcout(shift_srl_3Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92972),
            .ce(N__48238),
            .sr(_gnd_net_));
    defparam shift_srl_3_12_LC_1_8_2.C_ON=1'b0;
    defparam shift_srl_3_12_LC_1_8_2.SEQ_MODE=4'b1000;
    defparam shift_srl_3_12_LC_1_8_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_3_12_LC_1_8_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48202),
            .lcout(shift_srl_3Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92972),
            .ce(N__48238),
            .sr(_gnd_net_));
    defparam shift_srl_3_13_LC_1_8_3.C_ON=1'b0;
    defparam shift_srl_3_13_LC_1_8_3.SEQ_MODE=4'b1000;
    defparam shift_srl_3_13_LC_1_8_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_3_13_LC_1_8_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48196),
            .lcout(shift_srl_3Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92972),
            .ce(N__48238),
            .sr(_gnd_net_));
    defparam shift_srl_3_8_LC_1_8_4.C_ON=1'b0;
    defparam shift_srl_3_8_LC_1_8_4.SEQ_MODE=4'b1000;
    defparam shift_srl_3_8_LC_1_8_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_3_8_LC_1_8_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48166),
            .lcout(shift_srl_3Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92972),
            .ce(N__48238),
            .sr(_gnd_net_));
    defparam shift_srl_3_9_LC_1_8_6.C_ON=1'b0;
    defparam shift_srl_3_9_LC_1_8_6.SEQ_MODE=4'b1000;
    defparam shift_srl_3_9_LC_1_8_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_3_9_LC_1_8_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48190),
            .lcout(shift_srl_3Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92972),
            .ce(N__48238),
            .sr(_gnd_net_));
    defparam shift_srl_13_4_LC_1_9_1.C_ON=1'b0;
    defparam shift_srl_13_4_LC_1_9_1.SEQ_MODE=4'b1000;
    defparam shift_srl_13_4_LC_1_9_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_13_4_LC_1_9_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48655),
            .lcout(shift_srl_13Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92961),
            .ce(N__49573),
            .sr(_gnd_net_));
    defparam shift_srl_3_5_LC_1_10_0.C_ON=1'b0;
    defparam shift_srl_3_5_LC_1_10_0.SEQ_MODE=4'b1000;
    defparam shift_srl_3_5_LC_1_10_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_3_5_LC_1_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48280),
            .lcout(shift_srl_3Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92948),
            .ce(N__48234),
            .sr(_gnd_net_));
    defparam shift_srl_3_6_LC_1_10_1.C_ON=1'b0;
    defparam shift_srl_3_6_LC_1_10_1.SEQ_MODE=4'b1000;
    defparam shift_srl_3_6_LC_1_10_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_3_6_LC_1_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48178),
            .lcout(shift_srl_3Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92948),
            .ce(N__48234),
            .sr(_gnd_net_));
    defparam shift_srl_3_7_LC_1_10_2.C_ON=1'b0;
    defparam shift_srl_3_7_LC_1_10_2.SEQ_MODE=4'b1000;
    defparam shift_srl_3_7_LC_1_10_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_3_7_LC_1_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48172),
            .lcout(shift_srl_3Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92948),
            .ce(N__48234),
            .sr(_gnd_net_));
    defparam shift_srl_3_15_LC_1_10_3.C_ON=1'b0;
    defparam shift_srl_3_15_LC_1_10_3.SEQ_MODE=4'b1000;
    defparam shift_srl_3_15_LC_1_10_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_3_15_LC_1_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48292),
            .lcout(shift_srl_3Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92948),
            .ce(N__48234),
            .sr(_gnd_net_));
    defparam shift_srl_3_14_LC_1_10_4.C_ON=1'b0;
    defparam shift_srl_3_14_LC_1_10_4.SEQ_MODE=4'b1000;
    defparam shift_srl_3_14_LC_1_10_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_3_14_LC_1_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48301),
            .lcout(shift_srl_3Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92948),
            .ce(N__48234),
            .sr(_gnd_net_));
    defparam shift_srl_3_3_LC_1_10_5.C_ON=1'b0;
    defparam shift_srl_3_3_LC_1_10_5.SEQ_MODE=4'b1000;
    defparam shift_srl_3_3_LC_1_10_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_3_3_LC_1_10_5 (
            .in0(N__48244),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_3Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92948),
            .ce(N__48234),
            .sr(_gnd_net_));
    defparam shift_srl_3_4_LC_1_10_7.C_ON=1'b0;
    defparam shift_srl_3_4_LC_1_10_7.SEQ_MODE=4'b1000;
    defparam shift_srl_3_4_LC_1_10_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_3_4_LC_1_10_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48286),
            .lcout(shift_srl_3Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92948),
            .ce(N__48234),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNI2I4S_15_LC_1_11_0.C_ON=1'b0;
    defparam shift_srl_0_RNI2I4S_15_LC_1_11_0.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNI2I4S_15_LC_1_11_0.LUT_INIT=16'b0101010100000000;
    LogicCell40 shift_srl_0_RNI2I4S_15_LC_1_11_0 (
            .in0(N__53725),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__90040),
            .lcout(clk_en_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_3_RNI5UM81_15_LC_1_11_1.C_ON=1'b0;
    defparam shift_srl_3_RNI5UM81_15_LC_1_11_1.SEQ_MODE=4'b0000;
    defparam shift_srl_3_RNI5UM81_15_LC_1_11_1.LUT_INIT=16'b0011001100000000;
    LogicCell40 shift_srl_3_RNI5UM81_15_LC_1_11_1 (
            .in0(_gnd_net_),
            .in1(N__53724),
            .in2(_gnd_net_),
            .in3(N__49457),
            .lcout(rco_c_3),
            .ltout(rco_c_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNI0AH91_15_LC_1_11_2.C_ON=1'b0;
    defparam shift_srl_0_RNI0AH91_15_LC_1_11_2.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNI0AH91_15_LC_1_11_2.LUT_INIT=16'b1111000000000000;
    LogicCell40 shift_srl_0_RNI0AH91_15_LC_1_11_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__48259),
            .in3(N__90041),
            .lcout(clk_en_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_3_0_LC_1_11_3.C_ON=1'b0;
    defparam shift_srl_3_0_LC_1_11_3.SEQ_MODE=4'b1000;
    defparam shift_srl_3_0_LC_1_11_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_3_0_LC_1_11_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49458),
            .lcout(shift_srl_3Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92939),
            .ce(N__48233),
            .sr(_gnd_net_));
    defparam shift_srl_3_1_LC_1_11_4.C_ON=1'b0;
    defparam shift_srl_3_1_LC_1_11_4.SEQ_MODE=4'b1000;
    defparam shift_srl_3_1_LC_1_11_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_3_1_LC_1_11_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48256),
            .lcout(shift_srl_3Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92939),
            .ce(N__48233),
            .sr(_gnd_net_));
    defparam shift_srl_3_2_LC_1_11_5.C_ON=1'b0;
    defparam shift_srl_3_2_LC_1_11_5.SEQ_MODE=4'b1000;
    defparam shift_srl_3_2_LC_1_11_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_3_2_LC_1_11_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48250),
            .lcout(shift_srl_3Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92939),
            .ce(N__48233),
            .sr(_gnd_net_));
    defparam shift_srl_4_0_LC_1_12_0.C_ON=1'b0;
    defparam shift_srl_4_0_LC_1_12_0.SEQ_MODE=4'b1000;
    defparam shift_srl_4_0_LC_1_12_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_4_0_LC_1_12_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49310),
            .lcout(shift_srl_4Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92930),
            .ce(N__48726),
            .sr(_gnd_net_));
    defparam shift_srl_4_1_LC_1_12_1.C_ON=1'b0;
    defparam shift_srl_4_1_LC_1_12_1.SEQ_MODE=4'b1000;
    defparam shift_srl_4_1_LC_1_12_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_4_1_LC_1_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48343),
            .lcout(shift_srl_4Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92930),
            .ce(N__48726),
            .sr(_gnd_net_));
    defparam shift_srl_4_2_LC_1_12_2.C_ON=1'b0;
    defparam shift_srl_4_2_LC_1_12_2.SEQ_MODE=4'b1000;
    defparam shift_srl_4_2_LC_1_12_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_4_2_LC_1_12_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48337),
            .lcout(shift_srl_4Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92930),
            .ce(N__48726),
            .sr(_gnd_net_));
    defparam shift_srl_4_3_LC_1_12_3.C_ON=1'b0;
    defparam shift_srl_4_3_LC_1_12_3.SEQ_MODE=4'b1000;
    defparam shift_srl_4_3_LC_1_12_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_4_3_LC_1_12_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48331),
            .lcout(shift_srl_4Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92930),
            .ce(N__48726),
            .sr(_gnd_net_));
    defparam shift_srl_4_4_LC_1_12_4.C_ON=1'b0;
    defparam shift_srl_4_4_LC_1_12_4.SEQ_MODE=4'b1000;
    defparam shift_srl_4_4_LC_1_12_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_4_4_LC_1_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48325),
            .lcout(shift_srl_4Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92930),
            .ce(N__48726),
            .sr(_gnd_net_));
    defparam shift_srl_4_5_LC_1_12_5.C_ON=1'b0;
    defparam shift_srl_4_5_LC_1_12_5.SEQ_MODE=4'b1000;
    defparam shift_srl_4_5_LC_1_12_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_4_5_LC_1_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48319),
            .lcout(shift_srl_4Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92930),
            .ce(N__48726),
            .sr(_gnd_net_));
    defparam shift_srl_4_6_LC_1_12_6.C_ON=1'b0;
    defparam shift_srl_4_6_LC_1_12_6.SEQ_MODE=4'b1000;
    defparam shift_srl_4_6_LC_1_12_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_4_6_LC_1_12_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48313),
            .lcout(shift_srl_4Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92930),
            .ce(N__48726),
            .sr(_gnd_net_));
    defparam shift_srl_4_7_LC_1_12_7.C_ON=1'b0;
    defparam shift_srl_4_7_LC_1_12_7.SEQ_MODE=4'b1000;
    defparam shift_srl_4_7_LC_1_12_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_4_7_LC_1_12_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48307),
            .lcout(shift_srl_4Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92930),
            .ce(N__48726),
            .sr(_gnd_net_));
    defparam shift_srl_6_RNIUNNU_15_LC_1_13_0.C_ON=1'b0;
    defparam shift_srl_6_RNIUNNU_15_LC_1_13_0.SEQ_MODE=4'b0000;
    defparam shift_srl_6_RNIUNNU_15_LC_1_13_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_6_RNIUNNU_15_LC_1_13_0 (
            .in0(N__49336),
            .in1(N__49303),
            .in2(N__49368),
            .in3(N__49464),
            .lcout(rco_int_0_a2_out_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_6_15_LC_1_13_1.C_ON=1'b0;
    defparam shift_srl_6_15_LC_1_13_1.SEQ_MODE=4'b1000;
    defparam shift_srl_6_15_LC_1_13_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_6_15_LC_1_13_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48391),
            .lcout(shift_srl_6Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92922),
            .ce(N__48812),
            .sr(_gnd_net_));
    defparam shift_srl_6_14_LC_1_13_2.C_ON=1'b0;
    defparam shift_srl_6_14_LC_1_13_2.SEQ_MODE=4'b1000;
    defparam shift_srl_6_14_LC_1_13_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_6_14_LC_1_13_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48385),
            .lcout(shift_srl_6Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92922),
            .ce(N__48812),
            .sr(_gnd_net_));
    defparam shift_srl_6_13_LC_1_13_3.C_ON=1'b0;
    defparam shift_srl_6_13_LC_1_13_3.SEQ_MODE=4'b1000;
    defparam shift_srl_6_13_LC_1_13_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_6_13_LC_1_13_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48379),
            .lcout(shift_srl_6Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92922),
            .ce(N__48812),
            .sr(_gnd_net_));
    defparam shift_srl_6_12_LC_1_13_4.C_ON=1'b0;
    defparam shift_srl_6_12_LC_1_13_4.SEQ_MODE=4'b1000;
    defparam shift_srl_6_12_LC_1_13_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_6_12_LC_1_13_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48373),
            .lcout(shift_srl_6Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92922),
            .ce(N__48812),
            .sr(_gnd_net_));
    defparam shift_srl_6_11_LC_1_13_5.C_ON=1'b0;
    defparam shift_srl_6_11_LC_1_13_5.SEQ_MODE=4'b1000;
    defparam shift_srl_6_11_LC_1_13_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_6_11_LC_1_13_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48367),
            .lcout(shift_srl_6Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92922),
            .ce(N__48812),
            .sr(_gnd_net_));
    defparam shift_srl_6_10_LC_1_13_6.C_ON=1'b0;
    defparam shift_srl_6_10_LC_1_13_6.SEQ_MODE=4'b1000;
    defparam shift_srl_6_10_LC_1_13_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_6_10_LC_1_13_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48361),
            .lcout(shift_srl_6Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92922),
            .ce(N__48812),
            .sr(_gnd_net_));
    defparam shift_srl_6_9_LC_1_13_7.C_ON=1'b0;
    defparam shift_srl_6_9_LC_1_13_7.SEQ_MODE=4'b1000;
    defparam shift_srl_6_9_LC_1_13_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_6_9_LC_1_13_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48715),
            .lcout(shift_srl_6Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92922),
            .ce(N__48812),
            .sr(_gnd_net_));
    defparam shift_srl_5_10_LC_1_14_0.C_ON=1'b0;
    defparam shift_srl_5_10_LC_1_14_0.SEQ_MODE=4'b1000;
    defparam shift_srl_5_10_LC_1_14_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_5_10_LC_1_14_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48436),
            .lcout(shift_srl_5Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92916),
            .ce(N__48471),
            .sr(_gnd_net_));
    defparam shift_srl_5_11_LC_1_14_1.C_ON=1'b0;
    defparam shift_srl_5_11_LC_1_14_1.SEQ_MODE=4'b1000;
    defparam shift_srl_5_11_LC_1_14_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_5_11_LC_1_14_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48355),
            .lcout(shift_srl_5Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92916),
            .ce(N__48471),
            .sr(_gnd_net_));
    defparam shift_srl_5_12_LC_1_14_2.C_ON=1'b0;
    defparam shift_srl_5_12_LC_1_14_2.SEQ_MODE=4'b1000;
    defparam shift_srl_5_12_LC_1_14_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_5_12_LC_1_14_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48349),
            .lcout(shift_srl_5Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92916),
            .ce(N__48471),
            .sr(_gnd_net_));
    defparam shift_srl_5_13_LC_1_14_3.C_ON=1'b0;
    defparam shift_srl_5_13_LC_1_14_3.SEQ_MODE=4'b1000;
    defparam shift_srl_5_13_LC_1_14_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_5_13_LC_1_14_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48454),
            .lcout(shift_srl_5Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92916),
            .ce(N__48471),
            .sr(_gnd_net_));
    defparam shift_srl_5_14_LC_1_14_4.C_ON=1'b0;
    defparam shift_srl_5_14_LC_1_14_4.SEQ_MODE=4'b1000;
    defparam shift_srl_5_14_LC_1_14_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_5_14_LC_1_14_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48448),
            .lcout(shift_srl_5Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92916),
            .ce(N__48471),
            .sr(_gnd_net_));
    defparam shift_srl_5_15_LC_1_14_5.C_ON=1'b0;
    defparam shift_srl_5_15_LC_1_14_5.SEQ_MODE=4'b1000;
    defparam shift_srl_5_15_LC_1_14_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_5_15_LC_1_14_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48442),
            .lcout(shift_srl_5Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92916),
            .ce(N__48471),
            .sr(_gnd_net_));
    defparam shift_srl_5_9_LC_1_14_6.C_ON=1'b0;
    defparam shift_srl_5_9_LC_1_14_6.SEQ_MODE=4'b1000;
    defparam shift_srl_5_9_LC_1_14_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_5_9_LC_1_14_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48430),
            .lcout(shift_srl_5Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92916),
            .ce(N__48471),
            .sr(_gnd_net_));
    defparam shift_srl_5_8_LC_1_14_7.C_ON=1'b0;
    defparam shift_srl_5_8_LC_1_14_7.SEQ_MODE=4'b1000;
    defparam shift_srl_5_8_LC_1_14_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_5_8_LC_1_14_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48505),
            .lcout(shift_srl_5Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92916),
            .ce(N__48471),
            .sr(_gnd_net_));
    defparam shift_srl_5_RNI4Q2G1_15_LC_1_15_0.C_ON=1'b0;
    defparam shift_srl_5_RNI4Q2G1_15_LC_1_15_0.SEQ_MODE=4'b0000;
    defparam shift_srl_5_RNI4Q2G1_15_LC_1_15_0.LUT_INIT=16'b0100000000000000;
    LogicCell40 shift_srl_5_RNI4Q2G1_15_LC_1_15_0 (
            .in0(N__53728),
            .in1(N__49340),
            .in2(N__49318),
            .in3(N__49474),
            .lcout(rco_c_5),
            .ltout(rco_c_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIV5TG1_15_LC_1_15_1.C_ON=1'b0;
    defparam shift_srl_0_RNIV5TG1_15_LC_1_15_1.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIV5TG1_15_LC_1_15_1.LUT_INIT=16'b1111000000000000;
    LogicCell40 shift_srl_0_RNIV5TG1_15_LC_1_15_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__48409),
            .in3(N__89787),
            .lcout(clk_en_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_4_RNI4Q9A1_15_LC_1_15_2.C_ON=1'b0;
    defparam shift_srl_4_RNI4Q9A1_15_LC_1_15_2.SEQ_MODE=4'b0000;
    defparam shift_srl_4_RNI4Q9A1_15_LC_1_15_2.LUT_INIT=16'b0101000000000000;
    LogicCell40 shift_srl_4_RNI4Q9A1_15_LC_1_15_2 (
            .in0(N__53727),
            .in1(_gnd_net_),
            .in2(N__49317),
            .in3(N__49473),
            .lcout(rco_c_4),
            .ltout(rco_c_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIV54B1_15_LC_1_15_3.C_ON=1'b0;
    defparam shift_srl_0_RNIV54B1_15_LC_1_15_3.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIV54B1_15_LC_1_15_3.LUT_INIT=16'b1111000000000000;
    LogicCell40 shift_srl_0_RNIV54B1_15_LC_1_15_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__48394),
            .in3(N__89788),
            .lcout(clk_en_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_5_0_LC_1_15_4.C_ON=1'b0;
    defparam shift_srl_5_0_LC_1_15_4.SEQ_MODE=4'b1000;
    defparam shift_srl_5_0_LC_1_15_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_5_0_LC_1_15_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49341),
            .lcout(shift_srl_5Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92911),
            .ce(N__48470),
            .sr(_gnd_net_));
    defparam shift_srl_5_4_LC_1_16_0.C_ON=1'b0;
    defparam shift_srl_5_4_LC_1_16_0.SEQ_MODE=4'b1000;
    defparam shift_srl_5_4_LC_1_16_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_5_4_LC_1_16_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48496),
            .lcout(shift_srl_5Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92908),
            .ce(N__48472),
            .sr(_gnd_net_));
    defparam shift_srl_5_5_LC_1_16_1.C_ON=1'b0;
    defparam shift_srl_5_5_LC_1_16_1.SEQ_MODE=4'b1000;
    defparam shift_srl_5_5_LC_1_16_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_5_5_LC_1_16_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48523),
            .lcout(shift_srl_5Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92908),
            .ce(N__48472),
            .sr(_gnd_net_));
    defparam shift_srl_5_6_LC_1_16_2.C_ON=1'b0;
    defparam shift_srl_5_6_LC_1_16_2.SEQ_MODE=4'b1000;
    defparam shift_srl_5_6_LC_1_16_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_5_6_LC_1_16_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48517),
            .lcout(shift_srl_5Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92908),
            .ce(N__48472),
            .sr(_gnd_net_));
    defparam shift_srl_5_7_LC_1_16_3.C_ON=1'b0;
    defparam shift_srl_5_7_LC_1_16_3.SEQ_MODE=4'b1000;
    defparam shift_srl_5_7_LC_1_16_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_5_7_LC_1_16_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48511),
            .lcout(shift_srl_5Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92908),
            .ce(N__48472),
            .sr(_gnd_net_));
    defparam shift_srl_5_3_LC_1_16_4.C_ON=1'b0;
    defparam shift_srl_5_3_LC_1_16_4.SEQ_MODE=4'b1000;
    defparam shift_srl_5_3_LC_1_16_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_5_3_LC_1_16_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48478),
            .lcout(shift_srl_5Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92908),
            .ce(N__48472),
            .sr(_gnd_net_));
    defparam shift_srl_5_1_LC_1_16_6.C_ON=1'b0;
    defparam shift_srl_5_1_LC_1_16_6.SEQ_MODE=4'b1000;
    defparam shift_srl_5_1_LC_1_16_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_5_1_LC_1_16_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48490),
            .lcout(shift_srl_5Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92908),
            .ce(N__48472),
            .sr(_gnd_net_));
    defparam shift_srl_5_2_LC_1_16_7.C_ON=1'b0;
    defparam shift_srl_5_2_LC_1_16_7.SEQ_MODE=4'b1000;
    defparam shift_srl_5_2_LC_1_16_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_5_2_LC_1_16_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48484),
            .lcout(shift_srl_5Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92908),
            .ce(N__48472),
            .sr(_gnd_net_));
    defparam shift_srl_130_8_LC_1_18_0.C_ON=1'b0;
    defparam shift_srl_130_8_LC_1_18_0.SEQ_MODE=4'b1000;
    defparam shift_srl_130_8_LC_1_18_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_130_8_LC_1_18_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48559),
            .lcout(shift_srl_130Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92909),
            .ce(N__49882),
            .sr(_gnd_net_));
    defparam shift_srl_130_9_LC_1_18_1.C_ON=1'b0;
    defparam shift_srl_130_9_LC_1_18_1.SEQ_MODE=4'b1000;
    defparam shift_srl_130_9_LC_1_18_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_130_9_LC_1_18_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48571),
            .lcout(shift_srl_130Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92909),
            .ce(N__49882),
            .sr(_gnd_net_));
    defparam shift_srl_130_6_LC_1_18_2.C_ON=1'b0;
    defparam shift_srl_130_6_LC_1_18_2.SEQ_MODE=4'b1000;
    defparam shift_srl_130_6_LC_1_18_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_130_6_LC_1_18_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48916),
            .lcout(shift_srl_130Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92909),
            .ce(N__49882),
            .sr(_gnd_net_));
    defparam shift_srl_130_7_LC_1_18_4.C_ON=1'b0;
    defparam shift_srl_130_7_LC_1_18_4.SEQ_MODE=4'b1000;
    defparam shift_srl_130_7_LC_1_18_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_130_7_LC_1_18_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48565),
            .lcout(shift_srl_130Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92909),
            .ce(N__49882),
            .sr(_gnd_net_));
    defparam shift_srl_137_0_LC_1_19_0.C_ON=1'b0;
    defparam shift_srl_137_0_LC_1_19_0.SEQ_MODE=4'b1000;
    defparam shift_srl_137_0_LC_1_19_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_137_0_LC_1_19_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51268),
            .lcout(shift_srl_137Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92912),
            .ce(N__49986),
            .sr(_gnd_net_));
    defparam shift_srl_137_1_LC_1_19_1.C_ON=1'b0;
    defparam shift_srl_137_1_LC_1_19_1.SEQ_MODE=4'b1000;
    defparam shift_srl_137_1_LC_1_19_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_137_1_LC_1_19_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48553),
            .lcout(shift_srl_137Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92912),
            .ce(N__49986),
            .sr(_gnd_net_));
    defparam shift_srl_137_2_LC_1_19_2.C_ON=1'b0;
    defparam shift_srl_137_2_LC_1_19_2.SEQ_MODE=4'b1000;
    defparam shift_srl_137_2_LC_1_19_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_137_2_LC_1_19_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48547),
            .lcout(shift_srl_137Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92912),
            .ce(N__49986),
            .sr(_gnd_net_));
    defparam shift_srl_137_3_LC_1_19_3.C_ON=1'b0;
    defparam shift_srl_137_3_LC_1_19_3.SEQ_MODE=4'b1000;
    defparam shift_srl_137_3_LC_1_19_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_137_3_LC_1_19_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48541),
            .lcout(shift_srl_137Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92912),
            .ce(N__49986),
            .sr(_gnd_net_));
    defparam shift_srl_137_4_LC_1_19_4.C_ON=1'b0;
    defparam shift_srl_137_4_LC_1_19_4.SEQ_MODE=4'b1000;
    defparam shift_srl_137_4_LC_1_19_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_137_4_LC_1_19_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48535),
            .lcout(shift_srl_137Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92912),
            .ce(N__49986),
            .sr(_gnd_net_));
    defparam shift_srl_137_5_LC_1_19_5.C_ON=1'b0;
    defparam shift_srl_137_5_LC_1_19_5.SEQ_MODE=4'b1000;
    defparam shift_srl_137_5_LC_1_19_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_137_5_LC_1_19_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48529),
            .lcout(shift_srl_137Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92912),
            .ce(N__49986),
            .sr(_gnd_net_));
    defparam shift_srl_137_6_LC_1_19_6.C_ON=1'b0;
    defparam shift_srl_137_6_LC_1_19_6.SEQ_MODE=4'b1000;
    defparam shift_srl_137_6_LC_1_19_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_137_6_LC_1_19_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48613),
            .lcout(shift_srl_137Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92912),
            .ce(N__49986),
            .sr(_gnd_net_));
    defparam shift_srl_137_7_LC_1_19_7.C_ON=1'b0;
    defparam shift_srl_137_7_LC_1_19_7.SEQ_MODE=4'b1000;
    defparam shift_srl_137_7_LC_1_19_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_137_7_LC_1_19_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48607),
            .lcout(shift_srl_137Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92912),
            .ce(N__49986),
            .sr(_gnd_net_));
    defparam shift_srl_136_15_LC_1_20_3.C_ON=1'b0;
    defparam shift_srl_136_15_LC_1_20_3.SEQ_MODE=4'b1000;
    defparam shift_srl_136_15_LC_1_20_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_136_15_LC_1_20_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48964),
            .lcout(shift_srl_136Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92917),
            .ce(N__49954),
            .sr(_gnd_net_));
    defparam shift_srl_22_4_LC_2_7_3.C_ON=1'b0;
    defparam shift_srl_22_4_LC_2_7_3.SEQ_MODE=4'b1000;
    defparam shift_srl_22_4_LC_2_7_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_22_4_LC_2_7_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48601),
            .lcout(shift_srl_22Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93001),
            .ce(N__52207),
            .sr(_gnd_net_));
    defparam shift_srl_22_3_LC_2_7_4.C_ON=1'b0;
    defparam shift_srl_22_3_LC_2_7_4.SEQ_MODE=4'b1000;
    defparam shift_srl_22_3_LC_2_7_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_22_3_LC_2_7_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49060),
            .lcout(shift_srl_22Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93001),
            .ce(N__52207),
            .sr(_gnd_net_));
    defparam shift_srl_22_5_LC_2_7_6.C_ON=1'b0;
    defparam shift_srl_22_5_LC_2_7_6.SEQ_MODE=4'b1000;
    defparam shift_srl_22_5_LC_2_7_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_22_5_LC_2_7_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48595),
            .lcout(shift_srl_22Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93001),
            .ce(N__52207),
            .sr(_gnd_net_));
    defparam shift_srl_22_6_LC_2_7_7.C_ON=1'b0;
    defparam shift_srl_22_6_LC_2_7_7.SEQ_MODE=4'b1000;
    defparam shift_srl_22_6_LC_2_7_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_22_6_LC_2_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48589),
            .lcout(shift_srl_22Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93001),
            .ce(N__52207),
            .sr(_gnd_net_));
    defparam shift_srl_22_7_LC_2_8_0.C_ON=1'b0;
    defparam shift_srl_22_7_LC_2_8_0.SEQ_MODE=4'b1000;
    defparam shift_srl_22_7_LC_2_8_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_22_7_LC_2_8_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48583),
            .lcout(shift_srl_22Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92986),
            .ce(N__52201),
            .sr(_gnd_net_));
    defparam shift_srl_22_0_LC_2_8_1.C_ON=1'b0;
    defparam shift_srl_22_0_LC_2_8_1.SEQ_MODE=4'b1000;
    defparam shift_srl_22_0_LC_2_8_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_22_0_LC_2_8_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53433),
            .lcout(shift_srl_22Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92986),
            .ce(N__52201),
            .sr(_gnd_net_));
    defparam shift_srl_22_1_LC_2_8_3.C_ON=1'b0;
    defparam shift_srl_22_1_LC_2_8_3.SEQ_MODE=4'b1000;
    defparam shift_srl_22_1_LC_2_8_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_22_1_LC_2_8_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48577),
            .lcout(shift_srl_22Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92986),
            .ce(N__52201),
            .sr(_gnd_net_));
    defparam shift_srl_13_0_LC_2_9_0.C_ON=1'b0;
    defparam shift_srl_13_0_LC_2_9_0.SEQ_MODE=4'b1000;
    defparam shift_srl_13_0_LC_2_9_0.LUT_INIT=16'b1100110011001100;
    LogicCell40 shift_srl_13_0_LC_2_9_0 (
            .in0(_gnd_net_),
            .in1(N__50778),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_13Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92973),
            .ce(N__49569),
            .sr(_gnd_net_));
    defparam shift_srl_13_2_LC_2_9_2.C_ON=1'b0;
    defparam shift_srl_13_2_LC_2_9_2.SEQ_MODE=4'b1000;
    defparam shift_srl_13_2_LC_2_9_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_13_2_LC_2_9_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48643),
            .lcout(shift_srl_13Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92973),
            .ce(N__49569),
            .sr(_gnd_net_));
    defparam shift_srl_13_3_LC_2_9_3.C_ON=1'b0;
    defparam shift_srl_13_3_LC_2_9_3.SEQ_MODE=4'b1000;
    defparam shift_srl_13_3_LC_2_9_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_13_3_LC_2_9_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48661),
            .lcout(shift_srl_13Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92973),
            .ce(N__49569),
            .sr(_gnd_net_));
    defparam shift_srl_13_1_LC_2_9_4.C_ON=1'b0;
    defparam shift_srl_13_1_LC_2_9_4.SEQ_MODE=4'b1000;
    defparam shift_srl_13_1_LC_2_9_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_13_1_LC_2_9_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48649),
            .lcout(shift_srl_13Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92973),
            .ce(N__49569),
            .sr(_gnd_net_));
    defparam shift_srl_13_5_LC_2_9_5.C_ON=1'b0;
    defparam shift_srl_13_5_LC_2_9_5.SEQ_MODE=4'b1000;
    defparam shift_srl_13_5_LC_2_9_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_13_5_LC_2_9_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48637),
            .lcout(shift_srl_13Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92973),
            .ce(N__49569),
            .sr(_gnd_net_));
    defparam shift_srl_13_6_LC_2_9_6.C_ON=1'b0;
    defparam shift_srl_13_6_LC_2_9_6.SEQ_MODE=4'b1000;
    defparam shift_srl_13_6_LC_2_9_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_13_6_LC_2_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48631),
            .lcout(shift_srl_13Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92973),
            .ce(N__49569),
            .sr(_gnd_net_));
    defparam shift_srl_13_7_LC_2_9_7.C_ON=1'b0;
    defparam shift_srl_13_7_LC_2_9_7.SEQ_MODE=4'b1000;
    defparam shift_srl_13_7_LC_2_9_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_13_7_LC_2_9_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48625),
            .lcout(shift_srl_13Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92973),
            .ce(N__49569),
            .sr(_gnd_net_));
    defparam shift_srl_12_7_LC_2_10_0.C_ON=1'b0;
    defparam shift_srl_12_7_LC_2_10_0.SEQ_MODE=4'b1000;
    defparam shift_srl_12_7_LC_2_10_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_12_7_LC_2_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48703),
            .lcout(shift_srl_12Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92962),
            .ce(N__49395),
            .sr(_gnd_net_));
    defparam shift_srl_12_8_LC_2_10_1.C_ON=1'b0;
    defparam shift_srl_12_8_LC_2_10_1.SEQ_MODE=4'b1000;
    defparam shift_srl_12_8_LC_2_10_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_12_8_LC_2_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48619),
            .lcout(shift_srl_12Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92962),
            .ce(N__49395),
            .sr(_gnd_net_));
    defparam shift_srl_12_6_LC_2_10_2.C_ON=1'b0;
    defparam shift_srl_12_6_LC_2_10_2.SEQ_MODE=4'b1000;
    defparam shift_srl_12_6_LC_2_10_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_12_6_LC_2_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48667),
            .lcout(shift_srl_12Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92962),
            .ce(N__49395),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNI2HF43_15_LC_2_11_0.C_ON=1'b0;
    defparam shift_srl_0_RNI2HF43_15_LC_2_11_0.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNI2HF43_15_LC_2_11_0.LUT_INIT=16'b1010101000000000;
    LogicCell40 shift_srl_0_RNI2HF43_15_LC_2_11_0 (
            .in0(N__50373),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__89524),
            .lcout(clk_en_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_12_0_LC_2_11_1.C_ON=1'b0;
    defparam shift_srl_12_0_LC_2_11_1.SEQ_MODE=4'b1000;
    defparam shift_srl_12_0_LC_2_11_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_12_0_LC_2_11_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50815),
            .lcout(shift_srl_12Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92949),
            .ce(N__49394),
            .sr(_gnd_net_));
    defparam shift_srl_12_1_LC_2_11_2.C_ON=1'b0;
    defparam shift_srl_12_1_LC_2_11_2.SEQ_MODE=4'b1000;
    defparam shift_srl_12_1_LC_2_11_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_12_1_LC_2_11_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48697),
            .lcout(shift_srl_12Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92949),
            .ce(N__49394),
            .sr(_gnd_net_));
    defparam shift_srl_12_2_LC_2_11_3.C_ON=1'b0;
    defparam shift_srl_12_2_LC_2_11_3.SEQ_MODE=4'b1000;
    defparam shift_srl_12_2_LC_2_11_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_12_2_LC_2_11_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48691),
            .lcout(shift_srl_12Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92949),
            .ce(N__49394),
            .sr(_gnd_net_));
    defparam shift_srl_12_3_LC_2_11_4.C_ON=1'b0;
    defparam shift_srl_12_3_LC_2_11_4.SEQ_MODE=4'b1000;
    defparam shift_srl_12_3_LC_2_11_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_12_3_LC_2_11_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48685),
            .lcout(shift_srl_12Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92949),
            .ce(N__49394),
            .sr(_gnd_net_));
    defparam shift_srl_12_4_LC_2_11_5.C_ON=1'b0;
    defparam shift_srl_12_4_LC_2_11_5.SEQ_MODE=4'b1000;
    defparam shift_srl_12_4_LC_2_11_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_12_4_LC_2_11_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48679),
            .lcout(shift_srl_12Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92949),
            .ce(N__49394),
            .sr(_gnd_net_));
    defparam shift_srl_12_5_LC_2_11_6.C_ON=1'b0;
    defparam shift_srl_12_5_LC_2_11_6.SEQ_MODE=4'b1000;
    defparam shift_srl_12_5_LC_2_11_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_12_5_LC_2_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48673),
            .lcout(shift_srl_12Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92949),
            .ce(N__49394),
            .sr(_gnd_net_));
    defparam shift_srl_4_10_LC_2_12_0.C_ON=1'b0;
    defparam shift_srl_4_10_LC_2_12_0.SEQ_MODE=4'b1000;
    defparam shift_srl_4_10_LC_2_12_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_4_10_LC_2_12_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48745),
            .lcout(shift_srl_4Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92940),
            .ce(N__48727),
            .sr(_gnd_net_));
    defparam shift_srl_4_11_LC_2_12_1.C_ON=1'b0;
    defparam shift_srl_4_11_LC_2_12_1.SEQ_MODE=4'b1000;
    defparam shift_srl_4_11_LC_2_12_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_4_11_LC_2_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48775),
            .lcout(shift_srl_4Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92940),
            .ce(N__48727),
            .sr(_gnd_net_));
    defparam shift_srl_4_12_LC_2_12_2.C_ON=1'b0;
    defparam shift_srl_4_12_LC_2_12_2.SEQ_MODE=4'b1000;
    defparam shift_srl_4_12_LC_2_12_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_4_12_LC_2_12_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48769),
            .lcout(shift_srl_4Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92940),
            .ce(N__48727),
            .sr(_gnd_net_));
    defparam shift_srl_4_13_LC_2_12_3.C_ON=1'b0;
    defparam shift_srl_4_13_LC_2_12_3.SEQ_MODE=4'b1000;
    defparam shift_srl_4_13_LC_2_12_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_4_13_LC_2_12_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48763),
            .lcout(shift_srl_4Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92940),
            .ce(N__48727),
            .sr(_gnd_net_));
    defparam shift_srl_4_14_LC_2_12_4.C_ON=1'b0;
    defparam shift_srl_4_14_LC_2_12_4.SEQ_MODE=4'b1000;
    defparam shift_srl_4_14_LC_2_12_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_4_14_LC_2_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48757),
            .lcout(shift_srl_4Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92940),
            .ce(N__48727),
            .sr(_gnd_net_));
    defparam shift_srl_4_15_LC_2_12_5.C_ON=1'b0;
    defparam shift_srl_4_15_LC_2_12_5.SEQ_MODE=4'b1000;
    defparam shift_srl_4_15_LC_2_12_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_4_15_LC_2_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48751),
            .lcout(shift_srl_4Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92940),
            .ce(N__48727),
            .sr(_gnd_net_));
    defparam shift_srl_4_9_LC_2_12_6.C_ON=1'b0;
    defparam shift_srl_4_9_LC_2_12_6.SEQ_MODE=4'b1000;
    defparam shift_srl_4_9_LC_2_12_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_4_9_LC_2_12_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48733),
            .lcout(shift_srl_4Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92940),
            .ce(N__48727),
            .sr(_gnd_net_));
    defparam shift_srl_4_8_LC_2_12_7.C_ON=1'b0;
    defparam shift_srl_4_8_LC_2_12_7.SEQ_MODE=4'b1000;
    defparam shift_srl_4_8_LC_2_12_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_4_8_LC_2_12_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48739),
            .lcout(shift_srl_4Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92940),
            .ce(N__48727),
            .sr(_gnd_net_));
    defparam shift_srl_6_8_LC_2_13_0.C_ON=1'b0;
    defparam shift_srl_6_8_LC_2_13_0.SEQ_MODE=4'b1000;
    defparam shift_srl_6_8_LC_2_13_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_6_8_LC_2_13_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48709),
            .lcout(shift_srl_6Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92931),
            .ce(N__48816),
            .sr(_gnd_net_));
    defparam shift_srl_6_7_LC_2_13_6.C_ON=1'b0;
    defparam shift_srl_6_7_LC_2_13_6.SEQ_MODE=4'b1000;
    defparam shift_srl_6_7_LC_2_13_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_6_7_LC_2_13_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48826),
            .lcout(shift_srl_6Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92931),
            .ce(N__48816),
            .sr(_gnd_net_));
    defparam shift_srl_6_0_LC_2_14_0.C_ON=1'b0;
    defparam shift_srl_6_0_LC_2_14_0.SEQ_MODE=4'b1000;
    defparam shift_srl_6_0_LC_2_14_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_6_0_LC_2_14_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49367),
            .lcout(shift_srl_6Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92923),
            .ce(N__48820),
            .sr(_gnd_net_));
    defparam shift_srl_6_1_LC_2_14_1.C_ON=1'b0;
    defparam shift_srl_6_1_LC_2_14_1.SEQ_MODE=4'b1000;
    defparam shift_srl_6_1_LC_2_14_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_6_1_LC_2_14_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48862),
            .lcout(shift_srl_6Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92923),
            .ce(N__48820),
            .sr(_gnd_net_));
    defparam shift_srl_6_2_LC_2_14_2.C_ON=1'b0;
    defparam shift_srl_6_2_LC_2_14_2.SEQ_MODE=4'b1000;
    defparam shift_srl_6_2_LC_2_14_2.LUT_INIT=16'b1100110011001100;
    LogicCell40 shift_srl_6_2_LC_2_14_2 (
            .in0(_gnd_net_),
            .in1(N__48856),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_6Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92923),
            .ce(N__48820),
            .sr(_gnd_net_));
    defparam shift_srl_6_3_LC_2_14_3.C_ON=1'b0;
    defparam shift_srl_6_3_LC_2_14_3.SEQ_MODE=4'b1000;
    defparam shift_srl_6_3_LC_2_14_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_6_3_LC_2_14_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48850),
            .lcout(shift_srl_6Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92923),
            .ce(N__48820),
            .sr(_gnd_net_));
    defparam shift_srl_6_4_LC_2_14_4.C_ON=1'b0;
    defparam shift_srl_6_4_LC_2_14_4.SEQ_MODE=4'b1000;
    defparam shift_srl_6_4_LC_2_14_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_6_4_LC_2_14_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48844),
            .lcout(shift_srl_6Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92923),
            .ce(N__48820),
            .sr(_gnd_net_));
    defparam shift_srl_6_5_LC_2_14_5.C_ON=1'b0;
    defparam shift_srl_6_5_LC_2_14_5.SEQ_MODE=4'b1000;
    defparam shift_srl_6_5_LC_2_14_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_6_5_LC_2_14_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48838),
            .lcout(shift_srl_6Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92923),
            .ce(N__48820),
            .sr(_gnd_net_));
    defparam shift_srl_6_6_LC_2_14_6.C_ON=1'b0;
    defparam shift_srl_6_6_LC_2_14_6.SEQ_MODE=4'b1000;
    defparam shift_srl_6_6_LC_2_14_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_6_6_LC_2_14_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48832),
            .lcout(shift_srl_6Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92923),
            .ce(N__48820),
            .sr(_gnd_net_));
    defparam shift_srl_7_0_LC_2_15_0.C_ON=1'b0;
    defparam shift_srl_7_0_LC_2_15_0.SEQ_MODE=4'b1000;
    defparam shift_srl_7_0_LC_2_15_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_7_0_LC_2_15_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53762),
            .lcout(shift_srl_7Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92918),
            .ce(N__49675),
            .sr(_gnd_net_));
    defparam shift_srl_6_RNI5U1Q1_15_LC_2_15_1.C_ON=1'b0;
    defparam shift_srl_6_RNI5U1Q1_15_LC_2_15_1.SEQ_MODE=4'b0000;
    defparam shift_srl_6_RNI5U1Q1_15_LC_2_15_1.LUT_INIT=16'b0011001100000000;
    LogicCell40 shift_srl_6_RNI5U1Q1_15_LC_2_15_1 (
            .in0(_gnd_net_),
            .in1(N__53726),
            .in2(_gnd_net_),
            .in3(N__53639),
            .lcout(rco_c_6),
            .ltout(rco_c_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNI0ASQ1_15_LC_2_15_2.C_ON=1'b0;
    defparam shift_srl_0_RNI0ASQ1_15_LC_2_15_2.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNI0ASQ1_15_LC_2_15_2.LUT_INIT=16'b1111000000000000;
    LogicCell40 shift_srl_0_RNI0ASQ1_15_LC_2_15_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__48907),
            .in3(N__89525),
            .lcout(clk_en_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_7_1_LC_2_15_3.C_ON=1'b0;
    defparam shift_srl_7_1_LC_2_15_3.SEQ_MODE=4'b1000;
    defparam shift_srl_7_1_LC_2_15_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_7_1_LC_2_15_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48904),
            .lcout(shift_srl_7Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92918),
            .ce(N__49675),
            .sr(_gnd_net_));
    defparam shift_srl_7_2_LC_2_15_4.C_ON=1'b0;
    defparam shift_srl_7_2_LC_2_15_4.SEQ_MODE=4'b1000;
    defparam shift_srl_7_2_LC_2_15_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_7_2_LC_2_15_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48898),
            .lcout(shift_srl_7Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92918),
            .ce(N__49675),
            .sr(_gnd_net_));
    defparam shift_srl_7_3_LC_2_15_5.C_ON=1'b0;
    defparam shift_srl_7_3_LC_2_15_5.SEQ_MODE=4'b1000;
    defparam shift_srl_7_3_LC_2_15_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_7_3_LC_2_15_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48892),
            .lcout(shift_srl_7Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92918),
            .ce(N__49675),
            .sr(_gnd_net_));
    defparam shift_srl_7_4_LC_2_15_6.C_ON=1'b0;
    defparam shift_srl_7_4_LC_2_15_6.SEQ_MODE=4'b1000;
    defparam shift_srl_7_4_LC_2_15_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_7_4_LC_2_15_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48886),
            .lcout(shift_srl_7Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92918),
            .ce(N__49675),
            .sr(_gnd_net_));
    defparam shift_srl_7_6_LC_2_16_0.C_ON=1'b0;
    defparam shift_srl_7_6_LC_2_16_0.SEQ_MODE=4'b1000;
    defparam shift_srl_7_6_LC_2_16_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_7_6_LC_2_16_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48874),
            .lcout(shift_srl_7Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92913),
            .ce(N__49676),
            .sr(_gnd_net_));
    defparam shift_srl_7_5_LC_2_16_4.C_ON=1'b0;
    defparam shift_srl_7_5_LC_2_16_4.SEQ_MODE=4'b1000;
    defparam shift_srl_7_5_LC_2_16_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_7_5_LC_2_16_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48880),
            .lcout(shift_srl_7Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92913),
            .ce(N__49676),
            .sr(_gnd_net_));
    defparam shift_srl_129_8_LC_2_17_0.C_ON=1'b0;
    defparam shift_srl_129_8_LC_2_17_0.SEQ_MODE=4'b1000;
    defparam shift_srl_129_8_LC_2_17_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_129_8_LC_2_17_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49801),
            .lcout(shift_srl_129Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92907),
            .ce(N__53994),
            .sr(_gnd_net_));
    defparam shift_srl_129_9_LC_2_17_1.C_ON=1'b0;
    defparam shift_srl_129_9_LC_2_17_1.SEQ_MODE=4'b1000;
    defparam shift_srl_129_9_LC_2_17_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_129_9_LC_2_17_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48868),
            .lcout(shift_srl_129Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92907),
            .ce(N__53994),
            .sr(_gnd_net_));
    defparam shift_srl_130_0_LC_2_18_0.C_ON=1'b0;
    defparam shift_srl_130_0_LC_2_18_0.SEQ_MODE=4'b1000;
    defparam shift_srl_130_0_LC_2_18_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_130_0_LC_2_18_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52927),
            .lcout(shift_srl_130Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92914),
            .ce(N__49877),
            .sr(_gnd_net_));
    defparam shift_srl_130_1_LC_2_18_1.C_ON=1'b0;
    defparam shift_srl_130_1_LC_2_18_1.SEQ_MODE=4'b1000;
    defparam shift_srl_130_1_LC_2_18_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_130_1_LC_2_18_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48946),
            .lcout(shift_srl_130Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92914),
            .ce(N__49877),
            .sr(_gnd_net_));
    defparam shift_srl_130_2_LC_2_18_2.C_ON=1'b0;
    defparam shift_srl_130_2_LC_2_18_2.SEQ_MODE=4'b1000;
    defparam shift_srl_130_2_LC_2_18_2.LUT_INIT=16'b1100110011001100;
    LogicCell40 shift_srl_130_2_LC_2_18_2 (
            .in0(_gnd_net_),
            .in1(N__48940),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_130Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92914),
            .ce(N__49877),
            .sr(_gnd_net_));
    defparam shift_srl_130_3_LC_2_18_3.C_ON=1'b0;
    defparam shift_srl_130_3_LC_2_18_3.SEQ_MODE=4'b1000;
    defparam shift_srl_130_3_LC_2_18_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_130_3_LC_2_18_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48934),
            .lcout(shift_srl_130Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92914),
            .ce(N__49877),
            .sr(_gnd_net_));
    defparam shift_srl_130_4_LC_2_18_4.C_ON=1'b0;
    defparam shift_srl_130_4_LC_2_18_4.SEQ_MODE=4'b1000;
    defparam shift_srl_130_4_LC_2_18_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_130_4_LC_2_18_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48928),
            .lcout(shift_srl_130Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92914),
            .ce(N__49877),
            .sr(_gnd_net_));
    defparam shift_srl_130_5_LC_2_18_5.C_ON=1'b0;
    defparam shift_srl_130_5_LC_2_18_5.SEQ_MODE=4'b1000;
    defparam shift_srl_130_5_LC_2_18_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_130_5_LC_2_18_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48922),
            .lcout(shift_srl_130Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92914),
            .ce(N__49877),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIORHN01_15_LC_2_19_0.C_ON=1'b0;
    defparam shift_srl_0_RNIORHN01_15_LC_2_19_0.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIORHN01_15_LC_2_19_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNIORHN01_15_LC_2_19_0 (
            .in0(N__90420),
            .in1(N__65751),
            .in2(N__91374),
            .in3(N__57616),
            .lcout(clk_en_130),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_129_RNIDM4D_15_LC_2_19_1.C_ON=1'b0;
    defparam shift_srl_129_RNIDM4D_15_LC_2_19_1.SEQ_MODE=4'b0000;
    defparam shift_srl_129_RNIDM4D_15_LC_2_19_1.LUT_INIT=16'b1100110000000000;
    LogicCell40 shift_srl_129_RNIDM4D_15_LC_2_19_1 (
            .in0(_gnd_net_),
            .in1(N__91246),
            .in2(_gnd_net_),
            .in3(N__54234),
            .lcout(shift_srl_129_RNIDM4DZ0Z_15),
            .ltout(shift_srl_129_RNIDM4DZ0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_129_RNIVMDO2_15_LC_2_19_2.C_ON=1'b0;
    defparam shift_srl_129_RNIVMDO2_15_LC_2_19_2.SEQ_MODE=4'b0000;
    defparam shift_srl_129_RNIVMDO2_15_LC_2_19_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_129_RNIVMDO2_15_LC_2_19_2 (
            .in0(N__65567),
            .in1(N__65750),
            .in2(N__48910),
            .in3(N__65363),
            .lcout(g0_16_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_135_RNI46TQ_15_LC_2_19_3.C_ON=1'b0;
    defparam shift_srl_135_RNI46TQ_15_LC_2_19_3.SEQ_MODE=4'b0000;
    defparam shift_srl_135_RNI46TQ_15_LC_2_19_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_135_RNI46TQ_15_LC_2_19_3 (
            .in0(N__89786),
            .in1(N__53103),
            .in2(N__66257),
            .in3(N__52021),
            .lcout(),
            .ltout(g0_11_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_135_RNILIJH3_15_LC_2_19_4.C_ON=1'b0;
    defparam shift_srl_135_RNILIJH3_15_LC_2_19_4.SEQ_MODE=4'b0000;
    defparam shift_srl_135_RNILIJH3_15_LC_2_19_4.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_135_RNILIJH3_15_LC_2_19_4 (
            .in0(N__54433),
            .in1(N__56458),
            .in2(N__49000),
            .in3(N__49795),
            .lcout(),
            .ltout(g0_17_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_107_RNI6IDC21_15_LC_2_19_5.C_ON=1'b0;
    defparam shift_srl_107_RNI6IDC21_15_LC_2_19_5.SEQ_MODE=4'b0000;
    defparam shift_srl_107_RNI6IDC21_15_LC_2_19_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_107_RNI6IDC21_15_LC_2_19_5 (
            .in0(N__48997),
            .in1(N__64990),
            .in2(N__48991),
            .in3(N__79551),
            .lcout(clk_en_137),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_136_10_LC_2_20_0.C_ON=1'b0;
    defparam shift_srl_136_10_LC_2_20_0.SEQ_MODE=4'b1000;
    defparam shift_srl_136_10_LC_2_20_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_136_10_LC_2_20_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48958),
            .lcout(shift_srl_136Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92924),
            .ce(N__49953),
            .sr(_gnd_net_));
    defparam shift_srl_136_11_LC_2_20_1.C_ON=1'b0;
    defparam shift_srl_136_11_LC_2_20_1.SEQ_MODE=4'b1000;
    defparam shift_srl_136_11_LC_2_20_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_136_11_LC_2_20_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48988),
            .lcout(shift_srl_136Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92924),
            .ce(N__49953),
            .sr(_gnd_net_));
    defparam shift_srl_136_12_LC_2_20_2.C_ON=1'b0;
    defparam shift_srl_136_12_LC_2_20_2.SEQ_MODE=4'b1000;
    defparam shift_srl_136_12_LC_2_20_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_136_12_LC_2_20_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48982),
            .lcout(shift_srl_136Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92924),
            .ce(N__49953),
            .sr(_gnd_net_));
    defparam shift_srl_136_13_LC_2_20_3.C_ON=1'b0;
    defparam shift_srl_136_13_LC_2_20_3.SEQ_MODE=4'b1000;
    defparam shift_srl_136_13_LC_2_20_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_136_13_LC_2_20_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48976),
            .lcout(shift_srl_136Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92924),
            .ce(N__49953),
            .sr(_gnd_net_));
    defparam shift_srl_136_14_LC_2_20_4.C_ON=1'b0;
    defparam shift_srl_136_14_LC_2_20_4.SEQ_MODE=4'b1000;
    defparam shift_srl_136_14_LC_2_20_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_136_14_LC_2_20_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48970),
            .lcout(shift_srl_136Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92924),
            .ce(N__49953),
            .sr(_gnd_net_));
    defparam shift_srl_136_9_LC_2_20_6.C_ON=1'b0;
    defparam shift_srl_136_9_LC_2_20_6.SEQ_MODE=4'b1000;
    defparam shift_srl_136_9_LC_2_20_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_136_9_LC_2_20_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48952),
            .lcout(shift_srl_136Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92924),
            .ce(N__49953),
            .sr(_gnd_net_));
    defparam shift_srl_136_8_LC_2_20_7.C_ON=1'b0;
    defparam shift_srl_136_8_LC_2_20_7.SEQ_MODE=4'b1000;
    defparam shift_srl_136_8_LC_2_20_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_136_8_LC_2_20_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49006),
            .lcout(shift_srl_136Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92924),
            .ce(N__49953),
            .sr(_gnd_net_));
    defparam shift_srl_136_0_LC_2_21_0.C_ON=1'b0;
    defparam shift_srl_136_0_LC_2_21_0.SEQ_MODE=4'b1000;
    defparam shift_srl_136_0_LC_2_21_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_136_0_LC_2_21_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54460),
            .lcout(shift_srl_136Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92932),
            .ce(N__49952),
            .sr(_gnd_net_));
    defparam shift_srl_136_1_LC_2_21_1.C_ON=1'b0;
    defparam shift_srl_136_1_LC_2_21_1.SEQ_MODE=4'b1000;
    defparam shift_srl_136_1_LC_2_21_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_136_1_LC_2_21_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49048),
            .lcout(shift_srl_136Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92932),
            .ce(N__49952),
            .sr(_gnd_net_));
    defparam shift_srl_136_2_LC_2_21_2.C_ON=1'b0;
    defparam shift_srl_136_2_LC_2_21_2.SEQ_MODE=4'b1000;
    defparam shift_srl_136_2_LC_2_21_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_136_2_LC_2_21_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49042),
            .lcout(shift_srl_136Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92932),
            .ce(N__49952),
            .sr(_gnd_net_));
    defparam shift_srl_136_3_LC_2_21_3.C_ON=1'b0;
    defparam shift_srl_136_3_LC_2_21_3.SEQ_MODE=4'b1000;
    defparam shift_srl_136_3_LC_2_21_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_136_3_LC_2_21_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49036),
            .lcout(shift_srl_136Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92932),
            .ce(N__49952),
            .sr(_gnd_net_));
    defparam shift_srl_136_4_LC_2_21_4.C_ON=1'b0;
    defparam shift_srl_136_4_LC_2_21_4.SEQ_MODE=4'b1000;
    defparam shift_srl_136_4_LC_2_21_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_136_4_LC_2_21_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49030),
            .lcout(shift_srl_136Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92932),
            .ce(N__49952),
            .sr(_gnd_net_));
    defparam shift_srl_136_5_LC_2_21_5.C_ON=1'b0;
    defparam shift_srl_136_5_LC_2_21_5.SEQ_MODE=4'b1000;
    defparam shift_srl_136_5_LC_2_21_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_136_5_LC_2_21_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49024),
            .lcout(shift_srl_136Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92932),
            .ce(N__49952),
            .sr(_gnd_net_));
    defparam shift_srl_136_6_LC_2_21_6.C_ON=1'b0;
    defparam shift_srl_136_6_LC_2_21_6.SEQ_MODE=4'b1000;
    defparam shift_srl_136_6_LC_2_21_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_136_6_LC_2_21_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49018),
            .lcout(shift_srl_136Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92932),
            .ce(N__49952),
            .sr(_gnd_net_));
    defparam shift_srl_136_7_LC_2_21_7.C_ON=1'b0;
    defparam shift_srl_136_7_LC_2_21_7.SEQ_MODE=4'b1000;
    defparam shift_srl_136_7_LC_2_21_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_136_7_LC_2_21_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49012),
            .lcout(shift_srl_136Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92932),
            .ce(N__49952),
            .sr(_gnd_net_));
    defparam shift_srl_138_11_LC_2_22_0.C_ON=1'b0;
    defparam shift_srl_138_11_LC_2_22_0.SEQ_MODE=4'b1000;
    defparam shift_srl_138_11_LC_2_22_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_138_11_LC_2_22_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49072),
            .lcout(shift_srl_138Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92941),
            .ce(N__50038),
            .sr(_gnd_net_));
    defparam shift_srl_138_1_LC_2_22_1.C_ON=1'b0;
    defparam shift_srl_138_1_LC_2_22_1.SEQ_MODE=4'b1000;
    defparam shift_srl_138_1_LC_2_22_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_138_1_LC_2_22_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49078),
            .lcout(shift_srl_138Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92941),
            .ce(N__50038),
            .sr(_gnd_net_));
    defparam shift_srl_138_2_LC_2_22_2.C_ON=1'b0;
    defparam shift_srl_138_2_LC_2_22_2.SEQ_MODE=4'b1000;
    defparam shift_srl_138_2_LC_2_22_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_138_2_LC_2_22_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49102),
            .lcout(shift_srl_138Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92941),
            .ce(N__50038),
            .sr(_gnd_net_));
    defparam shift_srl_138_3_LC_2_22_3.C_ON=1'b0;
    defparam shift_srl_138_3_LC_2_22_3.SEQ_MODE=4'b1000;
    defparam shift_srl_138_3_LC_2_22_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_138_3_LC_2_22_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49096),
            .lcout(shift_srl_138Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92941),
            .ce(N__50038),
            .sr(_gnd_net_));
    defparam shift_srl_138_4_LC_2_22_4.C_ON=1'b0;
    defparam shift_srl_138_4_LC_2_22_4.SEQ_MODE=4'b1000;
    defparam shift_srl_138_4_LC_2_22_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_138_4_LC_2_22_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49090),
            .lcout(shift_srl_138Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92941),
            .ce(N__50038),
            .sr(_gnd_net_));
    defparam shift_srl_138_5_LC_2_22_5.C_ON=1'b0;
    defparam shift_srl_138_5_LC_2_22_5.SEQ_MODE=4'b1000;
    defparam shift_srl_138_5_LC_2_22_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_138_5_LC_2_22_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49084),
            .lcout(shift_srl_138Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92941),
            .ce(N__50038),
            .sr(_gnd_net_));
    defparam shift_srl_138_0_LC_2_22_6.C_ON=1'b0;
    defparam shift_srl_138_0_LC_2_22_6.SEQ_MODE=4'b1000;
    defparam shift_srl_138_0_LC_2_22_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_138_0_LC_2_22_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51324),
            .lcout(shift_srl_138Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92941),
            .ce(N__50038),
            .sr(_gnd_net_));
    defparam shift_srl_138_10_LC_2_22_7.C_ON=1'b0;
    defparam shift_srl_138_10_LC_2_22_7.SEQ_MODE=4'b1000;
    defparam shift_srl_138_10_LC_2_22_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_138_10_LC_2_22_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50092),
            .lcout(shift_srl_138Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92941),
            .ce(N__50038),
            .sr(_gnd_net_));
    defparam shift_srl_22_2_LC_3_7_1.C_ON=1'b0;
    defparam shift_srl_22_2_LC_3_7_1.SEQ_MODE=4'b1000;
    defparam shift_srl_22_2_LC_3_7_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_22_2_LC_3_7_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49066),
            .lcout(shift_srl_22Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93017),
            .ce(N__52202),
            .sr(_gnd_net_));
    defparam shift_srl_15_0_LC_3_9_0.C_ON=1'b0;
    defparam shift_srl_15_0_LC_3_9_0.SEQ_MODE=4'b1000;
    defparam shift_srl_15_0_LC_3_9_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_15_0_LC_3_9_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50546),
            .lcout(shift_srl_15Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92987),
            .ce(N__50118),
            .sr(_gnd_net_));
    defparam shift_srl_15_1_LC_3_9_1.C_ON=1'b0;
    defparam shift_srl_15_1_LC_3_9_1.SEQ_MODE=4'b1000;
    defparam shift_srl_15_1_LC_3_9_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_15_1_LC_3_9_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49054),
            .lcout(shift_srl_15Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92987),
            .ce(N__50118),
            .sr(_gnd_net_));
    defparam shift_srl_15_2_LC_3_9_2.C_ON=1'b0;
    defparam shift_srl_15_2_LC_3_9_2.SEQ_MODE=4'b1000;
    defparam shift_srl_15_2_LC_3_9_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_15_2_LC_3_9_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49150),
            .lcout(shift_srl_15Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92987),
            .ce(N__50118),
            .sr(_gnd_net_));
    defparam shift_srl_15_3_LC_3_9_3.C_ON=1'b0;
    defparam shift_srl_15_3_LC_3_9_3.SEQ_MODE=4'b1000;
    defparam shift_srl_15_3_LC_3_9_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_15_3_LC_3_9_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49144),
            .lcout(shift_srl_15Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92987),
            .ce(N__50118),
            .sr(_gnd_net_));
    defparam shift_srl_15_4_LC_3_9_4.C_ON=1'b0;
    defparam shift_srl_15_4_LC_3_9_4.SEQ_MODE=4'b1000;
    defparam shift_srl_15_4_LC_3_9_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_15_4_LC_3_9_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49138),
            .lcout(shift_srl_15Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92987),
            .ce(N__50118),
            .sr(_gnd_net_));
    defparam shift_srl_15_5_LC_3_9_5.C_ON=1'b0;
    defparam shift_srl_15_5_LC_3_9_5.SEQ_MODE=4'b1000;
    defparam shift_srl_15_5_LC_3_9_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_15_5_LC_3_9_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49132),
            .lcout(shift_srl_15Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92987),
            .ce(N__50118),
            .sr(_gnd_net_));
    defparam shift_srl_15_6_LC_3_9_6.C_ON=1'b0;
    defparam shift_srl_15_6_LC_3_9_6.SEQ_MODE=4'b1000;
    defparam shift_srl_15_6_LC_3_9_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_15_6_LC_3_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49126),
            .lcout(shift_srl_15Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92987),
            .ce(N__50118),
            .sr(_gnd_net_));
    defparam shift_srl_15_7_LC_3_9_7.C_ON=1'b0;
    defparam shift_srl_15_7_LC_3_9_7.SEQ_MODE=4'b1000;
    defparam shift_srl_15_7_LC_3_9_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_15_7_LC_3_9_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49120),
            .lcout(shift_srl_15Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92987),
            .ce(N__50118),
            .sr(_gnd_net_));
    defparam shift_srl_14_10_LC_3_10_0.C_ON=1'b0;
    defparam shift_srl_14_10_LC_3_10_0.SEQ_MODE=4'b1000;
    defparam shift_srl_14_10_LC_3_10_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_14_10_LC_3_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49186),
            .lcout(shift_srl_14Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92974),
            .ce(N__50202),
            .sr(_gnd_net_));
    defparam shift_srl_14_11_LC_3_10_1.C_ON=1'b0;
    defparam shift_srl_14_11_LC_3_10_1.SEQ_MODE=4'b1000;
    defparam shift_srl_14_11_LC_3_10_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_14_11_LC_3_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49114),
            .lcout(shift_srl_14Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92974),
            .ce(N__50202),
            .sr(_gnd_net_));
    defparam shift_srl_14_12_LC_3_10_2.C_ON=1'b0;
    defparam shift_srl_14_12_LC_3_10_2.SEQ_MODE=4'b1000;
    defparam shift_srl_14_12_LC_3_10_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_14_12_LC_3_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49108),
            .lcout(shift_srl_14Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92974),
            .ce(N__50202),
            .sr(_gnd_net_));
    defparam shift_srl_14_5_LC_3_10_3.C_ON=1'b0;
    defparam shift_srl_14_5_LC_3_10_3.SEQ_MODE=4'b1000;
    defparam shift_srl_14_5_LC_3_10_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_14_5_LC_3_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50227),
            .lcout(shift_srl_14Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92974),
            .ce(N__50202),
            .sr(_gnd_net_));
    defparam shift_srl_14_6_LC_3_10_4.C_ON=1'b0;
    defparam shift_srl_14_6_LC_3_10_4.SEQ_MODE=4'b1000;
    defparam shift_srl_14_6_LC_3_10_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_14_6_LC_3_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49198),
            .lcout(shift_srl_14Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92974),
            .ce(N__50202),
            .sr(_gnd_net_));
    defparam shift_srl_14_7_LC_3_10_5.C_ON=1'b0;
    defparam shift_srl_14_7_LC_3_10_5.SEQ_MODE=4'b1000;
    defparam shift_srl_14_7_LC_3_10_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_14_7_LC_3_10_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49192),
            .lcout(shift_srl_14Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92974),
            .ce(N__50202),
            .sr(_gnd_net_));
    defparam shift_srl_14_9_LC_3_10_6.C_ON=1'b0;
    defparam shift_srl_14_9_LC_3_10_6.SEQ_MODE=4'b1000;
    defparam shift_srl_14_9_LC_3_10_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_14_9_LC_3_10_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49174),
            .lcout(shift_srl_14Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92974),
            .ce(N__50202),
            .sr(_gnd_net_));
    defparam shift_srl_14_8_LC_3_10_7.C_ON=1'b0;
    defparam shift_srl_14_8_LC_3_10_7.SEQ_MODE=4'b1000;
    defparam shift_srl_14_8_LC_3_10_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_14_8_LC_3_10_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49180),
            .lcout(shift_srl_14Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92974),
            .ce(N__50202),
            .sr(_gnd_net_));
    defparam shift_srl_13_10_LC_3_11_0.C_ON=1'b0;
    defparam shift_srl_13_10_LC_3_11_0.SEQ_MODE=4'b1000;
    defparam shift_srl_13_10_LC_3_11_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_13_10_LC_3_11_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49237),
            .lcout(shift_srl_13Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92963),
            .ce(N__49568),
            .sr(_gnd_net_));
    defparam shift_srl_13_11_LC_3_11_1.C_ON=1'b0;
    defparam shift_srl_13_11_LC_3_11_1.SEQ_MODE=4'b1000;
    defparam shift_srl_13_11_LC_3_11_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_13_11_LC_3_11_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49168),
            .lcout(shift_srl_13Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92963),
            .ce(N__49568),
            .sr(_gnd_net_));
    defparam shift_srl_13_12_LC_3_11_2.C_ON=1'b0;
    defparam shift_srl_13_12_LC_3_11_2.SEQ_MODE=4'b1000;
    defparam shift_srl_13_12_LC_3_11_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_13_12_LC_3_11_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49162),
            .lcout(shift_srl_13Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92963),
            .ce(N__49568),
            .sr(_gnd_net_));
    defparam shift_srl_13_13_LC_3_11_3.C_ON=1'b0;
    defparam shift_srl_13_13_LC_3_11_3.SEQ_MODE=4'b1000;
    defparam shift_srl_13_13_LC_3_11_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_13_13_LC_3_11_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49156),
            .lcout(shift_srl_13Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92963),
            .ce(N__49568),
            .sr(_gnd_net_));
    defparam shift_srl_13_14_LC_3_11_4.C_ON=1'b0;
    defparam shift_srl_13_14_LC_3_11_4.SEQ_MODE=4'b1000;
    defparam shift_srl_13_14_LC_3_11_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_13_14_LC_3_11_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49249),
            .lcout(shift_srl_13Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92963),
            .ce(N__49568),
            .sr(_gnd_net_));
    defparam shift_srl_13_15_LC_3_11_5.C_ON=1'b0;
    defparam shift_srl_13_15_LC_3_11_5.SEQ_MODE=4'b1000;
    defparam shift_srl_13_15_LC_3_11_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_13_15_LC_3_11_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49243),
            .lcout(shift_srl_13Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92963),
            .ce(N__49568),
            .sr(_gnd_net_));
    defparam shift_srl_13_9_LC_3_11_6.C_ON=1'b0;
    defparam shift_srl_13_9_LC_3_11_6.SEQ_MODE=4'b1000;
    defparam shift_srl_13_9_LC_3_11_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_13_9_LC_3_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49222),
            .lcout(shift_srl_13Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92963),
            .ce(N__49568),
            .sr(_gnd_net_));
    defparam shift_srl_13_8_LC_3_11_7.C_ON=1'b0;
    defparam shift_srl_13_8_LC_3_11_7.SEQ_MODE=4'b1000;
    defparam shift_srl_13_8_LC_3_11_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_13_8_LC_3_11_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49231),
            .lcout(shift_srl_13Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92963),
            .ce(N__49568),
            .sr(_gnd_net_));
    defparam shift_srl_12_RNIV3PN3_15_LC_3_12_0.C_ON=1'b0;
    defparam shift_srl_12_RNIV3PN3_15_LC_3_12_0.SEQ_MODE=4'b0000;
    defparam shift_srl_12_RNIV3PN3_15_LC_3_12_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_12_RNIV3PN3_15_LC_3_12_0 (
            .in0(N__50366),
            .in1(N__50767),
            .in2(N__90579),
            .in3(N__50814),
            .lcout(clk_en_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_12_15_LC_3_12_1.C_ON=1'b0;
    defparam shift_srl_12_15_LC_3_12_1.SEQ_MODE=4'b1000;
    defparam shift_srl_12_15_LC_3_12_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_12_15_LC_3_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49216),
            .lcout(shift_srl_12Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92950),
            .ce(N__49399),
            .sr(_gnd_net_));
    defparam shift_srl_12_14_LC_3_12_2.C_ON=1'b0;
    defparam shift_srl_12_14_LC_3_12_2.SEQ_MODE=4'b1000;
    defparam shift_srl_12_14_LC_3_12_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_12_14_LC_3_12_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49210),
            .lcout(shift_srl_12Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92950),
            .ce(N__49399),
            .sr(_gnd_net_));
    defparam shift_srl_12_13_LC_3_12_3.C_ON=1'b0;
    defparam shift_srl_12_13_LC_3_12_3.SEQ_MODE=4'b1000;
    defparam shift_srl_12_13_LC_3_12_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_12_13_LC_3_12_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49204),
            .lcout(shift_srl_12Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92950),
            .ce(N__49399),
            .sr(_gnd_net_));
    defparam shift_srl_12_12_LC_3_12_4.C_ON=1'b0;
    defparam shift_srl_12_12_LC_3_12_4.SEQ_MODE=4'b1000;
    defparam shift_srl_12_12_LC_3_12_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_12_12_LC_3_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49426),
            .lcout(shift_srl_12Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92950),
            .ce(N__49399),
            .sr(_gnd_net_));
    defparam shift_srl_12_11_LC_3_12_5.C_ON=1'b0;
    defparam shift_srl_12_11_LC_3_12_5.SEQ_MODE=4'b1000;
    defparam shift_srl_12_11_LC_3_12_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_12_11_LC_3_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49420),
            .lcout(shift_srl_12Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92950),
            .ce(N__49399),
            .sr(_gnd_net_));
    defparam shift_srl_12_10_LC_3_12_6.C_ON=1'b0;
    defparam shift_srl_12_10_LC_3_12_6.SEQ_MODE=4'b1000;
    defparam shift_srl_12_10_LC_3_12_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_12_10_LC_3_12_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49405),
            .lcout(shift_srl_12Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92950),
            .ce(N__49399),
            .sr(_gnd_net_));
    defparam shift_srl_12_9_LC_3_12_7.C_ON=1'b0;
    defparam shift_srl_12_9_LC_3_12_7.SEQ_MODE=4'b1000;
    defparam shift_srl_12_9_LC_3_12_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_12_9_LC_3_12_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49414),
            .lcout(shift_srl_12Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92950),
            .ce(N__49399),
            .sr(_gnd_net_));
    defparam shift_srl_15_RNI07RB4_15_LC_3_13_0.C_ON=1'b0;
    defparam shift_srl_15_RNI07RB4_15_LC_3_13_0.SEQ_MODE=4'b0000;
    defparam shift_srl_15_RNI07RB4_15_LC_3_13_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_15_RNI07RB4_15_LC_3_13_0 (
            .in0(N__50557),
            .in1(N__90404),
            .in2(N__49272),
            .in3(N__50508),
            .lcout(clk_en_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_6_RNI00BH_15_LC_3_13_1.C_ON=1'b0;
    defparam shift_srl_6_RNI00BH_15_LC_3_13_1.SEQ_MODE=4'b0000;
    defparam shift_srl_6_RNI00BH_15_LC_3_13_1.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_6_RNI00BH_15_LC_3_13_1 (
            .in0(N__49369),
            .in1(N__49345),
            .in2(_gnd_net_),
            .in3(N__49304),
            .lcout(shift_srl_6_RNI00BHZ0Z_15),
            .ltout(shift_srl_6_RNI00BHZ0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_7_RNI00TC1_15_LC_3_13_2.C_ON=1'b0;
    defparam shift_srl_7_RNI00TC1_15_LC_3_13_2.SEQ_MODE=4'b0000;
    defparam shift_srl_7_RNI00TC1_15_LC_3_13_2.LUT_INIT=16'b1010000000000000;
    LogicCell40 shift_srl_7_RNI00TC1_15_LC_3_13_2 (
            .in0(N__49477),
            .in1(_gnd_net_),
            .in2(N__49282),
            .in3(N__53761),
            .lcout(shift_srl_7_RNI00TC1Z0Z_15),
            .ltout(shift_srl_7_RNI00TC1Z0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_11_RNI4OUM3_15_LC_3_13_3.C_ON=1'b0;
    defparam shift_srl_11_RNI4OUM3_15_LC_3_13_3.SEQ_MODE=4'b0000;
    defparam shift_srl_11_RNI4OUM3_15_LC_3_13_3.LUT_INIT=16'b0000000000100000;
    LogicCell40 shift_srl_11_RNI4OUM3_15_LC_3_13_3 (
            .in0(N__53803),
            .in1(N__50731),
            .in2(N__49279),
            .in3(N__53703),
            .lcout(rco_c_13),
            .ltout(rco_c_13_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_15_RNIN2BJ4_15_LC_3_13_4.C_ON=1'b0;
    defparam shift_srl_15_RNIN2BJ4_15_LC_3_13_4.SEQ_MODE=4'b0000;
    defparam shift_srl_15_RNIN2BJ4_15_LC_3_13_4.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_15_RNIN2BJ4_15_LC_3_13_4 (
            .in0(N__50556),
            .in1(N__50507),
            .in2(N__49255),
            .in3(N__50428),
            .lcout(rco_c_16),
            .ltout(rco_c_16_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_18_RNIP9C15_15_LC_3_13_5.C_ON=1'b0;
    defparam shift_srl_18_RNIP9C15_15_LC_3_13_5.SEQ_MODE=4'b0000;
    defparam shift_srl_18_RNIP9C15_15_LC_3_13_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_18_RNIP9C15_15_LC_3_13_5 (
            .in0(N__90405),
            .in1(N__52440),
            .in2(N__49252),
            .in3(N__50695),
            .lcout(clk_en_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_19_LC_3_13_6.C_ON=1'b0;
    defparam rco_obuf_RNO_19_LC_3_13_6.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_19_LC_3_13_6.LUT_INIT=16'b1000000000000000;
    LogicCell40 rco_obuf_RNO_19_LC_3_13_6 (
            .in0(N__49596),
            .in1(N__52560),
            .in2(N__50710),
            .in3(N__52438),
            .lcout(rco_c_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_11_RNI75L33_15_LC_3_13_7.C_ON=1'b0;
    defparam shift_srl_11_RNI75L33_15_LC_3_13_7.SEQ_MODE=4'b0000;
    defparam shift_srl_11_RNI75L33_15_LC_3_13_7.LUT_INIT=16'b0000000000001000;
    LogicCell40 shift_srl_11_RNI75L33_15_LC_3_13_7 (
            .in0(N__53802),
            .in1(N__49488),
            .in2(N__49504),
            .in3(N__53702),
            .lcout(rco_c_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_11_RNILS6B3_15_LC_3_14_0.C_ON=1'b0;
    defparam shift_srl_11_RNILS6B3_15_LC_3_14_0.SEQ_MODE=4'b0000;
    defparam shift_srl_11_RNILS6B3_15_LC_3_14_0.LUT_INIT=16'b0000000000100000;
    LogicCell40 shift_srl_11_RNILS6B3_15_LC_3_14_0 (
            .in0(N__53804),
            .in1(N__53723),
            .in2(N__53644),
            .in3(N__49534),
            .lcout(rco_c_12),
            .ltout(rco_c_12_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIG81C3_15_LC_3_14_1.C_ON=1'b0;
    defparam shift_srl_0_RNIG81C3_15_LC_3_14_1.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIG81C3_15_LC_3_14_1.LUT_INIT=16'b1111000000000000;
    LogicCell40 shift_srl_0_RNIG81C3_15_LC_3_14_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__49576),
            .in3(N__90461),
            .lcout(clk_en_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_11_RNI92881_15_LC_3_14_2.C_ON=1'b0;
    defparam shift_srl_11_RNI92881_15_LC_3_14_2.SEQ_MODE=4'b0000;
    defparam shift_srl_11_RNI92881_15_LC_3_14_2.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_11_RNI92881_15_LC_3_14_2 (
            .in0(N__51371),
            .in1(N__55724),
            .in2(N__53766),
            .in3(N__50818),
            .lcout(rco_int_0_a2_sx_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_13_RNIF3N74_15_LC_3_14_3.C_ON=1'b0;
    defparam shift_srl_13_RNIF3N74_15_LC_3_14_3.SEQ_MODE=4'b0000;
    defparam shift_srl_13_RNIF3N74_15_LC_3_14_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_13_RNIF3N74_15_LC_3_14_3 (
            .in0(N__50777),
            .in1(N__90462),
            .in2(N__49521),
            .in3(N__50509),
            .lcout(clk_en_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_7_15_LC_3_14_4.C_ON=1'b0;
    defparam shift_srl_7_15_LC_3_14_4.SEQ_MODE=4'b1000;
    defparam shift_srl_7_15_LC_3_14_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_7_15_LC_3_14_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49711),
            .lcout(shift_srl_7Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92933),
            .ce(N__49677),
            .sr(_gnd_net_));
    defparam shift_srl_11_RNIP23E1_15_LC_3_14_5.C_ON=1'b0;
    defparam shift_srl_11_RNIP23E1_15_LC_3_14_5.SEQ_MODE=4'b0000;
    defparam shift_srl_11_RNIP23E1_15_LC_3_14_5.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_11_RNIP23E1_15_LC_3_14_5 (
            .in0(N__49475),
            .in1(N__53756),
            .in2(N__55730),
            .in3(N__51370),
            .lcout(rco_int_0_a2_sx_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_7_RNI76782_15_LC_3_14_6.C_ON=1'b0;
    defparam shift_srl_7_RNI76782_15_LC_3_14_6.SEQ_MODE=4'b0000;
    defparam shift_srl_7_RNI76782_15_LC_3_14_6.LUT_INIT=16'b0010000000000000;
    LogicCell40 shift_srl_7_RNI76782_15_LC_3_14_6 (
            .in0(N__53760),
            .in1(N__53722),
            .in2(N__49492),
            .in3(N__49476),
            .lcout(rco_c_7),
            .ltout(rco_c_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_8_RNIAIIA2_15_LC_3_14_7.C_ON=1'b0;
    defparam shift_srl_8_RNIAIIA2_15_LC_3_14_7.SEQ_MODE=4'b0000;
    defparam shift_srl_8_RNIAIIA2_15_LC_3_14_7.LUT_INIT=16'b1111000000000000;
    LogicCell40 shift_srl_8_RNIAIIA2_15_LC_3_14_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__49648),
            .in3(N__53830),
            .lcout(rco_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_21_10_LC_3_15_0.C_ON=1'b0;
    defparam shift_srl_21_10_LC_3_15_0.SEQ_MODE=4'b1000;
    defparam shift_srl_21_10_LC_3_15_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_21_10_LC_3_15_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49615),
            .lcout(shift_srl_21Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92925),
            .ce(N__50920),
            .sr(_gnd_net_));
    defparam shift_srl_21_11_LC_3_15_1.C_ON=1'b0;
    defparam shift_srl_21_11_LC_3_15_1.SEQ_MODE=4'b1000;
    defparam shift_srl_21_11_LC_3_15_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_21_11_LC_3_15_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49645),
            .lcout(shift_srl_21Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92925),
            .ce(N__50920),
            .sr(_gnd_net_));
    defparam shift_srl_21_12_LC_3_15_2.C_ON=1'b0;
    defparam shift_srl_21_12_LC_3_15_2.SEQ_MODE=4'b1000;
    defparam shift_srl_21_12_LC_3_15_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_21_12_LC_3_15_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49639),
            .lcout(shift_srl_21Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92925),
            .ce(N__50920),
            .sr(_gnd_net_));
    defparam shift_srl_21_13_LC_3_15_3.C_ON=1'b0;
    defparam shift_srl_21_13_LC_3_15_3.SEQ_MODE=4'b1000;
    defparam shift_srl_21_13_LC_3_15_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_21_13_LC_3_15_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49633),
            .lcout(shift_srl_21Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92925),
            .ce(N__50920),
            .sr(_gnd_net_));
    defparam shift_srl_21_14_LC_3_15_4.C_ON=1'b0;
    defparam shift_srl_21_14_LC_3_15_4.SEQ_MODE=4'b1000;
    defparam shift_srl_21_14_LC_3_15_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_21_14_LC_3_15_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49627),
            .lcout(shift_srl_21Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92925),
            .ce(N__50920),
            .sr(_gnd_net_));
    defparam shift_srl_21_15_LC_3_15_5.C_ON=1'b0;
    defparam shift_srl_21_15_LC_3_15_5.SEQ_MODE=4'b1000;
    defparam shift_srl_21_15_LC_3_15_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_21_15_LC_3_15_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49621),
            .lcout(shift_srl_21Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92925),
            .ce(N__50920),
            .sr(_gnd_net_));
    defparam shift_srl_21_9_LC_3_15_6.C_ON=1'b0;
    defparam shift_srl_21_9_LC_3_15_6.SEQ_MODE=4'b1000;
    defparam shift_srl_21_9_LC_3_15_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_21_9_LC_3_15_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49609),
            .lcout(shift_srl_21Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92925),
            .ce(N__50920),
            .sr(_gnd_net_));
    defparam shift_srl_21_8_LC_3_15_7.C_ON=1'b0;
    defparam shift_srl_21_8_LC_3_15_7.SEQ_MODE=4'b1000;
    defparam shift_srl_21_8_LC_3_15_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_21_8_LC_3_15_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50926),
            .lcout(shift_srl_21Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92925),
            .ce(N__50920),
            .sr(_gnd_net_));
    defparam shift_srl_7_10_LC_3_16_0.C_ON=1'b0;
    defparam shift_srl_7_10_LC_3_16_0.SEQ_MODE=4'b1000;
    defparam shift_srl_7_10_LC_3_16_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_7_10_LC_3_16_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49702),
            .lcout(shift_srl_7Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92919),
            .ce(N__49678),
            .sr(_gnd_net_));
    defparam shift_srl_7_11_LC_3_16_1.C_ON=1'b0;
    defparam shift_srl_7_11_LC_3_16_1.SEQ_MODE=4'b1000;
    defparam shift_srl_7_11_LC_3_16_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_7_11_LC_3_16_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49735),
            .lcout(shift_srl_7Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92919),
            .ce(N__49678),
            .sr(_gnd_net_));
    defparam shift_srl_7_12_LC_3_16_2.C_ON=1'b0;
    defparam shift_srl_7_12_LC_3_16_2.SEQ_MODE=4'b1000;
    defparam shift_srl_7_12_LC_3_16_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_7_12_LC_3_16_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49729),
            .lcout(shift_srl_7Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92919),
            .ce(N__49678),
            .sr(_gnd_net_));
    defparam shift_srl_7_13_LC_3_16_3.C_ON=1'b0;
    defparam shift_srl_7_13_LC_3_16_3.SEQ_MODE=4'b1000;
    defparam shift_srl_7_13_LC_3_16_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_7_13_LC_3_16_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49723),
            .lcout(shift_srl_7Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92919),
            .ce(N__49678),
            .sr(_gnd_net_));
    defparam shift_srl_7_14_LC_3_16_4.C_ON=1'b0;
    defparam shift_srl_7_14_LC_3_16_4.SEQ_MODE=4'b1000;
    defparam shift_srl_7_14_LC_3_16_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_7_14_LC_3_16_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49717),
            .lcout(shift_srl_7Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92919),
            .ce(N__49678),
            .sr(_gnd_net_));
    defparam shift_srl_7_9_LC_3_16_5.C_ON=1'b0;
    defparam shift_srl_7_9_LC_3_16_5.SEQ_MODE=4'b1000;
    defparam shift_srl_7_9_LC_3_16_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_7_9_LC_3_16_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49696),
            .lcout(shift_srl_7Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92919),
            .ce(N__49678),
            .sr(_gnd_net_));
    defparam shift_srl_7_8_LC_3_16_6.C_ON=1'b0;
    defparam shift_srl_7_8_LC_3_16_6.SEQ_MODE=4'b1000;
    defparam shift_srl_7_8_LC_3_16_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_7_8_LC_3_16_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49684),
            .lcout(shift_srl_7Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92919),
            .ce(N__49678),
            .sr(_gnd_net_));
    defparam shift_srl_7_7_LC_3_16_7.C_ON=1'b0;
    defparam shift_srl_7_7_LC_3_16_7.SEQ_MODE=4'b1000;
    defparam shift_srl_7_7_LC_3_16_7.LUT_INIT=16'b1100110011001100;
    LogicCell40 shift_srl_7_7_LC_3_16_7 (
            .in0(_gnd_net_),
            .in1(N__49690),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_7Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92919),
            .ce(N__49678),
            .sr(_gnd_net_));
    defparam shift_srl_18_10_LC_3_17_0.C_ON=1'b0;
    defparam shift_srl_18_10_LC_3_17_0.SEQ_MODE=4'b1000;
    defparam shift_srl_18_10_LC_3_17_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_18_10_LC_3_17_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49759),
            .lcout(shift_srl_18Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92910),
            .ce(N__50854),
            .sr(_gnd_net_));
    defparam shift_srl_18_11_LC_3_17_1.C_ON=1'b0;
    defparam shift_srl_18_11_LC_3_17_1.SEQ_MODE=4'b1000;
    defparam shift_srl_18_11_LC_3_17_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_18_11_LC_3_17_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49654),
            .lcout(shift_srl_18Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92910),
            .ce(N__50854),
            .sr(_gnd_net_));
    defparam shift_srl_18_12_LC_3_17_2.C_ON=1'b0;
    defparam shift_srl_18_12_LC_3_17_2.SEQ_MODE=4'b1000;
    defparam shift_srl_18_12_LC_3_17_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_18_12_LC_3_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49783),
            .lcout(shift_srl_18Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92910),
            .ce(N__50854),
            .sr(_gnd_net_));
    defparam shift_srl_18_13_LC_3_17_3.C_ON=1'b0;
    defparam shift_srl_18_13_LC_3_17_3.SEQ_MODE=4'b1000;
    defparam shift_srl_18_13_LC_3_17_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_18_13_LC_3_17_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49777),
            .lcout(shift_srl_18Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92910),
            .ce(N__50854),
            .sr(_gnd_net_));
    defparam shift_srl_18_14_LC_3_17_4.C_ON=1'b0;
    defparam shift_srl_18_14_LC_3_17_4.SEQ_MODE=4'b1000;
    defparam shift_srl_18_14_LC_3_17_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_18_14_LC_3_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49771),
            .lcout(shift_srl_18Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92910),
            .ce(N__50854),
            .sr(_gnd_net_));
    defparam shift_srl_18_15_LC_3_17_5.C_ON=1'b0;
    defparam shift_srl_18_15_LC_3_17_5.SEQ_MODE=4'b1000;
    defparam shift_srl_18_15_LC_3_17_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_18_15_LC_3_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49765),
            .lcout(shift_srl_18Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92910),
            .ce(N__50854),
            .sr(_gnd_net_));
    defparam shift_srl_18_9_LC_3_17_6.C_ON=1'b0;
    defparam shift_srl_18_9_LC_3_17_6.SEQ_MODE=4'b1000;
    defparam shift_srl_18_9_LC_3_17_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_18_9_LC_3_17_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49753),
            .lcout(shift_srl_18Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92910),
            .ce(N__50854),
            .sr(_gnd_net_));
    defparam shift_srl_18_8_LC_3_17_7.C_ON=1'b0;
    defparam shift_srl_18_8_LC_3_17_7.SEQ_MODE=4'b1000;
    defparam shift_srl_18_8_LC_3_17_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_18_8_LC_3_17_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50860),
            .lcout(shift_srl_18Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92910),
            .ce(N__50854),
            .sr(_gnd_net_));
    defparam shift_srl_129_0_LC_3_18_0.C_ON=1'b0;
    defparam shift_srl_129_0_LC_3_18_0.SEQ_MODE=4'b1000;
    defparam shift_srl_129_0_LC_3_18_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_129_0_LC_3_18_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54235),
            .lcout(shift_srl_129Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92920),
            .ce(N__53987),
            .sr(_gnd_net_));
    defparam shift_srl_129_1_LC_3_18_1.C_ON=1'b0;
    defparam shift_srl_129_1_LC_3_18_1.SEQ_MODE=4'b1000;
    defparam shift_srl_129_1_LC_3_18_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_129_1_LC_3_18_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49747),
            .lcout(shift_srl_129Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92920),
            .ce(N__53987),
            .sr(_gnd_net_));
    defparam shift_srl_129_2_LC_3_18_2.C_ON=1'b0;
    defparam shift_srl_129_2_LC_3_18_2.SEQ_MODE=4'b1000;
    defparam shift_srl_129_2_LC_3_18_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_129_2_LC_3_18_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49741),
            .lcout(shift_srl_129Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92920),
            .ce(N__53987),
            .sr(_gnd_net_));
    defparam shift_srl_129_3_LC_3_18_3.C_ON=1'b0;
    defparam shift_srl_129_3_LC_3_18_3.SEQ_MODE=4'b1000;
    defparam shift_srl_129_3_LC_3_18_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_129_3_LC_3_18_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49831),
            .lcout(shift_srl_129Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92920),
            .ce(N__53987),
            .sr(_gnd_net_));
    defparam shift_srl_129_4_LC_3_18_4.C_ON=1'b0;
    defparam shift_srl_129_4_LC_3_18_4.SEQ_MODE=4'b1000;
    defparam shift_srl_129_4_LC_3_18_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_129_4_LC_3_18_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49825),
            .lcout(shift_srl_129Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92920),
            .ce(N__53987),
            .sr(_gnd_net_));
    defparam shift_srl_129_5_LC_3_18_5.C_ON=1'b0;
    defparam shift_srl_129_5_LC_3_18_5.SEQ_MODE=4'b1000;
    defparam shift_srl_129_5_LC_3_18_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_129_5_LC_3_18_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49819),
            .lcout(shift_srl_129Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92920),
            .ce(N__53987),
            .sr(_gnd_net_));
    defparam shift_srl_129_6_LC_3_18_6.C_ON=1'b0;
    defparam shift_srl_129_6_LC_3_18_6.SEQ_MODE=4'b1000;
    defparam shift_srl_129_6_LC_3_18_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_129_6_LC_3_18_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49813),
            .lcout(shift_srl_129Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92920),
            .ce(N__53987),
            .sr(_gnd_net_));
    defparam shift_srl_129_7_LC_3_18_7.C_ON=1'b0;
    defparam shift_srl_129_7_LC_3_18_7.SEQ_MODE=4'b1000;
    defparam shift_srl_129_7_LC_3_18_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_129_7_LC_3_18_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49807),
            .lcout(shift_srl_129Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92920),
            .ce(N__53987),
            .sr(_gnd_net_));
    defparam shift_srl_132_RNI4MAQ_15_LC_3_19_0.C_ON=1'b0;
    defparam shift_srl_132_RNI4MAQ_15_LC_3_19_0.SEQ_MODE=4'b0000;
    defparam shift_srl_132_RNI4MAQ_15_LC_3_19_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_132_RNI4MAQ_15_LC_3_19_0 (
            .in0(N__54369),
            .in1(N__54308),
            .in2(N__66462),
            .in3(N__52913),
            .lcout(g0_8_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_130_15_LC_3_19_1.C_ON=1'b0;
    defparam shift_srl_130_15_LC_3_19_1.SEQ_MODE=4'b1000;
    defparam shift_srl_130_15_LC_3_19_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_130_15_LC_3_19_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49789),
            .lcout(shift_srl_130Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92926),
            .ce(N__49881),
            .sr(_gnd_net_));
    defparam shift_srl_130_RNIQP2E_15_LC_3_19_2.C_ON=1'b0;
    defparam shift_srl_130_RNIQP2E_15_LC_3_19_2.SEQ_MODE=4'b0000;
    defparam shift_srl_130_RNIQP2E_15_LC_3_19_2.LUT_INIT=16'b1100110000000000;
    LogicCell40 shift_srl_130_RNIQP2E_15_LC_3_19_2 (
            .in0(_gnd_net_),
            .in1(N__90413),
            .in2(_gnd_net_),
            .in3(N__52912),
            .lcout(g0_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_130_14_LC_3_19_3.C_ON=1'b0;
    defparam shift_srl_130_14_LC_3_19_3.SEQ_MODE=4'b1000;
    defparam shift_srl_130_14_LC_3_19_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_130_14_LC_3_19_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49918),
            .lcout(shift_srl_130Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92926),
            .ce(N__49881),
            .sr(_gnd_net_));
    defparam shift_srl_130_13_LC_3_19_4.C_ON=1'b0;
    defparam shift_srl_130_13_LC_3_19_4.SEQ_MODE=4'b1000;
    defparam shift_srl_130_13_LC_3_19_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_130_13_LC_3_19_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49912),
            .lcout(shift_srl_130Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92926),
            .ce(N__49881),
            .sr(_gnd_net_));
    defparam shift_srl_130_12_LC_3_19_5.C_ON=1'b0;
    defparam shift_srl_130_12_LC_3_19_5.SEQ_MODE=4'b1000;
    defparam shift_srl_130_12_LC_3_19_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_130_12_LC_3_19_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49906),
            .lcout(shift_srl_130Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92926),
            .ce(N__49881),
            .sr(_gnd_net_));
    defparam shift_srl_130_11_LC_3_19_6.C_ON=1'b0;
    defparam shift_srl_130_11_LC_3_19_6.SEQ_MODE=4'b1000;
    defparam shift_srl_130_11_LC_3_19_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_130_11_LC_3_19_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49888),
            .lcout(shift_srl_130Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92926),
            .ce(N__49881),
            .sr(_gnd_net_));
    defparam shift_srl_130_10_LC_3_19_7.C_ON=1'b0;
    defparam shift_srl_130_10_LC_3_19_7.SEQ_MODE=4'b1000;
    defparam shift_srl_130_10_LC_3_19_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_130_10_LC_3_19_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49900),
            .lcout(shift_srl_130Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92926),
            .ce(N__49881),
            .sr(_gnd_net_));
    defparam shift_srl_137_10_LC_3_20_0.C_ON=1'b0;
    defparam shift_srl_137_10_LC_3_20_0.SEQ_MODE=4'b1000;
    defparam shift_srl_137_10_LC_3_20_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_137_10_LC_3_20_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50014),
            .lcout(shift_srl_137Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92934),
            .ce(N__49990),
            .sr(_gnd_net_));
    defparam shift_srl_137_11_LC_3_20_1.C_ON=1'b0;
    defparam shift_srl_137_11_LC_3_20_1.SEQ_MODE=4'b1000;
    defparam shift_srl_137_11_LC_3_20_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_137_11_LC_3_20_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49855),
            .lcout(shift_srl_137Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92934),
            .ce(N__49990),
            .sr(_gnd_net_));
    defparam shift_srl_137_12_LC_3_20_2.C_ON=1'b0;
    defparam shift_srl_137_12_LC_3_20_2.SEQ_MODE=4'b1000;
    defparam shift_srl_137_12_LC_3_20_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_137_12_LC_3_20_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49849),
            .lcout(shift_srl_137Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92934),
            .ce(N__49990),
            .sr(_gnd_net_));
    defparam shift_srl_137_13_LC_3_20_3.C_ON=1'b0;
    defparam shift_srl_137_13_LC_3_20_3.SEQ_MODE=4'b1000;
    defparam shift_srl_137_13_LC_3_20_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_137_13_LC_3_20_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49843),
            .lcout(shift_srl_137Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92934),
            .ce(N__49990),
            .sr(_gnd_net_));
    defparam shift_srl_137_14_LC_3_20_4.C_ON=1'b0;
    defparam shift_srl_137_14_LC_3_20_4.SEQ_MODE=4'b1000;
    defparam shift_srl_137_14_LC_3_20_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_137_14_LC_3_20_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49837),
            .lcout(shift_srl_137Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92934),
            .ce(N__49990),
            .sr(_gnd_net_));
    defparam shift_srl_137_15_LC_3_20_5.C_ON=1'b0;
    defparam shift_srl_137_15_LC_3_20_5.SEQ_MODE=4'b1000;
    defparam shift_srl_137_15_LC_3_20_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_137_15_LC_3_20_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50020),
            .lcout(shift_srl_137Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92934),
            .ce(N__49990),
            .sr(_gnd_net_));
    defparam shift_srl_137_9_LC_3_20_6.C_ON=1'b0;
    defparam shift_srl_137_9_LC_3_20_6.SEQ_MODE=4'b1000;
    defparam shift_srl_137_9_LC_3_20_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_137_9_LC_3_20_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49996),
            .lcout(shift_srl_137Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92934),
            .ce(N__49990),
            .sr(_gnd_net_));
    defparam shift_srl_137_8_LC_3_20_7.C_ON=1'b0;
    defparam shift_srl_137_8_LC_3_20_7.SEQ_MODE=4'b1000;
    defparam shift_srl_137_8_LC_3_20_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_137_8_LC_3_20_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50008),
            .lcout(shift_srl_137Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92934),
            .ce(N__49990),
            .sr(_gnd_net_));
    defparam shift_srl_132_RNI1837_15_LC_3_21_0.C_ON=1'b0;
    defparam shift_srl_132_RNI1837_15_LC_3_21_0.SEQ_MODE=4'b0000;
    defparam shift_srl_132_RNI1837_15_LC_3_21_0.LUT_INIT=16'b1100110000000000;
    LogicCell40 shift_srl_132_RNI1837_15_LC_3_21_0 (
            .in0(_gnd_net_),
            .in1(N__54365),
            .in2(_gnd_net_),
            .in3(N__54309),
            .lcout(),
            .ltout(g0_4_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_116_RNIKQMQ1_15_LC_3_21_1.C_ON=1'b0;
    defparam shift_srl_116_RNIKQMQ1_15_LC_3_21_1.SEQ_MODE=4'b0000;
    defparam shift_srl_116_RNIKQMQ1_15_LC_3_21_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_116_RNIKQMQ1_15_LC_3_21_1 (
            .in0(N__51100),
            .in1(N__58800),
            .in2(N__49969),
            .in3(N__63818),
            .lcout(g0_15_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_120_RNIID991_15_LC_3_21_2.C_ON=1'b0;
    defparam shift_srl_120_RNIID991_15_LC_3_21_2.SEQ_MODE=4'b0000;
    defparam shift_srl_120_RNIID991_15_LC_3_21_2.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_120_RNIID991_15_LC_3_21_2 (
            .in0(N__65752),
            .in1(N__65614),
            .in2(_gnd_net_),
            .in3(N__65866),
            .lcout(),
            .ltout(g0_13_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_135_RNIP0HR2_15_LC_3_21_3.C_ON=1'b0;
    defparam shift_srl_135_RNIP0HR2_15_LC_3_21_3.SEQ_MODE=4'b0000;
    defparam shift_srl_135_RNIP0HR2_15_LC_3_21_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_135_RNIP0HR2_15_LC_3_21_3 (
            .in0(N__53104),
            .in1(N__52015),
            .in2(N__49966),
            .in3(N__65364),
            .lcout(),
            .ltout(g0_16_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_116_RNI1C0621_15_LC_3_21_4.C_ON=1'b0;
    defparam shift_srl_116_RNI1C0621_15_LC_3_21_4.SEQ_MODE=4'b0000;
    defparam shift_srl_116_RNI1C0621_15_LC_3_21_4.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_116_RNI1C0621_15_LC_3_21_4 (
            .in0(N__49963),
            .in1(N__56473),
            .in2(N__49957),
            .in3(N__62004),
            .lcout(clk_en_136),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_132_RNIAGTV_15_LC_3_21_5.C_ON=1'b0;
    defparam shift_srl_132_RNIAGTV_15_LC_3_21_5.SEQ_MODE=4'b0000;
    defparam shift_srl_132_RNIAGTV_15_LC_3_21_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_132_RNIAGTV_15_LC_3_21_5 (
            .in0(N__54310),
            .in1(N__90518),
            .in2(N__54370),
            .in3(N__65753),
            .lcout(),
            .ltout(g0_8_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_132_RNICS0N21_15_LC_3_21_6.C_ON=1'b0;
    defparam shift_srl_132_RNICS0N21_15_LC_3_21_6.SEQ_MODE=4'b0000;
    defparam shift_srl_132_RNICS0N21_15_LC_3_21_6.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_132_RNICS0N21_15_LC_3_21_6 (
            .in0(N__51244),
            .in1(N__51094),
            .in2(N__50095),
            .in3(N__57612),
            .lcout(clk_en_138),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_138_9_LC_3_22_0.C_ON=1'b0;
    defparam shift_srl_138_9_LC_3_22_0.SEQ_MODE=4'b1000;
    defparam shift_srl_138_9_LC_3_22_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_138_9_LC_3_22_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50044),
            .lcout(shift_srl_138Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92951),
            .ce(N__50037),
            .sr(_gnd_net_));
    defparam shift_srl_138_12_LC_3_22_1.C_ON=1'b0;
    defparam shift_srl_138_12_LC_3_22_1.SEQ_MODE=4'b1000;
    defparam shift_srl_138_12_LC_3_22_1.LUT_INIT=16'b1100110011001100;
    LogicCell40 shift_srl_138_12_LC_3_22_1 (
            .in0(_gnd_net_),
            .in1(N__50086),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_138Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92951),
            .ce(N__50037),
            .sr(_gnd_net_));
    defparam shift_srl_138_7_LC_3_22_2.C_ON=1'b0;
    defparam shift_srl_138_7_LC_3_22_2.SEQ_MODE=4'b1000;
    defparam shift_srl_138_7_LC_3_22_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_138_7_LC_3_22_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50056),
            .lcout(shift_srl_138Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92951),
            .ce(N__50037),
            .sr(_gnd_net_));
    defparam shift_srl_138_13_LC_3_22_3.C_ON=1'b0;
    defparam shift_srl_138_13_LC_3_22_3.SEQ_MODE=4'b1000;
    defparam shift_srl_138_13_LC_3_22_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_138_13_LC_3_22_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50080),
            .lcout(shift_srl_138Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92951),
            .ce(N__50037),
            .sr(_gnd_net_));
    defparam shift_srl_138_14_LC_3_22_4.C_ON=1'b0;
    defparam shift_srl_138_14_LC_3_22_4.SEQ_MODE=4'b1000;
    defparam shift_srl_138_14_LC_3_22_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_138_14_LC_3_22_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50074),
            .lcout(shift_srl_138Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92951),
            .ce(N__50037),
            .sr(_gnd_net_));
    defparam shift_srl_138_15_LC_3_22_5.C_ON=1'b0;
    defparam shift_srl_138_15_LC_3_22_5.SEQ_MODE=4'b1000;
    defparam shift_srl_138_15_LC_3_22_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_138_15_LC_3_22_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50068),
            .lcout(shift_srl_138Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92951),
            .ce(N__50037),
            .sr(_gnd_net_));
    defparam shift_srl_138_6_LC_3_22_6.C_ON=1'b0;
    defparam shift_srl_138_6_LC_3_22_6.SEQ_MODE=4'b1000;
    defparam shift_srl_138_6_LC_3_22_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_138_6_LC_3_22_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50062),
            .lcout(shift_srl_138Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92951),
            .ce(N__50037),
            .sr(_gnd_net_));
    defparam shift_srl_138_8_LC_3_22_7.C_ON=1'b0;
    defparam shift_srl_138_8_LC_3_22_7.SEQ_MODE=4'b1000;
    defparam shift_srl_138_8_LC_3_22_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_138_8_LC_3_22_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50050),
            .lcout(shift_srl_138Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92951),
            .ce(N__50037),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_124_LC_3_24_5.C_ON=1'b0;
    defparam rco_obuf_RNO_124_LC_3_24_5.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_124_LC_3_24_5.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_124_LC_3_24_5 (
            .in0(N__65458),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57624),
            .lcout(rco_c_124),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_15_10_LC_4_9_0.C_ON=1'b0;
    defparam shift_srl_15_10_LC_4_9_0.SEQ_MODE=4'b1000;
    defparam shift_srl_15_10_LC_4_9_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_15_10_LC_4_9_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50137),
            .lcout(shift_srl_15Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93002),
            .ce(N__50119),
            .sr(_gnd_net_));
    defparam shift_srl_15_11_LC_4_9_1.C_ON=1'b0;
    defparam shift_srl_15_11_LC_4_9_1.SEQ_MODE=4'b1000;
    defparam shift_srl_15_11_LC_4_9_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_15_11_LC_4_9_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50167),
            .lcout(shift_srl_15Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93002),
            .ce(N__50119),
            .sr(_gnd_net_));
    defparam shift_srl_15_12_LC_4_9_2.C_ON=1'b0;
    defparam shift_srl_15_12_LC_4_9_2.SEQ_MODE=4'b1000;
    defparam shift_srl_15_12_LC_4_9_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_15_12_LC_4_9_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50161),
            .lcout(shift_srl_15Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93002),
            .ce(N__50119),
            .sr(_gnd_net_));
    defparam shift_srl_15_13_LC_4_9_3.C_ON=1'b0;
    defparam shift_srl_15_13_LC_4_9_3.SEQ_MODE=4'b1000;
    defparam shift_srl_15_13_LC_4_9_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_15_13_LC_4_9_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50155),
            .lcout(shift_srl_15Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93002),
            .ce(N__50119),
            .sr(_gnd_net_));
    defparam shift_srl_15_14_LC_4_9_4.C_ON=1'b0;
    defparam shift_srl_15_14_LC_4_9_4.SEQ_MODE=4'b1000;
    defparam shift_srl_15_14_LC_4_9_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_15_14_LC_4_9_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50149),
            .lcout(shift_srl_15Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93002),
            .ce(N__50119),
            .sr(_gnd_net_));
    defparam shift_srl_15_15_LC_4_9_5.C_ON=1'b0;
    defparam shift_srl_15_15_LC_4_9_5.SEQ_MODE=4'b1000;
    defparam shift_srl_15_15_LC_4_9_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_15_15_LC_4_9_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50143),
            .lcout(shift_srl_15Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93002),
            .ce(N__50119),
            .sr(_gnd_net_));
    defparam shift_srl_15_9_LC_4_9_6.C_ON=1'b0;
    defparam shift_srl_15_9_LC_4_9_6.SEQ_MODE=4'b1000;
    defparam shift_srl_15_9_LC_4_9_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_15_9_LC_4_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50125),
            .lcout(shift_srl_15Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93002),
            .ce(N__50119),
            .sr(_gnd_net_));
    defparam shift_srl_15_8_LC_4_9_7.C_ON=1'b0;
    defparam shift_srl_15_8_LC_4_9_7.SEQ_MODE=4'b1000;
    defparam shift_srl_15_8_LC_4_9_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_15_8_LC_4_9_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50131),
            .lcout(shift_srl_15Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93002),
            .ce(N__50119),
            .sr(_gnd_net_));
    defparam shift_srl_14_0_LC_4_10_0.C_ON=1'b0;
    defparam shift_srl_14_0_LC_4_10_0.SEQ_MODE=4'b1000;
    defparam shift_srl_14_0_LC_4_10_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_14_0_LC_4_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50501),
            .lcout(shift_srl_14Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92988),
            .ce(N__50203),
            .sr(_gnd_net_));
    defparam shift_srl_14_1_LC_4_10_1.C_ON=1'b0;
    defparam shift_srl_14_1_LC_4_10_1.SEQ_MODE=4'b1000;
    defparam shift_srl_14_1_LC_4_10_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_14_1_LC_4_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50251),
            .lcout(shift_srl_14Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92988),
            .ce(N__50203),
            .sr(_gnd_net_));
    defparam shift_srl_14_2_LC_4_10_2.C_ON=1'b0;
    defparam shift_srl_14_2_LC_4_10_2.SEQ_MODE=4'b1000;
    defparam shift_srl_14_2_LC_4_10_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_14_2_LC_4_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50245),
            .lcout(shift_srl_14Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92988),
            .ce(N__50203),
            .sr(_gnd_net_));
    defparam shift_srl_14_3_LC_4_10_3.C_ON=1'b0;
    defparam shift_srl_14_3_LC_4_10_3.SEQ_MODE=4'b1000;
    defparam shift_srl_14_3_LC_4_10_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_14_3_LC_4_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50239),
            .lcout(shift_srl_14Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92988),
            .ce(N__50203),
            .sr(_gnd_net_));
    defparam shift_srl_14_4_LC_4_10_4.C_ON=1'b0;
    defparam shift_srl_14_4_LC_4_10_4.SEQ_MODE=4'b1000;
    defparam shift_srl_14_4_LC_4_10_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_14_4_LC_4_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50233),
            .lcout(shift_srl_14Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92988),
            .ce(N__50203),
            .sr(_gnd_net_));
    defparam shift_srl_14_13_LC_4_10_5.C_ON=1'b0;
    defparam shift_srl_14_13_LC_4_10_5.SEQ_MODE=4'b1000;
    defparam shift_srl_14_13_LC_4_10_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_14_13_LC_4_10_5 (
            .in0(N__50221),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_14Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92988),
            .ce(N__50203),
            .sr(_gnd_net_));
    defparam shift_srl_14_14_LC_4_10_6.C_ON=1'b0;
    defparam shift_srl_14_14_LC_4_10_6.SEQ_MODE=4'b1000;
    defparam shift_srl_14_14_LC_4_10_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_14_14_LC_4_10_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50215),
            .lcout(shift_srl_14Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92988),
            .ce(N__50203),
            .sr(_gnd_net_));
    defparam shift_srl_14_15_LC_4_10_7.C_ON=1'b0;
    defparam shift_srl_14_15_LC_4_10_7.SEQ_MODE=4'b1000;
    defparam shift_srl_14_15_LC_4_10_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_14_15_LC_4_10_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50209),
            .lcout(shift_srl_14Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92988),
            .ce(N__50203),
            .sr(_gnd_net_));
    defparam shift_srl_11_RNI264O_15_LC_4_11_0.C_ON=1'b0;
    defparam shift_srl_11_RNI264O_15_LC_4_11_0.SEQ_MODE=4'b0000;
    defparam shift_srl_11_RNI264O_15_LC_4_11_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_11_RNI264O_15_LC_4_11_0 (
            .in0(N__50547),
            .in1(N__50486),
            .in2(N__50718),
            .in3(N__51348),
            .lcout(rco_int_0_a2_21_m6_0_a2_s_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_11_15_LC_4_11_1.C_ON=1'b0;
    defparam shift_srl_11_15_LC_4_11_1.SEQ_MODE=4'b1000;
    defparam shift_srl_11_15_LC_4_11_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_11_15_LC_4_11_1 (
            .in0(N__50299),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_11Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92975),
            .ce(N__51460),
            .sr(_gnd_net_));
    defparam shift_srl_11_14_LC_4_11_2.C_ON=1'b0;
    defparam shift_srl_11_14_LC_4_11_2.SEQ_MODE=4'b1000;
    defparam shift_srl_11_14_LC_4_11_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_11_14_LC_4_11_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50293),
            .lcout(shift_srl_11Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92975),
            .ce(N__51460),
            .sr(_gnd_net_));
    defparam shift_srl_11_13_LC_4_11_3.C_ON=1'b0;
    defparam shift_srl_11_13_LC_4_11_3.SEQ_MODE=4'b1000;
    defparam shift_srl_11_13_LC_4_11_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_11_13_LC_4_11_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50287),
            .lcout(shift_srl_11Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92975),
            .ce(N__51460),
            .sr(_gnd_net_));
    defparam shift_srl_11_12_LC_4_11_4.C_ON=1'b0;
    defparam shift_srl_11_12_LC_4_11_4.SEQ_MODE=4'b1000;
    defparam shift_srl_11_12_LC_4_11_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_11_12_LC_4_11_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50281),
            .lcout(shift_srl_11Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92975),
            .ce(N__51460),
            .sr(_gnd_net_));
    defparam shift_srl_11_11_LC_4_11_5.C_ON=1'b0;
    defparam shift_srl_11_11_LC_4_11_5.SEQ_MODE=4'b1000;
    defparam shift_srl_11_11_LC_4_11_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_11_11_LC_4_11_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50275),
            .lcout(shift_srl_11Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92975),
            .ce(N__51460),
            .sr(_gnd_net_));
    defparam shift_srl_11_10_LC_4_11_6.C_ON=1'b0;
    defparam shift_srl_11_10_LC_4_11_6.SEQ_MODE=4'b1000;
    defparam shift_srl_11_10_LC_4_11_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_11_10_LC_4_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50269),
            .lcout(shift_srl_11Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92975),
            .ce(N__51460),
            .sr(_gnd_net_));
    defparam shift_srl_11_9_LC_4_11_7.C_ON=1'b0;
    defparam shift_srl_11_9_LC_4_11_7.SEQ_MODE=4'b1000;
    defparam shift_srl_11_9_LC_4_11_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_11_9_LC_4_11_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51478),
            .lcout(shift_srl_11Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92975),
            .ce(N__51460),
            .sr(_gnd_net_));
    defparam shift_srl_16_10_LC_4_12_0.C_ON=1'b0;
    defparam shift_srl_16_10_LC_4_12_0.SEQ_MODE=4'b1000;
    defparam shift_srl_16_10_LC_4_12_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_16_10_LC_4_12_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51556),
            .lcout(shift_srl_16Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92964),
            .ce(N__51549),
            .sr(_gnd_net_));
    defparam shift_srl_16_11_LC_4_12_1.C_ON=1'b0;
    defparam shift_srl_16_11_LC_4_12_1.SEQ_MODE=4'b1000;
    defparam shift_srl_16_11_LC_4_12_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_16_11_LC_4_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50263),
            .lcout(shift_srl_16Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92964),
            .ce(N__51549),
            .sr(_gnd_net_));
    defparam shift_srl_16_12_LC_4_12_2.C_ON=1'b0;
    defparam shift_srl_16_12_LC_4_12_2.SEQ_MODE=4'b1000;
    defparam shift_srl_16_12_LC_4_12_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_16_12_LC_4_12_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50257),
            .lcout(shift_srl_16Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92964),
            .ce(N__51549),
            .sr(_gnd_net_));
    defparam shift_srl_16_13_LC_4_12_3.C_ON=1'b0;
    defparam shift_srl_16_13_LC_4_12_3.SEQ_MODE=4'b1000;
    defparam shift_srl_16_13_LC_4_12_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_16_13_LC_4_12_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50395),
            .lcout(shift_srl_16Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92964),
            .ce(N__51549),
            .sr(_gnd_net_));
    defparam shift_srl_16_14_LC_4_12_4.C_ON=1'b0;
    defparam shift_srl_16_14_LC_4_12_4.SEQ_MODE=4'b1000;
    defparam shift_srl_16_14_LC_4_12_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_16_14_LC_4_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50389),
            .lcout(shift_srl_16Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92964),
            .ce(N__51549),
            .sr(_gnd_net_));
    defparam shift_srl_16_15_LC_4_12_5.C_ON=1'b0;
    defparam shift_srl_16_15_LC_4_12_5.SEQ_MODE=4'b1000;
    defparam shift_srl_16_15_LC_4_12_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_16_15_LC_4_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50383),
            .lcout(shift_srl_16Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92964),
            .ce(N__51549),
            .sr(_gnd_net_));
    defparam shift_srl_16_0_LC_4_12_6.C_ON=1'b0;
    defparam shift_srl_16_0_LC_4_12_6.SEQ_MODE=4'b1000;
    defparam shift_srl_16_0_LC_4_12_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_16_0_LC_4_12_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50429),
            .lcout(shift_srl_16Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92964),
            .ce(N__51549),
            .sr(_gnd_net_));
    defparam shift_srl_16_2_LC_4_12_7.C_ON=1'b0;
    defparam shift_srl_16_2_LC_4_12_7.SEQ_MODE=4'b1000;
    defparam shift_srl_16_2_LC_4_12_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_16_2_LC_4_12_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51604),
            .lcout(shift_srl_16Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92964),
            .ce(N__51549),
            .sr(_gnd_net_));
    defparam shift_srl_12_RNIKNS64_15_LC_4_13_0.C_ON=1'b0;
    defparam shift_srl_12_RNIKNS64_15_LC_4_13_0.SEQ_MODE=4'b0000;
    defparam shift_srl_12_RNIKNS64_15_LC_4_13_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_12_RNIKNS64_15_LC_4_13_0 (
            .in0(N__50805),
            .in1(N__50365),
            .in2(N__50779),
            .in3(N__50503),
            .lcout(rco_c_14),
            .ltout(rco_c_14_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_15_RNIAERV4_15_LC_4_13_1.C_ON=1'b0;
    defparam shift_srl_15_RNIAERV4_15_LC_4_13_1.SEQ_MODE=4'b0000;
    defparam shift_srl_15_RNIAERV4_15_LC_4_13_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_15_RNIAERV4_15_LC_4_13_1 (
            .in0(N__50421),
            .in1(N__52431),
            .in2(N__50344),
            .in3(N__50549),
            .lcout(rco_c_17),
            .ltout(rco_c_17_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_20_LC_4_13_2.C_ON=1'b0;
    defparam rco_obuf_RNO_20_LC_4_13_2.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_20_LC_4_13_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 rco_obuf_RNO_20_LC_4_13_2 (
            .in0(N__50717),
            .in1(N__51746),
            .in2(N__50341),
            .in3(N__52559),
            .lcout(rco_c_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_19_RNIET865_15_LC_4_13_3.C_ON=1'b0;
    defparam shift_srl_19_RNIET865_15_LC_4_13_3.SEQ_MODE=4'b0000;
    defparam shift_srl_19_RNIET865_15_LC_4_13_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_19_RNIET865_15_LC_4_13_3 (
            .in0(N__52558),
            .in1(N__50310),
            .in2(N__50719),
            .in3(N__90403),
            .lcout(clk_en_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_15_RNIIE5K4_15_LC_4_13_4.C_ON=1'b0;
    defparam shift_srl_15_RNIIE5K4_15_LC_4_13_4.SEQ_MODE=4'b0000;
    defparam shift_srl_15_RNIIE5K4_15_LC_4_13_4.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_15_RNIIE5K4_15_LC_4_13_4 (
            .in0(N__50550),
            .in1(N__50592),
            .in2(N__90519),
            .in3(N__50422),
            .lcout(clk_en_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_12_RNI26481_15_LC_4_13_5.C_ON=1'b0;
    defparam shift_srl_12_RNI26481_15_LC_4_13_5.SEQ_MODE=4'b0000;
    defparam shift_srl_12_RNI26481_15_LC_4_13_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_12_RNI26481_15_LC_4_13_5 (
            .in0(N__50420),
            .in1(N__50771),
            .in2(N__52439),
            .in3(N__50804),
            .lcout(),
            .ltout(rco_int_0_a2_21_m6_0_a2_s_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_21_RNII6642_15_LC_4_13_6.C_ON=1'b0;
    defparam shift_srl_21_RNII6642_15_LC_4_13_6.SEQ_MODE=4'b0000;
    defparam shift_srl_21_RNII6642_15_LC_4_13_6.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_21_RNII6642_15_LC_4_13_6 (
            .in0(N__50644),
            .in1(N__51745),
            .in2(N__50581),
            .in3(N__52557),
            .lcout(rco_int_0_a2_21_m6_0_a2_s_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_17_15_LC_4_13_7.C_ON=1'b0;
    defparam shift_srl_17_15_LC_4_13_7.SEQ_MODE=4'b1000;
    defparam shift_srl_17_15_LC_4_13_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_17_15_LC_4_13_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52708),
            .lcout(shift_srl_17Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92952),
            .ce(N__52676),
            .sr(_gnd_net_));
    defparam shift_srl_18_RNIUTH05_15_LC_4_14_0.C_ON=1'b0;
    defparam shift_srl_18_RNIUTH05_15_LC_4_14_0.SEQ_MODE=4'b0000;
    defparam shift_srl_18_RNIUTH05_15_LC_4_14_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_18_RNIUTH05_15_LC_4_14_0 (
            .in0(N__50702),
            .in1(N__52429),
            .in2(N__50451),
            .in3(N__50430),
            .lcout(rco_c_18),
            .ltout(rco_c_18_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_20_RNIRHOF5_15_LC_4_14_1.C_ON=1'b0;
    defparam shift_srl_20_RNIRHOF5_15_LC_4_14_1.SEQ_MODE=4'b0000;
    defparam shift_srl_20_RNIRHOF5_15_LC_4_14_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_20_RNIRHOF5_15_LC_4_14_1 (
            .in0(N__90464),
            .in1(N__51751),
            .in2(N__50560),
            .in3(N__52561),
            .lcout(clk_en_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_11_RNIMLQ51_0_15_LC_4_14_2.C_ON=1'b0;
    defparam shift_srl_11_RNIMLQ51_0_15_LC_4_14_2.SEQ_MODE=4'b0000;
    defparam shift_srl_11_RNIMLQ51_0_15_LC_4_14_2.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_11_RNIMLQ51_0_15_LC_4_14_2 (
            .in0(N__55731),
            .in1(N__50775),
            .in2(N__51372),
            .in3(N__50816),
            .lcout(),
            .ltout(rco_int_0_a2_sx_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_15_RNI5R0B4_15_LC_4_14_3.C_ON=1'b0;
    defparam shift_srl_15_RNI5R0B4_15_LC_4_14_3.SEQ_MODE=4'b0000;
    defparam shift_srl_15_RNI5R0B4_15_LC_4_14_3.LUT_INIT=16'b0000100000000000;
    LogicCell40 shift_srl_15_RNI5R0B4_15_LC_4_14_3 (
            .in0(N__69178),
            .in1(N__50548),
            .in2(N__50512),
            .in3(N__50502),
            .lcout(rco_c_15),
            .ltout(rco_c_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_16_RNI5QL05_15_LC_4_14_4.C_ON=1'b0;
    defparam shift_srl_16_RNI5QL05_15_LC_4_14_4.SEQ_MODE=4'b0000;
    defparam shift_srl_16_RNI5QL05_15_LC_4_14_4.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_16_RNI5QL05_15_LC_4_14_4 (
            .in0(N__90463),
            .in1(N__52430),
            .in2(N__50434),
            .in3(N__50431),
            .lcout(clk_en_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_11_RNIMLQ51_15_LC_4_14_5.C_ON=1'b0;
    defparam shift_srl_11_RNIMLQ51_15_LC_4_14_5.SEQ_MODE=4'b0000;
    defparam shift_srl_11_RNIMLQ51_15_LC_4_14_5.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_11_RNIMLQ51_15_LC_4_14_5 (
            .in0(N__50817),
            .in1(N__55732),
            .in2(N__51373),
            .in3(N__50776),
            .lcout(rco_int_0_a2_sx_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_18_0_LC_4_14_6.C_ON=1'b0;
    defparam shift_srl_18_0_LC_4_14_6.SEQ_MODE=4'b1000;
    defparam shift_srl_18_0_LC_4_14_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_18_0_LC_4_14_6 (
            .in0(N__50703),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_18Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92942),
            .ce(N__50852),
            .sr(_gnd_net_));
    defparam shift_srl_18_1_LC_4_14_7.C_ON=1'b0;
    defparam shift_srl_18_1_LC_4_14_7.SEQ_MODE=4'b1000;
    defparam shift_srl_18_1_LC_4_14_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_18_1_LC_4_14_7 (
            .in0(N__50650),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_18Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92942),
            .ce(N__50852),
            .sr(_gnd_net_));
    defparam shift_srl_21_0_LC_4_15_0.C_ON=1'b0;
    defparam shift_srl_21_0_LC_4_15_0.SEQ_MODE=4'b1000;
    defparam shift_srl_21_0_LC_4_15_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_21_0_LC_4_15_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50643),
            .lcout(shift_srl_21Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92935),
            .ce(N__50919),
            .sr(_gnd_net_));
    defparam shift_srl_21_1_LC_4_15_1.C_ON=1'b0;
    defparam shift_srl_21_1_LC_4_15_1.SEQ_MODE=4'b1000;
    defparam shift_srl_21_1_LC_4_15_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_21_1_LC_4_15_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50629),
            .lcout(shift_srl_21Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92935),
            .ce(N__50919),
            .sr(_gnd_net_));
    defparam shift_srl_21_2_LC_4_15_2.C_ON=1'b0;
    defparam shift_srl_21_2_LC_4_15_2.SEQ_MODE=4'b1000;
    defparam shift_srl_21_2_LC_4_15_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_21_2_LC_4_15_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50623),
            .lcout(shift_srl_21Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92935),
            .ce(N__50919),
            .sr(_gnd_net_));
    defparam shift_srl_21_3_LC_4_15_3.C_ON=1'b0;
    defparam shift_srl_21_3_LC_4_15_3.SEQ_MODE=4'b1000;
    defparam shift_srl_21_3_LC_4_15_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_21_3_LC_4_15_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50617),
            .lcout(shift_srl_21Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92935),
            .ce(N__50919),
            .sr(_gnd_net_));
    defparam shift_srl_21_4_LC_4_15_4.C_ON=1'b0;
    defparam shift_srl_21_4_LC_4_15_4.SEQ_MODE=4'b1000;
    defparam shift_srl_21_4_LC_4_15_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_21_4_LC_4_15_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50611),
            .lcout(shift_srl_21Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92935),
            .ce(N__50919),
            .sr(_gnd_net_));
    defparam shift_srl_21_5_LC_4_15_5.C_ON=1'b0;
    defparam shift_srl_21_5_LC_4_15_5.SEQ_MODE=4'b1000;
    defparam shift_srl_21_5_LC_4_15_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_21_5_LC_4_15_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50605),
            .lcout(shift_srl_21Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92935),
            .ce(N__50919),
            .sr(_gnd_net_));
    defparam shift_srl_21_6_LC_4_15_6.C_ON=1'b0;
    defparam shift_srl_21_6_LC_4_15_6.SEQ_MODE=4'b1000;
    defparam shift_srl_21_6_LC_4_15_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_21_6_LC_4_15_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50938),
            .lcout(shift_srl_21Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92935),
            .ce(N__50919),
            .sr(_gnd_net_));
    defparam shift_srl_21_7_LC_4_15_7.C_ON=1'b0;
    defparam shift_srl_21_7_LC_4_15_7.SEQ_MODE=4'b1000;
    defparam shift_srl_21_7_LC_4_15_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_21_7_LC_4_15_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50932),
            .lcout(shift_srl_21Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92935),
            .ce(N__50919),
            .sr(_gnd_net_));
    defparam shift_srl_18_2_LC_4_16_0.C_ON=1'b0;
    defparam shift_srl_18_2_LC_4_16_0.SEQ_MODE=4'b1000;
    defparam shift_srl_18_2_LC_4_16_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_18_2_LC_4_16_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50899),
            .lcout(shift_srl_18Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92927),
            .ce(N__50853),
            .sr(_gnd_net_));
    defparam shift_srl_18_3_LC_4_16_1.C_ON=1'b0;
    defparam shift_srl_18_3_LC_4_16_1.SEQ_MODE=4'b1000;
    defparam shift_srl_18_3_LC_4_16_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_18_3_LC_4_16_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50890),
            .lcout(shift_srl_18Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92927),
            .ce(N__50853),
            .sr(_gnd_net_));
    defparam shift_srl_18_4_LC_4_16_2.C_ON=1'b0;
    defparam shift_srl_18_4_LC_4_16_2.SEQ_MODE=4'b1000;
    defparam shift_srl_18_4_LC_4_16_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_18_4_LC_4_16_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50884),
            .lcout(shift_srl_18Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92927),
            .ce(N__50853),
            .sr(_gnd_net_));
    defparam shift_srl_18_5_LC_4_16_3.C_ON=1'b0;
    defparam shift_srl_18_5_LC_4_16_3.SEQ_MODE=4'b1000;
    defparam shift_srl_18_5_LC_4_16_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_18_5_LC_4_16_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50878),
            .lcout(shift_srl_18Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92927),
            .ce(N__50853),
            .sr(_gnd_net_));
    defparam shift_srl_18_6_LC_4_16_4.C_ON=1'b0;
    defparam shift_srl_18_6_LC_4_16_4.SEQ_MODE=4'b1000;
    defparam shift_srl_18_6_LC_4_16_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_18_6_LC_4_16_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50872),
            .lcout(shift_srl_18Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92927),
            .ce(N__50853),
            .sr(_gnd_net_));
    defparam shift_srl_18_7_LC_4_16_5.C_ON=1'b0;
    defparam shift_srl_18_7_LC_4_16_5.SEQ_MODE=4'b1000;
    defparam shift_srl_18_7_LC_4_16_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_18_7_LC_4_16_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50866),
            .lcout(shift_srl_18Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92927),
            .ce(N__50853),
            .sr(_gnd_net_));
    defparam shift_srl_134_RNIVHU51_15_LC_4_17_0.C_ON=1'b0;
    defparam shift_srl_134_RNIVHU51_15_LC_4_17_0.SEQ_MODE=4'b0000;
    defparam shift_srl_134_RNIVHU51_15_LC_4_17_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_134_RNIVHU51_15_LC_4_17_0 (
            .in0(N__90399),
            .in1(N__52020),
            .in2(N__66237),
            .in3(N__52930),
            .lcout(g0_11_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_133_15_LC_4_17_1.C_ON=1'b0;
    defparam shift_srl_133_15_LC_4_17_1.SEQ_MODE=4'b1000;
    defparam shift_srl_133_15_LC_4_17_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_133_15_LC_4_17_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51285),
            .lcout(shift_srl_133Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92915),
            .ce(N__55375),
            .sr(_gnd_net_));
    defparam shift_srl_133_14_LC_4_17_2.C_ON=1'b0;
    defparam shift_srl_133_14_LC_4_17_2.SEQ_MODE=4'b1000;
    defparam shift_srl_133_14_LC_4_17_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_133_14_LC_4_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50968),
            .lcout(shift_srl_133Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92915),
            .ce(N__55375),
            .sr(_gnd_net_));
    defparam shift_srl_133_13_LC_4_17_3.C_ON=1'b0;
    defparam shift_srl_133_13_LC_4_17_3.SEQ_MODE=4'b1000;
    defparam shift_srl_133_13_LC_4_17_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_133_13_LC_4_17_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50962),
            .lcout(shift_srl_133Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92915),
            .ce(N__55375),
            .sr(_gnd_net_));
    defparam shift_srl_133_12_LC_4_17_4.C_ON=1'b0;
    defparam shift_srl_133_12_LC_4_17_4.SEQ_MODE=4'b1000;
    defparam shift_srl_133_12_LC_4_17_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_133_12_LC_4_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50956),
            .lcout(shift_srl_133Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92915),
            .ce(N__55375),
            .sr(_gnd_net_));
    defparam shift_srl_133_11_LC_4_17_5.C_ON=1'b0;
    defparam shift_srl_133_11_LC_4_17_5.SEQ_MODE=4'b1000;
    defparam shift_srl_133_11_LC_4_17_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_133_11_LC_4_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51859),
            .lcout(shift_srl_133Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92915),
            .ce(N__55375),
            .sr(_gnd_net_));
    defparam shift_srl_131_0_LC_4_18_0.C_ON=1'b0;
    defparam shift_srl_131_0_LC_4_18_0.SEQ_MODE=4'b1000;
    defparam shift_srl_131_0_LC_4_18_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_131_0_LC_4_18_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54297),
            .lcout(shift_srl_131Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92928),
            .ce(N__51888),
            .sr(_gnd_net_));
    defparam shift_srl_131_8_LC_4_18_1.C_ON=1'b0;
    defparam shift_srl_131_8_LC_4_18_1.SEQ_MODE=4'b1000;
    defparam shift_srl_131_8_LC_4_18_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_131_8_LC_4_18_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51034),
            .lcout(shift_srl_131Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92928),
            .ce(N__51888),
            .sr(_gnd_net_));
    defparam shift_srl_131_2_LC_4_18_2.C_ON=1'b0;
    defparam shift_srl_131_2_LC_4_18_2.SEQ_MODE=4'b1000;
    defparam shift_srl_131_2_LC_4_18_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_131_2_LC_4_18_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51895),
            .lcout(shift_srl_131Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92928),
            .ce(N__51888),
            .sr(_gnd_net_));
    defparam shift_srl_131_3_LC_4_18_3.C_ON=1'b0;
    defparam shift_srl_131_3_LC_4_18_3.SEQ_MODE=4'b1000;
    defparam shift_srl_131_3_LC_4_18_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_131_3_LC_4_18_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50950),
            .lcout(shift_srl_131Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92928),
            .ce(N__51888),
            .sr(_gnd_net_));
    defparam shift_srl_131_4_LC_4_18_4.C_ON=1'b0;
    defparam shift_srl_131_4_LC_4_18_4.SEQ_MODE=4'b1000;
    defparam shift_srl_131_4_LC_4_18_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_131_4_LC_4_18_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50944),
            .lcout(shift_srl_131Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92928),
            .ce(N__51888),
            .sr(_gnd_net_));
    defparam shift_srl_131_5_LC_4_18_5.C_ON=1'b0;
    defparam shift_srl_131_5_LC_4_18_5.SEQ_MODE=4'b1000;
    defparam shift_srl_131_5_LC_4_18_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_131_5_LC_4_18_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51052),
            .lcout(shift_srl_131Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92928),
            .ce(N__51888),
            .sr(_gnd_net_));
    defparam shift_srl_131_6_LC_4_18_6.C_ON=1'b0;
    defparam shift_srl_131_6_LC_4_18_6.SEQ_MODE=4'b1000;
    defparam shift_srl_131_6_LC_4_18_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_131_6_LC_4_18_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51046),
            .lcout(shift_srl_131Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92928),
            .ce(N__51888),
            .sr(_gnd_net_));
    defparam shift_srl_131_7_LC_4_18_7.C_ON=1'b0;
    defparam shift_srl_131_7_LC_4_18_7.SEQ_MODE=4'b1000;
    defparam shift_srl_131_7_LC_4_18_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_131_7_LC_4_18_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51040),
            .lcout(shift_srl_131Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92928),
            .ce(N__51888),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_0_131_LC_4_19_0.C_ON=1'b0;
    defparam rco_obuf_RNO_0_131_LC_4_19_0.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_0_131_LC_4_19_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 rco_obuf_RNO_0_131_LC_4_19_0 (
            .in0(N__54229),
            .in1(N__91249),
            .in2(N__52931),
            .in3(N__54298),
            .lcout(),
            .ltout(rco_obuf_RNO_0Z0Z_131_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_131_LC_4_19_1.C_ON=1'b0;
    defparam rco_obuf_RNO_131_LC_4_19_1.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_131_LC_4_19_1.LUT_INIT=16'b1010000010100000;
    LogicCell40 rco_obuf_RNO_131_LC_4_19_1 (
            .in0(N__91336),
            .in1(_gnd_net_),
            .in2(N__51028),
            .in3(_gnd_net_),
            .lcout(rco_c_131),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_130_LC_4_19_2.C_ON=1'b0;
    defparam rco_obuf_RNO_130_LC_4_19_2.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_130_LC_4_19_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 rco_obuf_RNO_130_LC_4_19_2 (
            .in0(N__54230),
            .in1(N__91335),
            .in2(N__52932),
            .in3(N__91250),
            .lcout(rco_c_130),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_129_RNI7G7R_15_LC_4_19_3.C_ON=1'b0;
    defparam shift_srl_129_RNI7G7R_15_LC_4_19_3.SEQ_MODE=4'b0000;
    defparam shift_srl_129_RNI7G7R_15_LC_4_19_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_129_RNI7G7R_15_LC_4_19_3 (
            .in0(N__91247),
            .in1(N__52917),
            .in2(N__90530),
            .in3(N__54228),
            .lcout(g0_2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_118_RNI2TIHV_15_LC_4_19_4.C_ON=1'b0;
    defparam shift_srl_118_RNI2TIHV_15_LC_4_19_4.SEQ_MODE=4'b0000;
    defparam shift_srl_118_RNI2TIHV_15_LC_4_19_4.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_118_RNI2TIHV_15_LC_4_19_4 (
            .in0(N__58738),
            .in1(N__65341),
            .in2(N__65566),
            .in3(N__79389),
            .lcout(rco_c_123),
            .ltout(rco_c_123_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_132_RNIOHTB11_15_LC_4_19_5.C_ON=1'b0;
    defparam shift_srl_132_RNIOHTB11_15_LC_4_19_5.SEQ_MODE=4'b0000;
    defparam shift_srl_132_RNIOHTB11_15_LC_4_19_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_132_RNIOHTB11_15_LC_4_19_5 (
            .in0(N__54151),
            .in1(N__50989),
            .in2(N__50983),
            .in3(N__65742),
            .lcout(clk_en_133),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_129_RNIN9Q411_15_LC_4_19_6.C_ON=1'b0;
    defparam shift_srl_129_RNIN9Q411_15_LC_4_19_6.SEQ_MODE=4'b0000;
    defparam shift_srl_129_RNIN9Q411_15_LC_4_19_6.LUT_INIT=16'b1010000000000000;
    LogicCell40 shift_srl_129_RNIN9Q411_15_LC_4_19_6 (
            .in0(N__57577),
            .in1(_gnd_net_),
            .in2(N__65754),
            .in3(N__51106),
            .lcout(clk_en_131),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_128_RNIHESE01_15_LC_4_19_7.C_ON=1'b0;
    defparam shift_srl_128_RNIHESE01_15_LC_4_19_7.SEQ_MODE=4'b0000;
    defparam shift_srl_128_RNIHESE01_15_LC_4_19_7.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_128_RNIHESE01_15_LC_4_19_7 (
            .in0(N__91248),
            .in1(N__65746),
            .in2(N__90531),
            .in3(N__57576),
            .lcout(clk_en_129),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_133_RNIEU741_15_LC_4_20_0.C_ON=1'b0;
    defparam shift_srl_133_RNIEU741_15_LC_4_20_0.SEQ_MODE=4'b0000;
    defparam shift_srl_133_RNIEU741_15_LC_4_20_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_133_RNIEU741_15_LC_4_20_0 (
            .in0(N__91266),
            .in1(N__52910),
            .in2(N__54232),
            .in3(N__66242),
            .lcout(g0_11_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_136_RNIHAQ01_15_LC_4_20_2.C_ON=1'b0;
    defparam shift_srl_136_RNIHAQ01_15_LC_4_20_2.SEQ_MODE=4'b0000;
    defparam shift_srl_136_RNIHAQ01_15_LC_4_20_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_136_RNIHAQ01_15_LC_4_20_2 (
            .in0(N__91267),
            .in1(N__54468),
            .in2(N__54233),
            .in3(N__52911),
            .lcout(g0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_129_14_LC_4_20_3.C_ON=1'b0;
    defparam shift_srl_129_14_LC_4_20_3.SEQ_MODE=4'b1000;
    defparam shift_srl_129_14_LC_4_20_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_129_14_LC_4_20_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51088),
            .lcout(shift_srl_129Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92943),
            .ce(N__53986),
            .sr(_gnd_net_));
    defparam shift_srl_129_13_LC_4_20_4.C_ON=1'b0;
    defparam shift_srl_129_13_LC_4_20_4.SEQ_MODE=4'b1000;
    defparam shift_srl_129_13_LC_4_20_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_129_13_LC_4_20_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51082),
            .lcout(shift_srl_129Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92943),
            .ce(N__53986),
            .sr(_gnd_net_));
    defparam shift_srl_129_12_LC_4_20_5.C_ON=1'b0;
    defparam shift_srl_129_12_LC_4_20_5.SEQ_MODE=4'b1000;
    defparam shift_srl_129_12_LC_4_20_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_129_12_LC_4_20_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51076),
            .lcout(shift_srl_129Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92943),
            .ce(N__53986),
            .sr(_gnd_net_));
    defparam shift_srl_129_11_LC_4_20_6.C_ON=1'b0;
    defparam shift_srl_129_11_LC_4_20_6.SEQ_MODE=4'b1000;
    defparam shift_srl_129_11_LC_4_20_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_129_11_LC_4_20_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51058),
            .lcout(shift_srl_129Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92943),
            .ce(N__53986),
            .sr(_gnd_net_));
    defparam shift_srl_129_10_LC_4_20_7.C_ON=1'b0;
    defparam shift_srl_129_10_LC_4_20_7.SEQ_MODE=4'b1000;
    defparam shift_srl_129_10_LC_4_20_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_129_10_LC_4_20_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51070),
            .lcout(shift_srl_129Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92943),
            .ce(N__53986),
            .sr(_gnd_net_));
    defparam shift_srl_134_10_LC_4_21_0.C_ON=1'b0;
    defparam shift_srl_134_10_LC_4_21_0.SEQ_MODE=4'b1000;
    defparam shift_srl_134_10_LC_4_21_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_134_10_LC_4_21_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51136),
            .lcout(shift_srl_134Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92953),
            .ce(N__53003),
            .sr(_gnd_net_));
    defparam shift_srl_134_11_LC_4_21_1.C_ON=1'b0;
    defparam shift_srl_134_11_LC_4_21_1.SEQ_MODE=4'b1000;
    defparam shift_srl_134_11_LC_4_21_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_134_11_LC_4_21_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51166),
            .lcout(shift_srl_134Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92953),
            .ce(N__53003),
            .sr(_gnd_net_));
    defparam shift_srl_134_12_LC_4_21_2.C_ON=1'b0;
    defparam shift_srl_134_12_LC_4_21_2.SEQ_MODE=4'b1000;
    defparam shift_srl_134_12_LC_4_21_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_134_12_LC_4_21_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51160),
            .lcout(shift_srl_134Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92953),
            .ce(N__53003),
            .sr(_gnd_net_));
    defparam shift_srl_134_13_LC_4_21_3.C_ON=1'b0;
    defparam shift_srl_134_13_LC_4_21_3.SEQ_MODE=4'b1000;
    defparam shift_srl_134_13_LC_4_21_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_134_13_LC_4_21_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51154),
            .lcout(shift_srl_134Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92953),
            .ce(N__53003),
            .sr(_gnd_net_));
    defparam shift_srl_134_14_LC_4_21_4.C_ON=1'b0;
    defparam shift_srl_134_14_LC_4_21_4.SEQ_MODE=4'b1000;
    defparam shift_srl_134_14_LC_4_21_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_134_14_LC_4_21_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51148),
            .lcout(shift_srl_134Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92953),
            .ce(N__53003),
            .sr(_gnd_net_));
    defparam shift_srl_134_15_LC_4_21_5.C_ON=1'b0;
    defparam shift_srl_134_15_LC_4_21_5.SEQ_MODE=4'b1000;
    defparam shift_srl_134_15_LC_4_21_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_134_15_LC_4_21_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51142),
            .lcout(shift_srl_134Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92953),
            .ce(N__53003),
            .sr(_gnd_net_));
    defparam shift_srl_134_9_LC_4_21_6.C_ON=1'b0;
    defparam shift_srl_134_9_LC_4_21_6.SEQ_MODE=4'b1000;
    defparam shift_srl_134_9_LC_4_21_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_134_9_LC_4_21_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51130),
            .lcout(shift_srl_134Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92953),
            .ce(N__53003),
            .sr(_gnd_net_));
    defparam shift_srl_134_8_LC_4_21_7.C_ON=1'b0;
    defparam shift_srl_134_8_LC_4_21_7.SEQ_MODE=4'b1000;
    defparam shift_srl_134_8_LC_4_21_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_134_8_LC_4_21_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53017),
            .lcout(shift_srl_134Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92953),
            .ce(N__53003),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_137_LC_4_22_0.C_ON=1'b0;
    defparam rco_obuf_RNO_137_LC_4_22_0.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_137_LC_4_22_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 rco_obuf_RNO_137_LC_4_22_0 (
            .in0(N__66302),
            .in1(N__51264),
            .in2(N__51217),
            .in3(N__54474),
            .lcout(rco_c_137),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_133_fast_RNIML0I_15_LC_4_22_1.C_ON=1'b0;
    defparam shift_srl_133_fast_RNIML0I_15_LC_4_22_1.SEQ_MODE=4'b0000;
    defparam shift_srl_133_fast_RNIML0I_15_LC_4_22_1.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_133_fast_RNIML0I_15_LC_4_22_1 (
            .in0(N__53085),
            .in1(N__52006),
            .in2(_gnd_net_),
            .in3(N__51274),
            .lcout(shift_srl_133_fast_RNIML0IZ0Z_15),
            .ltout(shift_srl_133_fast_RNIML0IZ0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_138_RNI8KQH1_15_LC_4_22_2.C_ON=1'b0;
    defparam shift_srl_138_RNI8KQH1_15_LC_4_22_2.SEQ_MODE=4'b0000;
    defparam shift_srl_138_RNI8KQH1_15_LC_4_22_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_138_RNI8KQH1_15_LC_4_22_2 (
            .in0(N__51325),
            .in1(N__51262),
            .in2(N__51310),
            .in3(N__54472),
            .lcout(rco_int_0_a3_0_a2_0_138),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_136_LC_4_22_3.C_ON=1'b0;
    defparam rco_obuf_RNO_136_LC_4_22_3.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_136_LC_4_22_3.LUT_INIT=16'b1000100000000000;
    LogicCell40 rco_obuf_RNO_136_LC_4_22_3 (
            .in0(N__54473),
            .in1(N__66301),
            .in2(_gnd_net_),
            .in3(N__51212),
            .lcout(rco_c_136),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_133_fast_15_LC_4_22_4.C_ON=1'b0;
    defparam shift_srl_133_fast_15_LC_4_22_4.SEQ_MODE=4'b1000;
    defparam shift_srl_133_fast_15_LC_4_22_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_133_fast_15_LC_4_22_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51289),
            .lcout(shift_srl_133_fastZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92965),
            .ce(N__55377),
            .sr(_gnd_net_));
    defparam shift_srl_137_RNIF4M41_15_LC_4_22_6.C_ON=1'b0;
    defparam shift_srl_137_RNIF4M41_15_LC_4_22_6.SEQ_MODE=4'b0000;
    defparam shift_srl_137_RNIF4M41_15_LC_4_22_6.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_137_RNIF4M41_15_LC_4_22_6 (
            .in0(N__52007),
            .in1(N__51263),
            .in2(N__53099),
            .in3(N__66243),
            .lcout(g0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_134_LC_4_22_7.C_ON=1'b0;
    defparam rco_obuf_RNO_134_LC_4_22_7.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_134_LC_4_22_7.LUT_INIT=16'b1000100000000000;
    LogicCell40 rco_obuf_RNO_134_LC_4_22_7 (
            .in0(N__66244),
            .in1(N__66300),
            .in2(_gnd_net_),
            .in3(N__52008),
            .lcout(rco_c_134),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_135_LC_4_23_5.C_ON=1'b0;
    defparam rco_obuf_RNO_135_LC_4_23_5.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_135_LC_4_23_5.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_135_LC_4_23_5 (
            .in0(N__51216),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66299),
            .lcout(rco_c_135),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_125_LC_4_24_0.C_ON=1'b0;
    defparam rco_obuf_RNO_125_LC_4_24_0.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_125_LC_4_24_0.LUT_INIT=16'b1000100000000000;
    LogicCell40 rco_obuf_RNO_125_LC_4_24_0 (
            .in0(N__66037),
            .in1(N__65457),
            .in2(_gnd_net_),
            .in3(N__57617),
            .lcout(rco_c_125),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_22_10_LC_5_8_0.C_ON=1'b0;
    defparam shift_srl_22_10_LC_5_8_0.SEQ_MODE=4'b1000;
    defparam shift_srl_22_10_LC_5_8_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_22_10_LC_5_8_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51379),
            .lcout(shift_srl_22Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93032),
            .ce(N__52206),
            .sr(_gnd_net_));
    defparam shift_srl_22_11_LC_5_8_1.C_ON=1'b0;
    defparam shift_srl_22_11_LC_5_8_1.SEQ_MODE=4'b1000;
    defparam shift_srl_22_11_LC_5_8_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_22_11_LC_5_8_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51424),
            .lcout(shift_srl_22Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93032),
            .ce(N__52206),
            .sr(_gnd_net_));
    defparam shift_srl_22_12_LC_5_8_2.C_ON=1'b0;
    defparam shift_srl_22_12_LC_5_8_2.SEQ_MODE=4'b1000;
    defparam shift_srl_22_12_LC_5_8_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_22_12_LC_5_8_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51418),
            .lcout(shift_srl_22Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93032),
            .ce(N__52206),
            .sr(_gnd_net_));
    defparam shift_srl_22_14_LC_5_8_4.C_ON=1'b0;
    defparam shift_srl_22_14_LC_5_8_4.SEQ_MODE=4'b1000;
    defparam shift_srl_22_14_LC_5_8_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_22_14_LC_5_8_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51406),
            .lcout(shift_srl_22Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93032),
            .ce(N__52206),
            .sr(_gnd_net_));
    defparam shift_srl_22_13_LC_5_8_6.C_ON=1'b0;
    defparam shift_srl_22_13_LC_5_8_6.SEQ_MODE=4'b1000;
    defparam shift_srl_22_13_LC_5_8_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_22_13_LC_5_8_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51412),
            .lcout(shift_srl_22Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93032),
            .ce(N__52206),
            .sr(_gnd_net_));
    defparam shift_srl_22_8_LC_5_8_7.C_ON=1'b0;
    defparam shift_srl_22_8_LC_5_8_7.SEQ_MODE=4'b1000;
    defparam shift_srl_22_8_LC_5_8_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_22_8_LC_5_8_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51400),
            .lcout(shift_srl_22Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93032),
            .ce(N__52206),
            .sr(_gnd_net_));
    defparam shift_srl_22_15_LC_5_9_1.C_ON=1'b0;
    defparam shift_srl_22_15_LC_5_9_1.SEQ_MODE=4'b1000;
    defparam shift_srl_22_15_LC_5_9_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_22_15_LC_5_9_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51391),
            .lcout(shift_srl_22Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93018),
            .ce(N__52197),
            .sr(_gnd_net_));
    defparam shift_srl_22_9_LC_5_9_3.C_ON=1'b0;
    defparam shift_srl_22_9_LC_5_9_3.SEQ_MODE=4'b1000;
    defparam shift_srl_22_9_LC_5_9_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_22_9_LC_5_9_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51385),
            .lcout(shift_srl_22Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93018),
            .ce(N__52197),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNILT313_15_LC_5_10_0.C_ON=1'b0;
    defparam shift_srl_0_RNILT313_15_LC_5_10_0.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNILT313_15_LC_5_10_0.LUT_INIT=16'b1100110000000000;
    LogicCell40 shift_srl_0_RNILT313_15_LC_5_10_0 (
            .in0(_gnd_net_),
            .in1(N__90044),
            .in2(_gnd_net_),
            .in3(N__52311),
            .lcout(clk_en_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_11_0_LC_5_10_1.C_ON=1'b0;
    defparam shift_srl_11_0_LC_5_10_1.SEQ_MODE=4'b1000;
    defparam shift_srl_11_0_LC_5_10_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_11_0_LC_5_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51358),
            .lcout(shift_srl_11Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93003),
            .ce(N__51449),
            .sr(_gnd_net_));
    defparam shift_srl_11_1_LC_5_10_2.C_ON=1'b0;
    defparam shift_srl_11_1_LC_5_10_2.SEQ_MODE=4'b1000;
    defparam shift_srl_11_1_LC_5_10_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_11_1_LC_5_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51514),
            .lcout(shift_srl_11Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93003),
            .ce(N__51449),
            .sr(_gnd_net_));
    defparam shift_srl_11_2_LC_5_10_3.C_ON=1'b0;
    defparam shift_srl_11_2_LC_5_10_3.SEQ_MODE=4'b1000;
    defparam shift_srl_11_2_LC_5_10_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_11_2_LC_5_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51508),
            .lcout(shift_srl_11Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93003),
            .ce(N__51449),
            .sr(_gnd_net_));
    defparam shift_srl_11_3_LC_5_10_4.C_ON=1'b0;
    defparam shift_srl_11_3_LC_5_10_4.SEQ_MODE=4'b1000;
    defparam shift_srl_11_3_LC_5_10_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_11_3_LC_5_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51502),
            .lcout(shift_srl_11Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93003),
            .ce(N__51449),
            .sr(_gnd_net_));
    defparam shift_srl_11_4_LC_5_10_5.C_ON=1'b0;
    defparam shift_srl_11_4_LC_5_10_5.SEQ_MODE=4'b1000;
    defparam shift_srl_11_4_LC_5_10_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_11_4_LC_5_10_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51496),
            .lcout(shift_srl_11Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93003),
            .ce(N__51449),
            .sr(_gnd_net_));
    defparam shift_srl_11_5_LC_5_10_6.C_ON=1'b0;
    defparam shift_srl_11_5_LC_5_10_6.SEQ_MODE=4'b1000;
    defparam shift_srl_11_5_LC_5_10_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_11_5_LC_5_10_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51490),
            .lcout(shift_srl_11Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93003),
            .ce(N__51449),
            .sr(_gnd_net_));
    defparam shift_srl_11_7_LC_5_11_0.C_ON=1'b0;
    defparam shift_srl_11_7_LC_5_11_0.SEQ_MODE=4'b1000;
    defparam shift_srl_11_7_LC_5_11_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_11_7_LC_5_11_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51466),
            .lcout(shift_srl_11Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92989),
            .ce(N__51456),
            .sr(_gnd_net_));
    defparam shift_srl_11_8_LC_5_11_1.C_ON=1'b0;
    defparam shift_srl_11_8_LC_5_11_1.SEQ_MODE=4'b1000;
    defparam shift_srl_11_8_LC_5_11_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_11_8_LC_5_11_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51484),
            .lcout(shift_srl_11Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92989),
            .ce(N__51456),
            .sr(_gnd_net_));
    defparam shift_srl_11_6_LC_5_11_6.C_ON=1'b0;
    defparam shift_srl_11_6_LC_5_11_6.SEQ_MODE=4'b1000;
    defparam shift_srl_11_6_LC_5_11_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_11_6_LC_5_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51472),
            .lcout(shift_srl_11Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92989),
            .ce(N__51456),
            .sr(_gnd_net_));
    defparam shift_srl_16_7_LC_5_12_0.C_ON=1'b0;
    defparam shift_srl_16_7_LC_5_12_0.SEQ_MODE=4'b1000;
    defparam shift_srl_16_7_LC_5_12_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_16_7_LC_5_12_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51568),
            .lcout(shift_srl_16Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92976),
            .ce(N__51550),
            .sr(_gnd_net_));
    defparam shift_srl_16_1_LC_5_12_1.C_ON=1'b0;
    defparam shift_srl_16_1_LC_5_12_1.SEQ_MODE=4'b1000;
    defparam shift_srl_16_1_LC_5_12_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_16_1_LC_5_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51430),
            .lcout(shift_srl_16Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92976),
            .ce(N__51550),
            .sr(_gnd_net_));
    defparam shift_srl_16_8_LC_5_12_2.C_ON=1'b0;
    defparam shift_srl_16_8_LC_5_12_2.SEQ_MODE=4'b1000;
    defparam shift_srl_16_8_LC_5_12_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_16_8_LC_5_12_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51598),
            .lcout(shift_srl_16Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92976),
            .ce(N__51550),
            .sr(_gnd_net_));
    defparam shift_srl_16_3_LC_5_12_3.C_ON=1'b0;
    defparam shift_srl_16_3_LC_5_12_3.SEQ_MODE=4'b1000;
    defparam shift_srl_16_3_LC_5_12_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_16_3_LC_5_12_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51592),
            .lcout(shift_srl_16Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92976),
            .ce(N__51550),
            .sr(_gnd_net_));
    defparam shift_srl_16_4_LC_5_12_4.C_ON=1'b0;
    defparam shift_srl_16_4_LC_5_12_4.SEQ_MODE=4'b1000;
    defparam shift_srl_16_4_LC_5_12_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_16_4_LC_5_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51586),
            .lcout(shift_srl_16Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92976),
            .ce(N__51550),
            .sr(_gnd_net_));
    defparam shift_srl_16_5_LC_5_12_5.C_ON=1'b0;
    defparam shift_srl_16_5_LC_5_12_5.SEQ_MODE=4'b1000;
    defparam shift_srl_16_5_LC_5_12_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_16_5_LC_5_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51580),
            .lcout(shift_srl_16Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92976),
            .ce(N__51550),
            .sr(_gnd_net_));
    defparam shift_srl_16_6_LC_5_12_6.C_ON=1'b0;
    defparam shift_srl_16_6_LC_5_12_6.SEQ_MODE=4'b1000;
    defparam shift_srl_16_6_LC_5_12_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_16_6_LC_5_12_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51574),
            .lcout(shift_srl_16Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92976),
            .ce(N__51550),
            .sr(_gnd_net_));
    defparam shift_srl_16_9_LC_5_12_7.C_ON=1'b0;
    defparam shift_srl_16_9_LC_5_12_7.SEQ_MODE=4'b1000;
    defparam shift_srl_16_9_LC_5_12_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_16_9_LC_5_12_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51562),
            .lcout(shift_srl_16Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92976),
            .ce(N__51550),
            .sr(_gnd_net_));
    defparam shift_srl_20_3_LC_5_13_0.C_ON=1'b0;
    defparam shift_srl_20_3_LC_5_13_0.SEQ_MODE=4'b1000;
    defparam shift_srl_20_3_LC_5_13_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_20_3_LC_5_13_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51652),
            .lcout(shift_srl_20Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92966),
            .ce(N__51702),
            .sr(_gnd_net_));
    defparam shift_srl_20_1_LC_5_13_1.C_ON=1'b0;
    defparam shift_srl_20_1_LC_5_13_1.SEQ_MODE=4'b1000;
    defparam shift_srl_20_1_LC_5_13_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_20_1_LC_5_13_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51646),
            .lcout(shift_srl_20Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92966),
            .ce(N__51702),
            .sr(_gnd_net_));
    defparam shift_srl_20_2_LC_5_13_2.C_ON=1'b0;
    defparam shift_srl_20_2_LC_5_13_2.SEQ_MODE=4'b1000;
    defparam shift_srl_20_2_LC_5_13_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_20_2_LC_5_13_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51520),
            .lcout(shift_srl_20Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92966),
            .ce(N__51702),
            .sr(_gnd_net_));
    defparam shift_srl_20_0_LC_5_13_3.C_ON=1'b0;
    defparam shift_srl_20_0_LC_5_13_3.SEQ_MODE=4'b1000;
    defparam shift_srl_20_0_LC_5_13_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_20_0_LC_5_13_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51750),
            .lcout(shift_srl_20Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92966),
            .ce(N__51702),
            .sr(_gnd_net_));
    defparam shift_srl_20_4_LC_5_13_4.C_ON=1'b0;
    defparam shift_srl_20_4_LC_5_13_4.SEQ_MODE=4'b1000;
    defparam shift_srl_20_4_LC_5_13_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_20_4_LC_5_13_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51640),
            .lcout(shift_srl_20Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92966),
            .ce(N__51702),
            .sr(_gnd_net_));
    defparam shift_srl_20_5_LC_5_13_5.C_ON=1'b0;
    defparam shift_srl_20_5_LC_5_13_5.SEQ_MODE=4'b1000;
    defparam shift_srl_20_5_LC_5_13_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_20_5_LC_5_13_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51634),
            .lcout(shift_srl_20Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92966),
            .ce(N__51702),
            .sr(_gnd_net_));
    defparam shift_srl_20_6_LC_5_13_6.C_ON=1'b0;
    defparam shift_srl_20_6_LC_5_13_6.SEQ_MODE=4'b1000;
    defparam shift_srl_20_6_LC_5_13_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_20_6_LC_5_13_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51628),
            .lcout(shift_srl_20Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92966),
            .ce(N__51702),
            .sr(_gnd_net_));
    defparam shift_srl_20_7_LC_5_13_7.C_ON=1'b0;
    defparam shift_srl_20_7_LC_5_13_7.SEQ_MODE=4'b1000;
    defparam shift_srl_20_7_LC_5_13_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_20_7_LC_5_13_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51622),
            .lcout(shift_srl_20Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92966),
            .ce(N__51702),
            .sr(_gnd_net_));
    defparam shift_srl_20_10_LC_5_14_0.C_ON=1'b0;
    defparam shift_srl_20_10_LC_5_14_0.SEQ_MODE=4'b1000;
    defparam shift_srl_20_10_LC_5_14_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_20_10_LC_5_14_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51610),
            .lcout(shift_srl_20Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92954),
            .ce(N__51703),
            .sr(_gnd_net_));
    defparam shift_srl_20_11_LC_5_14_1.C_ON=1'b0;
    defparam shift_srl_20_11_LC_5_14_1.SEQ_MODE=4'b1000;
    defparam shift_srl_20_11_LC_5_14_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_20_11_LC_5_14_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51616),
            .lcout(shift_srl_20Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92954),
            .ce(N__51703),
            .sr(_gnd_net_));
    defparam shift_srl_20_13_LC_5_14_2.C_ON=1'b0;
    defparam shift_srl_20_13_LC_5_14_2.SEQ_MODE=4'b1000;
    defparam shift_srl_20_13_LC_5_14_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_20_13_LC_5_14_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51721),
            .lcout(shift_srl_20Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92954),
            .ce(N__51703),
            .sr(_gnd_net_));
    defparam shift_srl_20_9_LC_5_14_3.C_ON=1'b0;
    defparam shift_srl_20_9_LC_5_14_3.SEQ_MODE=4'b1000;
    defparam shift_srl_20_9_LC_5_14_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_20_9_LC_5_14_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51709),
            .lcout(shift_srl_20Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92954),
            .ce(N__51703),
            .sr(_gnd_net_));
    defparam shift_srl_20_14_LC_5_14_4.C_ON=1'b0;
    defparam shift_srl_20_14_LC_5_14_4.SEQ_MODE=4'b1000;
    defparam shift_srl_20_14_LC_5_14_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_20_14_LC_5_14_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51763),
            .lcout(shift_srl_20Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92954),
            .ce(N__51703),
            .sr(_gnd_net_));
    defparam shift_srl_20_15_LC_5_14_5.C_ON=1'b0;
    defparam shift_srl_20_15_LC_5_14_5.SEQ_MODE=4'b1000;
    defparam shift_srl_20_15_LC_5_14_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_20_15_LC_5_14_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51757),
            .lcout(shift_srl_20Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92954),
            .ce(N__51703),
            .sr(_gnd_net_));
    defparam shift_srl_20_12_LC_5_14_6.C_ON=1'b0;
    defparam shift_srl_20_12_LC_5_14_6.SEQ_MODE=4'b1000;
    defparam shift_srl_20_12_LC_5_14_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_20_12_LC_5_14_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51727),
            .lcout(shift_srl_20Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92954),
            .ce(N__51703),
            .sr(_gnd_net_));
    defparam shift_srl_20_8_LC_5_14_7.C_ON=1'b0;
    defparam shift_srl_20_8_LC_5_14_7.SEQ_MODE=4'b1000;
    defparam shift_srl_20_8_LC_5_14_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_20_8_LC_5_14_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51715),
            .lcout(shift_srl_20Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92954),
            .ce(N__51703),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNI2I192_15_LC_5_15_0.C_ON=1'b0;
    defparam shift_srl_0_RNI2I192_15_LC_5_15_0.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNI2I192_15_LC_5_15_0.LUT_INIT=16'b1100110000000000;
    LogicCell40 shift_srl_0_RNI2I192_15_LC_5_15_0 (
            .in0(_gnd_net_),
            .in1(N__51691),
            .in2(_gnd_net_),
            .in3(N__90421),
            .lcout(clk_en_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_8_0_LC_5_15_1.C_ON=1'b0;
    defparam shift_srl_8_0_LC_5_15_1.SEQ_MODE=4'b1000;
    defparam shift_srl_8_0_LC_5_15_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_8_0_LC_5_15_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53826),
            .lcout(shift_srl_8Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92944),
            .ce(N__52829),
            .sr(_gnd_net_));
    defparam shift_srl_8_1_LC_5_15_2.C_ON=1'b0;
    defparam shift_srl_8_1_LC_5_15_2.SEQ_MODE=4'b1000;
    defparam shift_srl_8_1_LC_5_15_2.LUT_INIT=16'b1100110011001100;
    LogicCell40 shift_srl_8_1_LC_5_15_2 (
            .in0(_gnd_net_),
            .in1(N__51670),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_8Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92944),
            .ce(N__52829),
            .sr(_gnd_net_));
    defparam shift_srl_8_2_LC_5_15_3.C_ON=1'b0;
    defparam shift_srl_8_2_LC_5_15_3.SEQ_MODE=4'b1000;
    defparam shift_srl_8_2_LC_5_15_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_8_2_LC_5_15_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51664),
            .lcout(shift_srl_8Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92944),
            .ce(N__52829),
            .sr(_gnd_net_));
    defparam shift_srl_8_3_LC_5_15_4.C_ON=1'b0;
    defparam shift_srl_8_3_LC_5_15_4.SEQ_MODE=4'b1000;
    defparam shift_srl_8_3_LC_5_15_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_8_3_LC_5_15_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51658),
            .lcout(shift_srl_8Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92944),
            .ce(N__52829),
            .sr(_gnd_net_));
    defparam shift_srl_8_4_LC_5_15_5.C_ON=1'b0;
    defparam shift_srl_8_4_LC_5_15_5.SEQ_MODE=4'b1000;
    defparam shift_srl_8_4_LC_5_15_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_8_4_LC_5_15_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51811),
            .lcout(shift_srl_8Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92944),
            .ce(N__52829),
            .sr(_gnd_net_));
    defparam shift_srl_8_7_LC_5_16_0.C_ON=1'b0;
    defparam shift_srl_8_7_LC_5_16_0.SEQ_MODE=4'b1000;
    defparam shift_srl_8_7_LC_5_16_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_8_7_LC_5_16_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51805),
            .lcout(shift_srl_8Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92936),
            .ce(N__52836),
            .sr(_gnd_net_));
    defparam shift_srl_8_6_LC_5_16_1.C_ON=1'b0;
    defparam shift_srl_8_6_LC_5_16_1.SEQ_MODE=4'b1000;
    defparam shift_srl_8_6_LC_5_16_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_8_6_LC_5_16_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51793),
            .lcout(shift_srl_8Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92936),
            .ce(N__52836),
            .sr(_gnd_net_));
    defparam shift_srl_8_5_LC_5_16_4.C_ON=1'b0;
    defparam shift_srl_8_5_LC_5_16_4.SEQ_MODE=4'b1000;
    defparam shift_srl_8_5_LC_5_16_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_8_5_LC_5_16_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51799),
            .lcout(shift_srl_8Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92936),
            .ce(N__52836),
            .sr(_gnd_net_));
    defparam shift_srl_8_8_LC_5_16_5.C_ON=1'b0;
    defparam shift_srl_8_8_LC_5_16_5.SEQ_MODE=4'b1000;
    defparam shift_srl_8_8_LC_5_16_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_8_8_LC_5_16_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51787),
            .lcout(shift_srl_8Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92936),
            .ce(N__52836),
            .sr(_gnd_net_));
    defparam shift_srl_133_4_LC_5_17_0.C_ON=1'b0;
    defparam shift_srl_133_4_LC_5_17_0.SEQ_MODE=4'b1000;
    defparam shift_srl_133_4_LC_5_17_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_133_4_LC_5_17_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55393),
            .lcout(shift_srl_133Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92921),
            .ce(N__55376),
            .sr(_gnd_net_));
    defparam shift_srl_133_5_LC_5_17_1.C_ON=1'b0;
    defparam shift_srl_133_5_LC_5_17_1.SEQ_MODE=4'b1000;
    defparam shift_srl_133_5_LC_5_17_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_133_5_LC_5_17_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51781),
            .lcout(shift_srl_133Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92921),
            .ce(N__55376),
            .sr(_gnd_net_));
    defparam shift_srl_133_6_LC_5_17_2.C_ON=1'b0;
    defparam shift_srl_133_6_LC_5_17_2.SEQ_MODE=4'b1000;
    defparam shift_srl_133_6_LC_5_17_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_133_6_LC_5_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51775),
            .lcout(shift_srl_133Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92921),
            .ce(N__55376),
            .sr(_gnd_net_));
    defparam shift_srl_133_7_LC_5_17_3.C_ON=1'b0;
    defparam shift_srl_133_7_LC_5_17_3.SEQ_MODE=4'b1000;
    defparam shift_srl_133_7_LC_5_17_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_133_7_LC_5_17_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51769),
            .lcout(shift_srl_133Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92921),
            .ce(N__55376),
            .sr(_gnd_net_));
    defparam shift_srl_133_8_LC_5_17_4.C_ON=1'b0;
    defparam shift_srl_133_8_LC_5_17_4.SEQ_MODE=4'b1000;
    defparam shift_srl_133_8_LC_5_17_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_133_8_LC_5_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51865),
            .lcout(shift_srl_133Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92921),
            .ce(N__55376),
            .sr(_gnd_net_));
    defparam shift_srl_133_10_LC_5_17_6.C_ON=1'b0;
    defparam shift_srl_133_10_LC_5_17_6.SEQ_MODE=4'b1000;
    defparam shift_srl_133_10_LC_5_17_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_133_10_LC_5_17_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51847),
            .lcout(shift_srl_133Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92921),
            .ce(N__55376),
            .sr(_gnd_net_));
    defparam shift_srl_133_9_LC_5_17_7.C_ON=1'b0;
    defparam shift_srl_133_9_LC_5_17_7.SEQ_MODE=4'b1000;
    defparam shift_srl_133_9_LC_5_17_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_133_9_LC_5_17_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51853),
            .lcout(shift_srl_133Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92921),
            .ce(N__55376),
            .sr(_gnd_net_));
    defparam shift_srl_132_10_LC_5_18_0.C_ON=1'b0;
    defparam shift_srl_132_10_LC_5_18_0.SEQ_MODE=4'b1000;
    defparam shift_srl_132_10_LC_5_18_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_132_10_LC_5_18_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51817),
            .lcout(shift_srl_132Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92937),
            .ce(N__52954),
            .sr(_gnd_net_));
    defparam shift_srl_132_11_LC_5_18_1.C_ON=1'b0;
    defparam shift_srl_132_11_LC_5_18_1.SEQ_MODE=4'b1000;
    defparam shift_srl_132_11_LC_5_18_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_132_11_LC_5_18_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51841),
            .lcout(shift_srl_132Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92937),
            .ce(N__52954),
            .sr(_gnd_net_));
    defparam shift_srl_132_12_LC_5_18_2.C_ON=1'b0;
    defparam shift_srl_132_12_LC_5_18_2.SEQ_MODE=4'b1000;
    defparam shift_srl_132_12_LC_5_18_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_132_12_LC_5_18_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51835),
            .lcout(shift_srl_132Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92937),
            .ce(N__52954),
            .sr(_gnd_net_));
    defparam shift_srl_132_13_LC_5_18_3.C_ON=1'b0;
    defparam shift_srl_132_13_LC_5_18_3.SEQ_MODE=4'b1000;
    defparam shift_srl_132_13_LC_5_18_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_132_13_LC_5_18_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51829),
            .lcout(shift_srl_132Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92937),
            .ce(N__52954),
            .sr(_gnd_net_));
    defparam shift_srl_132_14_LC_5_18_4.C_ON=1'b0;
    defparam shift_srl_132_14_LC_5_18_4.SEQ_MODE=4'b1000;
    defparam shift_srl_132_14_LC_5_18_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_132_14_LC_5_18_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51823),
            .lcout(shift_srl_132Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92937),
            .ce(N__52954),
            .sr(_gnd_net_));
    defparam shift_srl_132_9_LC_5_18_5.C_ON=1'b0;
    defparam shift_srl_132_9_LC_5_18_5.SEQ_MODE=4'b1000;
    defparam shift_srl_132_9_LC_5_18_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_132_9_LC_5_18_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51949),
            .lcout(shift_srl_132Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92937),
            .ce(N__52954),
            .sr(_gnd_net_));
    defparam shift_srl_132_8_LC_5_18_6.C_ON=1'b0;
    defparam shift_srl_132_8_LC_5_18_6.SEQ_MODE=4'b1000;
    defparam shift_srl_132_8_LC_5_18_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_132_8_LC_5_18_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52969),
            .lcout(shift_srl_132Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92937),
            .ce(N__52954),
            .sr(_gnd_net_));
    defparam shift_srl_131_10_LC_5_19_0.C_ON=1'b0;
    defparam shift_srl_131_10_LC_5_19_0.SEQ_MODE=4'b1000;
    defparam shift_srl_131_10_LC_5_19_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_131_10_LC_5_19_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51907),
            .lcout(shift_srl_131Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92945),
            .ce(N__51889),
            .sr(_gnd_net_));
    defparam shift_srl_131_11_LC_5_19_1.C_ON=1'b0;
    defparam shift_srl_131_11_LC_5_19_1.SEQ_MODE=4'b1000;
    defparam shift_srl_131_11_LC_5_19_1.LUT_INIT=16'b1100110011001100;
    LogicCell40 shift_srl_131_11_LC_5_19_1 (
            .in0(_gnd_net_),
            .in1(N__51943),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_131Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92945),
            .ce(N__51889),
            .sr(_gnd_net_));
    defparam shift_srl_131_12_LC_5_19_2.C_ON=1'b0;
    defparam shift_srl_131_12_LC_5_19_2.SEQ_MODE=4'b1000;
    defparam shift_srl_131_12_LC_5_19_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_131_12_LC_5_19_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51937),
            .lcout(shift_srl_131Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92945),
            .ce(N__51889),
            .sr(_gnd_net_));
    defparam shift_srl_131_13_LC_5_19_3.C_ON=1'b0;
    defparam shift_srl_131_13_LC_5_19_3.SEQ_MODE=4'b1000;
    defparam shift_srl_131_13_LC_5_19_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_131_13_LC_5_19_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51931),
            .lcout(shift_srl_131Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92945),
            .ce(N__51889),
            .sr(_gnd_net_));
    defparam shift_srl_131_14_LC_5_19_4.C_ON=1'b0;
    defparam shift_srl_131_14_LC_5_19_4.SEQ_MODE=4'b1000;
    defparam shift_srl_131_14_LC_5_19_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_131_14_LC_5_19_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51925),
            .lcout(shift_srl_131Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92945),
            .ce(N__51889),
            .sr(_gnd_net_));
    defparam shift_srl_131_15_LC_5_19_5.C_ON=1'b0;
    defparam shift_srl_131_15_LC_5_19_5.SEQ_MODE=4'b1000;
    defparam shift_srl_131_15_LC_5_19_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_131_15_LC_5_19_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51919),
            .lcout(shift_srl_131Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92945),
            .ce(N__51889),
            .sr(_gnd_net_));
    defparam shift_srl_131_9_LC_5_19_6.C_ON=1'b0;
    defparam shift_srl_131_9_LC_5_19_6.SEQ_MODE=4'b1000;
    defparam shift_srl_131_9_LC_5_19_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_131_9_LC_5_19_6 (
            .in0(N__51913),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_131Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92945),
            .ce(N__51889),
            .sr(_gnd_net_));
    defparam shift_srl_131_1_LC_5_19_7.C_ON=1'b0;
    defparam shift_srl_131_1_LC_5_19_7.SEQ_MODE=4'b1000;
    defparam shift_srl_131_1_LC_5_19_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_131_1_LC_5_19_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51901),
            .lcout(shift_srl_131Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92945),
            .ce(N__51889),
            .sr(_gnd_net_));
    defparam shift_srl_134_0_LC_5_20_3.C_ON=1'b0;
    defparam shift_srl_134_0_LC_5_20_3.SEQ_MODE=4'b1000;
    defparam shift_srl_134_0_LC_5_20_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_134_0_LC_5_20_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52016),
            .lcout(shift_srl_134Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92955),
            .ce(N__53004),
            .sr(_gnd_net_));
    defparam shift_srl_133_RNI183N_15_LC_5_21_0.C_ON=1'b0;
    defparam shift_srl_133_RNI183N_15_LC_5_21_0.SEQ_MODE=4'b0000;
    defparam shift_srl_133_RNI183N_15_LC_5_21_0.LUT_INIT=16'b1100110000000000;
    LogicCell40 shift_srl_133_RNI183N_15_LC_5_21_0 (
            .in0(_gnd_net_),
            .in1(N__66241),
            .in2(_gnd_net_),
            .in3(N__52936),
            .lcout(),
            .ltout(g0_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_129_RNIIUCQ1_15_LC_5_21_1.C_ON=1'b0;
    defparam shift_srl_129_RNIIUCQ1_15_LC_5_21_1.SEQ_MODE=4'b0000;
    defparam shift_srl_129_RNIIUCQ1_15_LC_5_21_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_129_RNIIUCQ1_15_LC_5_21_1 (
            .in0(N__54502),
            .in1(N__91269),
            .in2(N__51976),
            .in3(N__54231),
            .lcout(),
            .ltout(g0_13_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_132_RNIQBOL11_15_LC_5_21_2.C_ON=1'b0;
    defparam shift_srl_132_RNIQBOL11_15_LC_5_21_2.SEQ_MODE=4'b0000;
    defparam shift_srl_132_RNIQBOL11_15_LC_5_21_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_132_RNIQBOL11_15_LC_5_21_2 (
            .in0(N__51961),
            .in1(N__51967),
            .in2(N__51973),
            .in3(N__61998),
            .lcout(clk_en_134),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_114_RNI00Q41_15_LC_5_21_3.C_ON=1'b0;
    defparam shift_srl_114_RNI00Q41_15_LC_5_21_3.SEQ_MODE=4'b0000;
    defparam shift_srl_114_RNI00Q41_15_LC_5_21_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_114_RNI00Q41_15_LC_5_21_3 (
            .in0(N__63813),
            .in1(N__58927),
            .in2(N__60535),
            .in3(N__60777),
            .lcout(),
            .ltout(g0_10_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_114_RNIEFPU2_15_LC_5_21_4.C_ON=1'b0;
    defparam shift_srl_114_RNIEFPU2_15_LC_5_21_4.SEQ_MODE=4'b0000;
    defparam shift_srl_114_RNIEFPU2_15_LC_5_21_4.LUT_INIT=16'b1100000000000000;
    LogicCell40 shift_srl_114_RNIEFPU2_15_LC_5_21_4 (
            .in0(_gnd_net_),
            .in1(N__65740),
            .in2(N__51970),
            .in3(N__65362),
            .lcout(g0_14_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_132_RNI8L5Q_15_LC_5_21_5.C_ON=1'b0;
    defparam shift_srl_132_RNI8L5Q_15_LC_5_21_5.SEQ_MODE=4'b0000;
    defparam shift_srl_132_RNI8L5Q_15_LC_5_21_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_132_RNI8L5Q_15_LC_5_21_5 (
            .in0(N__58801),
            .in1(N__54361),
            .in2(N__65572),
            .in3(N__54306),
            .lcout(g0_12_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_135_5_LC_5_22_0.C_ON=1'b0;
    defparam shift_srl_135_5_LC_5_22_0.SEQ_MODE=4'b1000;
    defparam shift_srl_135_5_LC_5_22_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_135_5_LC_5_22_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53212),
            .lcout(shift_srl_135Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92977),
            .ce(N__53176),
            .sr(_gnd_net_));
    defparam shift_srl_135_11_LC_5_22_1.C_ON=1'b0;
    defparam shift_srl_135_11_LC_5_22_1.SEQ_MODE=4'b1000;
    defparam shift_srl_135_11_LC_5_22_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_135_11_LC_5_22_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52033),
            .lcout(shift_srl_135Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92977),
            .ce(N__53176),
            .sr(_gnd_net_));
    defparam shift_srl_135_12_LC_5_22_2.C_ON=1'b0;
    defparam shift_srl_135_12_LC_5_22_2.SEQ_MODE=4'b1000;
    defparam shift_srl_135_12_LC_5_22_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_135_12_LC_5_22_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51955),
            .lcout(shift_srl_135Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92977),
            .ce(N__53176),
            .sr(_gnd_net_));
    defparam shift_srl_135_13_LC_5_22_3.C_ON=1'b0;
    defparam shift_srl_135_13_LC_5_22_3.SEQ_MODE=4'b1000;
    defparam shift_srl_135_13_LC_5_22_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_135_13_LC_5_22_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52057),
            .lcout(shift_srl_135Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92977),
            .ce(N__53176),
            .sr(_gnd_net_));
    defparam shift_srl_135_14_LC_5_22_4.C_ON=1'b0;
    defparam shift_srl_135_14_LC_5_22_4.SEQ_MODE=4'b1000;
    defparam shift_srl_135_14_LC_5_22_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_135_14_LC_5_22_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52051),
            .lcout(shift_srl_135Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92977),
            .ce(N__53176),
            .sr(_gnd_net_));
    defparam shift_srl_135_15_LC_5_22_5.C_ON=1'b0;
    defparam shift_srl_135_15_LC_5_22_5.SEQ_MODE=4'b1000;
    defparam shift_srl_135_15_LC_5_22_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_135_15_LC_5_22_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52045),
            .lcout(shift_srl_135Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92977),
            .ce(N__53176),
            .sr(_gnd_net_));
    defparam shift_srl_135_9_LC_5_22_6.C_ON=1'b0;
    defparam shift_srl_135_9_LC_5_22_6.SEQ_MODE=4'b1000;
    defparam shift_srl_135_9_LC_5_22_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_135_9_LC_5_22_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53110),
            .lcout(shift_srl_135Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92977),
            .ce(N__53176),
            .sr(_gnd_net_));
    defparam shift_srl_135_10_LC_5_22_7.C_ON=1'b0;
    defparam shift_srl_135_10_LC_5_22_7.SEQ_MODE=4'b1000;
    defparam shift_srl_135_10_LC_5_22_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_135_10_LC_5_22_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52039),
            .lcout(shift_srl_135Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92977),
            .ce(N__53176),
            .sr(_gnd_net_));
    defparam shift_srl_118_RNI944G_15_LC_5_23_2.C_ON=1'b0;
    defparam shift_srl_118_RNI944G_15_LC_5_23_2.SEQ_MODE=4'b0000;
    defparam shift_srl_118_RNI944G_15_LC_5_23_2.LUT_INIT=16'b1100110000000000;
    LogicCell40 shift_srl_118_RNI944G_15_LC_5_23_2 (
            .in0(_gnd_net_),
            .in1(N__60332),
            .in2(_gnd_net_),
            .in3(N__66443),
            .lcout(g0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_116_8_LC_5_24_0.C_ON=1'b0;
    defparam shift_srl_116_8_LC_5_24_0.SEQ_MODE=4'b1000;
    defparam shift_srl_116_8_LC_5_24_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_116_8_LC_5_24_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53266),
            .lcout(shift_srl_116Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93004),
            .ce(N__54577),
            .sr(_gnd_net_));
    defparam shift_srl_2_10_LC_6_7_0.C_ON=1'b0;
    defparam shift_srl_2_10_LC_6_7_0.SEQ_MODE=4'b1000;
    defparam shift_srl_2_10_LC_6_7_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_2_10_LC_6_7_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52087),
            .lcout(shift_srl_2Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93064),
            .ce(N__53333),
            .sr(_gnd_net_));
    defparam shift_srl_2_11_LC_6_7_1.C_ON=1'b0;
    defparam shift_srl_2_11_LC_6_7_1.SEQ_MODE=4'b1000;
    defparam shift_srl_2_11_LC_6_7_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_2_11_LC_6_7_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52027),
            .lcout(shift_srl_2Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93064),
            .ce(N__53333),
            .sr(_gnd_net_));
    defparam shift_srl_2_12_LC_6_7_2.C_ON=1'b0;
    defparam shift_srl_2_12_LC_6_7_2.SEQ_MODE=4'b1000;
    defparam shift_srl_2_12_LC_6_7_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_2_12_LC_6_7_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52105),
            .lcout(shift_srl_2Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93064),
            .ce(N__53333),
            .sr(_gnd_net_));
    defparam shift_srl_2_13_LC_6_7_3.C_ON=1'b0;
    defparam shift_srl_2_13_LC_6_7_3.SEQ_MODE=4'b1000;
    defparam shift_srl_2_13_LC_6_7_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_2_13_LC_6_7_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52099),
            .lcout(shift_srl_2Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93064),
            .ce(N__53333),
            .sr(_gnd_net_));
    defparam shift_srl_2_8_LC_6_7_4.C_ON=1'b0;
    defparam shift_srl_2_8_LC_6_7_4.SEQ_MODE=4'b1000;
    defparam shift_srl_2_8_LC_6_7_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_2_8_LC_6_7_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52213),
            .lcout(shift_srl_2Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93064),
            .ce(N__53333),
            .sr(_gnd_net_));
    defparam shift_srl_2_9_LC_6_7_5.C_ON=1'b0;
    defparam shift_srl_2_9_LC_6_7_5.SEQ_MODE=4'b1000;
    defparam shift_srl_2_9_LC_6_7_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_2_9_LC_6_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52093),
            .lcout(shift_srl_2Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93064),
            .ce(N__53333),
            .sr(_gnd_net_));
    defparam shift_srl_2_3_LC_6_7_6.C_ON=1'b0;
    defparam shift_srl_2_3_LC_6_7_6.SEQ_MODE=4'b1000;
    defparam shift_srl_2_3_LC_6_7_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_2_3_LC_6_7_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52081),
            .lcout(shift_srl_2Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93064),
            .ce(N__53333),
            .sr(_gnd_net_));
    defparam shift_srl_2_2_LC_6_7_7.C_ON=1'b0;
    defparam shift_srl_2_2_LC_6_7_7.SEQ_MODE=4'b1000;
    defparam shift_srl_2_2_LC_6_7_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_2_2_LC_6_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52069),
            .lcout(shift_srl_2Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93064),
            .ce(N__53333),
            .sr(_gnd_net_));
    defparam shift_srl_2_0_LC_6_8_0.C_ON=1'b0;
    defparam shift_srl_2_0_LC_6_8_0.SEQ_MODE=4'b1000;
    defparam shift_srl_2_0_LC_6_8_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_2_0_LC_6_8_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52300),
            .lcout(shift_srl_2Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93048),
            .ce(N__53338),
            .sr(_gnd_net_));
    defparam shift_srl_2_1_LC_6_8_1.C_ON=1'b0;
    defparam shift_srl_2_1_LC_6_8_1.SEQ_MODE=4'b1000;
    defparam shift_srl_2_1_LC_6_8_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_2_1_LC_6_8_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52075),
            .lcout(shift_srl_2Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93048),
            .ce(N__53338),
            .sr(_gnd_net_));
    defparam shift_srl_2_14_LC_6_8_2.C_ON=1'b0;
    defparam shift_srl_2_14_LC_6_8_2.SEQ_MODE=4'b1000;
    defparam shift_srl_2_14_LC_6_8_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_2_14_LC_6_8_2 (
            .in0(N__52063),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_2Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93048),
            .ce(N__53338),
            .sr(_gnd_net_));
    defparam shift_srl_2_5_LC_6_8_3.C_ON=1'b0;
    defparam shift_srl_2_5_LC_6_8_3.SEQ_MODE=4'b1000;
    defparam shift_srl_2_5_LC_6_8_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_2_5_LC_6_8_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52231),
            .lcout(shift_srl_2Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93048),
            .ce(N__53338),
            .sr(_gnd_net_));
    defparam shift_srl_2_4_LC_6_8_4.C_ON=1'b0;
    defparam shift_srl_2_4_LC_6_8_4.SEQ_MODE=4'b1000;
    defparam shift_srl_2_4_LC_6_8_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_2_4_LC_6_8_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52237),
            .lcout(shift_srl_2Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93048),
            .ce(N__53338),
            .sr(_gnd_net_));
    defparam shift_srl_2_6_LC_6_8_6.C_ON=1'b0;
    defparam shift_srl_2_6_LC_6_8_6.SEQ_MODE=4'b1000;
    defparam shift_srl_2_6_LC_6_8_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_2_6_LC_6_8_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52225),
            .lcout(shift_srl_2Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93048),
            .ce(N__53338),
            .sr(_gnd_net_));
    defparam shift_srl_2_7_LC_6_8_7.C_ON=1'b0;
    defparam shift_srl_2_7_LC_6_8_7.SEQ_MODE=4'b1000;
    defparam shift_srl_2_7_LC_6_8_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_2_7_LC_6_8_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52219),
            .lcout(shift_srl_2Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93048),
            .ce(N__53338),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNI9AET5_15_LC_6_9_0.C_ON=1'b0;
    defparam shift_srl_0_RNI9AET5_15_LC_6_9_0.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNI9AET5_15_LC_6_9_0.LUT_INIT=16'b1100110000000000;
    LogicCell40 shift_srl_0_RNI9AET5_15_LC_6_9_0 (
            .in0(_gnd_net_),
            .in1(N__90210),
            .in2(_gnd_net_),
            .in3(N__52130),
            .lcout(N_701),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_10_RNIQHCJ1_15_LC_6_9_1.C_ON=1'b0;
    defparam shift_srl_10_RNIQHCJ1_15_LC_6_9_1.SEQ_MODE=4'b0000;
    defparam shift_srl_10_RNIQHCJ1_15_LC_6_9_1.LUT_INIT=16'b0000000010001000;
    LogicCell40 shift_srl_10_RNIQHCJ1_15_LC_6_9_1 (
            .in0(N__53805),
            .in1(N__55719),
            .in2(_gnd_net_),
            .in3(N__53676),
            .lcout(),
            .ltout(shift_srl_10_RNIQHCJ1Z0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_10_RNIEUJS5_15_LC_6_9_2.C_ON=1'b0;
    defparam shift_srl_10_RNIEUJS5_15_LC_6_9_2.SEQ_MODE=4'b0000;
    defparam shift_srl_10_RNIEUJS5_15_LC_6_9_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_10_RNIEUJS5_15_LC_6_9_2 (
            .in0(N__52347),
            .in1(N__69272),
            .in2(N__52150),
            .in3(N__69231),
            .lcout(rco_c_21),
            .ltout(rco_c_21_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_22_RNIO6AV5_15_LC_6_9_3.C_ON=1'b0;
    defparam shift_srl_22_RNIO6AV5_15_LC_6_9_3.SEQ_MODE=4'b0000;
    defparam shift_srl_22_RNIO6AV5_15_LC_6_9_3.LUT_INIT=16'b1010000000000000;
    LogicCell40 shift_srl_22_RNIO6AV5_15_LC_6_9_3 (
            .in0(N__90211),
            .in1(_gnd_net_),
            .in2(N__52114),
            .in3(N__53419),
            .lcout(N_702),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_2_15_LC_6_9_4.C_ON=1'b0;
    defparam shift_srl_2_15_LC_6_9_4.SEQ_MODE=4'b1000;
    defparam shift_srl_2_15_LC_6_9_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_2_15_LC_6_9_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52111),
            .lcout(shift_srl_2Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93033),
            .ce(N__53337),
            .sr(_gnd_net_));
    defparam shift_srl_2_RNI76AR_15_LC_6_9_5.C_ON=1'b0;
    defparam shift_srl_2_RNI76AR_15_LC_6_9_5.SEQ_MODE=4'b0000;
    defparam shift_srl_2_RNI76AR_15_LC_6_9_5.LUT_INIT=16'b0111011111111111;
    LogicCell40 shift_srl_2_RNI76AR_15_LC_6_9_5 (
            .in0(N__57219),
            .in1(N__52298),
            .in2(_gnd_net_),
            .in3(N__57151),
            .lcout(N_453),
            .ltout(N_453_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_10_RNIQH903_15_LC_6_9_6.C_ON=1'b0;
    defparam shift_srl_10_RNIQH903_15_LC_6_9_6.SEQ_MODE=4'b0000;
    defparam shift_srl_10_RNIQH903_15_LC_6_9_6.LUT_INIT=16'b0000100000000000;
    LogicCell40 shift_srl_10_RNIQH903_15_LC_6_9_6 (
            .in0(N__55720),
            .in1(N__52348),
            .in2(N__52330),
            .in3(N__53806),
            .lcout(rco_c_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_2_LC_6_9_7.C_ON=1'b0;
    defparam rco_obuf_RNO_2_LC_6_9_7.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_2_LC_6_9_7.LUT_INIT=16'b1000100000000000;
    LogicCell40 rco_obuf_RNO_2_LC_6_9_7 (
            .in0(N__57218),
            .in1(N__52299),
            .in2(_gnd_net_),
            .in3(N__57152),
            .lcout(N_453_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_23_10_LC_6_10_0.C_ON=1'b0;
    defparam shift_srl_23_10_LC_6_10_0.SEQ_MODE=4'b1000;
    defparam shift_srl_23_10_LC_6_10_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_23_10_LC_6_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52243),
            .lcout(shift_srl_23Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93019),
            .ce(N__53579),
            .sr(_gnd_net_));
    defparam shift_srl_23_11_LC_6_10_1.C_ON=1'b0;
    defparam shift_srl_23_11_LC_6_10_1.SEQ_MODE=4'b1000;
    defparam shift_srl_23_11_LC_6_10_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_23_11_LC_6_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52267),
            .lcout(shift_srl_23Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93019),
            .ce(N__53579),
            .sr(_gnd_net_));
    defparam shift_srl_23_12_LC_6_10_2.C_ON=1'b0;
    defparam shift_srl_23_12_LC_6_10_2.SEQ_MODE=4'b1000;
    defparam shift_srl_23_12_LC_6_10_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_23_12_LC_6_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52261),
            .lcout(shift_srl_23Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93019),
            .ce(N__53579),
            .sr(_gnd_net_));
    defparam shift_srl_23_13_LC_6_10_3.C_ON=1'b0;
    defparam shift_srl_23_13_LC_6_10_3.SEQ_MODE=4'b1000;
    defparam shift_srl_23_13_LC_6_10_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_23_13_LC_6_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52255),
            .lcout(shift_srl_23Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93019),
            .ce(N__53579),
            .sr(_gnd_net_));
    defparam shift_srl_23_14_LC_6_10_4.C_ON=1'b0;
    defparam shift_srl_23_14_LC_6_10_4.SEQ_MODE=4'b1000;
    defparam shift_srl_23_14_LC_6_10_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_23_14_LC_6_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52249),
            .lcout(shift_srl_23Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93019),
            .ce(N__53579),
            .sr(_gnd_net_));
    defparam shift_srl_23_9_LC_6_10_5.C_ON=1'b0;
    defparam shift_srl_23_9_LC_6_10_5.SEQ_MODE=4'b1000;
    defparam shift_srl_23_9_LC_6_10_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_23_9_LC_6_10_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52396),
            .lcout(shift_srl_23Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93019),
            .ce(N__53579),
            .sr(_gnd_net_));
    defparam shift_srl_23_8_LC_6_10_6.C_ON=1'b0;
    defparam shift_srl_23_8_LC_6_10_6.SEQ_MODE=4'b1000;
    defparam shift_srl_23_8_LC_6_10_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_23_8_LC_6_10_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52390),
            .lcout(shift_srl_23Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93019),
            .ce(N__53579),
            .sr(_gnd_net_));
    defparam shift_srl_23_7_LC_6_10_7.C_ON=1'b0;
    defparam shift_srl_23_7_LC_6_10_7.SEQ_MODE=4'b1000;
    defparam shift_srl_23_7_LC_6_10_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_23_7_LC_6_10_7 (
            .in0(N__53587),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_23Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93019),
            .ce(N__53579),
            .sr(_gnd_net_));
    defparam shift_srl_19_10_LC_6_11_0.C_ON=1'b0;
    defparam shift_srl_19_10_LC_6_11_0.SEQ_MODE=4'b1000;
    defparam shift_srl_19_10_LC_6_11_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_19_10_LC_6_11_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52366),
            .lcout(shift_srl_19Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93005),
            .ce(N__52465),
            .sr(_gnd_net_));
    defparam shift_srl_19_11_LC_6_11_1.C_ON=1'b0;
    defparam shift_srl_19_11_LC_6_11_1.SEQ_MODE=4'b1000;
    defparam shift_srl_19_11_LC_6_11_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_19_11_LC_6_11_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52384),
            .lcout(shift_srl_19Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93005),
            .ce(N__52465),
            .sr(_gnd_net_));
    defparam shift_srl_19_6_LC_6_11_2.C_ON=1'b0;
    defparam shift_srl_19_6_LC_6_11_2.SEQ_MODE=4'b1000;
    defparam shift_srl_19_6_LC_6_11_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_19_6_LC_6_11_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52489),
            .lcout(shift_srl_19Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93005),
            .ce(N__52465),
            .sr(_gnd_net_));
    defparam shift_srl_19_7_LC_6_11_3.C_ON=1'b0;
    defparam shift_srl_19_7_LC_6_11_3.SEQ_MODE=4'b1000;
    defparam shift_srl_19_7_LC_6_11_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_19_7_LC_6_11_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52378),
            .lcout(shift_srl_19Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93005),
            .ce(N__52465),
            .sr(_gnd_net_));
    defparam shift_srl_19_14_LC_6_11_4.C_ON=1'b0;
    defparam shift_srl_19_14_LC_6_11_4.SEQ_MODE=4'b1000;
    defparam shift_srl_19_14_LC_6_11_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_19_14_LC_6_11_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52471),
            .lcout(shift_srl_19Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93005),
            .ce(N__52465),
            .sr(_gnd_net_));
    defparam shift_srl_19_15_LC_6_11_5.C_ON=1'b0;
    defparam shift_srl_19_15_LC_6_11_5.SEQ_MODE=4'b1000;
    defparam shift_srl_19_15_LC_6_11_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_19_15_LC_6_11_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52372),
            .lcout(shift_srl_19Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93005),
            .ce(N__52465),
            .sr(_gnd_net_));
    defparam shift_srl_19_9_LC_6_11_6.C_ON=1'b0;
    defparam shift_srl_19_9_LC_6_11_6.SEQ_MODE=4'b1000;
    defparam shift_srl_19_9_LC_6_11_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_19_9_LC_6_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52354),
            .lcout(shift_srl_19Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93005),
            .ce(N__52465),
            .sr(_gnd_net_));
    defparam shift_srl_19_8_LC_6_11_7.C_ON=1'b0;
    defparam shift_srl_19_8_LC_6_11_7.SEQ_MODE=4'b1000;
    defparam shift_srl_19_8_LC_6_11_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_19_8_LC_6_11_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52360),
            .lcout(shift_srl_19Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93005),
            .ce(N__52465),
            .sr(_gnd_net_));
    defparam shift_srl_19_0_LC_6_12_0.C_ON=1'b0;
    defparam shift_srl_19_0_LC_6_12_0.SEQ_MODE=4'b1000;
    defparam shift_srl_19_0_LC_6_12_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_19_0_LC_6_12_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52543),
            .lcout(shift_srl_19Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92990),
            .ce(N__52464),
            .sr(_gnd_net_));
    defparam shift_srl_19_1_LC_6_12_1.C_ON=1'b0;
    defparam shift_srl_19_1_LC_6_12_1.SEQ_MODE=4'b1000;
    defparam shift_srl_19_1_LC_6_12_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_19_1_LC_6_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52519),
            .lcout(shift_srl_19Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92990),
            .ce(N__52464),
            .sr(_gnd_net_));
    defparam shift_srl_19_2_LC_6_12_2.C_ON=1'b0;
    defparam shift_srl_19_2_LC_6_12_2.SEQ_MODE=4'b1000;
    defparam shift_srl_19_2_LC_6_12_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_19_2_LC_6_12_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52513),
            .lcout(shift_srl_19Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92990),
            .ce(N__52464),
            .sr(_gnd_net_));
    defparam shift_srl_19_3_LC_6_12_3.C_ON=1'b0;
    defparam shift_srl_19_3_LC_6_12_3.SEQ_MODE=4'b1000;
    defparam shift_srl_19_3_LC_6_12_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_19_3_LC_6_12_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52507),
            .lcout(shift_srl_19Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92990),
            .ce(N__52464),
            .sr(_gnd_net_));
    defparam shift_srl_19_4_LC_6_12_4.C_ON=1'b0;
    defparam shift_srl_19_4_LC_6_12_4.SEQ_MODE=4'b1000;
    defparam shift_srl_19_4_LC_6_12_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_19_4_LC_6_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52501),
            .lcout(shift_srl_19Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92990),
            .ce(N__52464),
            .sr(_gnd_net_));
    defparam shift_srl_19_5_LC_6_12_5.C_ON=1'b0;
    defparam shift_srl_19_5_LC_6_12_5.SEQ_MODE=4'b1000;
    defparam shift_srl_19_5_LC_6_12_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_19_5_LC_6_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52495),
            .lcout(shift_srl_19Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92990),
            .ce(N__52464),
            .sr(_gnd_net_));
    defparam shift_srl_19_12_LC_6_12_6.C_ON=1'b0;
    defparam shift_srl_19_12_LC_6_12_6.SEQ_MODE=4'b1000;
    defparam shift_srl_19_12_LC_6_12_6.LUT_INIT=16'b1100110011001100;
    LogicCell40 shift_srl_19_12_LC_6_12_6 (
            .in0(_gnd_net_),
            .in1(N__52483),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_19Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92990),
            .ce(N__52464),
            .sr(_gnd_net_));
    defparam shift_srl_19_13_LC_6_12_7.C_ON=1'b0;
    defparam shift_srl_19_13_LC_6_12_7.SEQ_MODE=4'b1000;
    defparam shift_srl_19_13_LC_6_12_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_19_13_LC_6_12_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52477),
            .lcout(shift_srl_19Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92990),
            .ce(N__52464),
            .sr(_gnd_net_));
    defparam shift_srl_17_0_LC_6_13_0.C_ON=1'b0;
    defparam shift_srl_17_0_LC_6_13_0.SEQ_MODE=4'b1000;
    defparam shift_srl_17_0_LC_6_13_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_17_0_LC_6_13_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52441),
            .lcout(shift_srl_17Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92978),
            .ce(N__52677),
            .sr(_gnd_net_));
    defparam shift_srl_17_1_LC_6_13_1.C_ON=1'b0;
    defparam shift_srl_17_1_LC_6_13_1.SEQ_MODE=4'b1000;
    defparam shift_srl_17_1_LC_6_13_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_17_1_LC_6_13_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52609),
            .lcout(shift_srl_17Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92978),
            .ce(N__52677),
            .sr(_gnd_net_));
    defparam shift_srl_17_2_LC_6_13_2.C_ON=1'b0;
    defparam shift_srl_17_2_LC_6_13_2.SEQ_MODE=4'b1000;
    defparam shift_srl_17_2_LC_6_13_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_17_2_LC_6_13_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52603),
            .lcout(shift_srl_17Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92978),
            .ce(N__52677),
            .sr(_gnd_net_));
    defparam shift_srl_17_3_LC_6_13_3.C_ON=1'b0;
    defparam shift_srl_17_3_LC_6_13_3.SEQ_MODE=4'b1000;
    defparam shift_srl_17_3_LC_6_13_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_17_3_LC_6_13_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52597),
            .lcout(shift_srl_17Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92978),
            .ce(N__52677),
            .sr(_gnd_net_));
    defparam shift_srl_17_4_LC_6_13_4.C_ON=1'b0;
    defparam shift_srl_17_4_LC_6_13_4.SEQ_MODE=4'b1000;
    defparam shift_srl_17_4_LC_6_13_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_17_4_LC_6_13_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52591),
            .lcout(shift_srl_17Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92978),
            .ce(N__52677),
            .sr(_gnd_net_));
    defparam shift_srl_17_5_LC_6_13_5.C_ON=1'b0;
    defparam shift_srl_17_5_LC_6_13_5.SEQ_MODE=4'b1000;
    defparam shift_srl_17_5_LC_6_13_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_17_5_LC_6_13_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52585),
            .lcout(shift_srl_17Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92978),
            .ce(N__52677),
            .sr(_gnd_net_));
    defparam shift_srl_17_6_LC_6_13_6.C_ON=1'b0;
    defparam shift_srl_17_6_LC_6_13_6.SEQ_MODE=4'b1000;
    defparam shift_srl_17_6_LC_6_13_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_17_6_LC_6_13_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52579),
            .lcout(shift_srl_17Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92978),
            .ce(N__52677),
            .sr(_gnd_net_));
    defparam shift_srl_17_7_LC_6_13_7.C_ON=1'b0;
    defparam shift_srl_17_7_LC_6_13_7.SEQ_MODE=4'b1000;
    defparam shift_srl_17_7_LC_6_13_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_17_7_LC_6_13_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52573),
            .lcout(shift_srl_17Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92978),
            .ce(N__52677),
            .sr(_gnd_net_));
    defparam shift_srl_17_10_LC_6_14_0.C_ON=1'b0;
    defparam shift_srl_17_10_LC_6_14_0.SEQ_MODE=4'b1000;
    defparam shift_srl_17_10_LC_6_14_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_17_10_LC_6_14_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52696),
            .lcout(shift_srl_17Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92967),
            .ce(N__52678),
            .sr(_gnd_net_));
    defparam shift_srl_17_11_LC_6_14_1.C_ON=1'b0;
    defparam shift_srl_17_11_LC_6_14_1.SEQ_MODE=4'b1000;
    defparam shift_srl_17_11_LC_6_14_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_17_11_LC_6_14_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52567),
            .lcout(shift_srl_17Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92967),
            .ce(N__52678),
            .sr(_gnd_net_));
    defparam shift_srl_17_12_LC_6_14_2.C_ON=1'b0;
    defparam shift_srl_17_12_LC_6_14_2.SEQ_MODE=4'b1000;
    defparam shift_srl_17_12_LC_6_14_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_17_12_LC_6_14_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52726),
            .lcout(shift_srl_17Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92967),
            .ce(N__52678),
            .sr(_gnd_net_));
    defparam shift_srl_17_13_LC_6_14_3.C_ON=1'b0;
    defparam shift_srl_17_13_LC_6_14_3.SEQ_MODE=4'b1000;
    defparam shift_srl_17_13_LC_6_14_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_17_13_LC_6_14_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52720),
            .lcout(shift_srl_17Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92967),
            .ce(N__52678),
            .sr(_gnd_net_));
    defparam shift_srl_17_14_LC_6_14_4.C_ON=1'b0;
    defparam shift_srl_17_14_LC_6_14_4.SEQ_MODE=4'b1000;
    defparam shift_srl_17_14_LC_6_14_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_17_14_LC_6_14_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52714),
            .lcout(shift_srl_17Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92967),
            .ce(N__52678),
            .sr(_gnd_net_));
    defparam shift_srl_17_9_LC_6_14_5.C_ON=1'b0;
    defparam shift_srl_17_9_LC_6_14_5.SEQ_MODE=4'b1000;
    defparam shift_srl_17_9_LC_6_14_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_17_9_LC_6_14_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52684),
            .lcout(shift_srl_17Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92967),
            .ce(N__52678),
            .sr(_gnd_net_));
    defparam shift_srl_17_8_LC_6_14_6.C_ON=1'b0;
    defparam shift_srl_17_8_LC_6_14_6.SEQ_MODE=4'b1000;
    defparam shift_srl_17_8_LC_6_14_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_17_8_LC_6_14_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52690),
            .lcout(shift_srl_17Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92967),
            .ce(N__52678),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNI5UCB2_15_LC_6_15_0.C_ON=1'b0;
    defparam shift_srl_0_RNI5UCB2_15_LC_6_15_0.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNI5UCB2_15_LC_6_15_0.LUT_INIT=16'b1100110000000000;
    LogicCell40 shift_srl_0_RNI5UCB2_15_LC_6_15_0 (
            .in0(_gnd_net_),
            .in1(N__90186),
            .in2(_gnd_net_),
            .in3(N__52642),
            .lcout(clk_en_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_9_0_LC_6_15_1.C_ON=1'b0;
    defparam shift_srl_9_0_LC_6_15_1.SEQ_MODE=4'b1000;
    defparam shift_srl_9_0_LC_6_15_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_9_0_LC_6_15_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53920),
            .lcout(shift_srl_9Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92956),
            .ce(N__54071),
            .sr(_gnd_net_));
    defparam shift_srl_9_1_LC_6_15_2.C_ON=1'b0;
    defparam shift_srl_9_1_LC_6_15_2.SEQ_MODE=4'b1000;
    defparam shift_srl_9_1_LC_6_15_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_9_1_LC_6_15_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52621),
            .lcout(shift_srl_9Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92956),
            .ce(N__54071),
            .sr(_gnd_net_));
    defparam shift_srl_9_2_LC_6_15_3.C_ON=1'b0;
    defparam shift_srl_9_2_LC_6_15_3.SEQ_MODE=4'b1000;
    defparam shift_srl_9_2_LC_6_15_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_9_2_LC_6_15_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52615),
            .lcout(shift_srl_9Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92956),
            .ce(N__54071),
            .sr(_gnd_net_));
    defparam shift_srl_9_3_LC_6_15_4.C_ON=1'b0;
    defparam shift_srl_9_3_LC_6_15_4.SEQ_MODE=4'b1000;
    defparam shift_srl_9_3_LC_6_15_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_9_3_LC_6_15_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52774),
            .lcout(shift_srl_9Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92956),
            .ce(N__54071),
            .sr(_gnd_net_));
    defparam shift_srl_9_4_LC_6_15_5.C_ON=1'b0;
    defparam shift_srl_9_4_LC_6_15_5.SEQ_MODE=4'b1000;
    defparam shift_srl_9_4_LC_6_15_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_9_4_LC_6_15_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52768),
            .lcout(shift_srl_9Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92956),
            .ce(N__54071),
            .sr(_gnd_net_));
    defparam shift_srl_9_5_LC_6_15_6.C_ON=1'b0;
    defparam shift_srl_9_5_LC_6_15_6.SEQ_MODE=4'b1000;
    defparam shift_srl_9_5_LC_6_15_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_9_5_LC_6_15_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52762),
            .lcout(shift_srl_9Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92956),
            .ce(N__54071),
            .sr(_gnd_net_));
    defparam shift_srl_9_6_LC_6_15_7.C_ON=1'b0;
    defparam shift_srl_9_6_LC_6_15_7.SEQ_MODE=4'b1000;
    defparam shift_srl_9_6_LC_6_15_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_9_6_LC_6_15_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52756),
            .lcout(shift_srl_9Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92956),
            .ce(N__54071),
            .sr(_gnd_net_));
    defparam shift_srl_8_10_LC_6_16_0.C_ON=1'b0;
    defparam shift_srl_8_10_LC_6_16_0.SEQ_MODE=4'b1000;
    defparam shift_srl_8_10_LC_6_16_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_8_10_LC_6_16_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52843),
            .lcout(shift_srl_8Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92946),
            .ce(N__52837),
            .sr(_gnd_net_));
    defparam shift_srl_8_11_LC_6_16_1.C_ON=1'b0;
    defparam shift_srl_8_11_LC_6_16_1.SEQ_MODE=4'b1000;
    defparam shift_srl_8_11_LC_6_16_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_8_11_LC_6_16_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52750),
            .lcout(shift_srl_8Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92946),
            .ce(N__52837),
            .sr(_gnd_net_));
    defparam shift_srl_8_12_LC_6_16_2.C_ON=1'b0;
    defparam shift_srl_8_12_LC_6_16_2.SEQ_MODE=4'b1000;
    defparam shift_srl_8_12_LC_6_16_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_8_12_LC_6_16_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52744),
            .lcout(shift_srl_8Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92946),
            .ce(N__52837),
            .sr(_gnd_net_));
    defparam shift_srl_8_13_LC_6_16_3.C_ON=1'b0;
    defparam shift_srl_8_13_LC_6_16_3.SEQ_MODE=4'b1000;
    defparam shift_srl_8_13_LC_6_16_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_8_13_LC_6_16_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52738),
            .lcout(shift_srl_8Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92946),
            .ce(N__52837),
            .sr(_gnd_net_));
    defparam shift_srl_8_14_LC_6_16_4.C_ON=1'b0;
    defparam shift_srl_8_14_LC_6_16_4.SEQ_MODE=4'b1000;
    defparam shift_srl_8_14_LC_6_16_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_8_14_LC_6_16_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52732),
            .lcout(shift_srl_8Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92946),
            .ce(N__52837),
            .sr(_gnd_net_));
    defparam shift_srl_8_15_LC_6_16_5.C_ON=1'b0;
    defparam shift_srl_8_15_LC_6_16_5.SEQ_MODE=4'b1000;
    defparam shift_srl_8_15_LC_6_16_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_8_15_LC_6_16_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52855),
            .lcout(shift_srl_8Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92946),
            .ce(N__52837),
            .sr(_gnd_net_));
    defparam shift_srl_8_9_LC_6_16_6.C_ON=1'b0;
    defparam shift_srl_8_9_LC_6_16_6.SEQ_MODE=4'b1000;
    defparam shift_srl_8_9_LC_6_16_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_8_9_LC_6_16_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52849),
            .lcout(shift_srl_8Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92946),
            .ce(N__52837),
            .sr(_gnd_net_));
    defparam shift_srl_128_8_LC_6_17_0.C_ON=1'b0;
    defparam shift_srl_128_8_LC_6_17_0.SEQ_MODE=4'b1000;
    defparam shift_srl_128_8_LC_6_17_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_128_8_LC_6_17_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52804),
            .lcout(shift_srl_128Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92929),
            .ce(N__56281),
            .sr(_gnd_net_));
    defparam shift_srl_128_7_LC_6_17_1.C_ON=1'b0;
    defparam shift_srl_128_7_LC_6_17_1.SEQ_MODE=4'b1000;
    defparam shift_srl_128_7_LC_6_17_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_128_7_LC_6_17_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54013),
            .lcout(shift_srl_128Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92929),
            .ce(N__56281),
            .sr(_gnd_net_));
    defparam shift_srl_132_0_LC_6_18_0.C_ON=1'b0;
    defparam shift_srl_132_0_LC_6_18_0.SEQ_MODE=4'b1000;
    defparam shift_srl_132_0_LC_6_18_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_132_0_LC_6_18_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54354),
            .lcout(shift_srl_132Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92947),
            .ce(N__52953),
            .sr(_gnd_net_));
    defparam shift_srl_132_1_LC_6_18_1.C_ON=1'b0;
    defparam shift_srl_132_1_LC_6_18_1.SEQ_MODE=4'b1000;
    defparam shift_srl_132_1_LC_6_18_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_132_1_LC_6_18_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52798),
            .lcout(shift_srl_132Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92947),
            .ce(N__52953),
            .sr(_gnd_net_));
    defparam shift_srl_132_2_LC_6_18_2.C_ON=1'b0;
    defparam shift_srl_132_2_LC_6_18_2.SEQ_MODE=4'b1000;
    defparam shift_srl_132_2_LC_6_18_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_132_2_LC_6_18_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52792),
            .lcout(shift_srl_132Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92947),
            .ce(N__52953),
            .sr(_gnd_net_));
    defparam shift_srl_132_3_LC_6_18_3.C_ON=1'b0;
    defparam shift_srl_132_3_LC_6_18_3.SEQ_MODE=4'b1000;
    defparam shift_srl_132_3_LC_6_18_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_132_3_LC_6_18_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52786),
            .lcout(shift_srl_132Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92947),
            .ce(N__52953),
            .sr(_gnd_net_));
    defparam shift_srl_132_4_LC_6_18_4.C_ON=1'b0;
    defparam shift_srl_132_4_LC_6_18_4.SEQ_MODE=4'b1000;
    defparam shift_srl_132_4_LC_6_18_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_132_4_LC_6_18_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52780),
            .lcout(shift_srl_132Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92947),
            .ce(N__52953),
            .sr(_gnd_net_));
    defparam shift_srl_132_5_LC_6_18_5.C_ON=1'b0;
    defparam shift_srl_132_5_LC_6_18_5.SEQ_MODE=4'b1000;
    defparam shift_srl_132_5_LC_6_18_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_132_5_LC_6_18_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52987),
            .lcout(shift_srl_132Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92947),
            .ce(N__52953),
            .sr(_gnd_net_));
    defparam shift_srl_132_6_LC_6_18_6.C_ON=1'b0;
    defparam shift_srl_132_6_LC_6_18_6.SEQ_MODE=4'b1000;
    defparam shift_srl_132_6_LC_6_18_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_132_6_LC_6_18_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52981),
            .lcout(shift_srl_132Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92947),
            .ce(N__52953),
            .sr(_gnd_net_));
    defparam shift_srl_132_7_LC_6_18_7.C_ON=1'b0;
    defparam shift_srl_132_7_LC_6_18_7.SEQ_MODE=4'b1000;
    defparam shift_srl_132_7_LC_6_18_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_132_7_LC_6_18_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52975),
            .lcout(shift_srl_132Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92947),
            .ce(N__52953),
            .sr(_gnd_net_));
    defparam shift_srl_132_15_LC_6_19_0.C_ON=1'b0;
    defparam shift_srl_132_15_LC_6_19_0.SEQ_MODE=4'b1000;
    defparam shift_srl_132_15_LC_6_19_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_132_15_LC_6_19_0 (
            .in0(N__52963),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_132Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92957),
            .ce(N__52952),
            .sr(_gnd_net_));
    defparam shift_srl_131_RNIJ56B1_15_LC_6_19_1.C_ON=1'b0;
    defparam shift_srl_131_RNIJ56B1_15_LC_6_19_1.SEQ_MODE=4'b0000;
    defparam shift_srl_131_RNIJ56B1_15_LC_6_19_1.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_131_RNIJ56B1_15_LC_6_19_1 (
            .in0(N__91214),
            .in1(N__54296),
            .in2(N__65755),
            .in3(N__52929),
            .lcout(),
            .ltout(g0_43_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_129_RNINR8611_15_LC_6_19_2.C_ON=1'b0;
    defparam shift_srl_129_RNINR8611_15_LC_6_19_2.SEQ_MODE=4'b0000;
    defparam shift_srl_129_RNINR8611_15_LC_6_19_2.LUT_INIT=16'b0000100000000000;
    LogicCell40 shift_srl_129_RNINR8611_15_LC_6_19_2 (
            .in0(N__54180),
            .in1(N__90183),
            .in2(N__52957),
            .in3(N__57605),
            .lcout(clk_en_132),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_132_RNI731T_15_LC_6_19_3.C_ON=1'b0;
    defparam shift_srl_132_RNI731T_15_LC_6_19_3.SEQ_MODE=4'b0000;
    defparam shift_srl_132_RNI731T_15_LC_6_19_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_132_RNI731T_15_LC_6_19_3 (
            .in0(N__54340),
            .in1(N__52928),
            .in2(N__54299),
            .in3(N__54179),
            .lcout(),
            .ltout(shift_srl_132_RNI731TZ0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_128_RNIDCG11_15_LC_6_19_4.C_ON=1'b0;
    defparam shift_srl_128_RNIDCG11_15_LC_6_19_4.SEQ_MODE=4'b0000;
    defparam shift_srl_128_RNIDCG11_15_LC_6_19_4.LUT_INIT=16'b1111000010101010;
    LogicCell40 shift_srl_128_RNIDCG11_15_LC_6_19_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__52861),
            .in3(N__91213),
            .lcout(rco_int_0_a3_0_a2_0_132),
            .ltout(rco_int_0_a3_0_a2_0_132_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_144_RNIM9VT1_15_LC_6_19_5.C_ON=1'b0;
    defparam shift_srl_144_RNIM9VT1_15_LC_6_19_5.SEQ_MODE=4'b0000;
    defparam shift_srl_144_RNIM9VT1_15_LC_6_19_5.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_144_RNIM9VT1_15_LC_6_19_5 (
            .in0(N__61820),
            .in1(N__61788),
            .in2(N__52858),
            .in3(N__63763),
            .lcout(rco_int_0_a2_0_a2_1_sx_sx_145),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_144_RNIM9VT1_0_15_LC_6_19_6.C_ON=1'b0;
    defparam shift_srl_144_RNIM9VT1_0_15_LC_6_19_6.SEQ_MODE=4'b0000;
    defparam shift_srl_144_RNIM9VT1_0_15_LC_6_19_6.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_144_RNIM9VT1_0_15_LC_6_19_6 (
            .in0(N__63764),
            .in1(N__62151),
            .in2(N__61792),
            .in3(N__61821),
            .lcout(rco_int_0_a2_0_a2_1_1_sx_145),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_134_1_LC_6_20_1.C_ON=1'b0;
    defparam shift_srl_134_1_LC_6_20_1.SEQ_MODE=4'b1000;
    defparam shift_srl_134_1_LC_6_20_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_134_1_LC_6_20_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53059),
            .lcout(shift_srl_134Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92968),
            .ce(N__53005),
            .sr(_gnd_net_));
    defparam shift_srl_134_2_LC_6_20_2.C_ON=1'b0;
    defparam shift_srl_134_2_LC_6_20_2.SEQ_MODE=4'b1000;
    defparam shift_srl_134_2_LC_6_20_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_134_2_LC_6_20_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53053),
            .lcout(shift_srl_134Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92968),
            .ce(N__53005),
            .sr(_gnd_net_));
    defparam shift_srl_134_3_LC_6_20_3.C_ON=1'b0;
    defparam shift_srl_134_3_LC_6_20_3.SEQ_MODE=4'b1000;
    defparam shift_srl_134_3_LC_6_20_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_134_3_LC_6_20_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53047),
            .lcout(shift_srl_134Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92968),
            .ce(N__53005),
            .sr(_gnd_net_));
    defparam shift_srl_134_4_LC_6_20_4.C_ON=1'b0;
    defparam shift_srl_134_4_LC_6_20_4.SEQ_MODE=4'b1000;
    defparam shift_srl_134_4_LC_6_20_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_134_4_LC_6_20_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53041),
            .lcout(shift_srl_134Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92968),
            .ce(N__53005),
            .sr(_gnd_net_));
    defparam shift_srl_134_5_LC_6_20_5.C_ON=1'b0;
    defparam shift_srl_134_5_LC_6_20_5.SEQ_MODE=4'b1000;
    defparam shift_srl_134_5_LC_6_20_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_134_5_LC_6_20_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53035),
            .lcout(shift_srl_134Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92968),
            .ce(N__53005),
            .sr(_gnd_net_));
    defparam shift_srl_134_6_LC_6_20_6.C_ON=1'b0;
    defparam shift_srl_134_6_LC_6_20_6.SEQ_MODE=4'b1000;
    defparam shift_srl_134_6_LC_6_20_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_134_6_LC_6_20_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53029),
            .lcout(shift_srl_134Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92968),
            .ce(N__53005),
            .sr(_gnd_net_));
    defparam shift_srl_134_7_LC_6_20_7.C_ON=1'b0;
    defparam shift_srl_134_7_LC_6_20_7.SEQ_MODE=4'b1000;
    defparam shift_srl_134_7_LC_6_20_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_134_7_LC_6_20_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53023),
            .lcout(shift_srl_134Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92968),
            .ce(N__53005),
            .sr(_gnd_net_));
    defparam shift_srl_115_RNID47DT_15_LC_6_21_0.C_ON=1'b0;
    defparam shift_srl_115_RNID47DT_15_LC_6_21_0.SEQ_MODE=4'b0000;
    defparam shift_srl_115_RNID47DT_15_LC_6_21_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_115_RNID47DT_15_LC_6_21_0 (
            .in0(N__63811),
            .in1(N__90395),
            .in2(N__62593),
            .in3(N__61999),
            .lcout(clk_en_116),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_115_15_LC_6_21_1.C_ON=1'b0;
    defparam shift_srl_115_15_LC_6_21_1.SEQ_MODE=4'b1000;
    defparam shift_srl_115_15_LC_6_21_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_115_15_LC_6_21_1 (
            .in0(N__64123),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_115Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92979),
            .ce(N__64084),
            .sr(_gnd_net_));
    defparam shift_srl_132_RNIEU7K_15_LC_6_21_2.C_ON=1'b0;
    defparam shift_srl_132_RNIEU7K_15_LC_6_21_2.SEQ_MODE=4'b0000;
    defparam shift_srl_132_RNIEU7K_15_LC_6_21_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_132_RNIEU7K_15_LC_6_21_2 (
            .in0(N__54205),
            .in1(N__54355),
            .in2(N__91268),
            .in3(N__54307),
            .lcout(g0_10_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_145_RNI57NS_15_LC_6_21_3.C_ON=1'b0;
    defparam shift_srl_145_RNI57NS_15_LC_6_21_3.SEQ_MODE=4'b0000;
    defparam shift_srl_145_RNI57NS_15_LC_6_21_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_145_RNI57NS_15_LC_6_21_3 (
            .in0(N__58785),
            .in1(N__63598),
            .in2(N__90517),
            .in3(N__63809),
            .lcout(g0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_116_RNI286T_15_LC_6_21_4.C_ON=1'b0;
    defparam shift_srl_116_RNI286T_15_LC_6_21_4.SEQ_MODE=4'b0000;
    defparam shift_srl_116_RNI286T_15_LC_6_21_4.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_116_RNI286T_15_LC_6_21_4 (
            .in0(N__63810),
            .in1(N__60534),
            .in2(N__60778),
            .in3(N__58786),
            .lcout(),
            .ltout(g0_9_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_116_RNIUVE13_15_LC_6_21_5.C_ON=1'b0;
    defparam shift_srl_116_RNIUVE13_15_LC_6_21_5.SEQ_MODE=4'b0000;
    defparam shift_srl_116_RNIUVE13_15_LC_6_21_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_116_RNIUVE13_15_LC_6_21_5 (
            .in0(N__53140),
            .in1(N__56443),
            .in2(N__53134),
            .in3(N__65568),
            .lcout(g0_16_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_123_RNIEFVP1_15_LC_6_21_6.C_ON=1'b0;
    defparam shift_srl_123_RNIEFVP1_15_LC_6_21_6.SEQ_MODE=4'b0000;
    defparam shift_srl_123_RNIEFVP1_15_LC_6_21_6.LUT_INIT=16'b1100110000000000;
    LogicCell40 shift_srl_123_RNIEFVP1_15_LC_6_21_6 (
            .in0(_gnd_net_),
            .in1(N__65728),
            .in2(_gnd_net_),
            .in3(N__65348),
            .lcout(),
            .ltout(g0_12_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_134_RNIT9P321_15_LC_6_21_7.C_ON=1'b0;
    defparam shift_srl_134_RNIT9P321_15_LC_6_21_7.SEQ_MODE=4'b0000;
    defparam shift_srl_134_RNIT9P321_15_LC_6_21_7.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_134_RNIT9P321_15_LC_6_21_7 (
            .in0(N__62000),
            .in1(N__53131),
            .in2(N__53119),
            .in3(N__53116),
            .lcout(clk_en_135),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_135_8_LC_6_22_0.C_ON=1'b0;
    defparam shift_srl_135_8_LC_6_22_0.SEQ_MODE=4'b1000;
    defparam shift_srl_135_8_LC_6_22_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_135_8_LC_6_22_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53182),
            .lcout(shift_srl_135Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92991),
            .ce(N__53175),
            .sr(_gnd_net_));
    defparam shift_srl_135_0_LC_6_22_1.C_ON=1'b0;
    defparam shift_srl_135_0_LC_6_22_1.SEQ_MODE=4'b1000;
    defparam shift_srl_135_0_LC_6_22_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_135_0_LC_6_22_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53095),
            .lcout(shift_srl_135Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92991),
            .ce(N__53175),
            .sr(_gnd_net_));
    defparam shift_srl_135_2_LC_6_22_2.C_ON=1'b0;
    defparam shift_srl_135_2_LC_6_22_2.SEQ_MODE=4'b1000;
    defparam shift_srl_135_2_LC_6_22_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_135_2_LC_6_22_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53200),
            .lcout(shift_srl_135Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92991),
            .ce(N__53175),
            .sr(_gnd_net_));
    defparam shift_srl_135_3_LC_6_22_3.C_ON=1'b0;
    defparam shift_srl_135_3_LC_6_22_3.SEQ_MODE=4'b1000;
    defparam shift_srl_135_3_LC_6_22_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_135_3_LC_6_22_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53224),
            .lcout(shift_srl_135Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92991),
            .ce(N__53175),
            .sr(_gnd_net_));
    defparam shift_srl_135_4_LC_6_22_4.C_ON=1'b0;
    defparam shift_srl_135_4_LC_6_22_4.SEQ_MODE=4'b1000;
    defparam shift_srl_135_4_LC_6_22_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_135_4_LC_6_22_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53218),
            .lcout(shift_srl_135Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92991),
            .ce(N__53175),
            .sr(_gnd_net_));
    defparam shift_srl_135_1_LC_6_22_5.C_ON=1'b0;
    defparam shift_srl_135_1_LC_6_22_5.SEQ_MODE=4'b1000;
    defparam shift_srl_135_1_LC_6_22_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_135_1_LC_6_22_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53206),
            .lcout(shift_srl_135Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92991),
            .ce(N__53175),
            .sr(_gnd_net_));
    defparam shift_srl_135_6_LC_6_22_6.C_ON=1'b0;
    defparam shift_srl_135_6_LC_6_22_6.SEQ_MODE=4'b1000;
    defparam shift_srl_135_6_LC_6_22_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_135_6_LC_6_22_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53194),
            .lcout(shift_srl_135Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92991),
            .ce(N__53175),
            .sr(_gnd_net_));
    defparam shift_srl_135_7_LC_6_22_7.C_ON=1'b0;
    defparam shift_srl_135_7_LC_6_22_7.SEQ_MODE=4'b1000;
    defparam shift_srl_135_7_LC_6_22_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_135_7_LC_6_22_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53188),
            .lcout(shift_srl_135Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92991),
            .ce(N__53175),
            .sr(_gnd_net_));
    defparam shift_srl_116_0_LC_6_23_0.C_ON=1'b0;
    defparam shift_srl_116_0_LC_6_23_0.SEQ_MODE=4'b1000;
    defparam shift_srl_116_0_LC_6_23_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_116_0_LC_6_23_0 (
            .in0(N__58802),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_116Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93006),
            .ce(N__54576),
            .sr(_gnd_net_));
    defparam shift_srl_116_1_LC_6_23_1.C_ON=1'b0;
    defparam shift_srl_116_1_LC_6_23_1.SEQ_MODE=4'b1000;
    defparam shift_srl_116_1_LC_6_23_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_116_1_LC_6_23_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53158),
            .lcout(shift_srl_116Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93006),
            .ce(N__54576),
            .sr(_gnd_net_));
    defparam shift_srl_116_2_LC_6_23_2.C_ON=1'b0;
    defparam shift_srl_116_2_LC_6_23_2.SEQ_MODE=4'b1000;
    defparam shift_srl_116_2_LC_6_23_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_116_2_LC_6_23_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53152),
            .lcout(shift_srl_116Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93006),
            .ce(N__54576),
            .sr(_gnd_net_));
    defparam shift_srl_116_3_LC_6_23_3.C_ON=1'b0;
    defparam shift_srl_116_3_LC_6_23_3.SEQ_MODE=4'b1000;
    defparam shift_srl_116_3_LC_6_23_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_116_3_LC_6_23_3 (
            .in0(N__53146),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_116Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93006),
            .ce(N__54576),
            .sr(_gnd_net_));
    defparam shift_srl_116_4_LC_6_23_4.C_ON=1'b0;
    defparam shift_srl_116_4_LC_6_23_4.SEQ_MODE=4'b1000;
    defparam shift_srl_116_4_LC_6_23_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_116_4_LC_6_23_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53290),
            .lcout(shift_srl_116Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93006),
            .ce(N__54576),
            .sr(_gnd_net_));
    defparam shift_srl_116_5_LC_6_23_5.C_ON=1'b0;
    defparam shift_srl_116_5_LC_6_23_5.SEQ_MODE=4'b1000;
    defparam shift_srl_116_5_LC_6_23_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_116_5_LC_6_23_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53284),
            .lcout(shift_srl_116Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93006),
            .ce(N__54576),
            .sr(_gnd_net_));
    defparam shift_srl_116_6_LC_6_23_6.C_ON=1'b0;
    defparam shift_srl_116_6_LC_6_23_6.SEQ_MODE=4'b1000;
    defparam shift_srl_116_6_LC_6_23_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_116_6_LC_6_23_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53278),
            .lcout(shift_srl_116Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93006),
            .ce(N__54576),
            .sr(_gnd_net_));
    defparam shift_srl_116_7_LC_6_23_7.C_ON=1'b0;
    defparam shift_srl_116_7_LC_6_23_7.SEQ_MODE=4'b1000;
    defparam shift_srl_116_7_LC_6_23_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_116_7_LC_6_23_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53272),
            .lcout(shift_srl_116Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93006),
            .ce(N__54576),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_113_LC_6_24_0.C_ON=1'b0;
    defparam rco_obuf_RNO_113_LC_6_24_0.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_113_LC_6_24_0.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_113_LC_6_24_0 (
            .in0(N__60451),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60354),
            .lcout(rco_c_113),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_107_0_LC_6_26_3.C_ON=1'b0;
    defparam shift_srl_107_0_LC_6_26_3.SEQ_MODE=4'b1000;
    defparam shift_srl_107_0_LC_6_26_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_107_0_LC_6_26_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62371),
            .lcout(shift_srl_107Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93047),
            .ce(N__56687),
            .sr(_gnd_net_));
    defparam shift_srl_107_1_LC_6_26_4.C_ON=1'b0;
    defparam shift_srl_107_1_LC_6_26_4.SEQ_MODE=4'b1000;
    defparam shift_srl_107_1_LC_6_26_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_107_1_LC_6_26_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53242),
            .lcout(shift_srl_107Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93047),
            .ce(N__56687),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_164_LC_7_2_5.C_ON=1'b0;
    defparam rco_obuf_RNO_164_LC_7_2_5.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_164_LC_7_2_5.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_164_LC_7_2_5 (
            .in0(N__82435),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87708),
            .lcout(rco_c_164),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_1_7_LC_7_6_0.C_ON=1'b0;
    defparam shift_srl_1_7_LC_7_6_0.SEQ_MODE=4'b1000;
    defparam shift_srl_1_7_LC_7_6_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_1_7_LC_7_6_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53356),
            .lcout(shift_srl_1Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93097),
            .ce(N__54669),
            .sr(_gnd_net_));
    defparam shift_srl_1_8_LC_7_6_1.C_ON=1'b0;
    defparam shift_srl_1_8_LC_7_6_1.SEQ_MODE=4'b1000;
    defparam shift_srl_1_8_LC_7_6_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_1_8_LC_7_6_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53362),
            .lcout(shift_srl_1Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93097),
            .ce(N__54669),
            .sr(_gnd_net_));
    defparam shift_srl_1_6_LC_7_6_3.C_ON=1'b0;
    defparam shift_srl_1_6_LC_7_6_3.SEQ_MODE=4'b1000;
    defparam shift_srl_1_6_LC_7_6_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_1_6_LC_7_6_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53350),
            .lcout(shift_srl_1Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93097),
            .ce(N__54669),
            .sr(_gnd_net_));
    defparam shift_srl_1_5_LC_7_6_4.C_ON=1'b0;
    defparam shift_srl_1_5_LC_7_6_4.SEQ_MODE=4'b1000;
    defparam shift_srl_1_5_LC_7_6_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_1_5_LC_7_6_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53344),
            .lcout(shift_srl_1Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93097),
            .ce(N__54669),
            .sr(_gnd_net_));
    defparam shift_srl_1_4_LC_7_6_6.C_ON=1'b0;
    defparam shift_srl_1_4_LC_7_6_6.SEQ_MODE=4'b1000;
    defparam shift_srl_1_4_LC_7_6_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_1_4_LC_7_6_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54685),
            .lcout(shift_srl_1Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93097),
            .ce(N__54669),
            .sr(_gnd_net_));
    defparam shift_srl_1_RNI5UTI_15_LC_7_7_0.C_ON=1'b0;
    defparam shift_srl_1_RNI5UTI_15_LC_7_7_0.SEQ_MODE=4'b0000;
    defparam shift_srl_1_RNI5UTI_15_LC_7_7_0.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_1_RNI5UTI_15_LC_7_7_0 (
            .in0(N__57220),
            .in1(N__89761),
            .in2(_gnd_net_),
            .in3(N__57153),
            .lcout(N_12_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_1_14_LC_7_7_2.C_ON=1'b0;
    defparam shift_srl_1_14_LC_7_7_2.SEQ_MODE=4'b1000;
    defparam shift_srl_1_14_LC_7_7_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_1_14_LC_7_7_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53308),
            .lcout(shift_srl_1Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93081),
            .ce(N__54657),
            .sr(_gnd_net_));
    defparam shift_srl_1_13_LC_7_7_3.C_ON=1'b0;
    defparam shift_srl_1_13_LC_7_7_3.SEQ_MODE=4'b1000;
    defparam shift_srl_1_13_LC_7_7_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_1_13_LC_7_7_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53302),
            .lcout(shift_srl_1Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93081),
            .ce(N__54657),
            .sr(_gnd_net_));
    defparam shift_srl_1_12_LC_7_7_4.C_ON=1'b0;
    defparam shift_srl_1_12_LC_7_7_4.SEQ_MODE=4'b1000;
    defparam shift_srl_1_12_LC_7_7_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_1_12_LC_7_7_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53296),
            .lcout(shift_srl_1Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93081),
            .ce(N__54657),
            .sr(_gnd_net_));
    defparam shift_srl_1_11_LC_7_7_5.C_ON=1'b0;
    defparam shift_srl_1_11_LC_7_7_5.SEQ_MODE=4'b1000;
    defparam shift_srl_1_11_LC_7_7_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_1_11_LC_7_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53458),
            .lcout(shift_srl_1Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93081),
            .ce(N__54657),
            .sr(_gnd_net_));
    defparam shift_srl_1_10_LC_7_7_6.C_ON=1'b0;
    defparam shift_srl_1_10_LC_7_7_6.SEQ_MODE=4'b1000;
    defparam shift_srl_1_10_LC_7_7_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_1_10_LC_7_7_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53446),
            .lcout(shift_srl_1Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93081),
            .ce(N__54657),
            .sr(_gnd_net_));
    defparam shift_srl_1_9_LC_7_7_7.C_ON=1'b0;
    defparam shift_srl_1_9_LC_7_7_7.SEQ_MODE=4'b1000;
    defparam shift_srl_1_9_LC_7_7_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_1_9_LC_7_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53452),
            .lcout(shift_srl_1Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93081),
            .ce(N__54657),
            .sr(_gnd_net_));
    defparam shift_srl_1_15_LC_7_8_4.C_ON=1'b0;
    defparam shift_srl_1_15_LC_7_8_4.SEQ_MODE=4'b1000;
    defparam shift_srl_1_15_LC_7_8_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_1_15_LC_7_8_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53440),
            .lcout(shift_srl_1Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93066),
            .ce(N__54673),
            .sr(_gnd_net_));
    defparam shift_srl_23_RNIBC3N_15_LC_7_9_0.C_ON=1'b0;
    defparam shift_srl_23_RNIBC3N_15_LC_7_9_0.SEQ_MODE=4'b0000;
    defparam shift_srl_23_RNIBC3N_15_LC_7_9_0.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_23_RNIBC3N_15_LC_7_9_0 (
            .in0(N__53388),
            .in1(N__53426),
            .in2(_gnd_net_),
            .in3(N__55710),
            .lcout(N_4016_i_0_a2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_23_15_LC_7_9_1.C_ON=1'b0;
    defparam shift_srl_23_15_LC_7_9_1.SEQ_MODE=4'b1000;
    defparam shift_srl_23_15_LC_7_9_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_23_15_LC_7_9_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53395),
            .lcout(shift_srl_23Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93050),
            .ce(N__53580),
            .sr(_gnd_net_));
    defparam shift_srl_23_0_LC_7_9_2.C_ON=1'b0;
    defparam shift_srl_23_0_LC_7_9_2.SEQ_MODE=4'b1000;
    defparam shift_srl_23_0_LC_7_9_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_23_0_LC_7_9_2 (
            .in0(N__53389),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_23Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93050),
            .ce(N__53580),
            .sr(_gnd_net_));
    defparam shift_srl_23_1_LC_7_9_3.C_ON=1'b0;
    defparam shift_srl_23_1_LC_7_9_3.SEQ_MODE=4'b1000;
    defparam shift_srl_23_1_LC_7_9_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_23_1_LC_7_9_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53380),
            .lcout(shift_srl_23Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93050),
            .ce(N__53580),
            .sr(_gnd_net_));
    defparam shift_srl_23_2_LC_7_9_4.C_ON=1'b0;
    defparam shift_srl_23_2_LC_7_9_4.SEQ_MODE=4'b1000;
    defparam shift_srl_23_2_LC_7_9_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_23_2_LC_7_9_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53374),
            .lcout(shift_srl_23Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93050),
            .ce(N__53580),
            .sr(_gnd_net_));
    defparam shift_srl_23_3_LC_7_9_5.C_ON=1'b0;
    defparam shift_srl_23_3_LC_7_9_5.SEQ_MODE=4'b1000;
    defparam shift_srl_23_3_LC_7_9_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_23_3_LC_7_9_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53368),
            .lcout(shift_srl_23Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93050),
            .ce(N__53580),
            .sr(_gnd_net_));
    defparam shift_srl_23_4_LC_7_9_6.C_ON=1'b0;
    defparam shift_srl_23_4_LC_7_9_6.SEQ_MODE=4'b1000;
    defparam shift_srl_23_4_LC_7_9_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_23_4_LC_7_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53605),
            .lcout(shift_srl_23Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93050),
            .ce(N__53580),
            .sr(_gnd_net_));
    defparam shift_srl_23_5_LC_7_9_7.C_ON=1'b0;
    defparam shift_srl_23_5_LC_7_9_7.SEQ_MODE=4'b1000;
    defparam shift_srl_23_5_LC_7_9_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_23_5_LC_7_9_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53599),
            .lcout(shift_srl_23Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93050),
            .ce(N__53580),
            .sr(_gnd_net_));
    defparam shift_srl_23_6_LC_7_10_0.C_ON=1'b0;
    defparam shift_srl_23_6_LC_7_10_0.SEQ_MODE=4'b1000;
    defparam shift_srl_23_6_LC_7_10_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_23_6_LC_7_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53593),
            .lcout(shift_srl_23Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93034),
            .ce(N__53581),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_155_LC_7_13_0.C_ON=1'b0;
    defparam rco_obuf_RNO_155_LC_7_13_0.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_155_LC_7_13_0.LUT_INIT=16'b1000100000000000;
    LogicCell40 rco_obuf_RNO_155_LC_7_13_0 (
            .in0(N__87905),
            .in1(N__77656),
            .in2(_gnd_net_),
            .in3(N__77606),
            .lcout(rco_c_155),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_154_LC_7_13_1.C_ON=1'b0;
    defparam rco_obuf_RNO_154_LC_7_13_1.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_154_LC_7_13_1.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_154_LC_7_13_1 (
            .in0(N__77605),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87904),
            .lcout(rco_c_154),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_156_LC_7_13_2.C_ON=1'b0;
    defparam rco_obuf_RNO_156_LC_7_13_2.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_156_LC_7_13_2.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_156_LC_7_13_2 (
            .in0(N__87906),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77557),
            .lcout(rco_c_156),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_159_LC_7_13_3.C_ON=1'b0;
    defparam rco_obuf_RNO_159_LC_7_13_3.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_159_LC_7_13_3.LUT_INIT=16'b1100110000000000;
    LogicCell40 rco_obuf_RNO_159_LC_7_13_3 (
            .in0(_gnd_net_),
            .in1(N__71656),
            .in2(_gnd_net_),
            .in3(N__87907),
            .lcout(rco_c_159),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_160_LC_7_13_4.C_ON=1'b0;
    defparam rco_obuf_RNO_160_LC_7_13_4.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_160_LC_7_13_4.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_160_LC_7_13_4 (
            .in0(N__87908),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69860),
            .lcout(rco_c_160),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_161_LC_7_13_5.C_ON=1'b0;
    defparam rco_obuf_RNO_161_LC_7_13_5.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_161_LC_7_13_5.LUT_INIT=16'b1000100000000000;
    LogicCell40 rco_obuf_RNO_161_LC_7_13_5 (
            .in0(N__69861),
            .in1(N__77369),
            .in2(_gnd_net_),
            .in3(N__87909),
            .lcout(rco_c_161),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_154_0_LC_7_13_6.C_ON=1'b0;
    defparam shift_srl_154_0_LC_7_13_6.SEQ_MODE=4'b1000;
    defparam shift_srl_154_0_LC_7_13_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_154_0_LC_7_13_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77604),
            .lcout(shift_srl_154Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92992),
            .ce(N__57341),
            .sr(_gnd_net_));
    defparam shift_srl_154_1_LC_7_13_7.C_ON=1'b0;
    defparam shift_srl_154_1_LC_7_13_7.SEQ_MODE=4'b1000;
    defparam shift_srl_154_1_LC_7_13_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_154_1_LC_7_13_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53866),
            .lcout(shift_srl_154Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92992),
            .ce(N__57341),
            .sr(_gnd_net_));
    defparam shift_srl_154_2_LC_7_14_0.C_ON=1'b0;
    defparam shift_srl_154_2_LC_7_14_0.SEQ_MODE=4'b1000;
    defparam shift_srl_154_2_LC_7_14_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_154_2_LC_7_14_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53860),
            .lcout(shift_srl_154Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92980),
            .ce(N__57355),
            .sr(_gnd_net_));
    defparam shift_srl_154_3_LC_7_14_1.C_ON=1'b0;
    defparam shift_srl_154_3_LC_7_14_1.SEQ_MODE=4'b1000;
    defparam shift_srl_154_3_LC_7_14_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_154_3_LC_7_14_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53854),
            .lcout(shift_srl_154Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92980),
            .ce(N__57355),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_26_LC_7_15_0.C_ON=1'b0;
    defparam rco_obuf_RNO_26_LC_7_15_0.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_26_LC_7_15_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 rco_obuf_RNO_26_LC_7_15_0 (
            .in0(N__83803),
            .in1(N__71542),
            .in2(N__71502),
            .in3(N__85116),
            .lcout(rco_c_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIBK2U6_15_LC_7_15_1.C_ON=1'b0;
    defparam shift_srl_0_RNIBK2U6_15_LC_7_15_1.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIBK2U6_15_LC_7_15_1.LUT_INIT=16'b1010101000000000;
    LogicCell40 shift_srl_0_RNIBK2U6_15_LC_7_15_1 (
            .in0(N__90185),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53933),
            .lcout(clk_en_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_9_RNI7SS8_15_LC_7_15_2.C_ON=1'b0;
    defparam shift_srl_9_RNI7SS8_15_LC_7_15_2.SEQ_MODE=4'b0000;
    defparam shift_srl_9_RNI7SS8_15_LC_7_15_2.LUT_INIT=16'b1100110000000000;
    LogicCell40 shift_srl_9_RNI7SS8_15_LC_7_15_2 (
            .in0(_gnd_net_),
            .in1(N__53919),
            .in2(_gnd_net_),
            .in3(N__53822),
            .lcout(rco_int_0_a2_0_9),
            .ltout(rco_int_0_a2_0_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_7_RNIE24H2_15_LC_7_15_3.C_ON=1'b0;
    defparam shift_srl_7_RNIE24H2_15_LC_7_15_3.SEQ_MODE=4'b0000;
    defparam shift_srl_7_RNIE24H2_15_LC_7_15_3.LUT_INIT=16'b0010000000000000;
    LogicCell40 shift_srl_7_RNIE24H2_15_LC_7_15_3 (
            .in0(N__53770),
            .in1(N__53701),
            .in2(N__53647),
            .in3(N__53643),
            .lcout(rco_c_9),
            .ltout(rco_c_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_23_RNIDRH46_15_LC_7_15_4.C_ON=1'b0;
    defparam shift_srl_23_RNIDRH46_15_LC_7_15_4.SEQ_MODE=4'b0000;
    defparam shift_srl_23_RNIDRH46_15_LC_7_15_4.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_23_RNIDRH46_15_LC_7_15_4 (
            .in0(N__69276),
            .in1(N__69294),
            .in2(N__53608),
            .in3(N__69227),
            .lcout(N_4016_i),
            .ltout(N_4016_i_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_25_RNIG88T6_15_LC_7_15_5.C_ON=1'b0;
    defparam shift_srl_25_RNIG88T6_15_LC_7_15_5.SEQ_MODE=4'b0000;
    defparam shift_srl_25_RNIG88T6_15_LC_7_15_5.LUT_INIT=16'b1100000000000000;
    LogicCell40 shift_srl_25_RNIG88T6_15_LC_7_15_5 (
            .in0(_gnd_net_),
            .in1(N__71492),
            .in2(N__53953),
            .in3(N__83802),
            .lcout(rco_c_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_26_RNIU0N07_15_LC_7_15_6.C_ON=1'b0;
    defparam shift_srl_26_RNIU0N07_15_LC_7_15_6.SEQ_MODE=4'b0000;
    defparam shift_srl_26_RNIU0N07_15_LC_7_15_6.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_26_RNIU0N07_15_LC_7_15_6 (
            .in0(N__53934),
            .in1(N__71541),
            .in2(_gnd_net_),
            .in3(N__90184),
            .lcout(clk_en_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_9_15_LC_7_15_7.C_ON=1'b0;
    defparam shift_srl_9_15_LC_7_15_7.SEQ_MODE=4'b1000;
    defparam shift_srl_9_15_LC_7_15_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_9_15_LC_7_15_7 (
            .in0(N__53884),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_9Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92969),
            .ce(N__54082),
            .sr(_gnd_net_));
    defparam shift_srl_9_10_LC_7_16_0.C_ON=1'b0;
    defparam shift_srl_9_10_LC_7_16_0.SEQ_MODE=4'b1000;
    defparam shift_srl_9_10_LC_7_16_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_9_10_LC_7_16_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53878),
            .lcout(shift_srl_9Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92958),
            .ce(N__54081),
            .sr(_gnd_net_));
    defparam shift_srl_9_11_LC_7_16_1.C_ON=1'b0;
    defparam shift_srl_9_11_LC_7_16_1.SEQ_MODE=4'b1000;
    defparam shift_srl_9_11_LC_7_16_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_9_11_LC_7_16_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53908),
            .lcout(shift_srl_9Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92958),
            .ce(N__54081),
            .sr(_gnd_net_));
    defparam shift_srl_9_12_LC_7_16_2.C_ON=1'b0;
    defparam shift_srl_9_12_LC_7_16_2.SEQ_MODE=4'b1000;
    defparam shift_srl_9_12_LC_7_16_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_9_12_LC_7_16_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53902),
            .lcout(shift_srl_9Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92958),
            .ce(N__54081),
            .sr(_gnd_net_));
    defparam shift_srl_9_13_LC_7_16_3.C_ON=1'b0;
    defparam shift_srl_9_13_LC_7_16_3.SEQ_MODE=4'b1000;
    defparam shift_srl_9_13_LC_7_16_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_9_13_LC_7_16_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53896),
            .lcout(shift_srl_9Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92958),
            .ce(N__54081),
            .sr(_gnd_net_));
    defparam shift_srl_9_14_LC_7_16_4.C_ON=1'b0;
    defparam shift_srl_9_14_LC_7_16_4.SEQ_MODE=4'b1000;
    defparam shift_srl_9_14_LC_7_16_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_9_14_LC_7_16_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53890),
            .lcout(shift_srl_9Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92958),
            .ce(N__54081),
            .sr(_gnd_net_));
    defparam shift_srl_9_9_LC_7_16_5.C_ON=1'b0;
    defparam shift_srl_9_9_LC_7_16_5.SEQ_MODE=4'b1000;
    defparam shift_srl_9_9_LC_7_16_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_9_9_LC_7_16_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53872),
            .lcout(shift_srl_9Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92958),
            .ce(N__54081),
            .sr(_gnd_net_));
    defparam shift_srl_9_8_LC_7_16_6.C_ON=1'b0;
    defparam shift_srl_9_8_LC_7_16_6.SEQ_MODE=4'b1000;
    defparam shift_srl_9_8_LC_7_16_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_9_8_LC_7_16_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54088),
            .lcout(shift_srl_9Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92958),
            .ce(N__54081),
            .sr(_gnd_net_));
    defparam shift_srl_9_7_LC_7_16_7.C_ON=1'b0;
    defparam shift_srl_9_7_LC_7_16_7.SEQ_MODE=4'b1000;
    defparam shift_srl_9_7_LC_7_16_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_9_7_LC_7_16_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54094),
            .lcout(shift_srl_9Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92958),
            .ce(N__54081),
            .sr(_gnd_net_));
    defparam shift_srl_128_0_LC_7_17_0.C_ON=1'b0;
    defparam shift_srl_128_0_LC_7_17_0.SEQ_MODE=4'b1000;
    defparam shift_srl_128_0_LC_7_17_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_128_0_LC_7_17_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__91256),
            .lcout(shift_srl_128Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92938),
            .ce(N__56280),
            .sr(_gnd_net_));
    defparam shift_srl_128_1_LC_7_17_1.C_ON=1'b0;
    defparam shift_srl_128_1_LC_7_17_1.SEQ_MODE=4'b1000;
    defparam shift_srl_128_1_LC_7_17_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_128_1_LC_7_17_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54049),
            .lcout(shift_srl_128Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92938),
            .ce(N__56280),
            .sr(_gnd_net_));
    defparam shift_srl_128_2_LC_7_17_2.C_ON=1'b0;
    defparam shift_srl_128_2_LC_7_17_2.SEQ_MODE=4'b1000;
    defparam shift_srl_128_2_LC_7_17_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_128_2_LC_7_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54043),
            .lcout(shift_srl_128Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92938),
            .ce(N__56280),
            .sr(_gnd_net_));
    defparam shift_srl_128_3_LC_7_17_3.C_ON=1'b0;
    defparam shift_srl_128_3_LC_7_17_3.SEQ_MODE=4'b1000;
    defparam shift_srl_128_3_LC_7_17_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_128_3_LC_7_17_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54037),
            .lcout(shift_srl_128Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92938),
            .ce(N__56280),
            .sr(_gnd_net_));
    defparam shift_srl_128_4_LC_7_17_4.C_ON=1'b0;
    defparam shift_srl_128_4_LC_7_17_4.SEQ_MODE=4'b1000;
    defparam shift_srl_128_4_LC_7_17_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_128_4_LC_7_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54031),
            .lcout(shift_srl_128Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92938),
            .ce(N__56280),
            .sr(_gnd_net_));
    defparam shift_srl_128_5_LC_7_17_5.C_ON=1'b0;
    defparam shift_srl_128_5_LC_7_17_5.SEQ_MODE=4'b1000;
    defparam shift_srl_128_5_LC_7_17_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_128_5_LC_7_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54025),
            .lcout(shift_srl_128Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92938),
            .ce(N__56280),
            .sr(_gnd_net_));
    defparam shift_srl_128_6_LC_7_17_6.C_ON=1'b0;
    defparam shift_srl_128_6_LC_7_17_6.SEQ_MODE=4'b1000;
    defparam shift_srl_128_6_LC_7_17_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_128_6_LC_7_17_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54019),
            .lcout(shift_srl_128Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92938),
            .ce(N__56280),
            .sr(_gnd_net_));
    defparam shift_srl_129_15_LC_7_18_4.C_ON=1'b0;
    defparam shift_srl_129_15_LC_7_18_4.SEQ_MODE=4'b1000;
    defparam shift_srl_129_15_LC_7_18_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_129_15_LC_7_18_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54007),
            .lcout(shift_srl_129Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92959),
            .ce(N__53995),
            .sr(_gnd_net_));
    defparam shift_srl_132_RNIEU7K_0_15_LC_7_19_0.C_ON=1'b0;
    defparam shift_srl_132_RNIEU7K_0_15_LC_7_19_0.SEQ_MODE=4'b0000;
    defparam shift_srl_132_RNIEU7K_0_15_LC_7_19_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_132_RNIEU7K_0_15_LC_7_19_0 (
            .in0(N__54341),
            .in1(N__54300),
            .in2(N__91245),
            .in3(N__54186),
            .lcout(g0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_128_15_LC_7_19_1.C_ON=1'b0;
    defparam shift_srl_128_15_LC_7_19_1.SEQ_MODE=4'b1000;
    defparam shift_srl_128_15_LC_7_19_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_128_15_LC_7_19_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54139),
            .lcout(shift_srl_128Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92970),
            .ce(N__56279),
            .sr(_gnd_net_));
    defparam shift_srl_128_14_LC_7_19_2.C_ON=1'b0;
    defparam shift_srl_128_14_LC_7_19_2.SEQ_MODE=4'b1000;
    defparam shift_srl_128_14_LC_7_19_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_128_14_LC_7_19_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54133),
            .lcout(shift_srl_128Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92970),
            .ce(N__56279),
            .sr(_gnd_net_));
    defparam shift_srl_128_13_LC_7_19_3.C_ON=1'b0;
    defparam shift_srl_128_13_LC_7_19_3.SEQ_MODE=4'b1000;
    defparam shift_srl_128_13_LC_7_19_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_128_13_LC_7_19_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54127),
            .lcout(shift_srl_128Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92970),
            .ce(N__56279),
            .sr(_gnd_net_));
    defparam shift_srl_128_12_LC_7_19_4.C_ON=1'b0;
    defparam shift_srl_128_12_LC_7_19_4.SEQ_MODE=4'b1000;
    defparam shift_srl_128_12_LC_7_19_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_128_12_LC_7_19_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54121),
            .lcout(shift_srl_128Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92970),
            .ce(N__56279),
            .sr(_gnd_net_));
    defparam shift_srl_128_11_LC_7_19_5.C_ON=1'b0;
    defparam shift_srl_128_11_LC_7_19_5.SEQ_MODE=4'b1000;
    defparam shift_srl_128_11_LC_7_19_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_128_11_LC_7_19_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54115),
            .lcout(shift_srl_128Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92970),
            .ce(N__56279),
            .sr(_gnd_net_));
    defparam shift_srl_128_10_LC_7_19_6.C_ON=1'b0;
    defparam shift_srl_128_10_LC_7_19_6.SEQ_MODE=4'b1000;
    defparam shift_srl_128_10_LC_7_19_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_128_10_LC_7_19_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54100),
            .lcout(shift_srl_128Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92970),
            .ce(N__56279),
            .sr(_gnd_net_));
    defparam shift_srl_128_9_LC_7_19_7.C_ON=1'b0;
    defparam shift_srl_128_9_LC_7_19_7.SEQ_MODE=4'b1000;
    defparam shift_srl_128_9_LC_7_19_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_128_9_LC_7_19_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54109),
            .lcout(shift_srl_128Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92970),
            .ce(N__56279),
            .sr(_gnd_net_));
    defparam shift_srl_113_RNI405M_15_LC_7_20_0.C_ON=1'b0;
    defparam shift_srl_113_RNI405M_15_LC_7_20_0.SEQ_MODE=4'b0000;
    defparam shift_srl_113_RNI405M_15_LC_7_20_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_113_RNI405M_15_LC_7_20_0 (
            .in0(N__60322),
            .in1(N__66461),
            .in2(N__90435),
            .in3(N__60450),
            .lcout(g0_9_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_144_RNILM4U4_15_LC_7_20_5.C_ON=1'b0;
    defparam shift_srl_144_RNILM4U4_15_LC_7_20_5.SEQ_MODE=4'b0000;
    defparam shift_srl_144_RNILM4U4_15_LC_7_20_5.LUT_INIT=16'b1111011111111111;
    LogicCell40 shift_srl_144_RNILM4U4_15_LC_7_20_5 (
            .in0(N__62130),
            .in1(N__65717),
            .in2(N__54490),
            .in3(N__66621),
            .lcout(rco_int_0_a2_0_a2_1_1_145),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_136_RNI96PM_15_LC_7_21_0.C_ON=1'b0;
    defparam shift_srl_136_RNI96PM_15_LC_7_21_0.SEQ_MODE=4'b0000;
    defparam shift_srl_136_RNI96PM_15_LC_7_21_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_136_RNI96PM_15_LC_7_21_0 (
            .in0(N__60529),
            .in1(N__63812),
            .in2(N__54481),
            .in3(N__58787),
            .lcout(g0_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_116_15_LC_7_21_1.C_ON=1'b0;
    defparam shift_srl_116_15_LC_7_21_1.SEQ_MODE=4'b1000;
    defparam shift_srl_116_15_LC_7_21_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_116_15_LC_7_21_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54418),
            .lcout(shift_srl_116Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92993),
            .ce(N__54569),
            .sr(_gnd_net_));
    defparam shift_srl_116_14_LC_7_21_2.C_ON=1'b0;
    defparam shift_srl_116_14_LC_7_21_2.SEQ_MODE=4'b1000;
    defparam shift_srl_116_14_LC_7_21_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_116_14_LC_7_21_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54412),
            .lcout(shift_srl_116Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92993),
            .ce(N__54569),
            .sr(_gnd_net_));
    defparam shift_srl_116_13_LC_7_21_3.C_ON=1'b0;
    defparam shift_srl_116_13_LC_7_21_3.SEQ_MODE=4'b1000;
    defparam shift_srl_116_13_LC_7_21_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_116_13_LC_7_21_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54406),
            .lcout(shift_srl_116Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92993),
            .ce(N__54569),
            .sr(_gnd_net_));
    defparam shift_srl_116_12_LC_7_21_4.C_ON=1'b0;
    defparam shift_srl_116_12_LC_7_21_4.SEQ_MODE=4'b1000;
    defparam shift_srl_116_12_LC_7_21_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_116_12_LC_7_21_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54400),
            .lcout(shift_srl_116Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92993),
            .ce(N__54569),
            .sr(_gnd_net_));
    defparam shift_srl_116_11_LC_7_21_5.C_ON=1'b0;
    defparam shift_srl_116_11_LC_7_21_5.SEQ_MODE=4'b1000;
    defparam shift_srl_116_11_LC_7_21_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_116_11_LC_7_21_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54394),
            .lcout(shift_srl_116Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92993),
            .ce(N__54569),
            .sr(_gnd_net_));
    defparam shift_srl_116_10_LC_7_21_6.C_ON=1'b0;
    defparam shift_srl_116_10_LC_7_21_6.SEQ_MODE=4'b1000;
    defparam shift_srl_116_10_LC_7_21_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_116_10_LC_7_21_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54376),
            .lcout(shift_srl_116Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92993),
            .ce(N__54569),
            .sr(_gnd_net_));
    defparam shift_srl_116_9_LC_7_21_7.C_ON=1'b0;
    defparam shift_srl_116_9_LC_7_21_7.SEQ_MODE=4'b1000;
    defparam shift_srl_116_9_LC_7_21_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_116_9_LC_7_21_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54388),
            .lcout(shift_srl_116Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92993),
            .ce(N__54569),
            .sr(_gnd_net_));
    defparam shift_srl_112_0_LC_7_22_0.C_ON=1'b0;
    defparam shift_srl_112_0_LC_7_22_0.SEQ_MODE=4'b1000;
    defparam shift_srl_112_0_LC_7_22_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_112_0_LC_7_22_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60528),
            .lcout(shift_srl_112Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93007),
            .ce(N__60169),
            .sr(_gnd_net_));
    defparam shift_srl_112_1_LC_7_22_1.C_ON=1'b0;
    defparam shift_srl_112_1_LC_7_22_1.SEQ_MODE=4'b1000;
    defparam shift_srl_112_1_LC_7_22_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_112_1_LC_7_22_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54544),
            .lcout(shift_srl_112Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93007),
            .ce(N__60169),
            .sr(_gnd_net_));
    defparam shift_srl_112_2_LC_7_22_2.C_ON=1'b0;
    defparam shift_srl_112_2_LC_7_22_2.SEQ_MODE=4'b1000;
    defparam shift_srl_112_2_LC_7_22_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_112_2_LC_7_22_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54538),
            .lcout(shift_srl_112Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93007),
            .ce(N__60169),
            .sr(_gnd_net_));
    defparam shift_srl_112_3_LC_7_22_3.C_ON=1'b0;
    defparam shift_srl_112_3_LC_7_22_3.SEQ_MODE=4'b1000;
    defparam shift_srl_112_3_LC_7_22_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_112_3_LC_7_22_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54532),
            .lcout(shift_srl_112Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93007),
            .ce(N__60169),
            .sr(_gnd_net_));
    defparam shift_srl_112_4_LC_7_22_4.C_ON=1'b0;
    defparam shift_srl_112_4_LC_7_22_4.SEQ_MODE=4'b1000;
    defparam shift_srl_112_4_LC_7_22_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_112_4_LC_7_22_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54526),
            .lcout(shift_srl_112Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93007),
            .ce(N__60169),
            .sr(_gnd_net_));
    defparam shift_srl_112_5_LC_7_22_5.C_ON=1'b0;
    defparam shift_srl_112_5_LC_7_22_5.SEQ_MODE=4'b1000;
    defparam shift_srl_112_5_LC_7_22_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_112_5_LC_7_22_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54520),
            .lcout(shift_srl_112Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93007),
            .ce(N__60169),
            .sr(_gnd_net_));
    defparam shift_srl_112_6_LC_7_22_6.C_ON=1'b0;
    defparam shift_srl_112_6_LC_7_22_6.SEQ_MODE=4'b1000;
    defparam shift_srl_112_6_LC_7_22_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_112_6_LC_7_22_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54514),
            .lcout(shift_srl_112Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93007),
            .ce(N__60169),
            .sr(_gnd_net_));
    defparam shift_srl_112_7_LC_7_22_7.C_ON=1'b0;
    defparam shift_srl_112_7_LC_7_22_7.SEQ_MODE=4'b1000;
    defparam shift_srl_112_7_LC_7_22_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_112_7_LC_7_22_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54508),
            .lcout(shift_srl_112Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93007),
            .ce(N__60169),
            .sr(_gnd_net_));
    defparam shift_srl_123_4_LC_7_23_0.C_ON=1'b0;
    defparam shift_srl_123_4_LC_7_23_0.SEQ_MODE=4'b1000;
    defparam shift_srl_123_4_LC_7_23_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_123_4_LC_7_23_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54607),
            .lcout(shift_srl_123Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93020),
            .ce(N__56206),
            .sr(_gnd_net_));
    defparam shift_srl_123_5_LC_7_23_1.C_ON=1'b0;
    defparam shift_srl_123_5_LC_7_23_1.SEQ_MODE=4'b1000;
    defparam shift_srl_123_5_LC_7_23_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_123_5_LC_7_23_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54619),
            .lcout(shift_srl_123Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93020),
            .ce(N__56206),
            .sr(_gnd_net_));
    defparam shift_srl_123_6_LC_7_23_2.C_ON=1'b0;
    defparam shift_srl_123_6_LC_7_23_2.SEQ_MODE=4'b1000;
    defparam shift_srl_123_6_LC_7_23_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_123_6_LC_7_23_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54613),
            .lcout(shift_srl_123Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93020),
            .ce(N__56206),
            .sr(_gnd_net_));
    defparam shift_srl_123_3_LC_7_23_6.C_ON=1'b0;
    defparam shift_srl_123_3_LC_7_23_6.SEQ_MODE=4'b1000;
    defparam shift_srl_123_3_LC_7_23_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_123_3_LC_7_23_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56218),
            .lcout(shift_srl_123Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93020),
            .ce(N__56206),
            .sr(_gnd_net_));
    defparam shift_srl_199_7_LC_7_24_0.C_ON=1'b0;
    defparam shift_srl_199_7_LC_7_24_0.SEQ_MODE=4'b1000;
    defparam shift_srl_199_7_LC_7_24_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_199_7_LC_7_24_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60862),
            .lcout(shift_srl_199Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93035),
            .ce(N__62731),
            .sr(_gnd_net_));
    defparam shift_srl_107_7_LC_7_25_4.C_ON=1'b0;
    defparam shift_srl_107_7_LC_7_25_4.SEQ_MODE=4'b1000;
    defparam shift_srl_107_7_LC_7_25_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_107_7_LC_7_25_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54583),
            .lcout(shift_srl_107Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93049),
            .ce(N__56692),
            .sr(_gnd_net_));
    defparam shift_srl_107_5_LC_7_26_0.C_ON=1'b0;
    defparam shift_srl_107_5_LC_7_26_0.SEQ_MODE=4'b1000;
    defparam shift_srl_107_5_LC_7_26_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_107_5_LC_7_26_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54595),
            .lcout(shift_srl_107Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93065),
            .ce(N__56691),
            .sr(_gnd_net_));
    defparam shift_srl_107_3_LC_7_26_1.C_ON=1'b0;
    defparam shift_srl_107_3_LC_7_26_1.SEQ_MODE=4'b1000;
    defparam shift_srl_107_3_LC_7_26_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_107_3_LC_7_26_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54718),
            .lcout(shift_srl_107Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93065),
            .ce(N__56691),
            .sr(_gnd_net_));
    defparam shift_srl_107_4_LC_7_26_2.C_ON=1'b0;
    defparam shift_srl_107_4_LC_7_26_2.SEQ_MODE=4'b1000;
    defparam shift_srl_107_4_LC_7_26_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_107_4_LC_7_26_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54601),
            .lcout(shift_srl_107Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93065),
            .ce(N__56691),
            .sr(_gnd_net_));
    defparam shift_srl_107_6_LC_7_26_3.C_ON=1'b0;
    defparam shift_srl_107_6_LC_7_26_3.SEQ_MODE=4'b1000;
    defparam shift_srl_107_6_LC_7_26_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_107_6_LC_7_26_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54589),
            .lcout(shift_srl_107Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93065),
            .ce(N__56691),
            .sr(_gnd_net_));
    defparam shift_srl_107_2_LC_7_26_4.C_ON=1'b0;
    defparam shift_srl_107_2_LC_7_26_4.SEQ_MODE=4'b1000;
    defparam shift_srl_107_2_LC_7_26_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_107_2_LC_7_26_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54724),
            .lcout(shift_srl_107Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93065),
            .ce(N__56691),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_151_LC_9_5_1.C_ON=1'b0;
    defparam rco_obuf_RNO_151_LC_9_5_1.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_151_LC_9_5_1.LUT_INIT=16'b1000100000000000;
    LogicCell40 rco_obuf_RNO_151_LC_9_5_1 (
            .in0(N__82222),
            .in1(N__66806),
            .in2(_gnd_net_),
            .in3(N__63427),
            .lcout(rco_c_151),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam en_in_ibuf_RNI9ETD_LC_9_7_0.C_ON=1'b0;
    defparam en_in_ibuf_RNI9ETD_LC_9_7_0.SEQ_MODE=4'b0000;
    defparam en_in_ibuf_RNI9ETD_LC_9_7_0.LUT_INIT=16'b1010101000000000;
    LogicCell40 en_in_ibuf_RNI9ETD_LC_9_7_0 (
            .in0(N__57234),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__89902),
            .lcout(N_10_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_1_0_LC_9_7_1.C_ON=1'b0;
    defparam shift_srl_1_0_LC_9_7_1.SEQ_MODE=4'b1000;
    defparam shift_srl_1_0_LC_9_7_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_1_0_LC_9_7_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57165),
            .lcout(shift_srl_1Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93116),
            .ce(N__54650),
            .sr(_gnd_net_));
    defparam shift_srl_1_1_LC_9_7_2.C_ON=1'b0;
    defparam shift_srl_1_1_LC_9_7_2.SEQ_MODE=4'b1000;
    defparam shift_srl_1_1_LC_9_7_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_1_1_LC_9_7_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54703),
            .lcout(shift_srl_1Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93116),
            .ce(N__54650),
            .sr(_gnd_net_));
    defparam shift_srl_1_2_LC_9_7_3.C_ON=1'b0;
    defparam shift_srl_1_2_LC_9_7_3.SEQ_MODE=4'b1000;
    defparam shift_srl_1_2_LC_9_7_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_1_2_LC_9_7_3 (
            .in0(N__54697),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_1Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93116),
            .ce(N__54650),
            .sr(_gnd_net_));
    defparam shift_srl_1_3_LC_9_7_4.C_ON=1'b0;
    defparam shift_srl_1_3_LC_9_7_4.SEQ_MODE=4'b1000;
    defparam shift_srl_1_3_LC_9_7_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_1_3_LC_9_7_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54691),
            .lcout(shift_srl_1Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93116),
            .ce(N__54650),
            .sr(_gnd_net_));
    defparam shift_srl_10_10_LC_9_9_0.C_ON=1'b0;
    defparam shift_srl_10_10_LC_9_9_0.SEQ_MODE=4'b1000;
    defparam shift_srl_10_10_LC_9_9_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_10_10_LC_9_9_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54754),
            .lcout(shift_srl_10Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93083),
            .ce(N__55645),
            .sr(_gnd_net_));
    defparam shift_srl_10_11_LC_9_9_1.C_ON=1'b0;
    defparam shift_srl_10_11_LC_9_9_1.SEQ_MODE=4'b1000;
    defparam shift_srl_10_11_LC_9_9_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_10_11_LC_9_9_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54625),
            .lcout(shift_srl_10Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93083),
            .ce(N__55645),
            .sr(_gnd_net_));
    defparam shift_srl_10_12_LC_9_9_2.C_ON=1'b0;
    defparam shift_srl_10_12_LC_9_9_2.SEQ_MODE=4'b1000;
    defparam shift_srl_10_12_LC_9_9_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_10_12_LC_9_9_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54778),
            .lcout(shift_srl_10Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93083),
            .ce(N__55645),
            .sr(_gnd_net_));
    defparam shift_srl_10_13_LC_9_9_3.C_ON=1'b0;
    defparam shift_srl_10_13_LC_9_9_3.SEQ_MODE=4'b1000;
    defparam shift_srl_10_13_LC_9_9_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_10_13_LC_9_9_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54772),
            .lcout(shift_srl_10Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93083),
            .ce(N__55645),
            .sr(_gnd_net_));
    defparam shift_srl_10_14_LC_9_9_4.C_ON=1'b0;
    defparam shift_srl_10_14_LC_9_9_4.SEQ_MODE=4'b1000;
    defparam shift_srl_10_14_LC_9_9_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_10_14_LC_9_9_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54766),
            .lcout(shift_srl_10Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93083),
            .ce(N__55645),
            .sr(_gnd_net_));
    defparam shift_srl_10_15_LC_9_9_5.C_ON=1'b0;
    defparam shift_srl_10_15_LC_9_9_5.SEQ_MODE=4'b1000;
    defparam shift_srl_10_15_LC_9_9_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_10_15_LC_9_9_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54760),
            .lcout(shift_srl_10Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93083),
            .ce(N__55645),
            .sr(_gnd_net_));
    defparam shift_srl_10_9_LC_9_9_6.C_ON=1'b0;
    defparam shift_srl_10_9_LC_9_9_6.SEQ_MODE=4'b1000;
    defparam shift_srl_10_9_LC_9_9_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_10_9_LC_9_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54748),
            .lcout(shift_srl_10Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93083),
            .ce(N__55645),
            .sr(_gnd_net_));
    defparam shift_srl_10_8_LC_9_9_7.C_ON=1'b0;
    defparam shift_srl_10_8_LC_9_9_7.SEQ_MODE=4'b1000;
    defparam shift_srl_10_8_LC_9_9_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_10_8_LC_9_9_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55552),
            .lcout(shift_srl_10Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93083),
            .ce(N__55645),
            .sr(_gnd_net_));
    defparam shift_srl_150_0_LC_9_10_0.C_ON=1'b0;
    defparam shift_srl_150_0_LC_9_10_0.SEQ_MODE=4'b1000;
    defparam shift_srl_150_0_LC_9_10_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_150_0_LC_9_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56088),
            .lcout(shift_srl_150Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93067),
            .ce(N__55615),
            .sr(_gnd_net_));
    defparam shift_srl_150_1_LC_9_10_1.C_ON=1'b0;
    defparam shift_srl_150_1_LC_9_10_1.SEQ_MODE=4'b1000;
    defparam shift_srl_150_1_LC_9_10_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_150_1_LC_9_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54742),
            .lcout(shift_srl_150Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93067),
            .ce(N__55615),
            .sr(_gnd_net_));
    defparam shift_srl_150_2_LC_9_10_2.C_ON=1'b0;
    defparam shift_srl_150_2_LC_9_10_2.SEQ_MODE=4'b1000;
    defparam shift_srl_150_2_LC_9_10_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_150_2_LC_9_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54736),
            .lcout(shift_srl_150Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93067),
            .ce(N__55615),
            .sr(_gnd_net_));
    defparam shift_srl_150_3_LC_9_10_3.C_ON=1'b0;
    defparam shift_srl_150_3_LC_9_10_3.SEQ_MODE=4'b1000;
    defparam shift_srl_150_3_LC_9_10_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_150_3_LC_9_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54730),
            .lcout(shift_srl_150Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93067),
            .ce(N__55615),
            .sr(_gnd_net_));
    defparam shift_srl_150_4_LC_9_10_4.C_ON=1'b0;
    defparam shift_srl_150_4_LC_9_10_4.SEQ_MODE=4'b1000;
    defparam shift_srl_150_4_LC_9_10_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_150_4_LC_9_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54826),
            .lcout(shift_srl_150Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93067),
            .ce(N__55615),
            .sr(_gnd_net_));
    defparam shift_srl_150_5_LC_9_10_5.C_ON=1'b0;
    defparam shift_srl_150_5_LC_9_10_5.SEQ_MODE=4'b1000;
    defparam shift_srl_150_5_LC_9_10_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_150_5_LC_9_10_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54820),
            .lcout(shift_srl_150Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93067),
            .ce(N__55615),
            .sr(_gnd_net_));
    defparam shift_srl_150_6_LC_9_10_6.C_ON=1'b0;
    defparam shift_srl_150_6_LC_9_10_6.SEQ_MODE=4'b1000;
    defparam shift_srl_150_6_LC_9_10_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_150_6_LC_9_10_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54814),
            .lcout(shift_srl_150Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93067),
            .ce(N__55615),
            .sr(_gnd_net_));
    defparam shift_srl_150_7_LC_9_10_7.C_ON=1'b0;
    defparam shift_srl_150_7_LC_9_10_7.SEQ_MODE=4'b1000;
    defparam shift_srl_150_7_LC_9_10_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_150_7_LC_9_10_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54808),
            .lcout(shift_srl_150Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93067),
            .ce(N__55615),
            .sr(_gnd_net_));
    defparam shift_srl_150_10_LC_9_11_0.C_ON=1'b0;
    defparam shift_srl_150_10_LC_9_11_0.SEQ_MODE=4'b1000;
    defparam shift_srl_150_10_LC_9_11_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_150_10_LC_9_11_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54862),
            .lcout(shift_srl_150Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93051),
            .ce(N__55614),
            .sr(_gnd_net_));
    defparam shift_srl_150_11_LC_9_11_1.C_ON=1'b0;
    defparam shift_srl_150_11_LC_9_11_1.SEQ_MODE=4'b1000;
    defparam shift_srl_150_11_LC_9_11_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_150_11_LC_9_11_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54802),
            .lcout(shift_srl_150Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93051),
            .ce(N__55614),
            .sr(_gnd_net_));
    defparam shift_srl_150_12_LC_9_11_2.C_ON=1'b0;
    defparam shift_srl_150_12_LC_9_11_2.SEQ_MODE=4'b1000;
    defparam shift_srl_150_12_LC_9_11_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_150_12_LC_9_11_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54796),
            .lcout(shift_srl_150Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93051),
            .ce(N__55614),
            .sr(_gnd_net_));
    defparam shift_srl_150_13_LC_9_11_3.C_ON=1'b0;
    defparam shift_srl_150_13_LC_9_11_3.SEQ_MODE=4'b1000;
    defparam shift_srl_150_13_LC_9_11_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_150_13_LC_9_11_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54790),
            .lcout(shift_srl_150Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93051),
            .ce(N__55614),
            .sr(_gnd_net_));
    defparam shift_srl_150_14_LC_9_11_4.C_ON=1'b0;
    defparam shift_srl_150_14_LC_9_11_4.SEQ_MODE=4'b1000;
    defparam shift_srl_150_14_LC_9_11_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_150_14_LC_9_11_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54784),
            .lcout(shift_srl_150Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93051),
            .ce(N__55614),
            .sr(_gnd_net_));
    defparam shift_srl_150_15_LC_9_11_5.C_ON=1'b0;
    defparam shift_srl_150_15_LC_9_11_5.SEQ_MODE=4'b1000;
    defparam shift_srl_150_15_LC_9_11_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_150_15_LC_9_11_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54868),
            .lcout(shift_srl_150Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93051),
            .ce(N__55614),
            .sr(_gnd_net_));
    defparam shift_srl_150_9_LC_9_11_6.C_ON=1'b0;
    defparam shift_srl_150_9_LC_9_11_6.SEQ_MODE=4'b1000;
    defparam shift_srl_150_9_LC_9_11_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_150_9_LC_9_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54850),
            .lcout(shift_srl_150Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93051),
            .ce(N__55614),
            .sr(_gnd_net_));
    defparam shift_srl_150_8_LC_9_11_7.C_ON=1'b0;
    defparam shift_srl_150_8_LC_9_11_7.SEQ_MODE=4'b1000;
    defparam shift_srl_150_8_LC_9_11_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_150_8_LC_9_11_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54856),
            .lcout(shift_srl_150Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93051),
            .ce(N__55614),
            .sr(_gnd_net_));
    defparam shift_srl_147_5_LC_9_12_1.C_ON=1'b0;
    defparam shift_srl_147_5_LC_9_12_1.SEQ_MODE=4'b1000;
    defparam shift_srl_147_5_LC_9_12_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_147_5_LC_9_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55864),
            .lcout(shift_srl_147Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93036),
            .ce(N__55836),
            .sr(_gnd_net_));
    defparam shift_srl_147_6_LC_9_12_3.C_ON=1'b0;
    defparam shift_srl_147_6_LC_9_12_3.SEQ_MODE=4'b1000;
    defparam shift_srl_147_6_LC_9_12_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_147_6_LC_9_12_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54844),
            .lcout(shift_srl_147Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93036),
            .ce(N__55836),
            .sr(_gnd_net_));
    defparam shift_srl_147_7_LC_9_12_7.C_ON=1'b0;
    defparam shift_srl_147_7_LC_9_12_7.SEQ_MODE=4'b1000;
    defparam shift_srl_147_7_LC_9_12_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_147_7_LC_9_12_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54838),
            .lcout(shift_srl_147Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93036),
            .ce(N__55836),
            .sr(_gnd_net_));
    defparam shift_srl_146_5_LC_9_13_0.C_ON=1'b0;
    defparam shift_srl_146_5_LC_9_13_0.SEQ_MODE=4'b1000;
    defparam shift_srl_146_5_LC_9_13_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_146_5_LC_9_13_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54922),
            .lcout(shift_srl_146Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93021),
            .ce(N__56157),
            .sr(_gnd_net_));
    defparam shift_srl_146_6_LC_9_13_1.C_ON=1'b0;
    defparam shift_srl_146_6_LC_9_13_1.SEQ_MODE=4'b1000;
    defparam shift_srl_146_6_LC_9_13_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_146_6_LC_9_13_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54832),
            .lcout(shift_srl_146Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93021),
            .ce(N__56157),
            .sr(_gnd_net_));
    defparam shift_srl_146_3_LC_9_13_2.C_ON=1'b0;
    defparam shift_srl_146_3_LC_9_13_2.SEQ_MODE=4'b1000;
    defparam shift_srl_146_3_LC_9_13_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_146_3_LC_9_13_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55804),
            .lcout(shift_srl_146Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93021),
            .ce(N__56157),
            .sr(_gnd_net_));
    defparam shift_srl_146_4_LC_9_13_5.C_ON=1'b0;
    defparam shift_srl_146_4_LC_9_13_5.SEQ_MODE=4'b1000;
    defparam shift_srl_146_4_LC_9_13_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_146_4_LC_9_13_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54928),
            .lcout(shift_srl_146Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93021),
            .ce(N__56157),
            .sr(_gnd_net_));
    defparam shift_srl_146_10_LC_9_14_0.C_ON=1'b0;
    defparam shift_srl_146_10_LC_9_14_0.SEQ_MODE=4'b1000;
    defparam shift_srl_146_10_LC_9_14_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_146_10_LC_9_14_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54892),
            .lcout(shift_srl_146Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93008),
            .ce(N__56153),
            .sr(_gnd_net_));
    defparam shift_srl_146_11_LC_9_14_1.C_ON=1'b0;
    defparam shift_srl_146_11_LC_9_14_1.SEQ_MODE=4'b1000;
    defparam shift_srl_146_11_LC_9_14_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_146_11_LC_9_14_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54916),
            .lcout(shift_srl_146Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93008),
            .ce(N__56153),
            .sr(_gnd_net_));
    defparam shift_srl_146_12_LC_9_14_2.C_ON=1'b0;
    defparam shift_srl_146_12_LC_9_14_2.SEQ_MODE=4'b1000;
    defparam shift_srl_146_12_LC_9_14_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_146_12_LC_9_14_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54910),
            .lcout(shift_srl_146Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93008),
            .ce(N__56153),
            .sr(_gnd_net_));
    defparam shift_srl_146_13_LC_9_14_3.C_ON=1'b0;
    defparam shift_srl_146_13_LC_9_14_3.SEQ_MODE=4'b1000;
    defparam shift_srl_146_13_LC_9_14_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_146_13_LC_9_14_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54904),
            .lcout(shift_srl_146Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93008),
            .ce(N__56153),
            .sr(_gnd_net_));
    defparam shift_srl_146_14_LC_9_14_4.C_ON=1'b0;
    defparam shift_srl_146_14_LC_9_14_4.SEQ_MODE=4'b1000;
    defparam shift_srl_146_14_LC_9_14_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_146_14_LC_9_14_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54898),
            .lcout(shift_srl_146Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93008),
            .ce(N__56153),
            .sr(_gnd_net_));
    defparam shift_srl_146_9_LC_9_14_5.C_ON=1'b0;
    defparam shift_srl_146_9_LC_9_14_5.SEQ_MODE=4'b1000;
    defparam shift_srl_146_9_LC_9_14_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_146_9_LC_9_14_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54886),
            .lcout(shift_srl_146Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93008),
            .ce(N__56153),
            .sr(_gnd_net_));
    defparam shift_srl_146_8_LC_9_14_6.C_ON=1'b0;
    defparam shift_srl_146_8_LC_9_14_6.SEQ_MODE=4'b1000;
    defparam shift_srl_146_8_LC_9_14_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_146_8_LC_9_14_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54874),
            .lcout(shift_srl_146Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93008),
            .ce(N__56153),
            .sr(_gnd_net_));
    defparam shift_srl_146_7_LC_9_14_7.C_ON=1'b0;
    defparam shift_srl_146_7_LC_9_14_7.SEQ_MODE=4'b1000;
    defparam shift_srl_146_7_LC_9_14_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_146_7_LC_9_14_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54880),
            .lcout(shift_srl_146Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93008),
            .ce(N__56153),
            .sr(_gnd_net_));
    defparam shift_srl_27_0_LC_9_15_0.C_ON=1'b0;
    defparam shift_srl_27_0_LC_9_15_0.SEQ_MODE=4'b1000;
    defparam shift_srl_27_0_LC_9_15_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_27_0_LC_9_15_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71421),
            .lcout(shift_srl_27Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92994),
            .ce(N__55005),
            .sr(_gnd_net_));
    defparam shift_srl_27_1_LC_9_15_1.C_ON=1'b0;
    defparam shift_srl_27_1_LC_9_15_1.SEQ_MODE=4'b1000;
    defparam shift_srl_27_1_LC_9_15_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_27_1_LC_9_15_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54976),
            .lcout(shift_srl_27Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92994),
            .ce(N__55005),
            .sr(_gnd_net_));
    defparam shift_srl_27_2_LC_9_15_2.C_ON=1'b0;
    defparam shift_srl_27_2_LC_9_15_2.SEQ_MODE=4'b1000;
    defparam shift_srl_27_2_LC_9_15_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_27_2_LC_9_15_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54970),
            .lcout(shift_srl_27Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92994),
            .ce(N__55005),
            .sr(_gnd_net_));
    defparam shift_srl_27_3_LC_9_15_3.C_ON=1'b0;
    defparam shift_srl_27_3_LC_9_15_3.SEQ_MODE=4'b1000;
    defparam shift_srl_27_3_LC_9_15_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_27_3_LC_9_15_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54964),
            .lcout(shift_srl_27Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92994),
            .ce(N__55005),
            .sr(_gnd_net_));
    defparam shift_srl_27_4_LC_9_15_4.C_ON=1'b0;
    defparam shift_srl_27_4_LC_9_15_4.SEQ_MODE=4'b1000;
    defparam shift_srl_27_4_LC_9_15_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_27_4_LC_9_15_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54958),
            .lcout(shift_srl_27Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92994),
            .ce(N__55005),
            .sr(_gnd_net_));
    defparam shift_srl_27_5_LC_9_15_5.C_ON=1'b0;
    defparam shift_srl_27_5_LC_9_15_5.SEQ_MODE=4'b1000;
    defparam shift_srl_27_5_LC_9_15_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_27_5_LC_9_15_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54952),
            .lcout(shift_srl_27Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92994),
            .ce(N__55005),
            .sr(_gnd_net_));
    defparam shift_srl_27_6_LC_9_15_6.C_ON=1'b0;
    defparam shift_srl_27_6_LC_9_15_6.SEQ_MODE=4'b1000;
    defparam shift_srl_27_6_LC_9_15_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_27_6_LC_9_15_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54946),
            .lcout(shift_srl_27Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92994),
            .ce(N__55005),
            .sr(_gnd_net_));
    defparam shift_srl_27_7_LC_9_15_7.C_ON=1'b0;
    defparam shift_srl_27_7_LC_9_15_7.SEQ_MODE=4'b1000;
    defparam shift_srl_27_7_LC_9_15_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_27_7_LC_9_15_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54940),
            .lcout(shift_srl_27Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92994),
            .ce(N__55005),
            .sr(_gnd_net_));
    defparam shift_srl_27_10_LC_9_16_0.C_ON=1'b0;
    defparam shift_srl_27_10_LC_9_16_0.SEQ_MODE=4'b1000;
    defparam shift_srl_27_10_LC_9_16_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_27_10_LC_9_16_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55015),
            .lcout(shift_srl_27Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92981),
            .ce(N__55009),
            .sr(_gnd_net_));
    defparam shift_srl_27_11_LC_9_16_1.C_ON=1'b0;
    defparam shift_srl_27_11_LC_9_16_1.SEQ_MODE=4'b1000;
    defparam shift_srl_27_11_LC_9_16_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_27_11_LC_9_16_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54934),
            .lcout(shift_srl_27Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92981),
            .ce(N__55009),
            .sr(_gnd_net_));
    defparam shift_srl_27_12_LC_9_16_2.C_ON=1'b0;
    defparam shift_srl_27_12_LC_9_16_2.SEQ_MODE=4'b1000;
    defparam shift_srl_27_12_LC_9_16_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_27_12_LC_9_16_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55051),
            .lcout(shift_srl_27Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92981),
            .ce(N__55009),
            .sr(_gnd_net_));
    defparam shift_srl_27_13_LC_9_16_3.C_ON=1'b0;
    defparam shift_srl_27_13_LC_9_16_3.SEQ_MODE=4'b1000;
    defparam shift_srl_27_13_LC_9_16_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_27_13_LC_9_16_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55045),
            .lcout(shift_srl_27Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92981),
            .ce(N__55009),
            .sr(_gnd_net_));
    defparam shift_srl_27_8_LC_9_16_4.C_ON=1'b0;
    defparam shift_srl_27_8_LC_9_16_4.SEQ_MODE=4'b1000;
    defparam shift_srl_27_8_LC_9_16_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_27_8_LC_9_16_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55039),
            .lcout(shift_srl_27Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92981),
            .ce(N__55009),
            .sr(_gnd_net_));
    defparam shift_srl_27_15_LC_9_16_5.C_ON=1'b0;
    defparam shift_srl_27_15_LC_9_16_5.SEQ_MODE=4'b1000;
    defparam shift_srl_27_15_LC_9_16_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_27_15_LC_9_16_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55027),
            .lcout(shift_srl_27Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92981),
            .ce(N__55009),
            .sr(_gnd_net_));
    defparam shift_srl_27_14_LC_9_16_6.C_ON=1'b0;
    defparam shift_srl_27_14_LC_9_16_6.SEQ_MODE=4'b1000;
    defparam shift_srl_27_14_LC_9_16_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_27_14_LC_9_16_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55033),
            .lcout(shift_srl_27Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92981),
            .ce(N__55009),
            .sr(_gnd_net_));
    defparam shift_srl_27_9_LC_9_16_7.C_ON=1'b0;
    defparam shift_srl_27_9_LC_9_16_7.SEQ_MODE=4'b1000;
    defparam shift_srl_27_9_LC_9_16_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_27_9_LC_9_16_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55021),
            .lcout(shift_srl_27Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92981),
            .ce(N__55009),
            .sr(_gnd_net_));
    defparam shift_srl_149_10_LC_9_17_0.C_ON=1'b0;
    defparam shift_srl_149_10_LC_9_17_0.SEQ_MODE=4'b1000;
    defparam shift_srl_149_10_LC_9_17_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_149_10_LC_9_17_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55081),
            .lcout(shift_srl_149Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92960),
            .ce(N__55977),
            .sr(_gnd_net_));
    defparam shift_srl_149_11_LC_9_17_1.C_ON=1'b0;
    defparam shift_srl_149_11_LC_9_17_1.SEQ_MODE=4'b1000;
    defparam shift_srl_149_11_LC_9_17_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_149_11_LC_9_17_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54988),
            .lcout(shift_srl_149Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92960),
            .ce(N__55977),
            .sr(_gnd_net_));
    defparam shift_srl_149_12_LC_9_17_2.C_ON=1'b0;
    defparam shift_srl_149_12_LC_9_17_2.SEQ_MODE=4'b1000;
    defparam shift_srl_149_12_LC_9_17_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_149_12_LC_9_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54982),
            .lcout(shift_srl_149Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92960),
            .ce(N__55977),
            .sr(_gnd_net_));
    defparam shift_srl_149_13_LC_9_17_3.C_ON=1'b0;
    defparam shift_srl_149_13_LC_9_17_3.SEQ_MODE=4'b1000;
    defparam shift_srl_149_13_LC_9_17_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_149_13_LC_9_17_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55099),
            .lcout(shift_srl_149Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92960),
            .ce(N__55977),
            .sr(_gnd_net_));
    defparam shift_srl_149_14_LC_9_17_4.C_ON=1'b0;
    defparam shift_srl_149_14_LC_9_17_4.SEQ_MODE=4'b1000;
    defparam shift_srl_149_14_LC_9_17_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_149_14_LC_9_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55093),
            .lcout(shift_srl_149Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92960),
            .ce(N__55977),
            .sr(_gnd_net_));
    defparam shift_srl_149_15_LC_9_17_5.C_ON=1'b0;
    defparam shift_srl_149_15_LC_9_17_5.SEQ_MODE=4'b1000;
    defparam shift_srl_149_15_LC_9_17_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_149_15_LC_9_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55087),
            .lcout(shift_srl_149Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92960),
            .ce(N__55977),
            .sr(_gnd_net_));
    defparam shift_srl_149_9_LC_9_17_6.C_ON=1'b0;
    defparam shift_srl_149_9_LC_9_17_6.SEQ_MODE=4'b1000;
    defparam shift_srl_149_9_LC_9_17_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_149_9_LC_9_17_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55075),
            .lcout(shift_srl_149Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92960),
            .ce(N__55977),
            .sr(_gnd_net_));
    defparam shift_srl_149_0_LC_9_17_7.C_ON=1'b0;
    defparam shift_srl_149_0_LC_9_17_7.SEQ_MODE=4'b1000;
    defparam shift_srl_149_0_LC_9_17_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_149_0_LC_9_17_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56115),
            .lcout(shift_srl_149Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92960),
            .ce(N__55977),
            .sr(_gnd_net_));
    defparam shift_srl_149_8_LC_9_18_0.C_ON=1'b0;
    defparam shift_srl_149_8_LC_9_18_0.SEQ_MODE=4'b1000;
    defparam shift_srl_149_8_LC_9_18_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_149_8_LC_9_18_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55129),
            .lcout(shift_srl_149Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92982),
            .ce(N__55978),
            .sr(_gnd_net_));
    defparam shift_srl_149_1_LC_9_18_1.C_ON=1'b0;
    defparam shift_srl_149_1_LC_9_18_1.SEQ_MODE=4'b1000;
    defparam shift_srl_149_1_LC_9_18_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_149_1_LC_9_18_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55069),
            .lcout(shift_srl_149Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92982),
            .ce(N__55978),
            .sr(_gnd_net_));
    defparam shift_srl_149_2_LC_9_18_2.C_ON=1'b0;
    defparam shift_srl_149_2_LC_9_18_2.SEQ_MODE=4'b1000;
    defparam shift_srl_149_2_LC_9_18_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_149_2_LC_9_18_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55063),
            .lcout(shift_srl_149Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92982),
            .ce(N__55978),
            .sr(_gnd_net_));
    defparam shift_srl_149_3_LC_9_18_3.C_ON=1'b0;
    defparam shift_srl_149_3_LC_9_18_3.SEQ_MODE=4'b1000;
    defparam shift_srl_149_3_LC_9_18_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_149_3_LC_9_18_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55057),
            .lcout(shift_srl_149Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92982),
            .ce(N__55978),
            .sr(_gnd_net_));
    defparam shift_srl_149_4_LC_9_18_4.C_ON=1'b0;
    defparam shift_srl_149_4_LC_9_18_4.SEQ_MODE=4'b1000;
    defparam shift_srl_149_4_LC_9_18_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_149_4_LC_9_18_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55153),
            .lcout(shift_srl_149Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92982),
            .ce(N__55978),
            .sr(_gnd_net_));
    defparam shift_srl_149_5_LC_9_18_5.C_ON=1'b0;
    defparam shift_srl_149_5_LC_9_18_5.SEQ_MODE=4'b1000;
    defparam shift_srl_149_5_LC_9_18_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_149_5_LC_9_18_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55147),
            .lcout(shift_srl_149Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92982),
            .ce(N__55978),
            .sr(_gnd_net_));
    defparam shift_srl_149_6_LC_9_18_6.C_ON=1'b0;
    defparam shift_srl_149_6_LC_9_18_6.SEQ_MODE=4'b1000;
    defparam shift_srl_149_6_LC_9_18_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_149_6_LC_9_18_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55141),
            .lcout(shift_srl_149Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92982),
            .ce(N__55978),
            .sr(_gnd_net_));
    defparam shift_srl_149_7_LC_9_18_7.C_ON=1'b0;
    defparam shift_srl_149_7_LC_9_18_7.SEQ_MODE=4'b1000;
    defparam shift_srl_149_7_LC_9_18_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_149_7_LC_9_18_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55135),
            .lcout(shift_srl_149Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92982),
            .ce(N__55978),
            .sr(_gnd_net_));
    defparam shift_srl_123_10_LC_9_19_0.C_ON=1'b0;
    defparam shift_srl_123_10_LC_9_19_0.SEQ_MODE=4'b1000;
    defparam shift_srl_123_10_LC_9_19_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_123_10_LC_9_19_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55195),
            .lcout(shift_srl_123Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92995),
            .ce(N__56198),
            .sr(_gnd_net_));
    defparam shift_srl_123_11_LC_9_19_1.C_ON=1'b0;
    defparam shift_srl_123_11_LC_9_19_1.SEQ_MODE=4'b1000;
    defparam shift_srl_123_11_LC_9_19_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_123_11_LC_9_19_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55123),
            .lcout(shift_srl_123Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92995),
            .ce(N__56198),
            .sr(_gnd_net_));
    defparam shift_srl_123_12_LC_9_19_2.C_ON=1'b0;
    defparam shift_srl_123_12_LC_9_19_2.SEQ_MODE=4'b1000;
    defparam shift_srl_123_12_LC_9_19_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_123_12_LC_9_19_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55117),
            .lcout(shift_srl_123Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92995),
            .ce(N__56198),
            .sr(_gnd_net_));
    defparam shift_srl_123_13_LC_9_19_3.C_ON=1'b0;
    defparam shift_srl_123_13_LC_9_19_3.SEQ_MODE=4'b1000;
    defparam shift_srl_123_13_LC_9_19_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_123_13_LC_9_19_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55111),
            .lcout(shift_srl_123Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92995),
            .ce(N__56198),
            .sr(_gnd_net_));
    defparam shift_srl_123_14_LC_9_19_4.C_ON=1'b0;
    defparam shift_srl_123_14_LC_9_19_4.SEQ_MODE=4'b1000;
    defparam shift_srl_123_14_LC_9_19_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_123_14_LC_9_19_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55105),
            .lcout(shift_srl_123Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92995),
            .ce(N__56198),
            .sr(_gnd_net_));
    defparam shift_srl_123_9_LC_9_19_5.C_ON=1'b0;
    defparam shift_srl_123_9_LC_9_19_5.SEQ_MODE=4'b1000;
    defparam shift_srl_123_9_LC_9_19_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_123_9_LC_9_19_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55189),
            .lcout(shift_srl_123Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92995),
            .ce(N__56198),
            .sr(_gnd_net_));
    defparam shift_srl_123_8_LC_9_19_6.C_ON=1'b0;
    defparam shift_srl_123_8_LC_9_19_6.SEQ_MODE=4'b1000;
    defparam shift_srl_123_8_LC_9_19_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_123_8_LC_9_19_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55171),
            .lcout(shift_srl_123Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92995),
            .ce(N__56198),
            .sr(_gnd_net_));
    defparam shift_srl_123_7_LC_9_19_7.C_ON=1'b0;
    defparam shift_srl_123_7_LC_9_19_7.SEQ_MODE=4'b1000;
    defparam shift_srl_123_7_LC_9_19_7.LUT_INIT=16'b1100110011001100;
    LogicCell40 shift_srl_123_7_LC_9_19_7 (
            .in0(_gnd_net_),
            .in1(N__55183),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_123Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92995),
            .ce(N__56198),
            .sr(_gnd_net_));
    defparam shift_srl_121_RNI3T2O_15_LC_9_20_0.C_ON=1'b0;
    defparam shift_srl_121_RNI3T2O_15_LC_9_20_0.SEQ_MODE=4'b0000;
    defparam shift_srl_121_RNI3T2O_15_LC_9_20_0.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_121_RNI3T2O_15_LC_9_20_0 (
            .in0(N__78447),
            .in1(N__60298),
            .in2(N__90406),
            .in3(N__66456),
            .lcout(),
            .ltout(clk_en_0_a3_0_a2_sx_123_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_122_RNISJS2V_15_LC_9_20_1.C_ON=1'b0;
    defparam shift_srl_122_RNISJS2V_15_LC_9_20_1.SEQ_MODE=4'b0000;
    defparam shift_srl_122_RNISJS2V_15_LC_9_20_1.LUT_INIT=16'b0000010000000000;
    LogicCell40 shift_srl_122_RNISJS2V_15_LC_9_20_1 (
            .in0(N__60651),
            .in1(N__60131),
            .in2(N__55165),
            .in3(N__79496),
            .lcout(clk_en_123),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_118_15_LC_9_20_2.C_ON=1'b0;
    defparam shift_srl_118_15_LC_9_20_2.SEQ_MODE=4'b1000;
    defparam shift_srl_118_15_LC_9_20_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_118_15_LC_9_20_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55159),
            .lcout(shift_srl_118Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93009),
            .ce(N__60810),
            .sr(_gnd_net_));
    defparam shift_srl_124_RNI69LK_15_LC_9_20_3.C_ON=1'b0;
    defparam shift_srl_124_RNI69LK_15_LC_9_20_3.SEQ_MODE=4'b0000;
    defparam shift_srl_124_RNI69LK_15_LC_9_20_3.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_124_RNI69LK_15_LC_9_20_3 (
            .in0(N__66455),
            .in1(N__90163),
            .in2(N__60323),
            .in3(N__65440),
            .lcout(),
            .ltout(clk_en_0_a3_0_a2_sx_125_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_124_RNIV14MV_15_LC_9_20_4.C_ON=1'b0;
    defparam shift_srl_124_RNIV14MV_15_LC_9_20_4.SEQ_MODE=4'b0000;
    defparam shift_srl_124_RNIV14MV_15_LC_9_20_4.LUT_INIT=16'b0000000000001000;
    LogicCell40 shift_srl_124_RNIV14MV_15_LC_9_20_4 (
            .in0(N__79497),
            .in1(N__65310),
            .in2(N__55162),
            .in3(N__60652),
            .lcout(clk_en_125),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_118_14_LC_9_20_5.C_ON=1'b0;
    defparam shift_srl_118_14_LC_9_20_5.SEQ_MODE=4'b1000;
    defparam shift_srl_118_14_LC_9_20_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_118_14_LC_9_20_5 (
            .in0(N__55249),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_118Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93009),
            .ce(N__60810),
            .sr(_gnd_net_));
    defparam shift_srl_118_13_LC_9_20_6.C_ON=1'b0;
    defparam shift_srl_118_13_LC_9_20_6.SEQ_MODE=4'b1000;
    defparam shift_srl_118_13_LC_9_20_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_118_13_LC_9_20_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55243),
            .lcout(shift_srl_118Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93009),
            .ce(N__60810),
            .sr(_gnd_net_));
    defparam shift_srl_118_12_LC_9_20_7.C_ON=1'b0;
    defparam shift_srl_118_12_LC_9_20_7.SEQ_MODE=4'b1000;
    defparam shift_srl_118_12_LC_9_20_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_118_12_LC_9_20_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55432),
            .lcout(shift_srl_118Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93009),
            .ce(N__60810),
            .sr(_gnd_net_));
    defparam shift_srl_125_0_LC_9_21_0.C_ON=1'b0;
    defparam shift_srl_125_0_LC_9_21_0.SEQ_MODE=4'b1000;
    defparam shift_srl_125_0_LC_9_21_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_125_0_LC_9_21_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66014),
            .lcout(shift_srl_125Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93022),
            .ce(N__56373),
            .sr(_gnd_net_));
    defparam shift_srl_125_1_LC_9_21_1.C_ON=1'b0;
    defparam shift_srl_125_1_LC_9_21_1.SEQ_MODE=4'b1000;
    defparam shift_srl_125_1_LC_9_21_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_125_1_LC_9_21_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55237),
            .lcout(shift_srl_125Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93022),
            .ce(N__56373),
            .sr(_gnd_net_));
    defparam shift_srl_125_2_LC_9_21_2.C_ON=1'b0;
    defparam shift_srl_125_2_LC_9_21_2.SEQ_MODE=4'b1000;
    defparam shift_srl_125_2_LC_9_21_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_125_2_LC_9_21_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55231),
            .lcout(shift_srl_125Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93022),
            .ce(N__56373),
            .sr(_gnd_net_));
    defparam shift_srl_125_3_LC_9_21_3.C_ON=1'b0;
    defparam shift_srl_125_3_LC_9_21_3.SEQ_MODE=4'b1000;
    defparam shift_srl_125_3_LC_9_21_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_125_3_LC_9_21_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55225),
            .lcout(shift_srl_125Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93022),
            .ce(N__56373),
            .sr(_gnd_net_));
    defparam shift_srl_125_4_LC_9_21_4.C_ON=1'b0;
    defparam shift_srl_125_4_LC_9_21_4.SEQ_MODE=4'b1000;
    defparam shift_srl_125_4_LC_9_21_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_125_4_LC_9_21_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55219),
            .lcout(shift_srl_125Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93022),
            .ce(N__56373),
            .sr(_gnd_net_));
    defparam shift_srl_125_5_LC_9_21_5.C_ON=1'b0;
    defparam shift_srl_125_5_LC_9_21_5.SEQ_MODE=4'b1000;
    defparam shift_srl_125_5_LC_9_21_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_125_5_LC_9_21_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55213),
            .lcout(shift_srl_125Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93022),
            .ce(N__56373),
            .sr(_gnd_net_));
    defparam shift_srl_125_6_LC_9_21_6.C_ON=1'b0;
    defparam shift_srl_125_6_LC_9_21_6.SEQ_MODE=4'b1000;
    defparam shift_srl_125_6_LC_9_21_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_125_6_LC_9_21_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55207),
            .lcout(shift_srl_125Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93022),
            .ce(N__56373),
            .sr(_gnd_net_));
    defparam shift_srl_125_7_LC_9_21_7.C_ON=1'b0;
    defparam shift_srl_125_7_LC_9_21_7.SEQ_MODE=4'b1000;
    defparam shift_srl_125_7_LC_9_21_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_125_7_LC_9_21_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55201),
            .lcout(shift_srl_125Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93022),
            .ce(N__56373),
            .sr(_gnd_net_));
    defparam shift_srl_113_7_LC_9_22_0.C_ON=1'b0;
    defparam shift_srl_113_7_LC_9_22_0.SEQ_MODE=4'b1000;
    defparam shift_srl_113_7_LC_9_22_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_113_7_LC_9_22_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55291),
            .lcout(shift_srl_113Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93037),
            .ce(N__57752),
            .sr(_gnd_net_));
    defparam shift_srl_113_8_LC_9_22_1.C_ON=1'b0;
    defparam shift_srl_113_8_LC_9_22_1.SEQ_MODE=4'b1000;
    defparam shift_srl_113_8_LC_9_22_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_113_8_LC_9_22_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55297),
            .lcout(shift_srl_113Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93037),
            .ce(N__57752),
            .sr(_gnd_net_));
    defparam shift_srl_113_6_LC_9_22_4.C_ON=1'b0;
    defparam shift_srl_113_6_LC_9_22_4.SEQ_MODE=4'b1000;
    defparam shift_srl_113_6_LC_9_22_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_113_6_LC_9_22_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55255),
            .lcout(shift_srl_113Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93037),
            .ce(N__57752),
            .sr(_gnd_net_));
    defparam shift_srl_113_0_LC_9_23_1.C_ON=1'b0;
    defparam shift_srl_113_0_LC_9_23_1.SEQ_MODE=4'b1000;
    defparam shift_srl_113_0_LC_9_23_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_113_0_LC_9_23_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60449),
            .lcout(shift_srl_113Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93052),
            .ce(N__57760),
            .sr(_gnd_net_));
    defparam shift_srl_113_1_LC_9_23_2.C_ON=1'b0;
    defparam shift_srl_113_1_LC_9_23_2.SEQ_MODE=4'b1000;
    defparam shift_srl_113_1_LC_9_23_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_113_1_LC_9_23_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55285),
            .lcout(shift_srl_113Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93052),
            .ce(N__57760),
            .sr(_gnd_net_));
    defparam shift_srl_113_2_LC_9_23_3.C_ON=1'b0;
    defparam shift_srl_113_2_LC_9_23_3.SEQ_MODE=4'b1000;
    defparam shift_srl_113_2_LC_9_23_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_113_2_LC_9_23_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55279),
            .lcout(shift_srl_113Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93052),
            .ce(N__57760),
            .sr(_gnd_net_));
    defparam shift_srl_113_3_LC_9_23_4.C_ON=1'b0;
    defparam shift_srl_113_3_LC_9_23_4.SEQ_MODE=4'b1000;
    defparam shift_srl_113_3_LC_9_23_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_113_3_LC_9_23_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55273),
            .lcout(shift_srl_113Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93052),
            .ce(N__57760),
            .sr(_gnd_net_));
    defparam shift_srl_113_4_LC_9_23_5.C_ON=1'b0;
    defparam shift_srl_113_4_LC_9_23_5.SEQ_MODE=4'b1000;
    defparam shift_srl_113_4_LC_9_23_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_113_4_LC_9_23_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55267),
            .lcout(shift_srl_113Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93052),
            .ce(N__57760),
            .sr(_gnd_net_));
    defparam shift_srl_113_5_LC_9_23_6.C_ON=1'b0;
    defparam shift_srl_113_5_LC_9_23_6.SEQ_MODE=4'b1000;
    defparam shift_srl_113_5_LC_9_23_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_113_5_LC_9_23_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55261),
            .lcout(shift_srl_113Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93052),
            .ce(N__57760),
            .sr(_gnd_net_));
    defparam shift_srl_110_10_LC_9_24_0.C_ON=1'b0;
    defparam shift_srl_110_10_LC_9_24_0.SEQ_MODE=4'b1000;
    defparam shift_srl_110_10_LC_9_24_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_110_10_LC_9_24_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55324),
            .lcout(shift_srl_110Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93068),
            .ce(N__62448),
            .sr(_gnd_net_));
    defparam shift_srl_110_11_LC_9_24_1.C_ON=1'b0;
    defparam shift_srl_110_11_LC_9_24_1.SEQ_MODE=4'b1000;
    defparam shift_srl_110_11_LC_9_24_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_110_11_LC_9_24_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55348),
            .lcout(shift_srl_110Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93068),
            .ce(N__62448),
            .sr(_gnd_net_));
    defparam shift_srl_110_12_LC_9_24_2.C_ON=1'b0;
    defparam shift_srl_110_12_LC_9_24_2.SEQ_MODE=4'b1000;
    defparam shift_srl_110_12_LC_9_24_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_110_12_LC_9_24_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55342),
            .lcout(shift_srl_110Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93068),
            .ce(N__62448),
            .sr(_gnd_net_));
    defparam shift_srl_110_13_LC_9_24_3.C_ON=1'b0;
    defparam shift_srl_110_13_LC_9_24_3.SEQ_MODE=4'b1000;
    defparam shift_srl_110_13_LC_9_24_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_110_13_LC_9_24_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55336),
            .lcout(shift_srl_110Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93068),
            .ce(N__62448),
            .sr(_gnd_net_));
    defparam shift_srl_110_14_LC_9_24_4.C_ON=1'b0;
    defparam shift_srl_110_14_LC_9_24_4.SEQ_MODE=4'b1000;
    defparam shift_srl_110_14_LC_9_24_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_110_14_LC_9_24_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55330),
            .lcout(shift_srl_110Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93068),
            .ce(N__62448),
            .sr(_gnd_net_));
    defparam shift_srl_110_9_LC_9_24_5.C_ON=1'b0;
    defparam shift_srl_110_9_LC_9_24_5.SEQ_MODE=4'b1000;
    defparam shift_srl_110_9_LC_9_24_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_110_9_LC_9_24_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56584),
            .lcout(shift_srl_110Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93068),
            .ce(N__62448),
            .sr(_gnd_net_));
    defparam shift_srl_110_6_LC_9_24_6.C_ON=1'b0;
    defparam shift_srl_110_6_LC_9_24_6.SEQ_MODE=4'b1000;
    defparam shift_srl_110_6_LC_9_24_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_110_6_LC_9_24_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56482),
            .lcout(shift_srl_110Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93068),
            .ce(N__62448),
            .sr(_gnd_net_));
    defparam shift_srl_118_RNIT53B11_15_LC_9_25_0.C_ON=1'b0;
    defparam shift_srl_118_RNIT53B11_15_LC_9_25_0.SEQ_MODE=4'b0000;
    defparam shift_srl_118_RNIT53B11_15_LC_9_25_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_118_RNIT53B11_15_LC_9_25_0 (
            .in0(N__78509),
            .in1(N__65741),
            .in2(N__65379),
            .in3(N__62180),
            .lcout(rco_c_132),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_122_LC_9_25_3.C_ON=1'b0;
    defparam rco_obuf_RNO_122_LC_9_25_3.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_122_LC_9_25_3.LUT_INIT=16'b1000100000000000;
    LogicCell40 rco_obuf_RNO_122_LC_9_25_3 (
            .in0(N__78474),
            .in1(N__60136),
            .in2(_gnd_net_),
            .in3(N__78508),
            .lcout(rco_c_122),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_133_0_LC_9_25_4.C_ON=1'b0;
    defparam shift_srl_133_0_LC_9_25_4.SEQ_MODE=4'b1000;
    defparam shift_srl_133_0_LC_9_25_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_133_0_LC_9_25_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66259),
            .lcout(shift_srl_133Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93082),
            .ce(N__55378),
            .sr(_gnd_net_));
    defparam shift_srl_133_1_LC_9_25_5.C_ON=1'b0;
    defparam shift_srl_133_1_LC_9_25_5.SEQ_MODE=4'b1000;
    defparam shift_srl_133_1_LC_9_25_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_133_1_LC_9_25_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55411),
            .lcout(shift_srl_133Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93082),
            .ce(N__55378),
            .sr(_gnd_net_));
    defparam shift_srl_133_2_LC_9_25_6.C_ON=1'b0;
    defparam shift_srl_133_2_LC_9_25_6.SEQ_MODE=4'b1000;
    defparam shift_srl_133_2_LC_9_25_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_133_2_LC_9_25_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55405),
            .lcout(shift_srl_133Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93082),
            .ce(N__55378),
            .sr(_gnd_net_));
    defparam shift_srl_133_3_LC_9_25_7.C_ON=1'b0;
    defparam shift_srl_133_3_LC_9_25_7.SEQ_MODE=4'b1000;
    defparam shift_srl_133_3_LC_9_25_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_133_3_LC_9_25_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55399),
            .lcout(shift_srl_133Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93082),
            .ce(N__55378),
            .sr(_gnd_net_));
    defparam shift_srl_105_7_LC_9_26_0.C_ON=1'b0;
    defparam shift_srl_105_7_LC_9_26_0.SEQ_MODE=4'b1000;
    defparam shift_srl_105_7_LC_9_26_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_105_7_LC_9_26_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55360),
            .lcout(shift_srl_105Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93098),
            .ce(N__58055),
            .sr(_gnd_net_));
    defparam shift_srl_105_6_LC_9_26_5.C_ON=1'b0;
    defparam shift_srl_105_6_LC_9_26_5.SEQ_MODE=4'b1000;
    defparam shift_srl_105_6_LC_9_26_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_105_6_LC_9_26_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55354),
            .lcout(shift_srl_105Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93098),
            .ce(N__58055),
            .sr(_gnd_net_));
    defparam shift_srl_105_5_LC_9_26_6.C_ON=1'b0;
    defparam shift_srl_105_5_LC_9_26_6.SEQ_MODE=4'b1000;
    defparam shift_srl_105_5_LC_9_26_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_105_5_LC_9_26_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57943),
            .lcout(shift_srl_105Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93098),
            .ce(N__58055),
            .sr(_gnd_net_));
    defparam shift_srl_106_0_LC_9_27_0.C_ON=1'b0;
    defparam shift_srl_106_0_LC_9_27_0.SEQ_MODE=4'b1000;
    defparam shift_srl_106_0_LC_9_27_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_106_0_LC_9_27_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59242),
            .lcout(shift_srl_106Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93115),
            .ce(N__56728),
            .sr(_gnd_net_));
    defparam shift_srl_106_4_LC_9_27_1.C_ON=1'b0;
    defparam shift_srl_106_4_LC_9_27_1.SEQ_MODE=4'b1000;
    defparam shift_srl_106_4_LC_9_27_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_106_4_LC_9_27_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55468),
            .lcout(shift_srl_106Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93115),
            .ce(N__56728),
            .sr(_gnd_net_));
    defparam shift_srl_106_2_LC_9_27_2.C_ON=1'b0;
    defparam shift_srl_106_2_LC_9_27_2.SEQ_MODE=4'b1000;
    defparam shift_srl_106_2_LC_9_27_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_106_2_LC_9_27_2 (
            .in0(N__56734),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_106Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93115),
            .ce(N__56728),
            .sr(_gnd_net_));
    defparam shift_srl_106_3_LC_9_27_3.C_ON=1'b0;
    defparam shift_srl_106_3_LC_9_27_3.SEQ_MODE=4'b1000;
    defparam shift_srl_106_3_LC_9_27_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_106_3_LC_9_27_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55474),
            .lcout(shift_srl_106Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93115),
            .ce(N__56728),
            .sr(_gnd_net_));
    defparam shift_srl_106_8_LC_9_27_4.C_ON=1'b0;
    defparam shift_srl_106_8_LC_9_27_4.SEQ_MODE=4'b1000;
    defparam shift_srl_106_8_LC_9_27_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_106_8_LC_9_27_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55444),
            .lcout(shift_srl_106Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93115),
            .ce(N__56728),
            .sr(_gnd_net_));
    defparam shift_srl_106_5_LC_9_27_5.C_ON=1'b0;
    defparam shift_srl_106_5_LC_9_27_5.SEQ_MODE=4'b1000;
    defparam shift_srl_106_5_LC_9_27_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_106_5_LC_9_27_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55462),
            .lcout(shift_srl_106Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93115),
            .ce(N__56728),
            .sr(_gnd_net_));
    defparam shift_srl_106_6_LC_9_27_6.C_ON=1'b0;
    defparam shift_srl_106_6_LC_9_27_6.SEQ_MODE=4'b1000;
    defparam shift_srl_106_6_LC_9_27_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_106_6_LC_9_27_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55456),
            .lcout(shift_srl_106Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93115),
            .ce(N__56728),
            .sr(_gnd_net_));
    defparam shift_srl_106_7_LC_9_27_7.C_ON=1'b0;
    defparam shift_srl_106_7_LC_9_27_7.SEQ_MODE=4'b1000;
    defparam shift_srl_106_7_LC_9_27_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_106_7_LC_9_27_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55450),
            .lcout(shift_srl_106Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93115),
            .ce(N__56728),
            .sr(_gnd_net_));
    defparam shift_srl_118_10_LC_9_28_0.C_ON=1'b0;
    defparam shift_srl_118_10_LC_9_28_0.SEQ_MODE=4'b1000;
    defparam shift_srl_118_10_LC_9_28_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_118_10_LC_9_28_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55423),
            .lcout(shift_srl_118Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93135),
            .ce(N__60811),
            .sr(_gnd_net_));
    defparam shift_srl_118_11_LC_9_28_1.C_ON=1'b0;
    defparam shift_srl_118_11_LC_9_28_1.SEQ_MODE=4'b1000;
    defparam shift_srl_118_11_LC_9_28_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_118_11_LC_9_28_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55438),
            .lcout(shift_srl_118Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93135),
            .ce(N__60811),
            .sr(_gnd_net_));
    defparam shift_srl_118_9_LC_9_28_2.C_ON=1'b0;
    defparam shift_srl_118_9_LC_9_28_2.SEQ_MODE=4'b1000;
    defparam shift_srl_118_9_LC_9_28_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_118_9_LC_9_28_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55417),
            .lcout(shift_srl_118Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93135),
            .ce(N__60811),
            .sr(_gnd_net_));
    defparam shift_srl_118_8_LC_9_28_3.C_ON=1'b0;
    defparam shift_srl_118_8_LC_9_28_3.SEQ_MODE=4'b1000;
    defparam shift_srl_118_8_LC_9_28_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_118_8_LC_9_28_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59053),
            .lcout(shift_srl_118Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93135),
            .ce(N__60811),
            .sr(_gnd_net_));
    defparam shift_srl_108_RNIG1NLR_15_LC_9_32_1.C_ON=1'b0;
    defparam shift_srl_108_RNIG1NLR_15_LC_9_32_1.SEQ_MODE=4'b0000;
    defparam shift_srl_108_RNIG1NLR_15_LC_9_32_1.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_108_RNIG1NLR_15_LC_9_32_1 (
            .in0(N__62308),
            .in1(N__62373),
            .in2(_gnd_net_),
            .in3(N__56634),
            .lcout(rco_c_108),
            .ltout(rco_c_108_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_109_LC_9_32_2.C_ON=1'b0;
    defparam rco_obuf_RNO_109_LC_9_32_2.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_109_LC_9_32_2.LUT_INIT=16'b1010000010100000;
    LogicCell40 rco_obuf_RNO_109_LC_9_32_2 (
            .in0(N__62410),
            .in1(_gnd_net_),
            .in2(N__55534),
            .in3(_gnd_net_),
            .lcout(rco_c_109),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_107_LC_9_32_7.C_ON=1'b0;
    defparam rco_obuf_RNO_107_LC_9_32_7.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_107_LC_9_32_7.LUT_INIT=16'b1100110000000000;
    LogicCell40 rco_obuf_RNO_107_LC_9_32_7 (
            .in0(_gnd_net_),
            .in1(N__56633),
            .in2(_gnd_net_),
            .in3(N__62372),
            .lcout(rco_c_107),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_0_LC_10_5_0.C_ON=1'b0;
    defparam shift_srl_0_0_LC_10_5_0.SEQ_MODE=4'b1000;
    defparam shift_srl_0_0_LC_10_5_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_0_0_LC_10_5_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__89331),
            .lcout(shift_srl_0Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93156),
            .ce(N__57235),
            .sr(_gnd_net_));
    defparam shift_srl_0_1_LC_10_5_1.C_ON=1'b0;
    defparam shift_srl_0_1_LC_10_5_1.SEQ_MODE=4'b1000;
    defparam shift_srl_0_1_LC_10_5_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_0_1_LC_10_5_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55504),
            .lcout(shift_srl_0Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93156),
            .ce(N__57235),
            .sr(_gnd_net_));
    defparam shift_srl_0_2_LC_10_5_2.C_ON=1'b0;
    defparam shift_srl_0_2_LC_10_5_2.SEQ_MODE=4'b1000;
    defparam shift_srl_0_2_LC_10_5_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_0_2_LC_10_5_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55498),
            .lcout(shift_srl_0Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93156),
            .ce(N__57235),
            .sr(_gnd_net_));
    defparam shift_srl_0_3_LC_10_5_3.C_ON=1'b0;
    defparam shift_srl_0_3_LC_10_5_3.SEQ_MODE=4'b1000;
    defparam shift_srl_0_3_LC_10_5_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_0_3_LC_10_5_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55492),
            .lcout(shift_srl_0Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93156),
            .ce(N__57235),
            .sr(_gnd_net_));
    defparam shift_srl_0_4_LC_10_5_4.C_ON=1'b0;
    defparam shift_srl_0_4_LC_10_5_4.SEQ_MODE=4'b1000;
    defparam shift_srl_0_4_LC_10_5_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_0_4_LC_10_5_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55486),
            .lcout(shift_srl_0Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93156),
            .ce(N__57235),
            .sr(_gnd_net_));
    defparam shift_srl_0_5_LC_10_5_5.C_ON=1'b0;
    defparam shift_srl_0_5_LC_10_5_5.SEQ_MODE=4'b1000;
    defparam shift_srl_0_5_LC_10_5_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_0_5_LC_10_5_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55480),
            .lcout(shift_srl_0Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93156),
            .ce(N__57235),
            .sr(_gnd_net_));
    defparam shift_srl_0_7_LC_10_6_1.C_ON=1'b0;
    defparam shift_srl_0_7_LC_10_6_1.SEQ_MODE=4'b1000;
    defparam shift_srl_0_7_LC_10_6_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_0_7_LC_10_6_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55591),
            .lcout(shift_srl_0Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93138),
            .ce(N__57245),
            .sr(_gnd_net_));
    defparam shift_srl_0_8_LC_10_6_3.C_ON=1'b0;
    defparam shift_srl_0_8_LC_10_6_3.SEQ_MODE=4'b1000;
    defparam shift_srl_0_8_LC_10_6_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_0_8_LC_10_6_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55603),
            .lcout(shift_srl_0Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93138),
            .ce(N__57245),
            .sr(_gnd_net_));
    defparam shift_srl_0_10_LC_10_6_4.C_ON=1'b0;
    defparam shift_srl_0_10_LC_10_6_4.SEQ_MODE=4'b1000;
    defparam shift_srl_0_10_LC_10_6_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_0_10_LC_10_6_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55579),
            .lcout(shift_srl_0Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93138),
            .ce(N__57245),
            .sr(_gnd_net_));
    defparam shift_srl_0_6_LC_10_6_5.C_ON=1'b0;
    defparam shift_srl_0_6_LC_10_6_5.SEQ_MODE=4'b1000;
    defparam shift_srl_0_6_LC_10_6_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_0_6_LC_10_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55597),
            .lcout(shift_srl_0Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93138),
            .ce(N__57245),
            .sr(_gnd_net_));
    defparam shift_srl_0_9_LC_10_6_7.C_ON=1'b0;
    defparam shift_srl_0_9_LC_10_6_7.SEQ_MODE=4'b1000;
    defparam shift_srl_0_9_LC_10_6_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_0_9_LC_10_6_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55585),
            .lcout(shift_srl_0Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93138),
            .ce(N__57245),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_152_LC_10_8_2.C_ON=1'b0;
    defparam rco_obuf_RNO_152_LC_10_8_2.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_152_LC_10_8_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 rco_obuf_RNO_152_LC_10_8_2 (
            .in0(N__82216),
            .in1(N__66805),
            .in2(N__63259),
            .in3(N__63423),
            .lcout(rco_c_152),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_10_4_LC_10_9_0.C_ON=1'b0;
    defparam shift_srl_10_4_LC_10_9_0.SEQ_MODE=4'b1000;
    defparam shift_srl_10_4_LC_10_9_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_10_4_LC_10_9_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55651),
            .lcout(shift_srl_10Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93086),
            .ce(N__55641),
            .sr(_gnd_net_));
    defparam shift_srl_10_5_LC_10_9_3.C_ON=1'b0;
    defparam shift_srl_10_5_LC_10_9_3.SEQ_MODE=4'b1000;
    defparam shift_srl_10_5_LC_10_9_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_10_5_LC_10_9_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55558),
            .lcout(shift_srl_10Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93086),
            .ce(N__55641),
            .sr(_gnd_net_));
    defparam shift_srl_10_7_LC_10_9_4.C_ON=1'b0;
    defparam shift_srl_10_7_LC_10_9_4.SEQ_MODE=4'b1000;
    defparam shift_srl_10_7_LC_10_9_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_10_7_LC_10_9_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55738),
            .lcout(shift_srl_10Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93086),
            .ce(N__55641),
            .sr(_gnd_net_));
    defparam shift_srl_10_6_LC_10_9_7.C_ON=1'b0;
    defparam shift_srl_10_6_LC_10_9_7.SEQ_MODE=4'b1000;
    defparam shift_srl_10_6_LC_10_9_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_10_6_LC_10_9_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55744),
            .lcout(shift_srl_10Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93086),
            .ce(N__55641),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNI9EUH2_15_LC_10_10_0.C_ON=1'b0;
    defparam shift_srl_0_RNI9EUH2_15_LC_10_10_0.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNI9EUH2_15_LC_10_10_0.LUT_INIT=16'b1100110000000000;
    LogicCell40 shift_srl_0_RNI9EUH2_15_LC_10_10_0 (
            .in0(_gnd_net_),
            .in1(N__89616),
            .in2(_gnd_net_),
            .in3(N__69188),
            .lcout(clk_en_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_10_0_LC_10_10_1.C_ON=1'b0;
    defparam shift_srl_10_0_LC_10_10_1.SEQ_MODE=4'b1000;
    defparam shift_srl_10_0_LC_10_10_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_10_0_LC_10_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55709),
            .lcout(shift_srl_10Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93070),
            .ce(N__55640),
            .sr(_gnd_net_));
    defparam shift_srl_10_1_LC_10_10_2.C_ON=1'b0;
    defparam shift_srl_10_1_LC_10_10_2.SEQ_MODE=4'b1000;
    defparam shift_srl_10_1_LC_10_10_2.LUT_INIT=16'b1100110011001100;
    LogicCell40 shift_srl_10_1_LC_10_10_2 (
            .in0(_gnd_net_),
            .in1(N__55669),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_10Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93070),
            .ce(N__55640),
            .sr(_gnd_net_));
    defparam shift_srl_10_2_LC_10_10_3.C_ON=1'b0;
    defparam shift_srl_10_2_LC_10_10_3.SEQ_MODE=4'b1000;
    defparam shift_srl_10_2_LC_10_10_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_10_2_LC_10_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55663),
            .lcout(shift_srl_10Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93070),
            .ce(N__55640),
            .sr(_gnd_net_));
    defparam shift_srl_10_3_LC_10_10_4.C_ON=1'b0;
    defparam shift_srl_10_3_LC_10_10_4.SEQ_MODE=4'b1000;
    defparam shift_srl_10_3_LC_10_10_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_10_3_LC_10_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55657),
            .lcout(shift_srl_10Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93070),
            .ce(N__55640),
            .sr(_gnd_net_));
    defparam shift_srl_147_15_LC_10_11_0.C_ON=1'b0;
    defparam shift_srl_147_15_LC_10_11_0.SEQ_MODE=4'b1000;
    defparam shift_srl_147_15_LC_10_11_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_147_15_LC_10_11_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55798),
            .lcout(shift_srl_147Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93054),
            .ce(N__55840),
            .sr(_gnd_net_));
    defparam shift_srl_149_RNIU42S_15_LC_10_11_1.C_ON=1'b0;
    defparam shift_srl_149_RNIU42S_15_LC_10_11_1.SEQ_MODE=4'b0000;
    defparam shift_srl_149_RNIU42S_15_LC_10_11_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_149_RNIU42S_15_LC_10_11_1 (
            .in0(N__56982),
            .in1(N__56119),
            .in2(N__70718),
            .in3(N__57019),
            .lcout(shift_srl_149_RNIU42SZ0Z_15),
            .ltout(shift_srl_149_RNIU42SZ0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNILB5P51_15_LC_10_11_2.C_ON=1'b0;
    defparam shift_srl_0_RNILB5P51_15_LC_10_11_2.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNILB5P51_15_LC_10_11_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNILB5P51_15_LC_10_11_2 (
            .in0(N__89618),
            .in1(N__77826),
            .in2(N__55618),
            .in3(N__79563),
            .lcout(clk_en_150),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_147_14_LC_10_11_3.C_ON=1'b0;
    defparam shift_srl_147_14_LC_10_11_3.SEQ_MODE=4'b1000;
    defparam shift_srl_147_14_LC_10_11_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_147_14_LC_10_11_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55792),
            .lcout(shift_srl_147Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93054),
            .ce(N__55840),
            .sr(_gnd_net_));
    defparam shift_srl_147_13_LC_10_11_4.C_ON=1'b0;
    defparam shift_srl_147_13_LC_10_11_4.SEQ_MODE=4'b1000;
    defparam shift_srl_147_13_LC_10_11_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_147_13_LC_10_11_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55786),
            .lcout(shift_srl_147Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93054),
            .ce(N__55840),
            .sr(_gnd_net_));
    defparam shift_srl_147_12_LC_10_11_5.C_ON=1'b0;
    defparam shift_srl_147_12_LC_10_11_5.SEQ_MODE=4'b1000;
    defparam shift_srl_147_12_LC_10_11_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_147_12_LC_10_11_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55780),
            .lcout(shift_srl_147Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93054),
            .ce(N__55840),
            .sr(_gnd_net_));
    defparam shift_srl_147_11_LC_10_11_6.C_ON=1'b0;
    defparam shift_srl_147_11_LC_10_11_6.SEQ_MODE=4'b1000;
    defparam shift_srl_147_11_LC_10_11_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_147_11_LC_10_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55774),
            .lcout(shift_srl_147Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93054),
            .ce(N__55840),
            .sr(_gnd_net_));
    defparam shift_srl_147_10_LC_10_11_7.C_ON=1'b0;
    defparam shift_srl_147_10_LC_10_11_7.SEQ_MODE=4'b1000;
    defparam shift_srl_147_10_LC_10_11_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_147_10_LC_10_11_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55858),
            .lcout(shift_srl_147Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93054),
            .ce(N__55840),
            .sr(_gnd_net_));
    defparam shift_srl_147_0_LC_10_12_0.C_ON=1'b0;
    defparam shift_srl_147_0_LC_10_12_0.SEQ_MODE=4'b1000;
    defparam shift_srl_147_0_LC_10_12_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_147_0_LC_10_12_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57023),
            .lcout(shift_srl_147Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93039),
            .ce(N__55832),
            .sr(_gnd_net_));
    defparam shift_srl_147_1_LC_10_12_1.C_ON=1'b0;
    defparam shift_srl_147_1_LC_10_12_1.SEQ_MODE=4'b1000;
    defparam shift_srl_147_1_LC_10_12_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_147_1_LC_10_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55768),
            .lcout(shift_srl_147Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93039),
            .ce(N__55832),
            .sr(_gnd_net_));
    defparam shift_srl_147_2_LC_10_12_2.C_ON=1'b0;
    defparam shift_srl_147_2_LC_10_12_2.SEQ_MODE=4'b1000;
    defparam shift_srl_147_2_LC_10_12_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_147_2_LC_10_12_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55762),
            .lcout(shift_srl_147Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93039),
            .ce(N__55832),
            .sr(_gnd_net_));
    defparam shift_srl_147_3_LC_10_12_3.C_ON=1'b0;
    defparam shift_srl_147_3_LC_10_12_3.SEQ_MODE=4'b1000;
    defparam shift_srl_147_3_LC_10_12_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_147_3_LC_10_12_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55756),
            .lcout(shift_srl_147Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93039),
            .ce(N__55832),
            .sr(_gnd_net_));
    defparam shift_srl_147_4_LC_10_12_4.C_ON=1'b0;
    defparam shift_srl_147_4_LC_10_12_4.SEQ_MODE=4'b1000;
    defparam shift_srl_147_4_LC_10_12_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_147_4_LC_10_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55750),
            .lcout(shift_srl_147Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93039),
            .ce(N__55832),
            .sr(_gnd_net_));
    defparam shift_srl_147_9_LC_10_12_5.C_ON=1'b0;
    defparam shift_srl_147_9_LC_10_12_5.SEQ_MODE=4'b1000;
    defparam shift_srl_147_9_LC_10_12_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_147_9_LC_10_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55846),
            .lcout(shift_srl_147Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93039),
            .ce(N__55832),
            .sr(_gnd_net_));
    defparam shift_srl_147_8_LC_10_12_7.C_ON=1'b0;
    defparam shift_srl_147_8_LC_10_12_7.SEQ_MODE=4'b1000;
    defparam shift_srl_147_8_LC_10_12_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_147_8_LC_10_12_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55852),
            .lcout(shift_srl_147Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93039),
            .ce(N__55832),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIV3TP61_15_LC_10_13_0.C_ON=1'b0;
    defparam shift_srl_0_RNIV3TP61_15_LC_10_13_0.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIV3TP61_15_LC_10_13_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNIV3TP61_15_LC_10_13_0 (
            .in0(N__79549),
            .in1(N__89613),
            .in2(N__77825),
            .in3(N__82288),
            .lcout(clk_en_154),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIN63T41_15_LC_10_13_1.C_ON=1'b0;
    defparam shift_srl_0_RNIN63T41_15_LC_10_13_1.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIN63T41_15_LC_10_13_1.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_0_RNIN63T41_15_LC_10_13_1 (
            .in0(N__89614),
            .in1(N__77805),
            .in2(_gnd_net_),
            .in3(N__79548),
            .lcout(clk_en_146),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_146_RNITHQT41_15_LC_10_13_2.C_ON=1'b0;
    defparam shift_srl_146_RNITHQT41_15_LC_10_13_2.SEQ_MODE=4'b0000;
    defparam shift_srl_146_RNITHQT41_15_LC_10_13_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_146_RNITHQT41_15_LC_10_13_2 (
            .in0(N__79550),
            .in1(N__89615),
            .in2(N__77824),
            .in3(N__70716),
            .lcout(clk_en_147),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_146_0_LC_10_13_3.C_ON=1'b0;
    defparam shift_srl_146_0_LC_10_13_3.SEQ_MODE=4'b1000;
    defparam shift_srl_146_0_LC_10_13_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_146_0_LC_10_13_3 (
            .in0(N__70717),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_146Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93024),
            .ce(N__56140),
            .sr(_gnd_net_));
    defparam shift_srl_146_1_LC_10_13_4.C_ON=1'b0;
    defparam shift_srl_146_1_LC_10_13_4.SEQ_MODE=4'b1000;
    defparam shift_srl_146_1_LC_10_13_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_146_1_LC_10_13_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55816),
            .lcout(shift_srl_146Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93024),
            .ce(N__56140),
            .sr(_gnd_net_));
    defparam shift_srl_146_2_LC_10_13_5.C_ON=1'b0;
    defparam shift_srl_146_2_LC_10_13_5.SEQ_MODE=4'b1000;
    defparam shift_srl_146_2_LC_10_13_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_146_2_LC_10_13_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55810),
            .lcout(shift_srl_146Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93024),
            .ce(N__56140),
            .sr(_gnd_net_));
    defparam shift_srl_160_10_LC_10_14_0.C_ON=1'b0;
    defparam shift_srl_160_10_LC_10_14_0.SEQ_MODE=4'b1000;
    defparam shift_srl_160_10_LC_10_14_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_160_10_LC_10_14_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55882),
            .lcout(shift_srl_160Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93011),
            .ce(N__57274),
            .sr(_gnd_net_));
    defparam shift_srl_160_11_LC_10_14_1.C_ON=1'b0;
    defparam shift_srl_160_11_LC_10_14_1.SEQ_MODE=4'b1000;
    defparam shift_srl_160_11_LC_10_14_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_160_11_LC_10_14_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55906),
            .lcout(shift_srl_160Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93011),
            .ce(N__57274),
            .sr(_gnd_net_));
    defparam shift_srl_160_4_LC_10_14_2.C_ON=1'b0;
    defparam shift_srl_160_4_LC_10_14_2.SEQ_MODE=4'b1000;
    defparam shift_srl_160_4_LC_10_14_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_160_4_LC_10_14_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55900),
            .lcout(shift_srl_160Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93011),
            .ce(N__57274),
            .sr(_gnd_net_));
    defparam shift_srl_160_3_LC_10_14_3.C_ON=1'b0;
    defparam shift_srl_160_3_LC_10_14_3.SEQ_MODE=4'b1000;
    defparam shift_srl_160_3_LC_10_14_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_160_3_LC_10_14_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55888),
            .lcout(shift_srl_160Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93011),
            .ce(N__57274),
            .sr(_gnd_net_));
    defparam shift_srl_160_1_LC_10_14_4.C_ON=1'b0;
    defparam shift_srl_160_1_LC_10_14_4.SEQ_MODE=4'b1000;
    defparam shift_srl_160_1_LC_10_14_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_160_1_LC_10_14_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55960),
            .lcout(shift_srl_160Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93011),
            .ce(N__57274),
            .sr(_gnd_net_));
    defparam shift_srl_160_2_LC_10_14_5.C_ON=1'b0;
    defparam shift_srl_160_2_LC_10_14_5.SEQ_MODE=4'b1000;
    defparam shift_srl_160_2_LC_10_14_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_160_2_LC_10_14_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55894),
            .lcout(shift_srl_160Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93011),
            .ce(N__57274),
            .sr(_gnd_net_));
    defparam shift_srl_160_9_LC_10_14_6.C_ON=1'b0;
    defparam shift_srl_160_9_LC_10_14_6.SEQ_MODE=4'b1000;
    defparam shift_srl_160_9_LC_10_14_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_160_9_LC_10_14_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55876),
            .lcout(shift_srl_160Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93011),
            .ce(N__57274),
            .sr(_gnd_net_));
    defparam shift_srl_160_8_LC_10_14_7.C_ON=1'b0;
    defparam shift_srl_160_8_LC_10_14_7.SEQ_MODE=4'b1000;
    defparam shift_srl_160_8_LC_10_14_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_160_8_LC_10_14_7 (
            .in0(N__55966),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_160Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93011),
            .ce(N__57274),
            .sr(_gnd_net_));
    defparam shift_srl_160_15_LC_10_15_0.C_ON=1'b0;
    defparam shift_srl_160_15_LC_10_15_0.SEQ_MODE=4'b1000;
    defparam shift_srl_160_15_LC_10_15_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_160_15_LC_10_15_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55870),
            .lcout(shift_srl_160Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92997),
            .ce(N__57270),
            .sr(_gnd_net_));
    defparam shift_srl_160_14_LC_10_15_1.C_ON=1'b0;
    defparam shift_srl_160_14_LC_10_15_1.SEQ_MODE=4'b1000;
    defparam shift_srl_160_14_LC_10_15_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_160_14_LC_10_15_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55924),
            .lcout(shift_srl_160Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92997),
            .ce(N__57270),
            .sr(_gnd_net_));
    defparam shift_srl_160_7_LC_10_15_2.C_ON=1'b0;
    defparam shift_srl_160_7_LC_10_15_2.SEQ_MODE=4'b1000;
    defparam shift_srl_160_7_LC_10_15_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_160_7_LC_10_15_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55936),
            .lcout(shift_srl_160Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92997),
            .ce(N__57270),
            .sr(_gnd_net_));
    defparam shift_srl_160_0_LC_10_15_3.C_ON=1'b0;
    defparam shift_srl_160_0_LC_10_15_3.SEQ_MODE=4'b1000;
    defparam shift_srl_160_0_LC_10_15_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_160_0_LC_10_15_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77420),
            .lcout(shift_srl_160Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92997),
            .ce(N__57270),
            .sr(_gnd_net_));
    defparam shift_srl_160_12_LC_10_15_4.C_ON=1'b0;
    defparam shift_srl_160_12_LC_10_15_4.SEQ_MODE=4'b1000;
    defparam shift_srl_160_12_LC_10_15_4.LUT_INIT=16'b1100110011001100;
    LogicCell40 shift_srl_160_12_LC_10_15_4 (
            .in0(_gnd_net_),
            .in1(N__55954),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_160Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92997),
            .ce(N__57270),
            .sr(_gnd_net_));
    defparam shift_srl_160_5_LC_10_15_5.C_ON=1'b0;
    defparam shift_srl_160_5_LC_10_15_5.SEQ_MODE=4'b1000;
    defparam shift_srl_160_5_LC_10_15_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_160_5_LC_10_15_5 (
            .in0(N__55948),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_160Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92997),
            .ce(N__57270),
            .sr(_gnd_net_));
    defparam shift_srl_160_6_LC_10_15_6.C_ON=1'b0;
    defparam shift_srl_160_6_LC_10_15_6.SEQ_MODE=4'b1000;
    defparam shift_srl_160_6_LC_10_15_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_160_6_LC_10_15_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55942),
            .lcout(shift_srl_160Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92997),
            .ce(N__57270),
            .sr(_gnd_net_));
    defparam shift_srl_160_13_LC_10_15_7.C_ON=1'b0;
    defparam shift_srl_160_13_LC_10_15_7.SEQ_MODE=4'b1000;
    defparam shift_srl_160_13_LC_10_15_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_160_13_LC_10_15_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55930),
            .lcout(shift_srl_160Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92997),
            .ce(N__57270),
            .sr(_gnd_net_));
    defparam shift_srl_161_10_LC_10_16_0.C_ON=1'b0;
    defparam shift_srl_161_10_LC_10_16_0.SEQ_MODE=4'b1000;
    defparam shift_srl_161_10_LC_10_16_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_161_10_LC_10_16_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56038),
            .lcout(shift_srl_161Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92984),
            .ce(N__57421),
            .sr(_gnd_net_));
    defparam shift_srl_161_11_LC_10_16_1.C_ON=1'b0;
    defparam shift_srl_161_11_LC_10_16_1.SEQ_MODE=4'b1000;
    defparam shift_srl_161_11_LC_10_16_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_161_11_LC_10_16_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55918),
            .lcout(shift_srl_161Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92984),
            .ce(N__57421),
            .sr(_gnd_net_));
    defparam shift_srl_161_12_LC_10_16_2.C_ON=1'b0;
    defparam shift_srl_161_12_LC_10_16_2.SEQ_MODE=4'b1000;
    defparam shift_srl_161_12_LC_10_16_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_161_12_LC_10_16_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55912),
            .lcout(shift_srl_161Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92984),
            .ce(N__57421),
            .sr(_gnd_net_));
    defparam shift_srl_161_13_LC_10_16_3.C_ON=1'b0;
    defparam shift_srl_161_13_LC_10_16_3.SEQ_MODE=4'b1000;
    defparam shift_srl_161_13_LC_10_16_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_161_13_LC_10_16_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56056),
            .lcout(shift_srl_161Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92984),
            .ce(N__57421),
            .sr(_gnd_net_));
    defparam shift_srl_161_14_LC_10_16_4.C_ON=1'b0;
    defparam shift_srl_161_14_LC_10_16_4.SEQ_MODE=4'b1000;
    defparam shift_srl_161_14_LC_10_16_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_161_14_LC_10_16_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56050),
            .lcout(shift_srl_161Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92984),
            .ce(N__57421),
            .sr(_gnd_net_));
    defparam shift_srl_161_15_LC_10_16_5.C_ON=1'b0;
    defparam shift_srl_161_15_LC_10_16_5.SEQ_MODE=4'b1000;
    defparam shift_srl_161_15_LC_10_16_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_161_15_LC_10_16_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56044),
            .lcout(shift_srl_161Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92984),
            .ce(N__57421),
            .sr(_gnd_net_));
    defparam shift_srl_161_9_LC_10_16_6.C_ON=1'b0;
    defparam shift_srl_161_9_LC_10_16_6.SEQ_MODE=4'b1000;
    defparam shift_srl_161_9_LC_10_16_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_161_9_LC_10_16_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56032),
            .lcout(shift_srl_161Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92984),
            .ce(N__57421),
            .sr(_gnd_net_));
    defparam shift_srl_161_8_LC_10_16_7.C_ON=1'b0;
    defparam shift_srl_161_8_LC_10_16_7.SEQ_MODE=4'b1000;
    defparam shift_srl_161_8_LC_10_16_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_161_8_LC_10_16_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57427),
            .lcout(shift_srl_161Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92984),
            .ce(N__57421),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_148_LC_10_17_0.C_ON=1'b0;
    defparam rco_obuf_RNO_148_LC_10_17_0.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_148_LC_10_17_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 rco_obuf_RNO_148_LC_10_17_0 (
            .in0(N__57027),
            .in1(N__70693),
            .in2(N__82212),
            .in3(N__56981),
            .lcout(rco_c_148),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_147_LC_10_17_1.C_ON=1'b0;
    defparam rco_obuf_RNO_147_LC_10_17_1.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_147_LC_10_17_1.LUT_INIT=16'b1000100000000000;
    LogicCell40 rco_obuf_RNO_147_LC_10_17_1 (
            .in0(N__70692),
            .in1(N__82194),
            .in2(_gnd_net_),
            .in3(N__57026),
            .lcout(rco_c_147),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_148_RNIGPIF_15_LC_10_17_2.C_ON=1'b0;
    defparam shift_srl_148_RNIGPIF_15_LC_10_17_2.SEQ_MODE=4'b0000;
    defparam shift_srl_148_RNIGPIF_15_LC_10_17_2.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_148_RNIGPIF_15_LC_10_17_2 (
            .in0(N__57025),
            .in1(N__70691),
            .in2(N__56989),
            .in3(N__89617),
            .lcout(),
            .ltout(clk_en_0_a3_0_a2_sx_149_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_148_RNICKRB51_15_LC_10_17_3.C_ON=1'b0;
    defparam shift_srl_148_RNICKRB51_15_LC_10_17_3.SEQ_MODE=4'b0000;
    defparam shift_srl_148_RNICKRB51_15_LC_10_17_3.LUT_INIT=16'b0000110000000000;
    LogicCell40 shift_srl_148_RNICKRB51_15_LC_10_17_3 (
            .in0(_gnd_net_),
            .in1(N__77774),
            .in2(N__55981),
            .in3(N__79511),
            .lcout(clk_en_149),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_146_15_LC_10_17_4.C_ON=1'b0;
    defparam shift_srl_146_15_LC_10_17_4.SEQ_MODE=4'b1000;
    defparam shift_srl_146_15_LC_10_17_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_146_15_LC_10_17_4 (
            .in0(N__56167),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_146Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92971),
            .ce(N__56158),
            .sr(_gnd_net_));
    defparam shift_srl_150_RNIPH7T_15_LC_10_17_5.C_ON=1'b0;
    defparam shift_srl_150_RNIPH7T_15_LC_10_17_5.SEQ_MODE=4'b0000;
    defparam shift_srl_150_RNIPH7T_15_LC_10_17_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_150_RNIPH7T_15_LC_10_17_5 (
            .in0(N__56980),
            .in1(N__56111),
            .in2(N__56095),
            .in3(N__57024),
            .lcout(),
            .ltout(shift_srl_150_RNIPH7TZ0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_146_RNIVSUT_15_LC_10_17_6.C_ON=1'b0;
    defparam shift_srl_146_RNIVSUT_15_LC_10_17_6.SEQ_MODE=4'b0000;
    defparam shift_srl_146_RNIVSUT_15_LC_10_17_6.LUT_INIT=16'b1111000010101010;
    LogicCell40 shift_srl_146_RNIVSUT_15_LC_10_17_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__56074),
            .in3(N__70690),
            .lcout(shift_srl_146_RNIVSUTZ0Z_15),
            .ltout(shift_srl_146_RNIVSUTZ0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_153_RNI8TPS1_15_LC_10_17_7.C_ON=1'b0;
    defparam shift_srl_153_RNI8TPS1_15_LC_10_17_7.SEQ_MODE=4'b0000;
    defparam shift_srl_153_RNI8TPS1_15_LC_10_17_7.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_153_RNI8TPS1_15_LC_10_17_7 (
            .in0(N__61645),
            .in1(N__63252),
            .in2(N__56071),
            .in3(N__63406),
            .lcout(rco_int_0_a2_0_a2_0_153),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_126_10_LC_10_18_0.C_ON=1'b0;
    defparam shift_srl_126_10_LC_10_18_0.SEQ_MODE=4'b1000;
    defparam shift_srl_126_10_LC_10_18_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_126_10_LC_10_18_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56302),
            .lcout(shift_srl_126Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92985),
            .ce(N__57547),
            .sr(_gnd_net_));
    defparam shift_srl_126_7_LC_10_18_1.C_ON=1'b0;
    defparam shift_srl_126_7_LC_10_18_1.SEQ_MODE=4'b1000;
    defparam shift_srl_126_7_LC_10_18_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_126_7_LC_10_18_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57664),
            .lcout(shift_srl_126Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92985),
            .ce(N__57547),
            .sr(_gnd_net_));
    defparam shift_srl_126_11_LC_10_18_2.C_ON=1'b0;
    defparam shift_srl_126_11_LC_10_18_2.SEQ_MODE=4'b1000;
    defparam shift_srl_126_11_LC_10_18_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_126_11_LC_10_18_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56068),
            .lcout(shift_srl_126Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92985),
            .ce(N__57547),
            .sr(_gnd_net_));
    defparam shift_srl_126_12_LC_10_18_3.C_ON=1'b0;
    defparam shift_srl_126_12_LC_10_18_3.SEQ_MODE=4'b1000;
    defparam shift_srl_126_12_LC_10_18_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_126_12_LC_10_18_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56062),
            .lcout(shift_srl_126Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92985),
            .ce(N__57547),
            .sr(_gnd_net_));
    defparam shift_srl_126_0_LC_10_18_4.C_ON=1'b0;
    defparam shift_srl_126_0_LC_10_18_4.SEQ_MODE=4'b1000;
    defparam shift_srl_126_0_LC_10_18_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_126_0_LC_10_18_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66061),
            .lcout(shift_srl_126Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92985),
            .ce(N__57547),
            .sr(_gnd_net_));
    defparam shift_srl_126_15_LC_10_18_5.C_ON=1'b0;
    defparam shift_srl_126_15_LC_10_18_5.SEQ_MODE=4'b1000;
    defparam shift_srl_126_15_LC_10_18_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_126_15_LC_10_18_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57652),
            .lcout(shift_srl_126Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92985),
            .ce(N__57547),
            .sr(_gnd_net_));
    defparam shift_srl_126_9_LC_10_18_6.C_ON=1'b0;
    defparam shift_srl_126_9_LC_10_18_6.SEQ_MODE=4'b1000;
    defparam shift_srl_126_9_LC_10_18_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_126_9_LC_10_18_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56290),
            .lcout(shift_srl_126Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92985),
            .ce(N__57547),
            .sr(_gnd_net_));
    defparam shift_srl_126_8_LC_10_18_7.C_ON=1'b0;
    defparam shift_srl_126_8_LC_10_18_7.SEQ_MODE=4'b1000;
    defparam shift_srl_126_8_LC_10_18_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_126_8_LC_10_18_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56296),
            .lcout(shift_srl_126Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92985),
            .ce(N__57547),
            .sr(_gnd_net_));
    defparam shift_srl_118_RNI43UI1_15_LC_10_19_0.C_ON=1'b0;
    defparam shift_srl_118_RNI43UI1_15_LC_10_19_0.SEQ_MODE=4'b0000;
    defparam shift_srl_118_RNI43UI1_15_LC_10_19_0.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_118_RNI43UI1_15_LC_10_19_0 (
            .in0(N__65301),
            .in1(N__60302),
            .in2(N__90077),
            .in3(N__66454),
            .lcout(),
            .ltout(clk_en_0_a2_0_a2_sx_128_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_118_RNIB5DA01_15_LC_10_19_1.C_ON=1'b0;
    defparam shift_srl_118_RNIB5DA01_15_LC_10_19_1.SEQ_MODE=4'b0000;
    defparam shift_srl_118_RNIB5DA01_15_LC_10_19_1.LUT_INIT=16'b0000010000000000;
    LogicCell40 shift_srl_118_RNIB5DA01_15_LC_10_19_1 (
            .in0(N__60650),
            .in1(N__65658),
            .in2(N__56284),
            .in3(N__79416),
            .lcout(clk_en_128),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_123_RNI0JV11_15_LC_10_19_2.C_ON=1'b0;
    defparam shift_srl_123_RNI0JV11_15_LC_10_19_2.SEQ_MODE=4'b0000;
    defparam shift_srl_123_RNI0JV11_15_LC_10_19_2.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_123_RNI0JV11_15_LC_10_19_2 (
            .in0(N__56238),
            .in1(N__60121),
            .in2(_gnd_net_),
            .in3(N__78446),
            .lcout(rco_int_0_a2_1_a2_0_123),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_123_15_LC_10_19_3.C_ON=1'b0;
    defparam shift_srl_123_15_LC_10_19_3.SEQ_MODE=4'b1000;
    defparam shift_srl_123_15_LC_10_19_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_123_15_LC_10_19_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56248),
            .lcout(shift_srl_123Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92998),
            .ce(N__56205),
            .sr(_gnd_net_));
    defparam shift_srl_123_0_LC_10_19_4.C_ON=1'b0;
    defparam shift_srl_123_0_LC_10_19_4.SEQ_MODE=4'b1000;
    defparam shift_srl_123_0_LC_10_19_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_123_0_LC_10_19_4 (
            .in0(N__56239),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_123Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92998),
            .ce(N__56205),
            .sr(_gnd_net_));
    defparam shift_srl_123_1_LC_10_19_5.C_ON=1'b0;
    defparam shift_srl_123_1_LC_10_19_5.SEQ_MODE=4'b1000;
    defparam shift_srl_123_1_LC_10_19_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_123_1_LC_10_19_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56230),
            .lcout(shift_srl_123Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92998),
            .ce(N__56205),
            .sr(_gnd_net_));
    defparam shift_srl_123_2_LC_10_19_6.C_ON=1'b0;
    defparam shift_srl_123_2_LC_10_19_6.SEQ_MODE=4'b1000;
    defparam shift_srl_123_2_LC_10_19_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_123_2_LC_10_19_6 (
            .in0(N__56224),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_123Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92998),
            .ce(N__56205),
            .sr(_gnd_net_));
    defparam shift_srl_121_10_LC_10_20_0.C_ON=1'b0;
    defparam shift_srl_121_10_LC_10_20_0.SEQ_MODE=4'b1000;
    defparam shift_srl_121_10_LC_10_20_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_121_10_LC_10_20_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56314),
            .lcout(shift_srl_121Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93012),
            .ce(N__59862),
            .sr(_gnd_net_));
    defparam shift_srl_121_11_LC_10_20_1.C_ON=1'b0;
    defparam shift_srl_121_11_LC_10_20_1.SEQ_MODE=4'b1000;
    defparam shift_srl_121_11_LC_10_20_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_121_11_LC_10_20_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56344),
            .lcout(shift_srl_121Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93012),
            .ce(N__59862),
            .sr(_gnd_net_));
    defparam shift_srl_121_12_LC_10_20_2.C_ON=1'b0;
    defparam shift_srl_121_12_LC_10_20_2.SEQ_MODE=4'b1000;
    defparam shift_srl_121_12_LC_10_20_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_121_12_LC_10_20_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56338),
            .lcout(shift_srl_121Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93012),
            .ce(N__59862),
            .sr(_gnd_net_));
    defparam shift_srl_121_13_LC_10_20_3.C_ON=1'b0;
    defparam shift_srl_121_13_LC_10_20_3.SEQ_MODE=4'b1000;
    defparam shift_srl_121_13_LC_10_20_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_121_13_LC_10_20_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56332),
            .lcout(shift_srl_121Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93012),
            .ce(N__59862),
            .sr(_gnd_net_));
    defparam shift_srl_121_14_LC_10_20_4.C_ON=1'b0;
    defparam shift_srl_121_14_LC_10_20_4.SEQ_MODE=4'b1000;
    defparam shift_srl_121_14_LC_10_20_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_121_14_LC_10_20_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56326),
            .lcout(shift_srl_121Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93012),
            .ce(N__59862),
            .sr(_gnd_net_));
    defparam shift_srl_121_15_LC_10_20_5.C_ON=1'b0;
    defparam shift_srl_121_15_LC_10_20_5.SEQ_MODE=4'b1000;
    defparam shift_srl_121_15_LC_10_20_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_121_15_LC_10_20_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56320),
            .lcout(shift_srl_121Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93012),
            .ce(N__59862),
            .sr(_gnd_net_));
    defparam shift_srl_121_9_LC_10_20_6.C_ON=1'b0;
    defparam shift_srl_121_9_LC_10_20_6.SEQ_MODE=4'b1000;
    defparam shift_srl_121_9_LC_10_20_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_121_9_LC_10_20_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56308),
            .lcout(shift_srl_121Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93012),
            .ce(N__59862),
            .sr(_gnd_net_));
    defparam shift_srl_121_8_LC_10_20_7.C_ON=1'b0;
    defparam shift_srl_121_8_LC_10_20_7.SEQ_MODE=4'b1000;
    defparam shift_srl_121_8_LC_10_20_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_121_8_LC_10_20_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59875),
            .lcout(shift_srl_121Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93012),
            .ce(N__59862),
            .sr(_gnd_net_));
    defparam shift_srl_125_10_LC_10_21_0.C_ON=1'b0;
    defparam shift_srl_125_10_LC_10_21_0.SEQ_MODE=4'b1000;
    defparam shift_srl_125_10_LC_10_21_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_125_10_LC_10_21_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56392),
            .lcout(shift_srl_125Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93025),
            .ce(N__56374),
            .sr(_gnd_net_));
    defparam shift_srl_125_11_LC_10_21_1.C_ON=1'b0;
    defparam shift_srl_125_11_LC_10_21_1.SEQ_MODE=4'b1000;
    defparam shift_srl_125_11_LC_10_21_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_125_11_LC_10_21_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56422),
            .lcout(shift_srl_125Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93025),
            .ce(N__56374),
            .sr(_gnd_net_));
    defparam shift_srl_125_12_LC_10_21_2.C_ON=1'b0;
    defparam shift_srl_125_12_LC_10_21_2.SEQ_MODE=4'b1000;
    defparam shift_srl_125_12_LC_10_21_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_125_12_LC_10_21_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56416),
            .lcout(shift_srl_125Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93025),
            .ce(N__56374),
            .sr(_gnd_net_));
    defparam shift_srl_125_13_LC_10_21_3.C_ON=1'b0;
    defparam shift_srl_125_13_LC_10_21_3.SEQ_MODE=4'b1000;
    defparam shift_srl_125_13_LC_10_21_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_125_13_LC_10_21_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56410),
            .lcout(shift_srl_125Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93025),
            .ce(N__56374),
            .sr(_gnd_net_));
    defparam shift_srl_125_14_LC_10_21_4.C_ON=1'b0;
    defparam shift_srl_125_14_LC_10_21_4.SEQ_MODE=4'b1000;
    defparam shift_srl_125_14_LC_10_21_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_125_14_LC_10_21_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56404),
            .lcout(shift_srl_125Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93025),
            .ce(N__56374),
            .sr(_gnd_net_));
    defparam shift_srl_125_15_LC_10_21_5.C_ON=1'b0;
    defparam shift_srl_125_15_LC_10_21_5.SEQ_MODE=4'b1000;
    defparam shift_srl_125_15_LC_10_21_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_125_15_LC_10_21_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56398),
            .lcout(shift_srl_125Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93025),
            .ce(N__56374),
            .sr(_gnd_net_));
    defparam shift_srl_125_9_LC_10_21_6.C_ON=1'b0;
    defparam shift_srl_125_9_LC_10_21_6.SEQ_MODE=4'b1000;
    defparam shift_srl_125_9_LC_10_21_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_125_9_LC_10_21_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56380),
            .lcout(shift_srl_125Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93025),
            .ce(N__56374),
            .sr(_gnd_net_));
    defparam shift_srl_125_8_LC_10_21_7.C_ON=1'b0;
    defparam shift_srl_125_8_LC_10_21_7.SEQ_MODE=4'b1000;
    defparam shift_srl_125_8_LC_10_21_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_125_8_LC_10_21_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56386),
            .lcout(shift_srl_125Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93025),
            .ce(N__56374),
            .sr(_gnd_net_));
    defparam shift_srl_112_RNIA81HS_15_LC_10_22_0.C_ON=1'b0;
    defparam shift_srl_112_RNIA81HS_15_LC_10_22_0.SEQ_MODE=4'b0000;
    defparam shift_srl_112_RNIA81HS_15_LC_10_22_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_112_RNIA81HS_15_LC_10_22_0 (
            .in0(N__60497),
            .in1(N__61991),
            .in2(N__60775),
            .in3(N__89794),
            .lcout(clk_en_113),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_112_15_LC_10_22_1.C_ON=1'b0;
    defparam shift_srl_112_15_LC_10_22_1.SEQ_MODE=4'b1000;
    defparam shift_srl_112_15_LC_10_22_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_112_15_LC_10_22_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57859),
            .lcout(shift_srl_112Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93040),
            .ce(N__60164),
            .sr(_gnd_net_));
    defparam shift_srl_114_RNIUNDS_15_LC_10_22_2.C_ON=1'b0;
    defparam shift_srl_114_RNIUNDS_15_LC_10_22_2.SEQ_MODE=4'b0000;
    defparam shift_srl_114_RNIUNDS_15_LC_10_22_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_114_RNIUNDS_15_LC_10_22_2 (
            .in0(N__58917),
            .in1(N__60415),
            .in2(N__60515),
            .in3(N__60732),
            .lcout(rco_int_0_a2_1_a2_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_114_RNIUNDS_0_15_LC_10_22_3.C_ON=1'b0;
    defparam shift_srl_114_RNIUNDS_0_15_LC_10_22_3.SEQ_MODE=4'b0000;
    defparam shift_srl_114_RNIUNDS_0_15_LC_10_22_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_114_RNIUNDS_0_15_LC_10_22_3 (
            .in0(N__60418),
            .in1(N__60496),
            .in2(N__60755),
            .in3(N__58920),
            .lcout(),
            .ltout(g0_9_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_118_RNI28CD1_15_LC_10_22_4.C_ON=1'b0;
    defparam shift_srl_118_RNI28CD1_15_LC_10_22_4.SEQ_MODE=4'b0000;
    defparam shift_srl_118_RNI28CD1_15_LC_10_22_4.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_118_RNI28CD1_15_LC_10_22_4 (
            .in0(N__60321),
            .in1(N__66447),
            .in2(N__56476),
            .in3(N__89793),
            .lcout(g0_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_114_RNI4GI51_15_LC_10_22_5.C_ON=1'b0;
    defparam shift_srl_114_RNI4GI51_15_LC_10_22_5.SEQ_MODE=4'b0000;
    defparam shift_srl_114_RNI4GI51_15_LC_10_22_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_114_RNI4GI51_15_LC_10_22_5 (
            .in0(N__60416),
            .in1(N__60319),
            .in2(N__60754),
            .in3(N__58918),
            .lcout(g0_9_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_114_RNIA8NU_15_LC_10_22_7.C_ON=1'b0;
    defparam shift_srl_114_RNIA8NU_15_LC_10_22_7.SEQ_MODE=4'b0000;
    defparam shift_srl_114_RNIA8NU_15_LC_10_22_7.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_114_RNIA8NU_15_LC_10_22_7 (
            .in0(N__60417),
            .in1(N__58919),
            .in2(N__66460),
            .in3(N__60320),
            .lcout(g0_8_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_108_RNIBDHMR_15_LC_10_23_0.C_ON=1'b0;
    defparam shift_srl_108_RNIBDHMR_15_LC_10_23_0.SEQ_MODE=4'b0000;
    defparam shift_srl_108_RNIBDHMR_15_LC_10_23_0.LUT_INIT=16'b0000100000000000;
    LogicCell40 shift_srl_108_RNIBDHMR_15_LC_10_23_0 (
            .in0(N__79595),
            .in1(N__62295),
            .in2(N__56596),
            .in3(N__79498),
            .lcout(clk_en_109),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_108_15_LC_10_23_1.C_ON=1'b0;
    defparam shift_srl_108_15_LC_10_23_1.SEQ_MODE=4'b1000;
    defparam shift_srl_108_15_LC_10_23_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_108_15_LC_10_23_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56530),
            .lcout(shift_srl_108Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93055),
            .ce(N__56926),
            .sr(_gnd_net_));
    defparam shift_srl_109_RNI3PIF_15_LC_10_23_2.C_ON=1'b0;
    defparam shift_srl_109_RNI3PIF_15_LC_10_23_2.SEQ_MODE=4'b0000;
    defparam shift_srl_109_RNI3PIF_15_LC_10_23_2.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_109_RNI3PIF_15_LC_10_23_2 (
            .in0(N__59290),
            .in1(N__59251),
            .in2(N__90076),
            .in3(N__62400),
            .lcout(),
            .ltout(clk_en_0_a3_0_a2_sx_110_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_109_RNIGGIQR_15_LC_10_23_3.C_ON=1'b0;
    defparam shift_srl_109_RNIGGIQR_15_LC_10_23_3.SEQ_MODE=4'b0000;
    defparam shift_srl_109_RNIGGIQR_15_LC_10_23_3.LUT_INIT=16'b0000010000000000;
    LogicCell40 shift_srl_109_RNIGGIQR_15_LC_10_23_3 (
            .in0(N__56428),
            .in1(N__79596),
            .in2(N__56431),
            .in3(N__79510),
            .lcout(clk_en_110),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_108_RNI7QFR_15_LC_10_23_4.C_ON=1'b0;
    defparam shift_srl_108_RNI7QFR_15_LC_10_23_4.SEQ_MODE=4'b0000;
    defparam shift_srl_108_RNI7QFR_15_LC_10_23_4.LUT_INIT=16'b0011001111111111;
    LogicCell40 shift_srl_108_RNI7QFR_15_LC_10_23_4 (
            .in0(_gnd_net_),
            .in1(N__62358),
            .in2(_gnd_net_),
            .in3(N__62294),
            .lcout(clk_en_0_a3_0_a2_1_110),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_108_14_LC_10_23_5.C_ON=1'b0;
    defparam shift_srl_108_14_LC_10_23_5.SEQ_MODE=4'b1000;
    defparam shift_srl_108_14_LC_10_23_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_108_14_LC_10_23_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56524),
            .lcout(shift_srl_108Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93055),
            .ce(N__56926),
            .sr(_gnd_net_));
    defparam shift_srl_108_13_LC_10_23_6.C_ON=1'b0;
    defparam shift_srl_108_13_LC_10_23_6.SEQ_MODE=4'b1000;
    defparam shift_srl_108_13_LC_10_23_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_108_13_LC_10_23_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56518),
            .lcout(shift_srl_108Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93055),
            .ce(N__56926),
            .sr(_gnd_net_));
    defparam shift_srl_108_12_LC_10_23_7.C_ON=1'b0;
    defparam shift_srl_108_12_LC_10_23_7.SEQ_MODE=4'b1000;
    defparam shift_srl_108_12_LC_10_23_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_108_12_LC_10_23_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56800),
            .lcout(shift_srl_108Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93055),
            .ce(N__56926),
            .sr(_gnd_net_));
    defparam shift_srl_110_0_LC_10_24_0.C_ON=1'b0;
    defparam shift_srl_110_0_LC_10_24_0.SEQ_MODE=4'b1000;
    defparam shift_srl_110_0_LC_10_24_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_110_0_LC_10_24_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62431),
            .lcout(shift_srl_110Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93071),
            .ce(N__62447),
            .sr(_gnd_net_));
    defparam shift_srl_110_1_LC_10_24_1.C_ON=1'b0;
    defparam shift_srl_110_1_LC_10_24_1.SEQ_MODE=4'b1000;
    defparam shift_srl_110_1_LC_10_24_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_110_1_LC_10_24_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56512),
            .lcout(shift_srl_110Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93071),
            .ce(N__62447),
            .sr(_gnd_net_));
    defparam shift_srl_110_2_LC_10_24_2.C_ON=1'b0;
    defparam shift_srl_110_2_LC_10_24_2.SEQ_MODE=4'b1000;
    defparam shift_srl_110_2_LC_10_24_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_110_2_LC_10_24_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56506),
            .lcout(shift_srl_110Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93071),
            .ce(N__62447),
            .sr(_gnd_net_));
    defparam shift_srl_110_3_LC_10_24_3.C_ON=1'b0;
    defparam shift_srl_110_3_LC_10_24_3.SEQ_MODE=4'b1000;
    defparam shift_srl_110_3_LC_10_24_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_110_3_LC_10_24_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56500),
            .lcout(shift_srl_110Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93071),
            .ce(N__62447),
            .sr(_gnd_net_));
    defparam shift_srl_110_4_LC_10_24_4.C_ON=1'b0;
    defparam shift_srl_110_4_LC_10_24_4.SEQ_MODE=4'b1000;
    defparam shift_srl_110_4_LC_10_24_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_110_4_LC_10_24_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56494),
            .lcout(shift_srl_110Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93071),
            .ce(N__62447),
            .sr(_gnd_net_));
    defparam shift_srl_110_5_LC_10_24_5.C_ON=1'b0;
    defparam shift_srl_110_5_LC_10_24_5.SEQ_MODE=4'b1000;
    defparam shift_srl_110_5_LC_10_24_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_110_5_LC_10_24_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56488),
            .lcout(shift_srl_110Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93071),
            .ce(N__62447),
            .sr(_gnd_net_));
    defparam shift_srl_110_8_LC_10_24_6.C_ON=1'b0;
    defparam shift_srl_110_8_LC_10_24_6.SEQ_MODE=4'b1000;
    defparam shift_srl_110_8_LC_10_24_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_110_8_LC_10_24_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56572),
            .lcout(shift_srl_110Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93071),
            .ce(N__62447),
            .sr(_gnd_net_));
    defparam shift_srl_110_7_LC_10_24_7.C_ON=1'b0;
    defparam shift_srl_110_7_LC_10_24_7.SEQ_MODE=4'b1000;
    defparam shift_srl_110_7_LC_10_24_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_110_7_LC_10_24_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56578),
            .lcout(shift_srl_110Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93071),
            .ce(N__62447),
            .sr(_gnd_net_));
    defparam shift_srl_107_10_LC_10_25_0.C_ON=1'b0;
    defparam shift_srl_107_10_LC_10_25_0.SEQ_MODE=4'b1000;
    defparam shift_srl_107_10_LC_10_25_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_107_10_LC_10_25_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56536),
            .lcout(shift_srl_107Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93085),
            .ce(N__56683),
            .sr(_gnd_net_));
    defparam shift_srl_107_11_LC_10_25_1.C_ON=1'b0;
    defparam shift_srl_107_11_LC_10_25_1.SEQ_MODE=4'b1000;
    defparam shift_srl_107_11_LC_10_25_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_107_11_LC_10_25_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56566),
            .lcout(shift_srl_107Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93085),
            .ce(N__56683),
            .sr(_gnd_net_));
    defparam shift_srl_107_12_LC_10_25_2.C_ON=1'b0;
    defparam shift_srl_107_12_LC_10_25_2.SEQ_MODE=4'b1000;
    defparam shift_srl_107_12_LC_10_25_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_107_12_LC_10_25_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56560),
            .lcout(shift_srl_107Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93085),
            .ce(N__56683),
            .sr(_gnd_net_));
    defparam shift_srl_107_13_LC_10_25_3.C_ON=1'b0;
    defparam shift_srl_107_13_LC_10_25_3.SEQ_MODE=4'b1000;
    defparam shift_srl_107_13_LC_10_25_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_107_13_LC_10_25_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56554),
            .lcout(shift_srl_107Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93085),
            .ce(N__56683),
            .sr(_gnd_net_));
    defparam shift_srl_107_14_LC_10_25_4.C_ON=1'b0;
    defparam shift_srl_107_14_LC_10_25_4.SEQ_MODE=4'b1000;
    defparam shift_srl_107_14_LC_10_25_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_107_14_LC_10_25_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56548),
            .lcout(shift_srl_107Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93085),
            .ce(N__56683),
            .sr(_gnd_net_));
    defparam shift_srl_107_15_LC_10_25_5.C_ON=1'b0;
    defparam shift_srl_107_15_LC_10_25_5.SEQ_MODE=4'b1000;
    defparam shift_srl_107_15_LC_10_25_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_107_15_LC_10_25_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56542),
            .lcout(shift_srl_107Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93085),
            .ce(N__56683),
            .sr(_gnd_net_));
    defparam shift_srl_107_9_LC_10_25_6.C_ON=1'b0;
    defparam shift_srl_107_9_LC_10_25_6.SEQ_MODE=4'b1000;
    defparam shift_srl_107_9_LC_10_25_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_107_9_LC_10_25_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56698),
            .lcout(shift_srl_107Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93085),
            .ce(N__56683),
            .sr(_gnd_net_));
    defparam shift_srl_107_8_LC_10_25_7.C_ON=1'b0;
    defparam shift_srl_107_8_LC_10_25_7.SEQ_MODE=4'b1000;
    defparam shift_srl_107_8_LC_10_25_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_107_8_LC_10_25_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56707),
            .lcout(shift_srl_107Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93085),
            .ce(N__56683),
            .sr(_gnd_net_));
    defparam shift_srl_105_RNI2SIJQ_15_LC_10_26_0.C_ON=1'b0;
    defparam shift_srl_105_RNI2SIJQ_15_LC_10_26_0.SEQ_MODE=4'b0000;
    defparam shift_srl_105_RNI2SIJQ_15_LC_10_26_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_105_RNI2SIJQ_15_LC_10_26_0 (
            .in0(N__59283),
            .in1(N__79585),
            .in2(N__90075),
            .in3(N__79544),
            .lcout(clk_en_106),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNI4J1RQ_15_LC_10_26_1.C_ON=1'b0;
    defparam shift_srl_0_RNI4J1RQ_15_LC_10_26_1.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNI4J1RQ_15_LC_10_26_1.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_0_RNI4J1RQ_15_LC_10_26_1 (
            .in0(N__79545),
            .in1(N__89799),
            .in2(_gnd_net_),
            .in3(N__56608),
            .lcout(clk_en_107),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_106_RNI977QQ_15_LC_10_26_2.C_ON=1'b0;
    defparam shift_srl_106_RNI977QQ_15_LC_10_26_2.SEQ_MODE=4'b0000;
    defparam shift_srl_106_RNI977QQ_15_LC_10_26_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_106_RNI977QQ_15_LC_10_26_2 (
            .in0(N__59284),
            .in1(N__79586),
            .in2(N__59246),
            .in3(N__79547),
            .lcout(rco_c_106),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_106_RNIPC6S1_15_LC_10_26_3.C_ON=1'b0;
    defparam shift_srl_106_RNIPC6S1_15_LC_10_26_3.SEQ_MODE=4'b0000;
    defparam shift_srl_106_RNIPC6S1_15_LC_10_26_3.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_106_RNIPC6S1_15_LC_10_26_3 (
            .in0(N__79584),
            .in1(N__59235),
            .in2(_gnd_net_),
            .in3(N__59282),
            .lcout(shift_srl_106_RNIPC6S1Z0Z_15),
            .ltout(shift_srl_106_RNIPC6S1Z0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_107_RNI7EM6R_15_LC_10_26_4.C_ON=1'b0;
    defparam shift_srl_107_RNI7EM6R_15_LC_10_26_4.SEQ_MODE=4'b0000;
    defparam shift_srl_107_RNI7EM6R_15_LC_10_26_4.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_107_RNI7EM6R_15_LC_10_26_4 (
            .in0(N__89798),
            .in1(N__62345),
            .in2(N__56602),
            .in3(N__79546),
            .lcout(clk_en_108),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_102_RNIM2FH1_15_LC_10_26_5.C_ON=1'b0;
    defparam shift_srl_102_RNIM2FH1_15_LC_10_26_5.SEQ_MODE=4'b0000;
    defparam shift_srl_102_RNIM2FH1_15_LC_10_26_5.LUT_INIT=16'b0011001100000000;
    LogicCell40 shift_srl_102_RNIM2FH1_15_LC_10_26_5 (
            .in0(_gnd_net_),
            .in1(N__60940),
            .in2(_gnd_net_),
            .in3(N__62704),
            .lcout(rco_int_0_a3_0_a2_out_0),
            .ltout(rco_int_0_a3_0_a2_out_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNI19AGQ_15_LC_10_26_6.C_ON=1'b0;
    defparam shift_srl_0_RNI19AGQ_15_LC_10_26_6.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNI19AGQ_15_LC_10_26_6.LUT_INIT=16'b1100000000000000;
    LogicCell40 shift_srl_0_RNI19AGQ_15_LC_10_26_6 (
            .in0(_gnd_net_),
            .in1(N__89792),
            .in2(N__56599),
            .in3(N__79543),
            .lcout(clk_en_105),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_106_RNI1H6N_15_LC_10_26_7.C_ON=1'b0;
    defparam shift_srl_106_RNI1H6N_15_LC_10_26_7.SEQ_MODE=4'b0000;
    defparam shift_srl_106_RNI1H6N_15_LC_10_26_7.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_106_RNI1H6N_15_LC_10_26_7 (
            .in0(N__62344),
            .in1(N__59234),
            .in2(N__90071),
            .in3(N__59281),
            .lcout(clk_en_0_a3_0_a2_sx_109),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_106_10_LC_10_27_0.C_ON=1'b0;
    defparam shift_srl_106_10_LC_10_27_0.SEQ_MODE=4'b1000;
    defparam shift_srl_106_10_LC_10_27_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_106_10_LC_10_27_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56746),
            .lcout(shift_srl_106Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93118),
            .ce(N__56724),
            .sr(_gnd_net_));
    defparam shift_srl_106_11_LC_10_27_1.C_ON=1'b0;
    defparam shift_srl_106_11_LC_10_27_1.SEQ_MODE=4'b1000;
    defparam shift_srl_106_11_LC_10_27_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_106_11_LC_10_27_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56782),
            .lcout(shift_srl_106Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93118),
            .ce(N__56724),
            .sr(_gnd_net_));
    defparam shift_srl_106_12_LC_10_27_2.C_ON=1'b0;
    defparam shift_srl_106_12_LC_10_27_2.SEQ_MODE=4'b1000;
    defparam shift_srl_106_12_LC_10_27_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_106_12_LC_10_27_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56776),
            .lcout(shift_srl_106Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93118),
            .ce(N__56724),
            .sr(_gnd_net_));
    defparam shift_srl_106_13_LC_10_27_3.C_ON=1'b0;
    defparam shift_srl_106_13_LC_10_27_3.SEQ_MODE=4'b1000;
    defparam shift_srl_106_13_LC_10_27_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_106_13_LC_10_27_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56770),
            .lcout(shift_srl_106Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93118),
            .ce(N__56724),
            .sr(_gnd_net_));
    defparam shift_srl_106_14_LC_10_27_4.C_ON=1'b0;
    defparam shift_srl_106_14_LC_10_27_4.SEQ_MODE=4'b1000;
    defparam shift_srl_106_14_LC_10_27_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_106_14_LC_10_27_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56764),
            .lcout(shift_srl_106Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93118),
            .ce(N__56724),
            .sr(_gnd_net_));
    defparam shift_srl_106_15_LC_10_27_5.C_ON=1'b0;
    defparam shift_srl_106_15_LC_10_27_5.SEQ_MODE=4'b1000;
    defparam shift_srl_106_15_LC_10_27_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_106_15_LC_10_27_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56758),
            .lcout(shift_srl_106Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93118),
            .ce(N__56724),
            .sr(_gnd_net_));
    defparam shift_srl_106_9_LC_10_27_6.C_ON=1'b0;
    defparam shift_srl_106_9_LC_10_27_6.SEQ_MODE=4'b1000;
    defparam shift_srl_106_9_LC_10_27_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_106_9_LC_10_27_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56752),
            .lcout(shift_srl_106Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93118),
            .ce(N__56724),
            .sr(_gnd_net_));
    defparam shift_srl_106_1_LC_10_27_7.C_ON=1'b0;
    defparam shift_srl_106_1_LC_10_27_7.SEQ_MODE=4'b1000;
    defparam shift_srl_106_1_LC_10_27_7.LUT_INIT=16'b1100110011001100;
    LogicCell40 shift_srl_106_1_LC_10_27_7 (
            .in0(_gnd_net_),
            .in1(N__56740),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_106Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93118),
            .ce(N__56724),
            .sr(_gnd_net_));
    defparam shift_srl_108_0_LC_10_28_0.C_ON=1'b0;
    defparam shift_srl_108_0_LC_10_28_0.SEQ_MODE=4'b1000;
    defparam shift_srl_108_0_LC_10_28_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_108_0_LC_10_28_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62304),
            .lcout(shift_srl_108Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93137),
            .ce(N__56921),
            .sr(_gnd_net_));
    defparam shift_srl_108_1_LC_10_28_1.C_ON=1'b0;
    defparam shift_srl_108_1_LC_10_28_1.SEQ_MODE=4'b1000;
    defparam shift_srl_108_1_LC_10_28_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_108_1_LC_10_28_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56848),
            .lcout(shift_srl_108Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93137),
            .ce(N__56921),
            .sr(_gnd_net_));
    defparam shift_srl_108_2_LC_10_28_2.C_ON=1'b0;
    defparam shift_srl_108_2_LC_10_28_2.SEQ_MODE=4'b1000;
    defparam shift_srl_108_2_LC_10_28_2.LUT_INIT=16'b1100110011001100;
    LogicCell40 shift_srl_108_2_LC_10_28_2 (
            .in0(_gnd_net_),
            .in1(N__56842),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_108Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93137),
            .ce(N__56921),
            .sr(_gnd_net_));
    defparam shift_srl_108_3_LC_10_28_3.C_ON=1'b0;
    defparam shift_srl_108_3_LC_10_28_3.SEQ_MODE=4'b1000;
    defparam shift_srl_108_3_LC_10_28_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_108_3_LC_10_28_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56836),
            .lcout(shift_srl_108Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93137),
            .ce(N__56921),
            .sr(_gnd_net_));
    defparam shift_srl_108_4_LC_10_28_4.C_ON=1'b0;
    defparam shift_srl_108_4_LC_10_28_4.SEQ_MODE=4'b1000;
    defparam shift_srl_108_4_LC_10_28_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_108_4_LC_10_28_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56830),
            .lcout(shift_srl_108Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93137),
            .ce(N__56921),
            .sr(_gnd_net_));
    defparam shift_srl_108_5_LC_10_28_5.C_ON=1'b0;
    defparam shift_srl_108_5_LC_10_28_5.SEQ_MODE=4'b1000;
    defparam shift_srl_108_5_LC_10_28_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_108_5_LC_10_28_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56824),
            .lcout(shift_srl_108Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93137),
            .ce(N__56921),
            .sr(_gnd_net_));
    defparam shift_srl_108_6_LC_10_28_6.C_ON=1'b0;
    defparam shift_srl_108_6_LC_10_28_6.SEQ_MODE=4'b1000;
    defparam shift_srl_108_6_LC_10_28_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_108_6_LC_10_28_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56818),
            .lcout(shift_srl_108Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93137),
            .ce(N__56921),
            .sr(_gnd_net_));
    defparam shift_srl_108_7_LC_10_28_7.C_ON=1'b0;
    defparam shift_srl_108_7_LC_10_28_7.SEQ_MODE=4'b1000;
    defparam shift_srl_108_7_LC_10_28_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_108_7_LC_10_28_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56812),
            .lcout(shift_srl_108Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93137),
            .ce(N__56921),
            .sr(_gnd_net_));
    defparam shift_srl_108_10_LC_10_29_0.C_ON=1'b0;
    defparam shift_srl_108_10_LC_10_29_0.SEQ_MODE=4'b1000;
    defparam shift_srl_108_10_LC_10_29_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_108_10_LC_10_29_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56788),
            .lcout(shift_srl_108Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93155),
            .ce(N__56925),
            .sr(_gnd_net_));
    defparam shift_srl_108_11_LC_10_29_1.C_ON=1'b0;
    defparam shift_srl_108_11_LC_10_29_1.SEQ_MODE=4'b1000;
    defparam shift_srl_108_11_LC_10_29_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_108_11_LC_10_29_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56806),
            .lcout(shift_srl_108Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93155),
            .ce(N__56925),
            .sr(_gnd_net_));
    defparam shift_srl_108_9_LC_10_29_2.C_ON=1'b0;
    defparam shift_srl_108_9_LC_10_29_2.SEQ_MODE=4'b1000;
    defparam shift_srl_108_9_LC_10_29_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_108_9_LC_10_29_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56932),
            .lcout(shift_srl_108Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93155),
            .ce(N__56925),
            .sr(_gnd_net_));
    defparam shift_srl_108_8_LC_10_29_3.C_ON=1'b0;
    defparam shift_srl_108_8_LC_10_29_3.SEQ_MODE=4'b1000;
    defparam shift_srl_108_8_LC_10_29_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_108_8_LC_10_29_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56938),
            .lcout(shift_srl_108Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93155),
            .ce(N__56925),
            .sr(_gnd_net_));
    defparam shift_srl_0_11_LC_11_6_1.C_ON=1'b0;
    defparam shift_srl_0_11_LC_11_6_1.SEQ_MODE=4'b1000;
    defparam shift_srl_0_11_LC_11_6_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_0_11_LC_11_6_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56890),
            .lcout(shift_srl_0Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93158),
            .ce(N__57246),
            .sr(_gnd_net_));
    defparam shift_srl_0_12_LC_11_6_2.C_ON=1'b0;
    defparam shift_srl_0_12_LC_11_6_2.SEQ_MODE=4'b1000;
    defparam shift_srl_0_12_LC_11_6_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_0_12_LC_11_6_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56884),
            .lcout(shift_srl_0Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93158),
            .ce(N__57246),
            .sr(_gnd_net_));
    defparam shift_srl_0_13_LC_11_6_3.C_ON=1'b0;
    defparam shift_srl_0_13_LC_11_6_3.SEQ_MODE=4'b1000;
    defparam shift_srl_0_13_LC_11_6_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_0_13_LC_11_6_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56878),
            .lcout(shift_srl_0Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93158),
            .ce(N__57246),
            .sr(_gnd_net_));
    defparam shift_srl_0_14_LC_11_6_4.C_ON=1'b0;
    defparam shift_srl_0_14_LC_11_6_4.SEQ_MODE=4'b1000;
    defparam shift_srl_0_14_LC_11_6_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_0_14_LC_11_6_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56872),
            .lcout(shift_srl_0Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93158),
            .ce(N__57246),
            .sr(_gnd_net_));
    defparam shift_srl_0_15_LC_11_6_5.C_ON=1'b0;
    defparam shift_srl_0_15_LC_11_6_5.SEQ_MODE=4'b1000;
    defparam shift_srl_0_15_LC_11_6_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_0_15_LC_11_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56866),
            .lcout(rco_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93158),
            .ce(N__57246),
            .sr(_gnd_net_));
    defparam shift_srl_148_10_LC_11_8_0.C_ON=1'b0;
    defparam shift_srl_148_10_LC_11_8_0.SEQ_MODE=4'b1000;
    defparam shift_srl_148_10_LC_11_8_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_148_10_LC_11_8_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57040),
            .lcout(shift_srl_148Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93120),
            .ce(N__58236),
            .sr(_gnd_net_));
    defparam shift_srl_148_11_LC_11_8_1.C_ON=1'b0;
    defparam shift_srl_148_11_LC_11_8_1.SEQ_MODE=4'b1000;
    defparam shift_srl_148_11_LC_11_8_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_148_11_LC_11_8_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56860),
            .lcout(shift_srl_148Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93120),
            .ce(N__58236),
            .sr(_gnd_net_));
    defparam shift_srl_148_12_LC_11_8_2.C_ON=1'b0;
    defparam shift_srl_148_12_LC_11_8_2.SEQ_MODE=4'b1000;
    defparam shift_srl_148_12_LC_11_8_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_148_12_LC_11_8_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56854),
            .lcout(shift_srl_148Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93120),
            .ce(N__58236),
            .sr(_gnd_net_));
    defparam shift_srl_148_13_LC_11_8_3.C_ON=1'b0;
    defparam shift_srl_148_13_LC_11_8_3.SEQ_MODE=4'b1000;
    defparam shift_srl_148_13_LC_11_8_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_148_13_LC_11_8_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57058),
            .lcout(shift_srl_148Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93120),
            .ce(N__58236),
            .sr(_gnd_net_));
    defparam shift_srl_148_14_LC_11_8_4.C_ON=1'b0;
    defparam shift_srl_148_14_LC_11_8_4.SEQ_MODE=4'b1000;
    defparam shift_srl_148_14_LC_11_8_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_148_14_LC_11_8_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57052),
            .lcout(shift_srl_148Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93120),
            .ce(N__58236),
            .sr(_gnd_net_));
    defparam shift_srl_148_15_LC_11_8_5.C_ON=1'b0;
    defparam shift_srl_148_15_LC_11_8_5.SEQ_MODE=4'b1000;
    defparam shift_srl_148_15_LC_11_8_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_148_15_LC_11_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57046),
            .lcout(shift_srl_148Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93120),
            .ce(N__58236),
            .sr(_gnd_net_));
    defparam shift_srl_148_9_LC_11_8_6.C_ON=1'b0;
    defparam shift_srl_148_9_LC_11_8_6.SEQ_MODE=4'b1000;
    defparam shift_srl_148_9_LC_11_8_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_148_9_LC_11_8_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57034),
            .lcout(shift_srl_148Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93120),
            .ce(N__58236),
            .sr(_gnd_net_));
    defparam shift_srl_148_8_LC_11_8_7.C_ON=1'b0;
    defparam shift_srl_148_8_LC_11_8_7.SEQ_MODE=4'b1000;
    defparam shift_srl_148_8_LC_11_8_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_148_8_LC_11_8_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58273),
            .lcout(shift_srl_148Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93120),
            .ce(N__58236),
            .sr(_gnd_net_));
    defparam shift_srl_147_RNI41O251_15_LC_11_9_0.C_ON=1'b0;
    defparam shift_srl_147_RNI41O251_15_LC_11_9_0.SEQ_MODE=4'b0000;
    defparam shift_srl_147_RNI41O251_15_LC_11_9_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_147_RNI41O251_15_LC_11_9_0 (
            .in0(N__70719),
            .in1(N__57028),
            .in2(N__89760),
            .in3(N__82185),
            .lcout(clk_en_148),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_148_0_LC_11_9_2.C_ON=1'b0;
    defparam shift_srl_148_0_LC_11_9_2.SEQ_MODE=4'b1000;
    defparam shift_srl_148_0_LC_11_9_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_148_0_LC_11_9_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56968),
            .lcout(shift_srl_148Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93101),
            .ce(N__58235),
            .sr(_gnd_net_));
    defparam shift_srl_148_1_LC_11_9_3.C_ON=1'b0;
    defparam shift_srl_148_1_LC_11_9_3.SEQ_MODE=4'b1000;
    defparam shift_srl_148_1_LC_11_9_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_148_1_LC_11_9_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56950),
            .lcout(shift_srl_148Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93101),
            .ce(N__58235),
            .sr(_gnd_net_));
    defparam shift_srl_148_2_LC_11_9_4.C_ON=1'b0;
    defparam shift_srl_148_2_LC_11_9_4.SEQ_MODE=4'b1000;
    defparam shift_srl_148_2_LC_11_9_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_148_2_LC_11_9_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56944),
            .lcout(shift_srl_148Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93101),
            .ce(N__58235),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_1_LC_11_10_3.C_ON=1'b0;
    defparam rco_obuf_RNO_1_LC_11_10_3.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_1_LC_11_10_3.LUT_INIT=16'b1100110000000000;
    LogicCell40 rco_obuf_RNO_1_LC_11_10_3 (
            .in0(_gnd_net_),
            .in1(N__57250),
            .in2(_gnd_net_),
            .in3(N__57169),
            .lcout(N_452_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_154_10_LC_11_13_0.C_ON=1'b0;
    defparam shift_srl_154_10_LC_11_13_0.SEQ_MODE=4'b1000;
    defparam shift_srl_154_10_LC_11_13_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_154_10_LC_11_13_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57106),
            .lcout(shift_srl_154Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93041),
            .ce(N__57340),
            .sr(_gnd_net_));
    defparam shift_srl_154_11_LC_11_13_1.C_ON=1'b0;
    defparam shift_srl_154_11_LC_11_13_1.SEQ_MODE=4'b1000;
    defparam shift_srl_154_11_LC_11_13_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_154_11_LC_11_13_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57112),
            .lcout(shift_srl_154Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93041),
            .ce(N__57340),
            .sr(_gnd_net_));
    defparam shift_srl_154_9_LC_11_13_2.C_ON=1'b0;
    defparam shift_srl_154_9_LC_11_13_2.SEQ_MODE=4'b1000;
    defparam shift_srl_154_9_LC_11_13_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_154_9_LC_11_13_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57100),
            .lcout(shift_srl_154Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93041),
            .ce(N__57340),
            .sr(_gnd_net_));
    defparam shift_srl_154_8_LC_11_13_3.C_ON=1'b0;
    defparam shift_srl_154_8_LC_11_13_3.SEQ_MODE=4'b1000;
    defparam shift_srl_154_8_LC_11_13_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_154_8_LC_11_13_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57094),
            .lcout(shift_srl_154Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93041),
            .ce(N__57340),
            .sr(_gnd_net_));
    defparam shift_srl_154_7_LC_11_13_4.C_ON=1'b0;
    defparam shift_srl_154_7_LC_11_13_4.SEQ_MODE=4'b1000;
    defparam shift_srl_154_7_LC_11_13_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_154_7_LC_11_13_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57088),
            .lcout(shift_srl_154Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93041),
            .ce(N__57340),
            .sr(_gnd_net_));
    defparam shift_srl_154_6_LC_11_13_5.C_ON=1'b0;
    defparam shift_srl_154_6_LC_11_13_5.SEQ_MODE=4'b1000;
    defparam shift_srl_154_6_LC_11_13_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_154_6_LC_11_13_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57082),
            .lcout(shift_srl_154Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93041),
            .ce(N__57340),
            .sr(_gnd_net_));
    defparam shift_srl_154_5_LC_11_13_6.C_ON=1'b0;
    defparam shift_srl_154_5_LC_11_13_6.SEQ_MODE=4'b1000;
    defparam shift_srl_154_5_LC_11_13_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_154_5_LC_11_13_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57064),
            .lcout(shift_srl_154Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93041),
            .ce(N__57340),
            .sr(_gnd_net_));
    defparam shift_srl_154_4_LC_11_13_7.C_ON=1'b0;
    defparam shift_srl_154_4_LC_11_13_7.SEQ_MODE=4'b1000;
    defparam shift_srl_154_4_LC_11_13_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_154_4_LC_11_13_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57076),
            .lcout(shift_srl_154Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93041),
            .ce(N__57340),
            .sr(_gnd_net_));
    defparam shift_srl_157_10_LC_11_14_0.C_ON=1'b0;
    defparam shift_srl_157_10_LC_11_14_0.SEQ_MODE=4'b1000;
    defparam shift_srl_157_10_LC_11_14_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_157_10_LC_11_14_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57286),
            .lcout(shift_srl_157Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93026),
            .ce(N__58413),
            .sr(_gnd_net_));
    defparam shift_srl_157_11_LC_11_14_1.C_ON=1'b0;
    defparam shift_srl_157_11_LC_11_14_1.SEQ_MODE=4'b1000;
    defparam shift_srl_157_11_LC_11_14_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_157_11_LC_11_14_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57304),
            .lcout(shift_srl_157Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93026),
            .ce(N__58413),
            .sr(_gnd_net_));
    defparam shift_srl_157_12_LC_11_14_2.C_ON=1'b0;
    defparam shift_srl_157_12_LC_11_14_2.SEQ_MODE=4'b1000;
    defparam shift_srl_157_12_LC_11_14_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_157_12_LC_11_14_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57298),
            .lcout(shift_srl_157Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93026),
            .ce(N__58413),
            .sr(_gnd_net_));
    defparam shift_srl_157_6_LC_11_14_3.C_ON=1'b0;
    defparam shift_srl_157_6_LC_11_14_3.SEQ_MODE=4'b1000;
    defparam shift_srl_157_6_LC_11_14_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_157_6_LC_11_14_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57292),
            .lcout(shift_srl_157Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93026),
            .ce(N__58413),
            .sr(_gnd_net_));
    defparam shift_srl_157_5_LC_11_14_4.C_ON=1'b0;
    defparam shift_srl_157_5_LC_11_14_4.SEQ_MODE=4'b1000;
    defparam shift_srl_157_5_LC_11_14_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_157_5_LC_11_14_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58450),
            .lcout(shift_srl_157Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93026),
            .ce(N__58413),
            .sr(_gnd_net_));
    defparam shift_srl_157_15_LC_11_14_5.C_ON=1'b0;
    defparam shift_srl_157_15_LC_11_14_5.SEQ_MODE=4'b1000;
    defparam shift_srl_157_15_LC_11_14_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_157_15_LC_11_14_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58432),
            .lcout(shift_srl_157Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93026),
            .ce(N__58413),
            .sr(_gnd_net_));
    defparam shift_srl_157_9_LC_11_14_6.C_ON=1'b0;
    defparam shift_srl_157_9_LC_11_14_6.SEQ_MODE=4'b1000;
    defparam shift_srl_157_9_LC_11_14_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_157_9_LC_11_14_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57280),
            .lcout(shift_srl_157Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93026),
            .ce(N__58413),
            .sr(_gnd_net_));
    defparam shift_srl_157_8_LC_11_14_7.C_ON=1'b0;
    defparam shift_srl_157_8_LC_11_14_7.SEQ_MODE=4'b1000;
    defparam shift_srl_157_8_LC_11_14_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_157_8_LC_11_14_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58420),
            .lcout(shift_srl_157Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93026),
            .ce(N__58413),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNICHO881_15_LC_11_15_0.C_ON=1'b0;
    defparam shift_srl_0_RNICHO881_15_LC_11_15_0.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNICHO881_15_LC_11_15_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNICHO881_15_LC_11_15_0 (
            .in0(N__82145),
            .in1(N__71649),
            .in2(N__90042),
            .in3(N__82292),
            .lcout(clk_en_160),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIEEVK81_15_LC_11_15_1.C_ON=1'b0;
    defparam shift_srl_0_RNIEEVK81_15_LC_11_15_1.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIEEVK81_15_LC_11_15_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNIEEVK81_15_LC_11_15_1 (
            .in0(N__82293),
            .in1(N__69865),
            .in2(N__90427),
            .in3(N__82146),
            .lcout(clk_en_161),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIH8FE71_15_LC_11_15_2.C_ON=1'b0;
    defparam shift_srl_0_RNIH8FE71_15_LC_11_15_2.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIH8FE71_15_LC_11_15_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNIH8FE71_15_LC_11_15_2 (
            .in0(N__82147),
            .in1(N__77552),
            .in2(N__90043),
            .in3(N__82295),
            .lcout(clk_en_157),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_154_RNI4CIS61_15_LC_11_15_3.C_ON=1'b0;
    defparam shift_srl_154_RNI4CIS61_15_LC_11_15_3.SEQ_MODE=4'b0000;
    defparam shift_srl_154_RNI4CIS61_15_LC_11_15_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_154_RNI4CIS61_15_LC_11_15_3 (
            .in0(N__82294),
            .in1(N__77581),
            .in2(N__90428),
            .in3(N__82148),
            .lcout(clk_en_155),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_154_15_LC_11_15_4.C_ON=1'b0;
    defparam shift_srl_154_15_LC_11_15_4.SEQ_MODE=4'b1000;
    defparam shift_srl_154_15_LC_11_15_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_154_15_LC_11_15_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57382),
            .lcout(shift_srl_154Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93013),
            .ce(N__57348),
            .sr(_gnd_net_));
    defparam shift_srl_154_14_LC_11_15_5.C_ON=1'b0;
    defparam shift_srl_154_14_LC_11_15_5.SEQ_MODE=4'b1000;
    defparam shift_srl_154_14_LC_11_15_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_154_14_LC_11_15_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57376),
            .lcout(shift_srl_154Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93013),
            .ce(N__57348),
            .sr(_gnd_net_));
    defparam shift_srl_154_13_LC_11_15_6.C_ON=1'b0;
    defparam shift_srl_154_13_LC_11_15_6.SEQ_MODE=4'b1000;
    defparam shift_srl_154_13_LC_11_15_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_154_13_LC_11_15_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57361),
            .lcout(shift_srl_154Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93013),
            .ce(N__57348),
            .sr(_gnd_net_));
    defparam shift_srl_154_12_LC_11_15_7.C_ON=1'b0;
    defparam shift_srl_154_12_LC_11_15_7.SEQ_MODE=4'b1000;
    defparam shift_srl_154_12_LC_11_15_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_154_12_LC_11_15_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57370),
            .lcout(shift_srl_154Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93013),
            .ce(N__57348),
            .sr(_gnd_net_));
    defparam shift_srl_161_0_LC_11_16_0.C_ON=1'b0;
    defparam shift_srl_161_0_LC_11_16_0.SEQ_MODE=4'b1000;
    defparam shift_srl_161_0_LC_11_16_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_161_0_LC_11_16_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77350),
            .lcout(shift_srl_161Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92999),
            .ce(N__57420),
            .sr(_gnd_net_));
    defparam shift_srl_161_1_LC_11_16_1.C_ON=1'b0;
    defparam shift_srl_161_1_LC_11_16_1.SEQ_MODE=4'b1000;
    defparam shift_srl_161_1_LC_11_16_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_161_1_LC_11_16_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57316),
            .lcout(shift_srl_161Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92999),
            .ce(N__57420),
            .sr(_gnd_net_));
    defparam shift_srl_161_2_LC_11_16_2.C_ON=1'b0;
    defparam shift_srl_161_2_LC_11_16_2.SEQ_MODE=4'b1000;
    defparam shift_srl_161_2_LC_11_16_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_161_2_LC_11_16_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57310),
            .lcout(shift_srl_161Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92999),
            .ce(N__57420),
            .sr(_gnd_net_));
    defparam shift_srl_161_3_LC_11_16_3.C_ON=1'b0;
    defparam shift_srl_161_3_LC_11_16_3.SEQ_MODE=4'b1000;
    defparam shift_srl_161_3_LC_11_16_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_161_3_LC_11_16_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57457),
            .lcout(shift_srl_161Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92999),
            .ce(N__57420),
            .sr(_gnd_net_));
    defparam shift_srl_161_4_LC_11_16_4.C_ON=1'b0;
    defparam shift_srl_161_4_LC_11_16_4.SEQ_MODE=4'b1000;
    defparam shift_srl_161_4_LC_11_16_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_161_4_LC_11_16_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57451),
            .lcout(shift_srl_161Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92999),
            .ce(N__57420),
            .sr(_gnd_net_));
    defparam shift_srl_161_5_LC_11_16_5.C_ON=1'b0;
    defparam shift_srl_161_5_LC_11_16_5.SEQ_MODE=4'b1000;
    defparam shift_srl_161_5_LC_11_16_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_161_5_LC_11_16_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57445),
            .lcout(shift_srl_161Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92999),
            .ce(N__57420),
            .sr(_gnd_net_));
    defparam shift_srl_161_6_LC_11_16_6.C_ON=1'b0;
    defparam shift_srl_161_6_LC_11_16_6.SEQ_MODE=4'b1000;
    defparam shift_srl_161_6_LC_11_16_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_161_6_LC_11_16_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57439),
            .lcout(shift_srl_161Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92999),
            .ce(N__57420),
            .sr(_gnd_net_));
    defparam shift_srl_161_7_LC_11_16_7.C_ON=1'b0;
    defparam shift_srl_161_7_LC_11_16_7.SEQ_MODE=4'b1000;
    defparam shift_srl_161_7_LC_11_16_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_161_7_LC_11_16_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57433),
            .lcout(shift_srl_161Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92999),
            .ce(N__57420),
            .sr(_gnd_net_));
    defparam shift_srl_124_10_LC_11_17_0.C_ON=1'b0;
    defparam shift_srl_124_10_LC_11_17_0.SEQ_MODE=4'b1000;
    defparam shift_srl_124_10_LC_11_17_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_124_10_LC_11_17_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57505),
            .lcout(shift_srl_124Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92983),
            .ce(N__58723),
            .sr(_gnd_net_));
    defparam shift_srl_124_11_LC_11_17_1.C_ON=1'b0;
    defparam shift_srl_124_11_LC_11_17_1.SEQ_MODE=4'b1000;
    defparam shift_srl_124_11_LC_11_17_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_124_11_LC_11_17_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57400),
            .lcout(shift_srl_124Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92983),
            .ce(N__58723),
            .sr(_gnd_net_));
    defparam shift_srl_124_12_LC_11_17_2.C_ON=1'b0;
    defparam shift_srl_124_12_LC_11_17_2.SEQ_MODE=4'b1000;
    defparam shift_srl_124_12_LC_11_17_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_124_12_LC_11_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57394),
            .lcout(shift_srl_124Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92983),
            .ce(N__58723),
            .sr(_gnd_net_));
    defparam shift_srl_124_13_LC_11_17_3.C_ON=1'b0;
    defparam shift_srl_124_13_LC_11_17_3.SEQ_MODE=4'b1000;
    defparam shift_srl_124_13_LC_11_17_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_124_13_LC_11_17_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57388),
            .lcout(shift_srl_124Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92983),
            .ce(N__58723),
            .sr(_gnd_net_));
    defparam shift_srl_124_14_LC_11_17_4.C_ON=1'b0;
    defparam shift_srl_124_14_LC_11_17_4.SEQ_MODE=4'b1000;
    defparam shift_srl_124_14_LC_11_17_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_124_14_LC_11_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57511),
            .lcout(shift_srl_124Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92983),
            .ce(N__58723),
            .sr(_gnd_net_));
    defparam shift_srl_124_9_LC_11_17_5.C_ON=1'b0;
    defparam shift_srl_124_9_LC_11_17_5.SEQ_MODE=4'b1000;
    defparam shift_srl_124_9_LC_11_17_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_124_9_LC_11_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57499),
            .lcout(shift_srl_124Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92983),
            .ce(N__58723),
            .sr(_gnd_net_));
    defparam shift_srl_124_8_LC_11_17_6.C_ON=1'b0;
    defparam shift_srl_124_8_LC_11_17_6.SEQ_MODE=4'b1000;
    defparam shift_srl_124_8_LC_11_17_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_124_8_LC_11_17_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58624),
            .lcout(shift_srl_124Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92983),
            .ce(N__58723),
            .sr(_gnd_net_));
    defparam shift_srl_126_13_LC_11_18_0.C_ON=1'b0;
    defparam shift_srl_126_13_LC_11_18_0.SEQ_MODE=4'b1000;
    defparam shift_srl_126_13_LC_11_18_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_126_13_LC_11_18_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57493),
            .lcout(shift_srl_126Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93000),
            .ce(N__57546),
            .sr(_gnd_net_));
    defparam shift_srl_126_1_LC_11_18_1.C_ON=1'b0;
    defparam shift_srl_126_1_LC_11_18_1.SEQ_MODE=4'b1000;
    defparam shift_srl_126_1_LC_11_18_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_126_1_LC_11_18_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57487),
            .lcout(shift_srl_126Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93000),
            .ce(N__57546),
            .sr(_gnd_net_));
    defparam shift_srl_126_2_LC_11_18_2.C_ON=1'b0;
    defparam shift_srl_126_2_LC_11_18_2.SEQ_MODE=4'b1000;
    defparam shift_srl_126_2_LC_11_18_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_126_2_LC_11_18_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57481),
            .lcout(shift_srl_126Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93000),
            .ce(N__57546),
            .sr(_gnd_net_));
    defparam shift_srl_126_3_LC_11_18_3.C_ON=1'b0;
    defparam shift_srl_126_3_LC_11_18_3.SEQ_MODE=4'b1000;
    defparam shift_srl_126_3_LC_11_18_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_126_3_LC_11_18_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57475),
            .lcout(shift_srl_126Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93000),
            .ce(N__57546),
            .sr(_gnd_net_));
    defparam shift_srl_126_4_LC_11_18_4.C_ON=1'b0;
    defparam shift_srl_126_4_LC_11_18_4.SEQ_MODE=4'b1000;
    defparam shift_srl_126_4_LC_11_18_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_126_4_LC_11_18_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57469),
            .lcout(shift_srl_126Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93000),
            .ce(N__57546),
            .sr(_gnd_net_));
    defparam shift_srl_126_5_LC_11_18_5.C_ON=1'b0;
    defparam shift_srl_126_5_LC_11_18_5.SEQ_MODE=4'b1000;
    defparam shift_srl_126_5_LC_11_18_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_126_5_LC_11_18_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57463),
            .lcout(shift_srl_126Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93000),
            .ce(N__57546),
            .sr(_gnd_net_));
    defparam shift_srl_126_6_LC_11_18_6.C_ON=1'b0;
    defparam shift_srl_126_6_LC_11_18_6.SEQ_MODE=4'b1000;
    defparam shift_srl_126_6_LC_11_18_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_126_6_LC_11_18_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57670),
            .lcout(shift_srl_126Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93000),
            .ce(N__57546),
            .sr(_gnd_net_));
    defparam shift_srl_126_14_LC_11_18_7.C_ON=1'b0;
    defparam shift_srl_126_14_LC_11_18_7.SEQ_MODE=4'b1000;
    defparam shift_srl_126_14_LC_11_18_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_126_14_LC_11_18_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57658),
            .lcout(shift_srl_126Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93000),
            .ce(N__57546),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_126_LC_11_19_0.C_ON=1'b0;
    defparam rco_obuf_RNO_126_LC_11_19_0.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_126_LC_11_19_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 rco_obuf_RNO_126_LC_11_19_0 (
            .in0(N__65412),
            .in1(N__66063),
            .in2(N__66028),
            .in3(N__57601),
            .lcout(rco_c_126),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_125_RNI2V0UV_15_LC_11_19_3.C_ON=1'b0;
    defparam shift_srl_125_RNI2V0UV_15_LC_11_19_3.SEQ_MODE=4'b0000;
    defparam shift_srl_125_RNI2V0UV_15_LC_11_19_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_125_RNI2V0UV_15_LC_11_19_3 (
            .in0(N__57600),
            .in1(N__65411),
            .in2(N__66029),
            .in3(N__89759),
            .lcout(clk_en_126),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_124_15_LC_11_19_4.C_ON=1'b0;
    defparam shift_srl_124_15_LC_11_19_4.SEQ_MODE=4'b1000;
    defparam shift_srl_124_15_LC_11_19_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_124_15_LC_11_19_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57535),
            .lcout(shift_srl_124Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93014),
            .ce(N__58722),
            .sr(_gnd_net_));
    defparam shift_srl_127_RNIESVN_15_LC_11_19_5.C_ON=1'b0;
    defparam shift_srl_127_RNIESVN_15_LC_11_19_5.SEQ_MODE=4'b0000;
    defparam shift_srl_127_RNIESVN_15_LC_11_19_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_127_RNIESVN_15_LC_11_19_5 (
            .in0(N__66062),
            .in1(N__66015),
            .in2(N__68092),
            .in3(N__65410),
            .lcout(rco_int_0_a2_1_a2_0_127),
            .ltout(rco_int_0_a2_1_a2_0_127_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_145_RNII9RO3_15_LC_11_19_6.C_ON=1'b0;
    defparam shift_srl_145_RNII9RO3_15_LC_11_19_6.SEQ_MODE=4'b0000;
    defparam shift_srl_145_RNII9RO3_15_LC_11_19_6.LUT_INIT=16'b1111111101111111;
    LogicCell40 shift_srl_145_RNII9RO3_15_LC_11_19_6 (
            .in0(N__63591),
            .in1(N__66607),
            .in2(N__57526),
            .in3(N__57523),
            .lcout(),
            .ltout(rco_int_0_a2_0_a2_1_sx_145_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_145_RNIC08UB_15_LC_11_19_7.C_ON=1'b0;
    defparam shift_srl_145_RNIC08UB_15_LC_11_19_7.SEQ_MODE=4'b0000;
    defparam shift_srl_145_RNIC08UB_15_LC_11_19_7.LUT_INIT=16'b0000100000000000;
    LogicCell40 shift_srl_145_RNIC08UB_15_LC_11_19_7 (
            .in0(N__62129),
            .in1(N__64976),
            .in2(N__57514),
            .in3(N__62236),
            .lcout(rco_int_0_a2_0_a2_1_145),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_122_10_LC_11_20_0.C_ON=1'b0;
    defparam shift_srl_122_10_LC_11_20_0.SEQ_MODE=4'b1000;
    defparam shift_srl_122_10_LC_11_20_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_122_10_LC_11_20_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57682),
            .lcout(shift_srl_122Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93027),
            .ce(N__60051),
            .sr(_gnd_net_));
    defparam shift_srl_122_11_LC_11_20_1.C_ON=1'b0;
    defparam shift_srl_122_11_LC_11_20_1.SEQ_MODE=4'b1000;
    defparam shift_srl_122_11_LC_11_20_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_122_11_LC_11_20_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57712),
            .lcout(shift_srl_122Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93027),
            .ce(N__60051),
            .sr(_gnd_net_));
    defparam shift_srl_122_12_LC_11_20_2.C_ON=1'b0;
    defparam shift_srl_122_12_LC_11_20_2.SEQ_MODE=4'b1000;
    defparam shift_srl_122_12_LC_11_20_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_122_12_LC_11_20_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57706),
            .lcout(shift_srl_122Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93027),
            .ce(N__60051),
            .sr(_gnd_net_));
    defparam shift_srl_122_13_LC_11_20_3.C_ON=1'b0;
    defparam shift_srl_122_13_LC_11_20_3.SEQ_MODE=4'b1000;
    defparam shift_srl_122_13_LC_11_20_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_122_13_LC_11_20_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57700),
            .lcout(shift_srl_122Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93027),
            .ce(N__60051),
            .sr(_gnd_net_));
    defparam shift_srl_122_14_LC_11_20_4.C_ON=1'b0;
    defparam shift_srl_122_14_LC_11_20_4.SEQ_MODE=4'b1000;
    defparam shift_srl_122_14_LC_11_20_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_122_14_LC_11_20_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57694),
            .lcout(shift_srl_122Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93027),
            .ce(N__60051),
            .sr(_gnd_net_));
    defparam shift_srl_122_15_LC_11_20_5.C_ON=1'b0;
    defparam shift_srl_122_15_LC_11_20_5.SEQ_MODE=4'b1000;
    defparam shift_srl_122_15_LC_11_20_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_122_15_LC_11_20_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57688),
            .lcout(shift_srl_122Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93027),
            .ce(N__60051),
            .sr(_gnd_net_));
    defparam shift_srl_122_9_LC_11_20_6.C_ON=1'b0;
    defparam shift_srl_122_9_LC_11_20_6.SEQ_MODE=4'b1000;
    defparam shift_srl_122_9_LC_11_20_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_122_9_LC_11_20_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57676),
            .lcout(shift_srl_122Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93027),
            .ce(N__60051),
            .sr(_gnd_net_));
    defparam shift_srl_122_8_LC_11_20_7.C_ON=1'b0;
    defparam shift_srl_122_8_LC_11_20_7.SEQ_MODE=4'b1000;
    defparam shift_srl_122_8_LC_11_20_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_122_8_LC_11_20_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60061),
            .lcout(shift_srl_122Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93027),
            .ce(N__60051),
            .sr(_gnd_net_));
    defparam shift_srl_114_RNI6OUT_15_LC_11_21_0.C_ON=1'b0;
    defparam shift_srl_114_RNI6OUT_15_LC_11_21_0.SEQ_MODE=4'b0000;
    defparam shift_srl_114_RNI6OUT_15_LC_11_21_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_114_RNI6OUT_15_LC_11_21_0 (
            .in0(N__63814),
            .in1(N__58903),
            .in2(N__58803),
            .in3(N__60414),
            .lcout(rco_int_0_a3_0_a2_138_m6_0_a2_7_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_113_15_LC_11_21_1.C_ON=1'b0;
    defparam shift_srl_113_15_LC_11_21_1.SEQ_MODE=4'b1000;
    defparam shift_srl_113_15_LC_11_21_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_113_15_LC_11_21_1 (
            .in0(N__57808),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_113Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93042),
            .ce(N__57759),
            .sr(_gnd_net_));
    defparam shift_srl_113_14_LC_11_21_2.C_ON=1'b0;
    defparam shift_srl_113_14_LC_11_21_2.SEQ_MODE=4'b1000;
    defparam shift_srl_113_14_LC_11_21_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_113_14_LC_11_21_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57802),
            .lcout(shift_srl_113Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93042),
            .ce(N__57759),
            .sr(_gnd_net_));
    defparam shift_srl_113_13_LC_11_21_3.C_ON=1'b0;
    defparam shift_srl_113_13_LC_11_21_3.SEQ_MODE=4'b1000;
    defparam shift_srl_113_13_LC_11_21_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_113_13_LC_11_21_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57796),
            .lcout(shift_srl_113Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93042),
            .ce(N__57759),
            .sr(_gnd_net_));
    defparam shift_srl_113_12_LC_11_21_4.C_ON=1'b0;
    defparam shift_srl_113_12_LC_11_21_4.SEQ_MODE=4'b1000;
    defparam shift_srl_113_12_LC_11_21_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_113_12_LC_11_21_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57790),
            .lcout(shift_srl_113Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93042),
            .ce(N__57759),
            .sr(_gnd_net_));
    defparam shift_srl_113_11_LC_11_21_5.C_ON=1'b0;
    defparam shift_srl_113_11_LC_11_21_5.SEQ_MODE=4'b1000;
    defparam shift_srl_113_11_LC_11_21_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_113_11_LC_11_21_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57784),
            .lcout(shift_srl_113Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93042),
            .ce(N__57759),
            .sr(_gnd_net_));
    defparam shift_srl_113_10_LC_11_21_6.C_ON=1'b0;
    defparam shift_srl_113_10_LC_11_21_6.SEQ_MODE=4'b1000;
    defparam shift_srl_113_10_LC_11_21_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_113_10_LC_11_21_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57766),
            .lcout(shift_srl_113Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93042),
            .ce(N__57759),
            .sr(_gnd_net_));
    defparam shift_srl_113_9_LC_11_21_7.C_ON=1'b0;
    defparam shift_srl_113_9_LC_11_21_7.SEQ_MODE=4'b1000;
    defparam shift_srl_113_9_LC_11_21_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_113_9_LC_11_21_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57778),
            .lcout(shift_srl_113Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93042),
            .ce(N__57759),
            .sr(_gnd_net_));
    defparam shift_srl_112_10_LC_11_22_0.C_ON=1'b0;
    defparam shift_srl_112_10_LC_11_22_0.SEQ_MODE=4'b1000;
    defparam shift_srl_112_10_LC_11_22_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_112_10_LC_11_22_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57853),
            .lcout(shift_srl_112Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93056),
            .ce(N__60165),
            .sr(_gnd_net_));
    defparam shift_srl_112_11_LC_11_22_1.C_ON=1'b0;
    defparam shift_srl_112_11_LC_11_22_1.SEQ_MODE=4'b1000;
    defparam shift_srl_112_11_LC_11_22_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_112_11_LC_11_22_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57724),
            .lcout(shift_srl_112Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93056),
            .ce(N__60165),
            .sr(_gnd_net_));
    defparam shift_srl_112_12_LC_11_22_2.C_ON=1'b0;
    defparam shift_srl_112_12_LC_11_22_2.SEQ_MODE=4'b1000;
    defparam shift_srl_112_12_LC_11_22_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_112_12_LC_11_22_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57718),
            .lcout(shift_srl_112Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93056),
            .ce(N__60165),
            .sr(_gnd_net_));
    defparam shift_srl_112_13_LC_11_22_3.C_ON=1'b0;
    defparam shift_srl_112_13_LC_11_22_3.SEQ_MODE=4'b1000;
    defparam shift_srl_112_13_LC_11_22_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_112_13_LC_11_22_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57871),
            .lcout(shift_srl_112Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93056),
            .ce(N__60165),
            .sr(_gnd_net_));
    defparam shift_srl_112_14_LC_11_22_4.C_ON=1'b0;
    defparam shift_srl_112_14_LC_11_22_4.SEQ_MODE=4'b1000;
    defparam shift_srl_112_14_LC_11_22_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_112_14_LC_11_22_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57865),
            .lcout(shift_srl_112Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93056),
            .ce(N__60165),
            .sr(_gnd_net_));
    defparam shift_srl_112_9_LC_11_22_5.C_ON=1'b0;
    defparam shift_srl_112_9_LC_11_22_5.SEQ_MODE=4'b1000;
    defparam shift_srl_112_9_LC_11_22_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_112_9_LC_11_22_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57838),
            .lcout(shift_srl_112Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93056),
            .ce(N__60165),
            .sr(_gnd_net_));
    defparam shift_srl_112_8_LC_11_22_6.C_ON=1'b0;
    defparam shift_srl_112_8_LC_11_22_6.SEQ_MODE=4'b1000;
    defparam shift_srl_112_8_LC_11_22_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_112_8_LC_11_22_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57847),
            .lcout(shift_srl_112Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93056),
            .ce(N__60165),
            .sr(_gnd_net_));
    defparam shift_srl_109_10_LC_11_23_0.C_ON=1'b0;
    defparam shift_srl_109_10_LC_11_23_0.SEQ_MODE=4'b1000;
    defparam shift_srl_109_10_LC_11_23_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_109_10_LC_11_23_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57919),
            .lcout(shift_srl_109Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93072),
            .ce(N__57999),
            .sr(_gnd_net_));
    defparam shift_srl_109_11_LC_11_23_1.C_ON=1'b0;
    defparam shift_srl_109_11_LC_11_23_1.SEQ_MODE=4'b1000;
    defparam shift_srl_109_11_LC_11_23_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_109_11_LC_11_23_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57832),
            .lcout(shift_srl_109Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93072),
            .ce(N__57999),
            .sr(_gnd_net_));
    defparam shift_srl_109_12_LC_11_23_2.C_ON=1'b0;
    defparam shift_srl_109_12_LC_11_23_2.SEQ_MODE=4'b1000;
    defparam shift_srl_109_12_LC_11_23_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_109_12_LC_11_23_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57826),
            .lcout(shift_srl_109Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93072),
            .ce(N__57999),
            .sr(_gnd_net_));
    defparam shift_srl_109_13_LC_11_23_3.C_ON=1'b0;
    defparam shift_srl_109_13_LC_11_23_3.SEQ_MODE=4'b1000;
    defparam shift_srl_109_13_LC_11_23_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_109_13_LC_11_23_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57820),
            .lcout(shift_srl_109Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93072),
            .ce(N__57999),
            .sr(_gnd_net_));
    defparam shift_srl_109_14_LC_11_23_4.C_ON=1'b0;
    defparam shift_srl_109_14_LC_11_23_4.SEQ_MODE=4'b1000;
    defparam shift_srl_109_14_LC_11_23_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_109_14_LC_11_23_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57814),
            .lcout(shift_srl_109Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93072),
            .ce(N__57999),
            .sr(_gnd_net_));
    defparam shift_srl_109_15_LC_11_23_5.C_ON=1'b0;
    defparam shift_srl_109_15_LC_11_23_5.SEQ_MODE=4'b1000;
    defparam shift_srl_109_15_LC_11_23_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_109_15_LC_11_23_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57925),
            .lcout(shift_srl_109Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93072),
            .ce(N__57999),
            .sr(_gnd_net_));
    defparam shift_srl_109_9_LC_11_23_6.C_ON=1'b0;
    defparam shift_srl_109_9_LC_11_23_6.SEQ_MODE=4'b1000;
    defparam shift_srl_109_9_LC_11_23_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_109_9_LC_11_23_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57913),
            .lcout(shift_srl_109Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93072),
            .ce(N__57999),
            .sr(_gnd_net_));
    defparam shift_srl_109_8_LC_11_23_7.C_ON=1'b0;
    defparam shift_srl_109_8_LC_11_23_7.SEQ_MODE=4'b1000;
    defparam shift_srl_109_8_LC_11_23_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_109_8_LC_11_23_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58009),
            .lcout(shift_srl_109Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93072),
            .ce(N__57999),
            .sr(_gnd_net_));
    defparam shift_srl_109_0_LC_11_24_0.C_ON=1'b0;
    defparam shift_srl_109_0_LC_11_24_0.SEQ_MODE=4'b1000;
    defparam shift_srl_109_0_LC_11_24_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_109_0_LC_11_24_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62401),
            .lcout(shift_srl_109Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93087),
            .ce(N__58003),
            .sr(_gnd_net_));
    defparam shift_srl_109_1_LC_11_24_1.C_ON=1'b0;
    defparam shift_srl_109_1_LC_11_24_1.SEQ_MODE=4'b1000;
    defparam shift_srl_109_1_LC_11_24_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_109_1_LC_11_24_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57907),
            .lcout(shift_srl_109Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93087),
            .ce(N__58003),
            .sr(_gnd_net_));
    defparam shift_srl_109_2_LC_11_24_2.C_ON=1'b0;
    defparam shift_srl_109_2_LC_11_24_2.SEQ_MODE=4'b1000;
    defparam shift_srl_109_2_LC_11_24_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_109_2_LC_11_24_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57901),
            .lcout(shift_srl_109Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93087),
            .ce(N__58003),
            .sr(_gnd_net_));
    defparam shift_srl_109_3_LC_11_24_3.C_ON=1'b0;
    defparam shift_srl_109_3_LC_11_24_3.SEQ_MODE=4'b1000;
    defparam shift_srl_109_3_LC_11_24_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_109_3_LC_11_24_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57895),
            .lcout(shift_srl_109Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93087),
            .ce(N__58003),
            .sr(_gnd_net_));
    defparam shift_srl_109_4_LC_11_24_4.C_ON=1'b0;
    defparam shift_srl_109_4_LC_11_24_4.SEQ_MODE=4'b1000;
    defparam shift_srl_109_4_LC_11_24_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_109_4_LC_11_24_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57889),
            .lcout(shift_srl_109Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93087),
            .ce(N__58003),
            .sr(_gnd_net_));
    defparam shift_srl_109_5_LC_11_24_5.C_ON=1'b0;
    defparam shift_srl_109_5_LC_11_24_5.SEQ_MODE=4'b1000;
    defparam shift_srl_109_5_LC_11_24_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_109_5_LC_11_24_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57883),
            .lcout(shift_srl_109Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93087),
            .ce(N__58003),
            .sr(_gnd_net_));
    defparam shift_srl_109_6_LC_11_24_6.C_ON=1'b0;
    defparam shift_srl_109_6_LC_11_24_6.SEQ_MODE=4'b1000;
    defparam shift_srl_109_6_LC_11_24_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_109_6_LC_11_24_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57877),
            .lcout(shift_srl_109Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93087),
            .ce(N__58003),
            .sr(_gnd_net_));
    defparam shift_srl_109_7_LC_11_24_7.C_ON=1'b0;
    defparam shift_srl_109_7_LC_11_24_7.SEQ_MODE=4'b1000;
    defparam shift_srl_109_7_LC_11_24_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_109_7_LC_11_24_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58015),
            .lcout(shift_srl_109Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93087),
            .ce(N__58003),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_105_LC_11_25_0.C_ON=1'b0;
    defparam rco_obuf_RNO_105_LC_11_25_0.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_105_LC_11_25_0.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_105_LC_11_25_0 (
            .in0(N__59289),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79252),
            .lcout(rco_c_105),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_105_0_LC_11_25_1.C_ON=1'b0;
    defparam shift_srl_105_0_LC_11_25_1.SEQ_MODE=4'b1000;
    defparam shift_srl_105_0_LC_11_25_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_105_0_LC_11_25_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59288),
            .lcout(shift_srl_105Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93100),
            .ce(N__58060),
            .sr(_gnd_net_));
    defparam shift_srl_105_1_LC_11_25_2.C_ON=1'b0;
    defparam shift_srl_105_1_LC_11_25_2.SEQ_MODE=4'b1000;
    defparam shift_srl_105_1_LC_11_25_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_105_1_LC_11_25_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57967),
            .lcout(shift_srl_105Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93100),
            .ce(N__58060),
            .sr(_gnd_net_));
    defparam shift_srl_105_2_LC_11_25_3.C_ON=1'b0;
    defparam shift_srl_105_2_LC_11_25_3.SEQ_MODE=4'b1000;
    defparam shift_srl_105_2_LC_11_25_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_105_2_LC_11_25_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57961),
            .lcout(shift_srl_105Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93100),
            .ce(N__58060),
            .sr(_gnd_net_));
    defparam shift_srl_105_3_LC_11_25_4.C_ON=1'b0;
    defparam shift_srl_105_3_LC_11_25_4.SEQ_MODE=4'b1000;
    defparam shift_srl_105_3_LC_11_25_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_105_3_LC_11_25_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57955),
            .lcout(shift_srl_105Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93100),
            .ce(N__58060),
            .sr(_gnd_net_));
    defparam shift_srl_105_4_LC_11_25_5.C_ON=1'b0;
    defparam shift_srl_105_4_LC_11_25_5.SEQ_MODE=4'b1000;
    defparam shift_srl_105_4_LC_11_25_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_105_4_LC_11_25_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57949),
            .lcout(shift_srl_105Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93100),
            .ce(N__58060),
            .sr(_gnd_net_));
    defparam shift_srl_105_10_LC_11_26_0.C_ON=1'b0;
    defparam shift_srl_105_10_LC_11_26_0.SEQ_MODE=4'b1000;
    defparam shift_srl_105_10_LC_11_26_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_105_10_LC_11_26_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58081),
            .lcout(shift_srl_105Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93119),
            .ce(N__58059),
            .sr(_gnd_net_));
    defparam shift_srl_105_11_LC_11_26_1.C_ON=1'b0;
    defparam shift_srl_105_11_LC_11_26_1.SEQ_MODE=4'b1000;
    defparam shift_srl_105_11_LC_11_26_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_105_11_LC_11_26_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57931),
            .lcout(shift_srl_105Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93119),
            .ce(N__58059),
            .sr(_gnd_net_));
    defparam shift_srl_105_12_LC_11_26_2.C_ON=1'b0;
    defparam shift_srl_105_12_LC_11_26_2.SEQ_MODE=4'b1000;
    defparam shift_srl_105_12_LC_11_26_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_105_12_LC_11_26_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58105),
            .lcout(shift_srl_105Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93119),
            .ce(N__58059),
            .sr(_gnd_net_));
    defparam shift_srl_105_13_LC_11_26_3.C_ON=1'b0;
    defparam shift_srl_105_13_LC_11_26_3.SEQ_MODE=4'b1000;
    defparam shift_srl_105_13_LC_11_26_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_105_13_LC_11_26_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58099),
            .lcout(shift_srl_105Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93119),
            .ce(N__58059),
            .sr(_gnd_net_));
    defparam shift_srl_105_14_LC_11_26_4.C_ON=1'b0;
    defparam shift_srl_105_14_LC_11_26_4.SEQ_MODE=4'b1000;
    defparam shift_srl_105_14_LC_11_26_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_105_14_LC_11_26_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58093),
            .lcout(shift_srl_105Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93119),
            .ce(N__58059),
            .sr(_gnd_net_));
    defparam shift_srl_105_15_LC_11_26_5.C_ON=1'b0;
    defparam shift_srl_105_15_LC_11_26_5.SEQ_MODE=4'b1000;
    defparam shift_srl_105_15_LC_11_26_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_105_15_LC_11_26_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58087),
            .lcout(shift_srl_105Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93119),
            .ce(N__58059),
            .sr(_gnd_net_));
    defparam shift_srl_105_9_LC_11_26_6.C_ON=1'b0;
    defparam shift_srl_105_9_LC_11_26_6.SEQ_MODE=4'b1000;
    defparam shift_srl_105_9_LC_11_26_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_105_9_LC_11_26_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58066),
            .lcout(shift_srl_105Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93119),
            .ce(N__58059),
            .sr(_gnd_net_));
    defparam shift_srl_105_8_LC_11_26_7.C_ON=1'b0;
    defparam shift_srl_105_8_LC_11_26_7.SEQ_MODE=4'b1000;
    defparam shift_srl_105_8_LC_11_26_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_105_8_LC_11_26_7 (
            .in0(N__58075),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_105Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93119),
            .ce(N__58059),
            .sr(_gnd_net_));
    defparam shift_srl_104_0_LC_11_27_0.C_ON=1'b0;
    defparam shift_srl_104_0_LC_11_27_0.SEQ_MODE=4'b1000;
    defparam shift_srl_104_0_LC_11_27_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_104_0_LC_11_27_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61000),
            .lcout(shift_srl_104Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93139),
            .ce(N__59307),
            .sr(_gnd_net_));
    defparam shift_srl_104_1_LC_11_27_1.C_ON=1'b0;
    defparam shift_srl_104_1_LC_11_27_1.SEQ_MODE=4'b1000;
    defparam shift_srl_104_1_LC_11_27_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_104_1_LC_11_27_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58027),
            .lcout(shift_srl_104Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93139),
            .ce(N__59307),
            .sr(_gnd_net_));
    defparam shift_srl_104_2_LC_11_27_2.C_ON=1'b0;
    defparam shift_srl_104_2_LC_11_27_2.SEQ_MODE=4'b1000;
    defparam shift_srl_104_2_LC_11_27_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_104_2_LC_11_27_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58021),
            .lcout(shift_srl_104Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93139),
            .ce(N__59307),
            .sr(_gnd_net_));
    defparam shift_srl_104_3_LC_11_27_3.C_ON=1'b0;
    defparam shift_srl_104_3_LC_11_27_3.SEQ_MODE=4'b1000;
    defparam shift_srl_104_3_LC_11_27_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_104_3_LC_11_27_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58153),
            .lcout(shift_srl_104Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93139),
            .ce(N__59307),
            .sr(_gnd_net_));
    defparam shift_srl_104_4_LC_11_27_4.C_ON=1'b0;
    defparam shift_srl_104_4_LC_11_27_4.SEQ_MODE=4'b1000;
    defparam shift_srl_104_4_LC_11_27_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_104_4_LC_11_27_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58147),
            .lcout(shift_srl_104Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93139),
            .ce(N__59307),
            .sr(_gnd_net_));
    defparam shift_srl_104_5_LC_11_27_5.C_ON=1'b0;
    defparam shift_srl_104_5_LC_11_27_5.SEQ_MODE=4'b1000;
    defparam shift_srl_104_5_LC_11_27_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_104_5_LC_11_27_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58141),
            .lcout(shift_srl_104Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93139),
            .ce(N__59307),
            .sr(_gnd_net_));
    defparam shift_srl_104_6_LC_11_27_6.C_ON=1'b0;
    defparam shift_srl_104_6_LC_11_27_6.SEQ_MODE=4'b1000;
    defparam shift_srl_104_6_LC_11_27_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_104_6_LC_11_27_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58135),
            .lcout(shift_srl_104Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93139),
            .ce(N__59307),
            .sr(_gnd_net_));
    defparam shift_srl_104_7_LC_11_27_7.C_ON=1'b0;
    defparam shift_srl_104_7_LC_11_27_7.SEQ_MODE=4'b1000;
    defparam shift_srl_104_7_LC_11_27_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_104_7_LC_11_27_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58129),
            .lcout(shift_srl_104Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93139),
            .ce(N__59307),
            .sr(_gnd_net_));
    defparam shift_srl_101_10_LC_11_28_0.C_ON=1'b0;
    defparam shift_srl_101_10_LC_11_28_0.SEQ_MODE=4'b1000;
    defparam shift_srl_101_10_LC_11_28_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_101_10_LC_11_28_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58204),
            .lcout(shift_srl_101Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93157),
            .ce(N__59205),
            .sr(_gnd_net_));
    defparam shift_srl_101_11_LC_11_28_1.C_ON=1'b0;
    defparam shift_srl_101_11_LC_11_28_1.SEQ_MODE=4'b1000;
    defparam shift_srl_101_11_LC_11_28_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_101_11_LC_11_28_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58123),
            .lcout(shift_srl_101Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93157),
            .ce(N__59205),
            .sr(_gnd_net_));
    defparam shift_srl_101_12_LC_11_28_2.C_ON=1'b0;
    defparam shift_srl_101_12_LC_11_28_2.SEQ_MODE=4'b1000;
    defparam shift_srl_101_12_LC_11_28_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_101_12_LC_11_28_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58117),
            .lcout(shift_srl_101Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93157),
            .ce(N__59205),
            .sr(_gnd_net_));
    defparam shift_srl_101_13_LC_11_28_3.C_ON=1'b0;
    defparam shift_srl_101_13_LC_11_28_3.SEQ_MODE=4'b1000;
    defparam shift_srl_101_13_LC_11_28_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_101_13_LC_11_28_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58111),
            .lcout(shift_srl_101Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93157),
            .ce(N__59205),
            .sr(_gnd_net_));
    defparam shift_srl_101_14_LC_11_28_4.C_ON=1'b0;
    defparam shift_srl_101_14_LC_11_28_4.SEQ_MODE=4'b1000;
    defparam shift_srl_101_14_LC_11_28_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_101_14_LC_11_28_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58210),
            .lcout(shift_srl_101Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93157),
            .ce(N__59205),
            .sr(_gnd_net_));
    defparam shift_srl_101_9_LC_11_28_5.C_ON=1'b0;
    defparam shift_srl_101_9_LC_11_28_5.SEQ_MODE=4'b1000;
    defparam shift_srl_101_9_LC_11_28_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_101_9_LC_11_28_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58198),
            .lcout(shift_srl_101Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93157),
            .ce(N__59205),
            .sr(_gnd_net_));
    defparam shift_srl_101_8_LC_11_28_6.C_ON=1'b0;
    defparam shift_srl_101_8_LC_11_28_6.SEQ_MODE=4'b1000;
    defparam shift_srl_101_8_LC_11_28_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_101_8_LC_11_28_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58192),
            .lcout(shift_srl_101Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93157),
            .ce(N__59205),
            .sr(_gnd_net_));
    defparam shift_srl_101_7_LC_11_28_7.C_ON=1'b0;
    defparam shift_srl_101_7_LC_11_28_7.SEQ_MODE=4'b1000;
    defparam shift_srl_101_7_LC_11_28_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_101_7_LC_11_28_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58318),
            .lcout(shift_srl_101Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93157),
            .ce(N__59205),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_101_LC_11_29_1.C_ON=1'b0;
    defparam rco_obuf_RNO_101_LC_11_29_1.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_101_LC_11_29_1.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_101_LC_11_29_1 (
            .in0(N__60985),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79642),
            .lcout(rco_c_101),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_101_0_LC_11_29_2.C_ON=1'b0;
    defparam shift_srl_101_0_LC_11_29_2.SEQ_MODE=4'b1000;
    defparam shift_srl_101_0_LC_11_29_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_101_0_LC_11_29_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60984),
            .lcout(shift_srl_101Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93177),
            .ce(N__59204),
            .sr(_gnd_net_));
    defparam shift_srl_101_1_LC_11_29_3.C_ON=1'b0;
    defparam shift_srl_101_1_LC_11_29_3.SEQ_MODE=4'b1000;
    defparam shift_srl_101_1_LC_11_29_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_101_1_LC_11_29_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58171),
            .lcout(shift_srl_101Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93177),
            .ce(N__59204),
            .sr(_gnd_net_));
    defparam shift_srl_101_2_LC_11_29_4.C_ON=1'b0;
    defparam shift_srl_101_2_LC_11_29_4.SEQ_MODE=4'b1000;
    defparam shift_srl_101_2_LC_11_29_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_101_2_LC_11_29_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58165),
            .lcout(shift_srl_101Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93177),
            .ce(N__59204),
            .sr(_gnd_net_));
    defparam shift_srl_101_3_LC_11_29_5.C_ON=1'b0;
    defparam shift_srl_101_3_LC_11_29_5.SEQ_MODE=4'b1000;
    defparam shift_srl_101_3_LC_11_29_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_101_3_LC_11_29_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58159),
            .lcout(shift_srl_101Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93177),
            .ce(N__59204),
            .sr(_gnd_net_));
    defparam shift_srl_101_4_LC_11_29_6.C_ON=1'b0;
    defparam shift_srl_101_4_LC_11_29_6.SEQ_MODE=4'b1000;
    defparam shift_srl_101_4_LC_11_29_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_101_4_LC_11_29_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58336),
            .lcout(shift_srl_101Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93177),
            .ce(N__59204),
            .sr(_gnd_net_));
    defparam shift_srl_101_5_LC_11_29_7.C_ON=1'b0;
    defparam shift_srl_101_5_LC_11_29_7.SEQ_MODE=4'b1000;
    defparam shift_srl_101_5_LC_11_29_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_101_5_LC_11_29_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58330),
            .lcout(shift_srl_101Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93177),
            .ce(N__59204),
            .sr(_gnd_net_));
    defparam shift_srl_101_6_LC_11_30_0.C_ON=1'b0;
    defparam shift_srl_101_6_LC_11_30_0.SEQ_MODE=4'b1000;
    defparam shift_srl_101_6_LC_11_30_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_101_6_LC_11_30_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58324),
            .lcout(shift_srl_101Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93199),
            .ce(N__59206),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_149_LC_12_4_1.C_ON=1'b0;
    defparam rco_obuf_RNO_149_LC_12_4_1.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_149_LC_12_4_1.LUT_INIT=16'b1100110000000000;
    LogicCell40 rco_obuf_RNO_149_LC_12_4_1 (
            .in0(_gnd_net_),
            .in1(N__58309),
            .in2(_gnd_net_),
            .in3(N__82198),
            .lcout(rco_c_149),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_148_6_LC_12_8_0.C_ON=1'b0;
    defparam shift_srl_148_6_LC_12_8_0.SEQ_MODE=4'b1000;
    defparam shift_srl_148_6_LC_12_8_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_148_6_LC_12_8_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58249),
            .lcout(shift_srl_148Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93141),
            .ce(N__58243),
            .sr(_gnd_net_));
    defparam shift_srl_148_7_LC_12_8_1.C_ON=1'b0;
    defparam shift_srl_148_7_LC_12_8_1.SEQ_MODE=4'b1000;
    defparam shift_srl_148_7_LC_12_8_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_148_7_LC_12_8_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58279),
            .lcout(shift_srl_148Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93141),
            .ce(N__58243),
            .sr(_gnd_net_));
    defparam shift_srl_148_4_LC_12_8_4.C_ON=1'b0;
    defparam shift_srl_148_4_LC_12_8_4.SEQ_MODE=4'b1000;
    defparam shift_srl_148_4_LC_12_8_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_148_4_LC_12_8_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58261),
            .lcout(shift_srl_148Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93141),
            .ce(N__58243),
            .sr(_gnd_net_));
    defparam shift_srl_148_3_LC_12_8_6.C_ON=1'b0;
    defparam shift_srl_148_3_LC_12_8_6.SEQ_MODE=4'b1000;
    defparam shift_srl_148_3_LC_12_8_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_148_3_LC_12_8_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58267),
            .lcout(shift_srl_148Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93141),
            .ce(N__58243),
            .sr(_gnd_net_));
    defparam shift_srl_148_5_LC_12_8_7.C_ON=1'b0;
    defparam shift_srl_148_5_LC_12_8_7.SEQ_MODE=4'b1000;
    defparam shift_srl_148_5_LC_12_8_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_148_5_LC_12_8_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58255),
            .lcout(shift_srl_148Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93141),
            .ce(N__58243),
            .sr(_gnd_net_));
    defparam shift_srl_25_3_LC_12_9_3.C_ON=1'b0;
    defparam shift_srl_25_3_LC_12_9_3.SEQ_MODE=4'b1000;
    defparam shift_srl_25_3_LC_12_9_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_25_3_LC_12_9_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58372),
            .lcout(shift_srl_25Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93122),
            .ce(N__59573),
            .sr(_gnd_net_));
    defparam shift_srl_25_4_LC_12_9_6.C_ON=1'b0;
    defparam shift_srl_25_4_LC_12_9_6.SEQ_MODE=4'b1000;
    defparam shift_srl_25_4_LC_12_9_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_25_4_LC_12_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58390),
            .lcout(shift_srl_25Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93122),
            .ce(N__59573),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIPBKF6_15_LC_12_10_0.C_ON=1'b0;
    defparam shift_srl_0_RNIPBKF6_15_LC_12_10_0.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIPBKF6_15_LC_12_10_0.LUT_INIT=16'b1100110000000000;
    LogicCell40 shift_srl_0_RNIPBKF6_15_LC_12_10_0 (
            .in0(_gnd_net_),
            .in1(N__89765),
            .in2(_gnd_net_),
            .in3(N__58359),
            .lcout(clk_en_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_25_0_LC_12_10_2.C_ON=1'b0;
    defparam shift_srl_25_0_LC_12_10_2.SEQ_MODE=4'b1000;
    defparam shift_srl_25_0_LC_12_10_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_25_0_LC_12_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71463),
            .lcout(shift_srl_25Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93102),
            .ce(N__59572),
            .sr(_gnd_net_));
    defparam shift_srl_25_1_LC_12_10_3.C_ON=1'b0;
    defparam shift_srl_25_1_LC_12_10_3.SEQ_MODE=4'b1000;
    defparam shift_srl_25_1_LC_12_10_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_25_1_LC_12_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58384),
            .lcout(shift_srl_25Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93102),
            .ce(N__59572),
            .sr(_gnd_net_));
    defparam shift_srl_25_2_LC_12_10_4.C_ON=1'b0;
    defparam shift_srl_25_2_LC_12_10_4.SEQ_MODE=4'b1000;
    defparam shift_srl_25_2_LC_12_10_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_25_2_LC_12_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58378),
            .lcout(shift_srl_25Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93102),
            .ce(N__59572),
            .sr(_gnd_net_));
    defparam shift_srl_24_RNIUVPE6_15_LC_12_11_5.C_ON=1'b0;
    defparam shift_srl_24_RNIUVPE6_15_LC_12_11_5.SEQ_MODE=4'b0000;
    defparam shift_srl_24_RNIUVPE6_15_LC_12_11_5.LUT_INIT=16'b1100110000000000;
    LogicCell40 shift_srl_24_RNIUVPE6_15_LC_12_11_5 (
            .in0(_gnd_net_),
            .in1(N__83796),
            .in2(_gnd_net_),
            .in3(N__85197),
            .lcout(rco_c_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_157_0_LC_12_14_0.C_ON=1'b0;
    defparam shift_srl_157_0_LC_12_14_0.SEQ_MODE=4'b1000;
    defparam shift_srl_157_0_LC_12_14_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_157_0_LC_12_14_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77871),
            .lcout(shift_srl_157Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93043),
            .ce(N__58414),
            .sr(_gnd_net_));
    defparam shift_srl_157_1_LC_12_14_1.C_ON=1'b0;
    defparam shift_srl_157_1_LC_12_14_1.SEQ_MODE=4'b1000;
    defparam shift_srl_157_1_LC_12_14_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_157_1_LC_12_14_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58348),
            .lcout(shift_srl_157Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93043),
            .ce(N__58414),
            .sr(_gnd_net_));
    defparam shift_srl_157_2_LC_12_14_2.C_ON=1'b0;
    defparam shift_srl_157_2_LC_12_14_2.SEQ_MODE=4'b1000;
    defparam shift_srl_157_2_LC_12_14_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_157_2_LC_12_14_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58342),
            .lcout(shift_srl_157Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93043),
            .ce(N__58414),
            .sr(_gnd_net_));
    defparam shift_srl_157_3_LC_12_14_3.C_ON=1'b0;
    defparam shift_srl_157_3_LC_12_14_3.SEQ_MODE=4'b1000;
    defparam shift_srl_157_3_LC_12_14_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_157_3_LC_12_14_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58462),
            .lcout(shift_srl_157Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93043),
            .ce(N__58414),
            .sr(_gnd_net_));
    defparam shift_srl_157_4_LC_12_14_4.C_ON=1'b0;
    defparam shift_srl_157_4_LC_12_14_4.SEQ_MODE=4'b1000;
    defparam shift_srl_157_4_LC_12_14_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_157_4_LC_12_14_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58456),
            .lcout(shift_srl_157Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93043),
            .ce(N__58414),
            .sr(_gnd_net_));
    defparam shift_srl_157_13_LC_12_14_5.C_ON=1'b0;
    defparam shift_srl_157_13_LC_12_14_5.SEQ_MODE=4'b1000;
    defparam shift_srl_157_13_LC_12_14_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_157_13_LC_12_14_5 (
            .in0(N__58444),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_157Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93043),
            .ce(N__58414),
            .sr(_gnd_net_));
    defparam shift_srl_157_14_LC_12_14_6.C_ON=1'b0;
    defparam shift_srl_157_14_LC_12_14_6.SEQ_MODE=4'b1000;
    defparam shift_srl_157_14_LC_12_14_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_157_14_LC_12_14_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58438),
            .lcout(shift_srl_157Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93043),
            .ce(N__58414),
            .sr(_gnd_net_));
    defparam shift_srl_157_7_LC_12_14_7.C_ON=1'b0;
    defparam shift_srl_157_7_LC_12_14_7.SEQ_MODE=4'b1000;
    defparam shift_srl_157_7_LC_12_14_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_157_7_LC_12_14_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58426),
            .lcout(shift_srl_157Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93043),
            .ce(N__58414),
            .sr(_gnd_net_));
    defparam shift_srl_155_0_LC_12_15_0.C_ON=1'b0;
    defparam shift_srl_155_0_LC_12_15_0.SEQ_MODE=4'b1000;
    defparam shift_srl_155_0_LC_12_15_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_155_0_LC_12_15_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77632),
            .lcout(shift_srl_155Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93028),
            .ce(N__58551),
            .sr(_gnd_net_));
    defparam shift_srl_155_1_LC_12_15_1.C_ON=1'b0;
    defparam shift_srl_155_1_LC_12_15_1.SEQ_MODE=4'b1000;
    defparam shift_srl_155_1_LC_12_15_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_155_1_LC_12_15_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58402),
            .lcout(shift_srl_155Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93028),
            .ce(N__58551),
            .sr(_gnd_net_));
    defparam shift_srl_155_2_LC_12_15_2.C_ON=1'b0;
    defparam shift_srl_155_2_LC_12_15_2.SEQ_MODE=4'b1000;
    defparam shift_srl_155_2_LC_12_15_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_155_2_LC_12_15_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58396),
            .lcout(shift_srl_155Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93028),
            .ce(N__58551),
            .sr(_gnd_net_));
    defparam shift_srl_155_7_LC_12_15_3.C_ON=1'b0;
    defparam shift_srl_155_7_LC_12_15_3.SEQ_MODE=4'b1000;
    defparam shift_srl_155_7_LC_12_15_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_155_7_LC_12_15_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58510),
            .lcout(shift_srl_155Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93028),
            .ce(N__58551),
            .sr(_gnd_net_));
    defparam shift_srl_155_6_LC_12_15_4.C_ON=1'b0;
    defparam shift_srl_155_6_LC_12_15_4.SEQ_MODE=4'b1000;
    defparam shift_srl_155_6_LC_12_15_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_155_6_LC_12_15_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58498),
            .lcout(shift_srl_155Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93028),
            .ce(N__58551),
            .sr(_gnd_net_));
    defparam shift_srl_155_9_LC_12_15_5.C_ON=1'b0;
    defparam shift_srl_155_9_LC_12_15_5.SEQ_MODE=4'b1000;
    defparam shift_srl_155_9_LC_12_15_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_155_9_LC_12_15_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58480),
            .lcout(shift_srl_155Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93028),
            .ce(N__58551),
            .sr(_gnd_net_));
    defparam shift_srl_155_10_LC_12_15_6.C_ON=1'b0;
    defparam shift_srl_155_10_LC_12_15_6.SEQ_MODE=4'b1000;
    defparam shift_srl_155_10_LC_12_15_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_155_10_LC_12_15_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58504),
            .lcout(shift_srl_155Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93028),
            .ce(N__58551),
            .sr(_gnd_net_));
    defparam shift_srl_155_5_LC_12_15_7.C_ON=1'b0;
    defparam shift_srl_155_5_LC_12_15_7.SEQ_MODE=4'b1000;
    defparam shift_srl_155_5_LC_12_15_7.LUT_INIT=16'b1100110011001100;
    LogicCell40 shift_srl_155_5_LC_12_15_7 (
            .in0(_gnd_net_),
            .in1(N__58492),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_155Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93028),
            .ce(N__58551),
            .sr(_gnd_net_));
    defparam shift_srl_155_4_LC_12_16_0.C_ON=1'b0;
    defparam shift_srl_155_4_LC_12_16_0.SEQ_MODE=4'b1000;
    defparam shift_srl_155_4_LC_12_16_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_155_4_LC_12_16_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58570),
            .lcout(shift_srl_155Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93015),
            .ce(N__58552),
            .sr(_gnd_net_));
    defparam shift_srl_155_8_LC_12_16_1.C_ON=1'b0;
    defparam shift_srl_155_8_LC_12_16_1.SEQ_MODE=4'b1000;
    defparam shift_srl_155_8_LC_12_16_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_155_8_LC_12_16_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58486),
            .lcout(shift_srl_155Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93015),
            .ce(N__58552),
            .sr(_gnd_net_));
    defparam shift_srl_155_12_LC_12_16_2.C_ON=1'b0;
    defparam shift_srl_155_12_LC_12_16_2.SEQ_MODE=4'b1000;
    defparam shift_srl_155_12_LC_12_16_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_155_12_LC_12_16_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58558),
            .lcout(shift_srl_155Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93015),
            .ce(N__58552),
            .sr(_gnd_net_));
    defparam shift_srl_155_13_LC_12_16_3.C_ON=1'b0;
    defparam shift_srl_155_13_LC_12_16_3.SEQ_MODE=4'b1000;
    defparam shift_srl_155_13_LC_12_16_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_155_13_LC_12_16_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58474),
            .lcout(shift_srl_155Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93015),
            .ce(N__58552),
            .sr(_gnd_net_));
    defparam shift_srl_155_14_LC_12_16_4.C_ON=1'b0;
    defparam shift_srl_155_14_LC_12_16_4.SEQ_MODE=4'b1000;
    defparam shift_srl_155_14_LC_12_16_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_155_14_LC_12_16_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58468),
            .lcout(shift_srl_155Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93015),
            .ce(N__58552),
            .sr(_gnd_net_));
    defparam shift_srl_155_15_LC_12_16_5.C_ON=1'b0;
    defparam shift_srl_155_15_LC_12_16_5.SEQ_MODE=4'b1000;
    defparam shift_srl_155_15_LC_12_16_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_155_15_LC_12_16_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58582),
            .lcout(shift_srl_155Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93015),
            .ce(N__58552),
            .sr(_gnd_net_));
    defparam shift_srl_155_3_LC_12_16_6.C_ON=1'b0;
    defparam shift_srl_155_3_LC_12_16_6.SEQ_MODE=4'b1000;
    defparam shift_srl_155_3_LC_12_16_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_155_3_LC_12_16_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58576),
            .lcout(shift_srl_155Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93015),
            .ce(N__58552),
            .sr(_gnd_net_));
    defparam shift_srl_155_11_LC_12_16_7.C_ON=1'b0;
    defparam shift_srl_155_11_LC_12_16_7.SEQ_MODE=4'b1000;
    defparam shift_srl_155_11_LC_12_16_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_155_11_LC_12_16_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58564),
            .lcout(shift_srl_155Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93015),
            .ce(N__58552),
            .sr(_gnd_net_));
    defparam shift_srl_124_0_LC_12_17_0.C_ON=1'b0;
    defparam shift_srl_124_0_LC_12_17_0.SEQ_MODE=4'b1000;
    defparam shift_srl_124_0_LC_12_17_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_124_0_LC_12_17_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65439),
            .lcout(shift_srl_124Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92996),
            .ce(N__58718),
            .sr(_gnd_net_));
    defparam shift_srl_124_1_LC_12_17_1.C_ON=1'b0;
    defparam shift_srl_124_1_LC_12_17_1.SEQ_MODE=4'b1000;
    defparam shift_srl_124_1_LC_12_17_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_124_1_LC_12_17_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58540),
            .lcout(shift_srl_124Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92996),
            .ce(N__58718),
            .sr(_gnd_net_));
    defparam shift_srl_124_2_LC_12_17_2.C_ON=1'b0;
    defparam shift_srl_124_2_LC_12_17_2.SEQ_MODE=4'b1000;
    defparam shift_srl_124_2_LC_12_17_2.LUT_INIT=16'b1100110011001100;
    LogicCell40 shift_srl_124_2_LC_12_17_2 (
            .in0(_gnd_net_),
            .in1(N__58534),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_124Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92996),
            .ce(N__58718),
            .sr(_gnd_net_));
    defparam shift_srl_124_3_LC_12_17_3.C_ON=1'b0;
    defparam shift_srl_124_3_LC_12_17_3.SEQ_MODE=4'b1000;
    defparam shift_srl_124_3_LC_12_17_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_124_3_LC_12_17_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58528),
            .lcout(shift_srl_124Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92996),
            .ce(N__58718),
            .sr(_gnd_net_));
    defparam shift_srl_124_4_LC_12_17_4.C_ON=1'b0;
    defparam shift_srl_124_4_LC_12_17_4.SEQ_MODE=4'b1000;
    defparam shift_srl_124_4_LC_12_17_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_124_4_LC_12_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58522),
            .lcout(shift_srl_124Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92996),
            .ce(N__58718),
            .sr(_gnd_net_));
    defparam shift_srl_124_5_LC_12_17_5.C_ON=1'b0;
    defparam shift_srl_124_5_LC_12_17_5.SEQ_MODE=4'b1000;
    defparam shift_srl_124_5_LC_12_17_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_124_5_LC_12_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58516),
            .lcout(shift_srl_124Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92996),
            .ce(N__58718),
            .sr(_gnd_net_));
    defparam shift_srl_124_6_LC_12_17_6.C_ON=1'b0;
    defparam shift_srl_124_6_LC_12_17_6.SEQ_MODE=4'b1000;
    defparam shift_srl_124_6_LC_12_17_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_124_6_LC_12_17_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58636),
            .lcout(shift_srl_124Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92996),
            .ce(N__58718),
            .sr(_gnd_net_));
    defparam shift_srl_124_7_LC_12_17_7.C_ON=1'b0;
    defparam shift_srl_124_7_LC_12_17_7.SEQ_MODE=4'b1000;
    defparam shift_srl_124_7_LC_12_17_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_124_7_LC_12_17_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58630),
            .lcout(shift_srl_124Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__92996),
            .ce(N__58718),
            .sr(_gnd_net_));
    defparam shift_srl_144_0_LC_12_18_0.C_ON=1'b0;
    defparam shift_srl_144_0_LC_12_18_0.SEQ_MODE=4'b1000;
    defparam shift_srl_144_0_LC_12_18_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_144_0_LC_12_18_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61819),
            .lcout(shift_srl_144Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93016),
            .ce(N__59989),
            .sr(_gnd_net_));
    defparam shift_srl_144_1_LC_12_18_1.C_ON=1'b0;
    defparam shift_srl_144_1_LC_12_18_1.SEQ_MODE=4'b1000;
    defparam shift_srl_144_1_LC_12_18_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_144_1_LC_12_18_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58618),
            .lcout(shift_srl_144Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93016),
            .ce(N__59989),
            .sr(_gnd_net_));
    defparam shift_srl_144_2_LC_12_18_2.C_ON=1'b0;
    defparam shift_srl_144_2_LC_12_18_2.SEQ_MODE=4'b1000;
    defparam shift_srl_144_2_LC_12_18_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_144_2_LC_12_18_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58612),
            .lcout(shift_srl_144Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93016),
            .ce(N__59989),
            .sr(_gnd_net_));
    defparam shift_srl_144_3_LC_12_18_3.C_ON=1'b0;
    defparam shift_srl_144_3_LC_12_18_3.SEQ_MODE=4'b1000;
    defparam shift_srl_144_3_LC_12_18_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_144_3_LC_12_18_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58606),
            .lcout(shift_srl_144Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93016),
            .ce(N__59989),
            .sr(_gnd_net_));
    defparam shift_srl_144_4_LC_12_18_4.C_ON=1'b0;
    defparam shift_srl_144_4_LC_12_18_4.SEQ_MODE=4'b1000;
    defparam shift_srl_144_4_LC_12_18_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_144_4_LC_12_18_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58600),
            .lcout(shift_srl_144Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93016),
            .ce(N__59989),
            .sr(_gnd_net_));
    defparam shift_srl_144_5_LC_12_18_5.C_ON=1'b0;
    defparam shift_srl_144_5_LC_12_18_5.SEQ_MODE=4'b1000;
    defparam shift_srl_144_5_LC_12_18_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_144_5_LC_12_18_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58594),
            .lcout(shift_srl_144Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93016),
            .ce(N__59989),
            .sr(_gnd_net_));
    defparam shift_srl_144_6_LC_12_18_6.C_ON=1'b0;
    defparam shift_srl_144_6_LC_12_18_6.SEQ_MODE=4'b1000;
    defparam shift_srl_144_6_LC_12_18_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_144_6_LC_12_18_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58588),
            .lcout(shift_srl_144Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93016),
            .ce(N__59989),
            .sr(_gnd_net_));
    defparam shift_srl_144_7_LC_12_18_7.C_ON=1'b0;
    defparam shift_srl_144_7_LC_12_18_7.SEQ_MODE=4'b1000;
    defparam shift_srl_144_7_LC_12_18_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_144_7_LC_12_18_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58690),
            .lcout(shift_srl_144Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93016),
            .ce(N__59989),
            .sr(_gnd_net_));
    defparam shift_srl_144_10_LC_12_19_0.C_ON=1'b0;
    defparam shift_srl_144_10_LC_12_19_0.SEQ_MODE=4'b1000;
    defparam shift_srl_144_10_LC_12_19_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_144_10_LC_12_19_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58654),
            .lcout(shift_srl_144Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93029),
            .ce(N__59988),
            .sr(_gnd_net_));
    defparam shift_srl_144_11_LC_12_19_1.C_ON=1'b0;
    defparam shift_srl_144_11_LC_12_19_1.SEQ_MODE=4'b1000;
    defparam shift_srl_144_11_LC_12_19_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_144_11_LC_12_19_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58684),
            .lcout(shift_srl_144Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93029),
            .ce(N__59988),
            .sr(_gnd_net_));
    defparam shift_srl_144_12_LC_12_19_2.C_ON=1'b0;
    defparam shift_srl_144_12_LC_12_19_2.SEQ_MODE=4'b1000;
    defparam shift_srl_144_12_LC_12_19_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_144_12_LC_12_19_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58678),
            .lcout(shift_srl_144Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93029),
            .ce(N__59988),
            .sr(_gnd_net_));
    defparam shift_srl_144_13_LC_12_19_3.C_ON=1'b0;
    defparam shift_srl_144_13_LC_12_19_3.SEQ_MODE=4'b1000;
    defparam shift_srl_144_13_LC_12_19_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_144_13_LC_12_19_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58672),
            .lcout(shift_srl_144Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93029),
            .ce(N__59988),
            .sr(_gnd_net_));
    defparam shift_srl_144_14_LC_12_19_4.C_ON=1'b0;
    defparam shift_srl_144_14_LC_12_19_4.SEQ_MODE=4'b1000;
    defparam shift_srl_144_14_LC_12_19_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_144_14_LC_12_19_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58666),
            .lcout(shift_srl_144Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93029),
            .ce(N__59988),
            .sr(_gnd_net_));
    defparam shift_srl_144_15_LC_12_19_5.C_ON=1'b0;
    defparam shift_srl_144_15_LC_12_19_5.SEQ_MODE=4'b1000;
    defparam shift_srl_144_15_LC_12_19_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_144_15_LC_12_19_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58660),
            .lcout(shift_srl_144Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93029),
            .ce(N__59988),
            .sr(_gnd_net_));
    defparam shift_srl_144_9_LC_12_19_6.C_ON=1'b0;
    defparam shift_srl_144_9_LC_12_19_6.SEQ_MODE=4'b1000;
    defparam shift_srl_144_9_LC_12_19_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_144_9_LC_12_19_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58642),
            .lcout(shift_srl_144Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93029),
            .ce(N__59988),
            .sr(_gnd_net_));
    defparam shift_srl_144_8_LC_12_19_7.C_ON=1'b0;
    defparam shift_srl_144_8_LC_12_19_7.SEQ_MODE=4'b1000;
    defparam shift_srl_144_8_LC_12_19_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_144_8_LC_12_19_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58648),
            .lcout(shift_srl_144Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93029),
            .ce(N__59988),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIG00FT_15_LC_12_20_0.C_ON=1'b0;
    defparam shift_srl_0_RNIG00FT_15_LC_12_20_0.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIG00FT_15_LC_12_20_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNIG00FT_15_LC_12_20_0 (
            .in0(N__79321),
            .in1(N__65882),
            .in2(N__90532),
            .in3(N__64986),
            .lcout(clk_en_117),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_116_RNI3CPB1_15_LC_12_20_1.C_ON=1'b0;
    defparam shift_srl_116_RNI3CPB1_15_LC_12_20_1.SEQ_MODE=4'b0000;
    defparam shift_srl_116_RNI3CPB1_15_LC_12_20_1.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_116_RNI3CPB1_15_LC_12_20_1 (
            .in0(N__62585),
            .in1(N__58809),
            .in2(_gnd_net_),
            .in3(N__63832),
            .lcout(rco_int_0_a2_1_a2_0_0_116),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_116_RNI5Q4G4_15_LC_12_20_2.C_ON=1'b0;
    defparam shift_srl_116_RNI5Q4G4_15_LC_12_20_2.SEQ_MODE=4'b0000;
    defparam shift_srl_116_RNI5Q4G4_15_LC_12_20_2.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_116_RNI5Q4G4_15_LC_12_20_2 (
            .in0(N__63833),
            .in1(N__62586),
            .in2(N__58813),
            .in3(N__64985),
            .lcout(),
            .ltout(rco_int_0_a2_1_a2_1_118_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_118_RNIUO9UT_15_LC_12_20_3.C_ON=1'b0;
    defparam shift_srl_118_RNIUO9UT_15_LC_12_20_3.SEQ_MODE=4'b0000;
    defparam shift_srl_118_RNIUO9UT_15_LC_12_20_3.LUT_INIT=16'b0000100000000000;
    LogicCell40 shift_srl_118_RNIUO9UT_15_LC_12_20_3 (
            .in0(N__60315),
            .in1(N__66392),
            .in2(N__58744),
            .in3(N__79320),
            .lcout(rco_c_118),
            .ltout(rco_c_118_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNITLDGU_15_LC_12_20_4.C_ON=1'b0;
    defparam shift_srl_0_RNITLDGU_15_LC_12_20_4.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNITLDGU_15_LC_12_20_4.LUT_INIT=16'b1010000000000000;
    LogicCell40 shift_srl_0_RNITLDGU_15_LC_12_20_4 (
            .in0(N__90439),
            .in1(_gnd_net_),
            .in2(N__58741),
            .in3(N__65551),
            .lcout(clk_en_121),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_118_RNIEU805_15_LC_12_20_5.C_ON=1'b0;
    defparam shift_srl_118_RNIEU805_15_LC_12_20_5.SEQ_MODE=4'b0000;
    defparam shift_srl_118_RNIEU805_15_LC_12_20_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_118_RNIEU805_15_LC_12_20_5 (
            .in0(N__64984),
            .in1(N__60314),
            .in2(N__65890),
            .in3(N__66391),
            .lcout(rco_int_0_a2_1_a2_1_123),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIT8DIV_15_LC_12_20_6.C_ON=1'b0;
    defparam shift_srl_0_RNIT8DIV_15_LC_12_20_6.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIT8DIV_15_LC_12_20_6.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNIT8DIV_15_LC_12_20_6 (
            .in0(N__65552),
            .in1(N__65370),
            .in2(N__90533),
            .in3(N__65947),
            .lcout(clk_en_124),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_121_RNIS2INU_15_LC_12_20_7.C_ON=1'b0;
    defparam shift_srl_121_RNIS2INU_15_LC_12_20_7.SEQ_MODE=4'b0000;
    defparam shift_srl_121_RNIS2INU_15_LC_12_20_7.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_121_RNIS2INU_15_LC_12_20_7 (
            .in0(N__65948),
            .in1(N__65553),
            .in2(N__78472),
            .in3(N__90443),
            .lcout(clk_en_122),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_118_RNI2AJFU_15_LC_12_21_0.C_ON=1'b0;
    defparam shift_srl_118_RNI2AJFU_15_LC_12_21_0.SEQ_MODE=4'b0000;
    defparam shift_srl_118_RNI2AJFU_15_LC_12_21_0.LUT_INIT=16'b0010000000000000;
    LogicCell40 shift_srl_118_RNI2AJFU_15_LC_12_21_0 (
            .in0(N__66415),
            .in1(N__60649),
            .in2(N__60334),
            .in3(N__79415),
            .lcout(rco_c_120),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_117_15_LC_12_21_2.C_ON=1'b0;
    defparam shift_srl_117_15_LC_12_21_2.SEQ_MODE=4'b1000;
    defparam shift_srl_117_15_LC_12_21_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_117_15_LC_12_21_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58861),
            .lcout(shift_srl_117Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93057),
            .ce(N__65060),
            .sr(_gnd_net_));
    defparam shift_srl_117_14_LC_12_21_3.C_ON=1'b0;
    defparam shift_srl_117_14_LC_12_21_3.SEQ_MODE=4'b1000;
    defparam shift_srl_117_14_LC_12_21_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_117_14_LC_12_21_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58855),
            .lcout(shift_srl_117Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93057),
            .ce(N__65060),
            .sr(_gnd_net_));
    defparam shift_srl_117_13_LC_12_21_4.C_ON=1'b0;
    defparam shift_srl_117_13_LC_12_21_4.SEQ_MODE=4'b1000;
    defparam shift_srl_117_13_LC_12_21_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_117_13_LC_12_21_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58849),
            .lcout(shift_srl_117Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93057),
            .ce(N__65060),
            .sr(_gnd_net_));
    defparam shift_srl_117_12_LC_12_21_5.C_ON=1'b0;
    defparam shift_srl_117_12_LC_12_21_5.SEQ_MODE=4'b1000;
    defparam shift_srl_117_12_LC_12_21_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_117_12_LC_12_21_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58843),
            .lcout(shift_srl_117Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93057),
            .ce(N__65060),
            .sr(_gnd_net_));
    defparam shift_srl_117_11_LC_12_21_6.C_ON=1'b0;
    defparam shift_srl_117_11_LC_12_21_6.SEQ_MODE=4'b1000;
    defparam shift_srl_117_11_LC_12_21_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_117_11_LC_12_21_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58837),
            .lcout(shift_srl_117Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93057),
            .ce(N__65060),
            .sr(_gnd_net_));
    defparam shift_srl_117_10_LC_12_21_7.C_ON=1'b0;
    defparam shift_srl_117_10_LC_12_21_7.SEQ_MODE=4'b1000;
    defparam shift_srl_117_10_LC_12_21_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_117_10_LC_12_21_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65083),
            .lcout(shift_srl_117Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93057),
            .ce(N__65060),
            .sr(_gnd_net_));
    defparam shift_srl_114_10_LC_12_22_0.C_ON=1'b0;
    defparam shift_srl_114_10_LC_12_22_0.SEQ_MODE=4'b1000;
    defparam shift_srl_114_10_LC_12_22_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_114_10_LC_12_22_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58939),
            .lcout(shift_srl_114Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93073),
            .ce(N__60382),
            .sr(_gnd_net_));
    defparam shift_srl_114_11_LC_12_22_1.C_ON=1'b0;
    defparam shift_srl_114_11_LC_12_22_1.SEQ_MODE=4'b1000;
    defparam shift_srl_114_11_LC_12_22_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_114_11_LC_12_22_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58831),
            .lcout(shift_srl_114Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93073),
            .ce(N__60382),
            .sr(_gnd_net_));
    defparam shift_srl_114_12_LC_12_22_2.C_ON=1'b0;
    defparam shift_srl_114_12_LC_12_22_2.SEQ_MODE=4'b1000;
    defparam shift_srl_114_12_LC_12_22_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_114_12_LC_12_22_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58825),
            .lcout(shift_srl_114Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93073),
            .ce(N__60382),
            .sr(_gnd_net_));
    defparam shift_srl_114_13_LC_12_22_3.C_ON=1'b0;
    defparam shift_srl_114_13_LC_12_22_3.SEQ_MODE=4'b1000;
    defparam shift_srl_114_13_LC_12_22_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_114_13_LC_12_22_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58819),
            .lcout(shift_srl_114Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93073),
            .ce(N__60382),
            .sr(_gnd_net_));
    defparam shift_srl_114_14_LC_12_22_4.C_ON=1'b0;
    defparam shift_srl_114_14_LC_12_22_4.SEQ_MODE=4'b1000;
    defparam shift_srl_114_14_LC_12_22_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_114_14_LC_12_22_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58951),
            .lcout(shift_srl_114Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93073),
            .ce(N__60382),
            .sr(_gnd_net_));
    defparam shift_srl_114_15_LC_12_22_5.C_ON=1'b0;
    defparam shift_srl_114_15_LC_12_22_5.SEQ_MODE=4'b1000;
    defparam shift_srl_114_15_LC_12_22_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_114_15_LC_12_22_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58945),
            .lcout(shift_srl_114Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93073),
            .ce(N__60382),
            .sr(_gnd_net_));
    defparam shift_srl_114_9_LC_12_22_6.C_ON=1'b0;
    defparam shift_srl_114_9_LC_12_22_6.SEQ_MODE=4'b1000;
    defparam shift_srl_114_9_LC_12_22_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_114_9_LC_12_22_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58933),
            .lcout(shift_srl_114Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93073),
            .ce(N__60382),
            .sr(_gnd_net_));
    defparam shift_srl_114_8_LC_12_22_7.C_ON=1'b0;
    defparam shift_srl_114_8_LC_12_22_7.SEQ_MODE=4'b1000;
    defparam shift_srl_114_8_LC_12_22_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_114_8_LC_12_22_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58987),
            .lcout(shift_srl_114Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93073),
            .ce(N__60382),
            .sr(_gnd_net_));
    defparam shift_srl_114_0_LC_12_23_0.C_ON=1'b0;
    defparam shift_srl_114_0_LC_12_23_0.SEQ_MODE=4'b1000;
    defparam shift_srl_114_0_LC_12_23_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_114_0_LC_12_23_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58916),
            .lcout(shift_srl_114Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93088),
            .ce(N__60375),
            .sr(_gnd_net_));
    defparam shift_srl_114_1_LC_12_23_1.C_ON=1'b0;
    defparam shift_srl_114_1_LC_12_23_1.SEQ_MODE=4'b1000;
    defparam shift_srl_114_1_LC_12_23_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_114_1_LC_12_23_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58885),
            .lcout(shift_srl_114Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93088),
            .ce(N__60375),
            .sr(_gnd_net_));
    defparam shift_srl_114_2_LC_12_23_2.C_ON=1'b0;
    defparam shift_srl_114_2_LC_12_23_2.SEQ_MODE=4'b1000;
    defparam shift_srl_114_2_LC_12_23_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_114_2_LC_12_23_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58879),
            .lcout(shift_srl_114Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93088),
            .ce(N__60375),
            .sr(_gnd_net_));
    defparam shift_srl_114_3_LC_12_23_3.C_ON=1'b0;
    defparam shift_srl_114_3_LC_12_23_3.SEQ_MODE=4'b1000;
    defparam shift_srl_114_3_LC_12_23_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_114_3_LC_12_23_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58873),
            .lcout(shift_srl_114Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93088),
            .ce(N__60375),
            .sr(_gnd_net_));
    defparam shift_srl_114_4_LC_12_23_4.C_ON=1'b0;
    defparam shift_srl_114_4_LC_12_23_4.SEQ_MODE=4'b1000;
    defparam shift_srl_114_4_LC_12_23_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_114_4_LC_12_23_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58867),
            .lcout(shift_srl_114Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93088),
            .ce(N__60375),
            .sr(_gnd_net_));
    defparam shift_srl_114_5_LC_12_23_5.C_ON=1'b0;
    defparam shift_srl_114_5_LC_12_23_5.SEQ_MODE=4'b1000;
    defparam shift_srl_114_5_LC_12_23_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_114_5_LC_12_23_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59005),
            .lcout(shift_srl_114Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93088),
            .ce(N__60375),
            .sr(_gnd_net_));
    defparam shift_srl_114_6_LC_12_23_6.C_ON=1'b0;
    defparam shift_srl_114_6_LC_12_23_6.SEQ_MODE=4'b1000;
    defparam shift_srl_114_6_LC_12_23_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_114_6_LC_12_23_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58999),
            .lcout(shift_srl_114Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93088),
            .ce(N__60375),
            .sr(_gnd_net_));
    defparam shift_srl_114_7_LC_12_23_7.C_ON=1'b0;
    defparam shift_srl_114_7_LC_12_23_7.SEQ_MODE=4'b1000;
    defparam shift_srl_114_7_LC_12_23_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_114_7_LC_12_23_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58993),
            .lcout(shift_srl_114Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93088),
            .ce(N__60375),
            .sr(_gnd_net_));
    defparam shift_srl_118_0_LC_12_24_0.C_ON=1'b0;
    defparam shift_srl_118_0_LC_12_24_0.SEQ_MODE=4'b1000;
    defparam shift_srl_118_0_LC_12_24_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_118_0_LC_12_24_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60328),
            .lcout(shift_srl_118Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93103),
            .ce(N__60800),
            .sr(_gnd_net_));
    defparam shift_srl_118_1_LC_12_24_1.C_ON=1'b0;
    defparam shift_srl_118_1_LC_12_24_1.SEQ_MODE=4'b1000;
    defparam shift_srl_118_1_LC_12_24_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_118_1_LC_12_24_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58981),
            .lcout(shift_srl_118Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93103),
            .ce(N__60800),
            .sr(_gnd_net_));
    defparam shift_srl_118_2_LC_12_24_2.C_ON=1'b0;
    defparam shift_srl_118_2_LC_12_24_2.SEQ_MODE=4'b1000;
    defparam shift_srl_118_2_LC_12_24_2.LUT_INIT=16'b1100110011001100;
    LogicCell40 shift_srl_118_2_LC_12_24_2 (
            .in0(_gnd_net_),
            .in1(N__58975),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_118Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93103),
            .ce(N__60800),
            .sr(_gnd_net_));
    defparam shift_srl_118_3_LC_12_24_3.C_ON=1'b0;
    defparam shift_srl_118_3_LC_12_24_3.SEQ_MODE=4'b1000;
    defparam shift_srl_118_3_LC_12_24_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_118_3_LC_12_24_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58969),
            .lcout(shift_srl_118Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93103),
            .ce(N__60800),
            .sr(_gnd_net_));
    defparam shift_srl_118_4_LC_12_24_4.C_ON=1'b0;
    defparam shift_srl_118_4_LC_12_24_4.SEQ_MODE=4'b1000;
    defparam shift_srl_118_4_LC_12_24_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_118_4_LC_12_24_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58963),
            .lcout(shift_srl_118Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93103),
            .ce(N__60800),
            .sr(_gnd_net_));
    defparam shift_srl_118_5_LC_12_24_5.C_ON=1'b0;
    defparam shift_srl_118_5_LC_12_24_5.SEQ_MODE=4'b1000;
    defparam shift_srl_118_5_LC_12_24_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_118_5_LC_12_24_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58957),
            .lcout(shift_srl_118Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93103),
            .ce(N__60800),
            .sr(_gnd_net_));
    defparam shift_srl_118_6_LC_12_24_6.C_ON=1'b0;
    defparam shift_srl_118_6_LC_12_24_6.SEQ_MODE=4'b1000;
    defparam shift_srl_118_6_LC_12_24_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_118_6_LC_12_24_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59065),
            .lcout(shift_srl_118Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93103),
            .ce(N__60800),
            .sr(_gnd_net_));
    defparam shift_srl_118_7_LC_12_24_7.C_ON=1'b0;
    defparam shift_srl_118_7_LC_12_24_7.SEQ_MODE=4'b1000;
    defparam shift_srl_118_7_LC_12_24_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_118_7_LC_12_24_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59059),
            .lcout(shift_srl_118Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93103),
            .ce(N__60800),
            .sr(_gnd_net_));
    defparam shift_srl_100_0_LC_12_25_0.C_ON=1'b0;
    defparam shift_srl_100_0_LC_12_25_0.SEQ_MODE=4'b1000;
    defparam shift_srl_100_0_LC_12_25_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_100_0_LC_12_25_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79689),
            .lcout(shift_srl_100Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93121),
            .ce(N__60890),
            .sr(_gnd_net_));
    defparam shift_srl_100_1_LC_12_25_1.C_ON=1'b0;
    defparam shift_srl_100_1_LC_12_25_1.SEQ_MODE=4'b1000;
    defparam shift_srl_100_1_LC_12_25_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_100_1_LC_12_25_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59041),
            .lcout(shift_srl_100Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93121),
            .ce(N__60890),
            .sr(_gnd_net_));
    defparam shift_srl_100_2_LC_12_25_2.C_ON=1'b0;
    defparam shift_srl_100_2_LC_12_25_2.SEQ_MODE=4'b1000;
    defparam shift_srl_100_2_LC_12_25_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_100_2_LC_12_25_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59035),
            .lcout(shift_srl_100Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93121),
            .ce(N__60890),
            .sr(_gnd_net_));
    defparam shift_srl_100_3_LC_12_25_3.C_ON=1'b0;
    defparam shift_srl_100_3_LC_12_25_3.SEQ_MODE=4'b1000;
    defparam shift_srl_100_3_LC_12_25_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_100_3_LC_12_25_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59029),
            .lcout(shift_srl_100Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93121),
            .ce(N__60890),
            .sr(_gnd_net_));
    defparam shift_srl_100_4_LC_12_25_4.C_ON=1'b0;
    defparam shift_srl_100_4_LC_12_25_4.SEQ_MODE=4'b1000;
    defparam shift_srl_100_4_LC_12_25_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_100_4_LC_12_25_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59023),
            .lcout(shift_srl_100Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93121),
            .ce(N__60890),
            .sr(_gnd_net_));
    defparam shift_srl_100_5_LC_12_25_5.C_ON=1'b0;
    defparam shift_srl_100_5_LC_12_25_5.SEQ_MODE=4'b1000;
    defparam shift_srl_100_5_LC_12_25_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_100_5_LC_12_25_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59017),
            .lcout(shift_srl_100Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93121),
            .ce(N__60890),
            .sr(_gnd_net_));
    defparam shift_srl_100_6_LC_12_25_6.C_ON=1'b0;
    defparam shift_srl_100_6_LC_12_25_6.SEQ_MODE=4'b1000;
    defparam shift_srl_100_6_LC_12_25_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_100_6_LC_12_25_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59011),
            .lcout(shift_srl_100Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93121),
            .ce(N__60890),
            .sr(_gnd_net_));
    defparam shift_srl_104_10_LC_12_26_0.C_ON=1'b0;
    defparam shift_srl_104_10_LC_12_26_0.SEQ_MODE=4'b1000;
    defparam shift_srl_104_10_LC_12_26_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_104_10_LC_12_26_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59083),
            .lcout(shift_srl_104Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93140),
            .ce(N__59308),
            .sr(_gnd_net_));
    defparam shift_srl_104_11_LC_12_26_1.C_ON=1'b0;
    defparam shift_srl_104_11_LC_12_26_1.SEQ_MODE=4'b1000;
    defparam shift_srl_104_11_LC_12_26_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_104_11_LC_12_26_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59113),
            .lcout(shift_srl_104Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93140),
            .ce(N__59308),
            .sr(_gnd_net_));
    defparam shift_srl_104_12_LC_12_26_2.C_ON=1'b0;
    defparam shift_srl_104_12_LC_12_26_2.SEQ_MODE=4'b1000;
    defparam shift_srl_104_12_LC_12_26_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_104_12_LC_12_26_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59107),
            .lcout(shift_srl_104Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93140),
            .ce(N__59308),
            .sr(_gnd_net_));
    defparam shift_srl_104_13_LC_12_26_3.C_ON=1'b0;
    defparam shift_srl_104_13_LC_12_26_3.SEQ_MODE=4'b1000;
    defparam shift_srl_104_13_LC_12_26_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_104_13_LC_12_26_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59101),
            .lcout(shift_srl_104Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93140),
            .ce(N__59308),
            .sr(_gnd_net_));
    defparam shift_srl_104_14_LC_12_26_4.C_ON=1'b0;
    defparam shift_srl_104_14_LC_12_26_4.SEQ_MODE=4'b1000;
    defparam shift_srl_104_14_LC_12_26_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_104_14_LC_12_26_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59095),
            .lcout(shift_srl_104Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93140),
            .ce(N__59308),
            .sr(_gnd_net_));
    defparam shift_srl_104_15_LC_12_26_5.C_ON=1'b0;
    defparam shift_srl_104_15_LC_12_26_5.SEQ_MODE=4'b1000;
    defparam shift_srl_104_15_LC_12_26_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_104_15_LC_12_26_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59089),
            .lcout(shift_srl_104Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93140),
            .ce(N__59308),
            .sr(_gnd_net_));
    defparam shift_srl_104_9_LC_12_26_6.C_ON=1'b0;
    defparam shift_srl_104_9_LC_12_26_6.SEQ_MODE=4'b1000;
    defparam shift_srl_104_9_LC_12_26_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_104_9_LC_12_26_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59071),
            .lcout(shift_srl_104Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93140),
            .ce(N__59308),
            .sr(_gnd_net_));
    defparam shift_srl_104_8_LC_12_26_7.C_ON=1'b0;
    defparam shift_srl_104_8_LC_12_26_7.SEQ_MODE=4'b1000;
    defparam shift_srl_104_8_LC_12_26_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_104_8_LC_12_26_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59077),
            .lcout(shift_srl_104Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93140),
            .ce(N__59308),
            .sr(_gnd_net_));
    defparam shift_srl_102_RNI73HLP_15_LC_12_27_0.C_ON=1'b0;
    defparam shift_srl_102_RNI73HLP_15_LC_12_27_0.SEQ_MODE=4'b0000;
    defparam shift_srl_102_RNI73HLP_15_LC_12_27_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_102_RNI73HLP_15_LC_12_27_0 (
            .in0(N__79530),
            .in1(N__62698),
            .in2(N__79688),
            .in3(N__60961),
            .lcout(rco_c_102),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_102_RNIN8GN_15_LC_12_27_1.C_ON=1'b0;
    defparam shift_srl_102_RNIN8GN_15_LC_12_27_1.SEQ_MODE=4'b0000;
    defparam shift_srl_102_RNIN8GN_15_LC_12_27_1.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_102_RNIN8GN_15_LC_12_27_1 (
            .in0(N__60960),
            .in1(N__62702),
            .in2(_gnd_net_),
            .in3(N__79678),
            .lcout(),
            .ltout(shift_srl_102_RNIN8GNZ0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_103_RNI1Q71Q_15_LC_12_27_2.C_ON=1'b0;
    defparam shift_srl_103_RNI1Q71Q_15_LC_12_27_2.SEQ_MODE=4'b0000;
    defparam shift_srl_103_RNI1Q71Q_15_LC_12_27_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_103_RNI1Q71Q_15_LC_12_27_2 (
            .in0(N__79529),
            .in1(N__90565),
            .in2(N__59311),
            .in3(N__61093),
            .lcout(clk_en_104),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_101_15_LC_12_27_3.C_ON=1'b0;
    defparam shift_srl_101_15_LC_12_27_3.SEQ_MODE=4'b1000;
    defparam shift_srl_101_15_LC_12_27_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_101_15_LC_12_27_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59296),
            .lcout(shift_srl_101Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93159),
            .ce(N__59194),
            .sr(_gnd_net_));
    defparam shift_srl_102_RNIUJTJ_15_LC_12_27_4.C_ON=1'b0;
    defparam shift_srl_102_RNIUJTJ_15_LC_12_27_4.SEQ_MODE=4'b0000;
    defparam shift_srl_102_RNIUJTJ_15_LC_12_27_4.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_102_RNIUJTJ_15_LC_12_27_4 (
            .in0(N__59280),
            .in1(N__62696),
            .in2(N__59250),
            .in3(N__60959),
            .lcout(rco_int_0_a2_0_a2_s_0_sx_110),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_100_RNI755DP_15_LC_12_27_5.C_ON=1'b0;
    defparam shift_srl_100_RNI755DP_15_LC_12_27_5.SEQ_MODE=4'b0000;
    defparam shift_srl_100_RNI755DP_15_LC_12_27_5.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_100_RNI755DP_15_LC_12_27_5 (
            .in0(N__90563),
            .in1(N__79677),
            .in2(_gnd_net_),
            .in3(N__79527),
            .lcout(clk_en_101),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_102_RNIIKAO_15_LC_12_27_6.C_ON=1'b0;
    defparam shift_srl_102_RNIIKAO_15_LC_12_27_6.SEQ_MODE=4'b0000;
    defparam shift_srl_102_RNIIKAO_15_LC_12_27_6.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_102_RNIIKAO_15_LC_12_27_6 (
            .in0(N__79676),
            .in1(N__62697),
            .in2(N__60983),
            .in3(N__90564),
            .lcout(),
            .ltout(clk_en_0_a3_0_a2_sx_103_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_102_RNI2FBMP_15_LC_12_27_7.C_ON=1'b0;
    defparam shift_srl_102_RNI2FBMP_15_LC_12_27_7.SEQ_MODE=4'b0000;
    defparam shift_srl_102_RNI2FBMP_15_LC_12_27_7.LUT_INIT=16'b0000111100000000;
    LogicCell40 shift_srl_102_RNI2FBMP_15_LC_12_27_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__59170),
            .in3(N__79528),
            .lcout(clk_en_103),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_103_LC_12_28_0.C_ON=1'b0;
    defparam rco_obuf_RNO_103_LC_12_28_0.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_103_LC_12_28_0.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_103_LC_12_28_0 (
            .in0(N__61095),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59151),
            .lcout(rco_c_103),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_103_0_LC_12_28_1.C_ON=1'b0;
    defparam shift_srl_103_0_LC_12_28_1.SEQ_MODE=4'b1000;
    defparam shift_srl_103_0_LC_12_28_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_103_0_LC_12_28_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61094),
            .lcout(shift_srl_103Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93178),
            .ce(N__61046),
            .sr(_gnd_net_));
    defparam shift_srl_103_1_LC_12_28_2.C_ON=1'b0;
    defparam shift_srl_103_1_LC_12_28_2.SEQ_MODE=4'b1000;
    defparam shift_srl_103_1_LC_12_28_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_103_1_LC_12_28_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59119),
            .lcout(shift_srl_103Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93178),
            .ce(N__61046),
            .sr(_gnd_net_));
    defparam shift_srl_103_2_LC_12_28_3.C_ON=1'b0;
    defparam shift_srl_103_2_LC_12_28_3.SEQ_MODE=4'b1000;
    defparam shift_srl_103_2_LC_12_28_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_103_2_LC_12_28_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59371),
            .lcout(shift_srl_103Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93178),
            .ce(N__61046),
            .sr(_gnd_net_));
    defparam shift_srl_103_3_LC_12_28_4.C_ON=1'b0;
    defparam shift_srl_103_3_LC_12_28_4.SEQ_MODE=4'b1000;
    defparam shift_srl_103_3_LC_12_28_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_103_3_LC_12_28_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59365),
            .lcout(shift_srl_103Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93178),
            .ce(N__61046),
            .sr(_gnd_net_));
    defparam shift_srl_103_4_LC_12_28_5.C_ON=1'b0;
    defparam shift_srl_103_4_LC_12_28_5.SEQ_MODE=4'b1000;
    defparam shift_srl_103_4_LC_12_28_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_103_4_LC_12_28_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59359),
            .lcout(shift_srl_103Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93178),
            .ce(N__61046),
            .sr(_gnd_net_));
    defparam shift_srl_103_5_LC_12_28_6.C_ON=1'b0;
    defparam shift_srl_103_5_LC_12_28_6.SEQ_MODE=4'b1000;
    defparam shift_srl_103_5_LC_12_28_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_103_5_LC_12_28_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59353),
            .lcout(shift_srl_103Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93178),
            .ce(N__61046),
            .sr(_gnd_net_));
    defparam shift_srl_103_6_LC_12_28_7.C_ON=1'b0;
    defparam shift_srl_103_6_LC_12_28_7.SEQ_MODE=4'b1000;
    defparam shift_srl_103_6_LC_12_28_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_103_6_LC_12_28_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59347),
            .lcout(shift_srl_103Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93178),
            .ce(N__61046),
            .sr(_gnd_net_));
    defparam shift_srl_100_10_LC_12_29_0.C_ON=1'b0;
    defparam shift_srl_100_10_LC_12_29_0.SEQ_MODE=4'b1000;
    defparam shift_srl_100_10_LC_12_29_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_100_10_LC_12_29_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59341),
            .lcout(shift_srl_100Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93200),
            .ce(N__60895),
            .sr(_gnd_net_));
    defparam shift_srl_100_9_LC_12_29_1.C_ON=1'b0;
    defparam shift_srl_100_9_LC_12_29_1.SEQ_MODE=4'b1000;
    defparam shift_srl_100_9_LC_12_29_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_100_9_LC_12_29_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59335),
            .lcout(shift_srl_100Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93200),
            .ce(N__60895),
            .sr(_gnd_net_));
    defparam shift_srl_100_8_LC_12_29_2.C_ON=1'b0;
    defparam shift_srl_100_8_LC_12_29_2.SEQ_MODE=4'b1000;
    defparam shift_srl_100_8_LC_12_29_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_100_8_LC_12_29_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59317),
            .lcout(shift_srl_100Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93200),
            .ce(N__60895),
            .sr(_gnd_net_));
    defparam shift_srl_100_7_LC_12_29_6.C_ON=1'b0;
    defparam shift_srl_100_7_LC_12_29_6.SEQ_MODE=4'b1000;
    defparam shift_srl_100_7_LC_12_29_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_100_7_LC_12_29_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59329),
            .lcout(shift_srl_100Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93200),
            .ce(N__60895),
            .sr(_gnd_net_));
    defparam shift_srl_103_7_LC_12_30_0.C_ON=1'b0;
    defparam shift_srl_103_7_LC_12_30_0.SEQ_MODE=4'b1000;
    defparam shift_srl_103_7_LC_12_30_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_103_7_LC_12_30_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59422),
            .lcout(shift_srl_103Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93221),
            .ce(N__61047),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_165_LC_13_4_3.C_ON=1'b0;
    defparam rco_obuf_RNO_165_LC_13_4_3.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_165_LC_13_4_3.LUT_INIT=16'b1000100000000000;
    LogicCell40 rco_obuf_RNO_165_LC_13_4_3 (
            .in0(N__87724),
            .in1(N__82428),
            .in2(_gnd_net_),
            .in3(N__83983),
            .lcout(rco_c_165),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_90_10_LC_13_5_0.C_ON=1'b0;
    defparam shift_srl_90_10_LC_13_5_0.SEQ_MODE=4'b1000;
    defparam shift_srl_90_10_LC_13_5_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_90_10_LC_13_5_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59401),
            .lcout(shift_srl_90Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93222),
            .ce(N__61228),
            .sr(_gnd_net_));
    defparam shift_srl_90_9_LC_13_5_1.C_ON=1'b0;
    defparam shift_srl_90_9_LC_13_5_1.SEQ_MODE=4'b1000;
    defparam shift_srl_90_9_LC_13_5_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_90_9_LC_13_5_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59395),
            .lcout(shift_srl_90Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93222),
            .ce(N__61228),
            .sr(_gnd_net_));
    defparam shift_srl_90_8_LC_13_5_2.C_ON=1'b0;
    defparam shift_srl_90_8_LC_13_5_2.SEQ_MODE=4'b1000;
    defparam shift_srl_90_8_LC_13_5_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_90_8_LC_13_5_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59383),
            .lcout(shift_srl_90Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93222),
            .ce(N__61228),
            .sr(_gnd_net_));
    defparam shift_srl_90_6_LC_13_5_5.C_ON=1'b0;
    defparam shift_srl_90_6_LC_13_5_5.SEQ_MODE=4'b1000;
    defparam shift_srl_90_6_LC_13_5_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_90_6_LC_13_5_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61156),
            .lcout(shift_srl_90Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93222),
            .ce(N__61228),
            .sr(_gnd_net_));
    defparam shift_srl_90_7_LC_13_5_6.C_ON=1'b0;
    defparam shift_srl_90_7_LC_13_5_6.SEQ_MODE=4'b1000;
    defparam shift_srl_90_7_LC_13_5_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_90_7_LC_13_5_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59389),
            .lcout(shift_srl_90Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93222),
            .ce(N__61228),
            .sr(_gnd_net_));
    defparam shift_srl_91_10_LC_13_6_0.C_ON=1'b0;
    defparam shift_srl_91_10_LC_13_6_0.SEQ_MODE=4'b1000;
    defparam shift_srl_91_10_LC_13_6_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_91_10_LC_13_6_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59452),
            .lcout(shift_srl_91Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93202),
            .ce(N__61146),
            .sr(_gnd_net_));
    defparam shift_srl_91_11_LC_13_6_1.C_ON=1'b0;
    defparam shift_srl_91_11_LC_13_6_1.SEQ_MODE=4'b1000;
    defparam shift_srl_91_11_LC_13_6_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_91_11_LC_13_6_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59377),
            .lcout(shift_srl_91Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93202),
            .ce(N__61146),
            .sr(_gnd_net_));
    defparam shift_srl_91_12_LC_13_6_2.C_ON=1'b0;
    defparam shift_srl_91_12_LC_13_6_2.SEQ_MODE=4'b1000;
    defparam shift_srl_91_12_LC_13_6_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_91_12_LC_13_6_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59476),
            .lcout(shift_srl_91Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93202),
            .ce(N__61146),
            .sr(_gnd_net_));
    defparam shift_srl_91_13_LC_13_6_3.C_ON=1'b0;
    defparam shift_srl_91_13_LC_13_6_3.SEQ_MODE=4'b1000;
    defparam shift_srl_91_13_LC_13_6_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_91_13_LC_13_6_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59470),
            .lcout(shift_srl_91Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93202),
            .ce(N__61146),
            .sr(_gnd_net_));
    defparam shift_srl_91_14_LC_13_6_4.C_ON=1'b0;
    defparam shift_srl_91_14_LC_13_6_4.SEQ_MODE=4'b1000;
    defparam shift_srl_91_14_LC_13_6_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_91_14_LC_13_6_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59464),
            .lcout(shift_srl_91Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93202),
            .ce(N__61146),
            .sr(_gnd_net_));
    defparam shift_srl_91_15_LC_13_6_5.C_ON=1'b0;
    defparam shift_srl_91_15_LC_13_6_5.SEQ_MODE=4'b1000;
    defparam shift_srl_91_15_LC_13_6_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_91_15_LC_13_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59458),
            .lcout(shift_srl_91Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93202),
            .ce(N__61146),
            .sr(_gnd_net_));
    defparam shift_srl_91_9_LC_13_6_6.C_ON=1'b0;
    defparam shift_srl_91_9_LC_13_6_6.SEQ_MODE=4'b1000;
    defparam shift_srl_91_9_LC_13_6_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_91_9_LC_13_6_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59446),
            .lcout(shift_srl_91Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93202),
            .ce(N__61146),
            .sr(_gnd_net_));
    defparam shift_srl_91_8_LC_13_6_7.C_ON=1'b0;
    defparam shift_srl_91_8_LC_13_6_7.SEQ_MODE=4'b1000;
    defparam shift_srl_91_8_LC_13_6_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_91_8_LC_13_6_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59506),
            .lcout(shift_srl_91Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93202),
            .ce(N__61146),
            .sr(_gnd_net_));
    defparam shift_srl_91_0_LC_13_7_0.C_ON=1'b0;
    defparam shift_srl_91_0_LC_13_7_0.SEQ_MODE=4'b1000;
    defparam shift_srl_91_0_LC_13_7_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_91_0_LC_13_7_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66938),
            .lcout(shift_srl_91Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93180),
            .ce(N__61150),
            .sr(_gnd_net_));
    defparam shift_srl_91_1_LC_13_7_1.C_ON=1'b0;
    defparam shift_srl_91_1_LC_13_7_1.SEQ_MODE=4'b1000;
    defparam shift_srl_91_1_LC_13_7_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_91_1_LC_13_7_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59440),
            .lcout(shift_srl_91Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93180),
            .ce(N__61150),
            .sr(_gnd_net_));
    defparam shift_srl_91_2_LC_13_7_2.C_ON=1'b0;
    defparam shift_srl_91_2_LC_13_7_2.SEQ_MODE=4'b1000;
    defparam shift_srl_91_2_LC_13_7_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_91_2_LC_13_7_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59434),
            .lcout(shift_srl_91Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93180),
            .ce(N__61150),
            .sr(_gnd_net_));
    defparam shift_srl_91_3_LC_13_7_3.C_ON=1'b0;
    defparam shift_srl_91_3_LC_13_7_3.SEQ_MODE=4'b1000;
    defparam shift_srl_91_3_LC_13_7_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_91_3_LC_13_7_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59428),
            .lcout(shift_srl_91Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93180),
            .ce(N__61150),
            .sr(_gnd_net_));
    defparam shift_srl_91_4_LC_13_7_4.C_ON=1'b0;
    defparam shift_srl_91_4_LC_13_7_4.SEQ_MODE=4'b1000;
    defparam shift_srl_91_4_LC_13_7_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_91_4_LC_13_7_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59530),
            .lcout(shift_srl_91Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93180),
            .ce(N__61150),
            .sr(_gnd_net_));
    defparam shift_srl_91_5_LC_13_7_5.C_ON=1'b0;
    defparam shift_srl_91_5_LC_13_7_5.SEQ_MODE=4'b1000;
    defparam shift_srl_91_5_LC_13_7_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_91_5_LC_13_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59524),
            .lcout(shift_srl_91Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93180),
            .ce(N__61150),
            .sr(_gnd_net_));
    defparam shift_srl_91_6_LC_13_7_6.C_ON=1'b0;
    defparam shift_srl_91_6_LC_13_7_6.SEQ_MODE=4'b1000;
    defparam shift_srl_91_6_LC_13_7_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_91_6_LC_13_7_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59518),
            .lcout(shift_srl_91Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93180),
            .ce(N__61150),
            .sr(_gnd_net_));
    defparam shift_srl_91_7_LC_13_7_7.C_ON=1'b0;
    defparam shift_srl_91_7_LC_13_7_7.SEQ_MODE=4'b1000;
    defparam shift_srl_91_7_LC_13_7_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_91_7_LC_13_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59512),
            .lcout(shift_srl_91Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93180),
            .ce(N__61150),
            .sr(_gnd_net_));
    defparam shift_srl_25_7_LC_13_9_1.C_ON=1'b0;
    defparam shift_srl_25_7_LC_13_9_1.SEQ_MODE=4'b1000;
    defparam shift_srl_25_7_LC_13_9_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_25_7_LC_13_9_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59488),
            .lcout(shift_srl_25Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93143),
            .ce(N__59581),
            .sr(_gnd_net_));
    defparam shift_srl_25_5_LC_13_9_2.C_ON=1'b0;
    defparam shift_srl_25_5_LC_13_9_2.SEQ_MODE=4'b1000;
    defparam shift_srl_25_5_LC_13_9_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_25_5_LC_13_9_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59500),
            .lcout(shift_srl_25Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93143),
            .ce(N__59581),
            .sr(_gnd_net_));
    defparam shift_srl_25_6_LC_13_9_4.C_ON=1'b0;
    defparam shift_srl_25_6_LC_13_9_4.SEQ_MODE=4'b1000;
    defparam shift_srl_25_6_LC_13_9_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_25_6_LC_13_9_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59494),
            .lcout(shift_srl_25Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93143),
            .ce(N__59581),
            .sr(_gnd_net_));
    defparam shift_srl_25_10_LC_13_10_0.C_ON=1'b0;
    defparam shift_srl_25_10_LC_13_10_0.SEQ_MODE=4'b1000;
    defparam shift_srl_25_10_LC_13_10_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_25_10_LC_13_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59599),
            .lcout(shift_srl_25Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93123),
            .ce(N__59574),
            .sr(_gnd_net_));
    defparam shift_srl_25_11_LC_13_10_1.C_ON=1'b0;
    defparam shift_srl_25_11_LC_13_10_1.SEQ_MODE=4'b1000;
    defparam shift_srl_25_11_LC_13_10_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_25_11_LC_13_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59482),
            .lcout(shift_srl_25Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93123),
            .ce(N__59574),
            .sr(_gnd_net_));
    defparam shift_srl_25_12_LC_13_10_2.C_ON=1'b0;
    defparam shift_srl_25_12_LC_13_10_2.SEQ_MODE=4'b1000;
    defparam shift_srl_25_12_LC_13_10_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_25_12_LC_13_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59623),
            .lcout(shift_srl_25Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93123),
            .ce(N__59574),
            .sr(_gnd_net_));
    defparam shift_srl_25_13_LC_13_10_3.C_ON=1'b0;
    defparam shift_srl_25_13_LC_13_10_3.SEQ_MODE=4'b1000;
    defparam shift_srl_25_13_LC_13_10_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_25_13_LC_13_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59617),
            .lcout(shift_srl_25Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93123),
            .ce(N__59574),
            .sr(_gnd_net_));
    defparam shift_srl_25_14_LC_13_10_4.C_ON=1'b0;
    defparam shift_srl_25_14_LC_13_10_4.SEQ_MODE=4'b1000;
    defparam shift_srl_25_14_LC_13_10_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_25_14_LC_13_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59611),
            .lcout(shift_srl_25Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93123),
            .ce(N__59574),
            .sr(_gnd_net_));
    defparam shift_srl_25_15_LC_13_10_5.C_ON=1'b0;
    defparam shift_srl_25_15_LC_13_10_5.SEQ_MODE=4'b1000;
    defparam shift_srl_25_15_LC_13_10_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_25_15_LC_13_10_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59605),
            .lcout(shift_srl_25Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93123),
            .ce(N__59574),
            .sr(_gnd_net_));
    defparam shift_srl_25_9_LC_13_10_6.C_ON=1'b0;
    defparam shift_srl_25_9_LC_13_10_6.SEQ_MODE=4'b1000;
    defparam shift_srl_25_9_LC_13_10_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_25_9_LC_13_10_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59587),
            .lcout(shift_srl_25Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93123),
            .ce(N__59574),
            .sr(_gnd_net_));
    defparam shift_srl_25_8_LC_13_10_7.C_ON=1'b0;
    defparam shift_srl_25_8_LC_13_10_7.SEQ_MODE=4'b1000;
    defparam shift_srl_25_8_LC_13_10_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_25_8_LC_13_10_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59593),
            .lcout(shift_srl_25Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93123),
            .ce(N__59574),
            .sr(_gnd_net_));
    defparam shift_srl_89_0_LC_13_11_0.C_ON=1'b0;
    defparam shift_srl_89_0_LC_13_11_0.SEQ_MODE=4'b1000;
    defparam shift_srl_89_0_LC_13_11_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_89_0_LC_13_11_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67011),
            .lcout(shift_srl_89Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93104),
            .ce(N__61429),
            .sr(_gnd_net_));
    defparam shift_srl_89_1_LC_13_11_1.C_ON=1'b0;
    defparam shift_srl_89_1_LC_13_11_1.SEQ_MODE=4'b1000;
    defparam shift_srl_89_1_LC_13_11_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_89_1_LC_13_11_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59542),
            .lcout(shift_srl_89Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93104),
            .ce(N__61429),
            .sr(_gnd_net_));
    defparam shift_srl_89_2_LC_13_11_2.C_ON=1'b0;
    defparam shift_srl_89_2_LC_13_11_2.SEQ_MODE=4'b1000;
    defparam shift_srl_89_2_LC_13_11_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_89_2_LC_13_11_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59536),
            .lcout(shift_srl_89Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93104),
            .ce(N__61429),
            .sr(_gnd_net_));
    defparam shift_srl_89_3_LC_13_11_3.C_ON=1'b0;
    defparam shift_srl_89_3_LC_13_11_3.SEQ_MODE=4'b1000;
    defparam shift_srl_89_3_LC_13_11_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_89_3_LC_13_11_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59671),
            .lcout(shift_srl_89Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93104),
            .ce(N__61429),
            .sr(_gnd_net_));
    defparam shift_srl_89_4_LC_13_11_4.C_ON=1'b0;
    defparam shift_srl_89_4_LC_13_11_4.SEQ_MODE=4'b1000;
    defparam shift_srl_89_4_LC_13_11_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_89_4_LC_13_11_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59665),
            .lcout(shift_srl_89Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93104),
            .ce(N__61429),
            .sr(_gnd_net_));
    defparam shift_srl_89_5_LC_13_11_5.C_ON=1'b0;
    defparam shift_srl_89_5_LC_13_11_5.SEQ_MODE=4'b1000;
    defparam shift_srl_89_5_LC_13_11_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_89_5_LC_13_11_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59659),
            .lcout(shift_srl_89Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93104),
            .ce(N__61429),
            .sr(_gnd_net_));
    defparam shift_srl_89_6_LC_13_11_6.C_ON=1'b0;
    defparam shift_srl_89_6_LC_13_11_6.SEQ_MODE=4'b1000;
    defparam shift_srl_89_6_LC_13_11_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_89_6_LC_13_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59653),
            .lcout(shift_srl_89Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93104),
            .ce(N__61429),
            .sr(_gnd_net_));
    defparam shift_srl_89_7_LC_13_11_7.C_ON=1'b0;
    defparam shift_srl_89_7_LC_13_11_7.SEQ_MODE=4'b1000;
    defparam shift_srl_89_7_LC_13_11_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_89_7_LC_13_11_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59647),
            .lcout(shift_srl_89Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93104),
            .ce(N__61429),
            .sr(_gnd_net_));
    defparam shift_srl_89_10_LC_13_12_0.C_ON=1'b0;
    defparam shift_srl_89_10_LC_13_12_0.SEQ_MODE=4'b1000;
    defparam shift_srl_89_10_LC_13_12_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_89_10_LC_13_12_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59707),
            .lcout(shift_srl_89Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93089),
            .ce(N__61428),
            .sr(_gnd_net_));
    defparam shift_srl_89_11_LC_13_12_1.C_ON=1'b0;
    defparam shift_srl_89_11_LC_13_12_1.SEQ_MODE=4'b1000;
    defparam shift_srl_89_11_LC_13_12_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_89_11_LC_13_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59641),
            .lcout(shift_srl_89Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93089),
            .ce(N__61428),
            .sr(_gnd_net_));
    defparam shift_srl_89_12_LC_13_12_2.C_ON=1'b0;
    defparam shift_srl_89_12_LC_13_12_2.SEQ_MODE=4'b1000;
    defparam shift_srl_89_12_LC_13_12_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_89_12_LC_13_12_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59635),
            .lcout(shift_srl_89Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93089),
            .ce(N__61428),
            .sr(_gnd_net_));
    defparam shift_srl_89_13_LC_13_12_3.C_ON=1'b0;
    defparam shift_srl_89_13_LC_13_12_3.SEQ_MODE=4'b1000;
    defparam shift_srl_89_13_LC_13_12_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_89_13_LC_13_12_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59629),
            .lcout(shift_srl_89Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93089),
            .ce(N__61428),
            .sr(_gnd_net_));
    defparam shift_srl_89_14_LC_13_12_4.C_ON=1'b0;
    defparam shift_srl_89_14_LC_13_12_4.SEQ_MODE=4'b1000;
    defparam shift_srl_89_14_LC_13_12_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_89_14_LC_13_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59713),
            .lcout(shift_srl_89Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93089),
            .ce(N__61428),
            .sr(_gnd_net_));
    defparam shift_srl_89_9_LC_13_12_5.C_ON=1'b0;
    defparam shift_srl_89_9_LC_13_12_5.SEQ_MODE=4'b1000;
    defparam shift_srl_89_9_LC_13_12_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_89_9_LC_13_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59695),
            .lcout(shift_srl_89Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93089),
            .ce(N__61428),
            .sr(_gnd_net_));
    defparam shift_srl_89_8_LC_13_12_6.C_ON=1'b0;
    defparam shift_srl_89_8_LC_13_12_6.SEQ_MODE=4'b1000;
    defparam shift_srl_89_8_LC_13_12_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_89_8_LC_13_12_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59701),
            .lcout(shift_srl_89Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93089),
            .ce(N__61428),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNI87C56_15_LC_13_13_0.C_ON=1'b0;
    defparam shift_srl_0_RNI87C56_15_LC_13_13_0.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNI87C56_15_LC_13_13_0.LUT_INIT=16'b1100110000000000;
    LogicCell40 shift_srl_0_RNI87C56_15_LC_13_13_0 (
            .in0(_gnd_net_),
            .in1(N__90426),
            .in2(_gnd_net_),
            .in3(N__85194),
            .lcout(clk_en_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_24_0_LC_13_13_1.C_ON=1'b0;
    defparam shift_srl_24_0_LC_13_13_1.SEQ_MODE=4'b1000;
    defparam shift_srl_24_0_LC_13_13_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_24_0_LC_13_13_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83790),
            .lcout(shift_srl_24Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93074),
            .ce(N__63150),
            .sr(_gnd_net_));
    defparam shift_srl_24_1_LC_13_13_2.C_ON=1'b0;
    defparam shift_srl_24_1_LC_13_13_2.SEQ_MODE=4'b1000;
    defparam shift_srl_24_1_LC_13_13_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_24_1_LC_13_13_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59689),
            .lcout(shift_srl_24Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93074),
            .ce(N__63150),
            .sr(_gnd_net_));
    defparam shift_srl_24_2_LC_13_13_3.C_ON=1'b0;
    defparam shift_srl_24_2_LC_13_13_3.SEQ_MODE=4'b1000;
    defparam shift_srl_24_2_LC_13_13_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_24_2_LC_13_13_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59683),
            .lcout(shift_srl_24Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93074),
            .ce(N__63150),
            .sr(_gnd_net_));
    defparam shift_srl_24_3_LC_13_13_4.C_ON=1'b0;
    defparam shift_srl_24_3_LC_13_13_4.SEQ_MODE=4'b1000;
    defparam shift_srl_24_3_LC_13_13_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_24_3_LC_13_13_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59677),
            .lcout(shift_srl_24Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93074),
            .ce(N__63150),
            .sr(_gnd_net_));
    defparam shift_srl_143_0_LC_13_14_0.C_ON=1'b0;
    defparam shift_srl_143_0_LC_13_14_0.SEQ_MODE=4'b1000;
    defparam shift_srl_143_0_LC_13_14_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_143_0_LC_13_14_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61781),
            .lcout(shift_srl_143Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93058),
            .ce(N__59974),
            .sr(_gnd_net_));
    defparam shift_srl_143_1_LC_13_14_1.C_ON=1'b0;
    defparam shift_srl_143_1_LC_13_14_1.SEQ_MODE=4'b1000;
    defparam shift_srl_143_1_LC_13_14_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_143_1_LC_13_14_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59767),
            .lcout(shift_srl_143Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93058),
            .ce(N__59974),
            .sr(_gnd_net_));
    defparam shift_srl_143_2_LC_13_14_2.C_ON=1'b0;
    defparam shift_srl_143_2_LC_13_14_2.SEQ_MODE=4'b1000;
    defparam shift_srl_143_2_LC_13_14_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_143_2_LC_13_14_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59761),
            .lcout(shift_srl_143Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93058),
            .ce(N__59974),
            .sr(_gnd_net_));
    defparam shift_srl_143_3_LC_13_14_3.C_ON=1'b0;
    defparam shift_srl_143_3_LC_13_14_3.SEQ_MODE=4'b1000;
    defparam shift_srl_143_3_LC_13_14_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_143_3_LC_13_14_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59755),
            .lcout(shift_srl_143Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93058),
            .ce(N__59974),
            .sr(_gnd_net_));
    defparam shift_srl_143_4_LC_13_14_4.C_ON=1'b0;
    defparam shift_srl_143_4_LC_13_14_4.SEQ_MODE=4'b1000;
    defparam shift_srl_143_4_LC_13_14_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_143_4_LC_13_14_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59749),
            .lcout(shift_srl_143Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93058),
            .ce(N__59974),
            .sr(_gnd_net_));
    defparam shift_srl_143_5_LC_13_14_5.C_ON=1'b0;
    defparam shift_srl_143_5_LC_13_14_5.SEQ_MODE=4'b1000;
    defparam shift_srl_143_5_LC_13_14_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_143_5_LC_13_14_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59743),
            .lcout(shift_srl_143Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93058),
            .ce(N__59974),
            .sr(_gnd_net_));
    defparam shift_srl_143_6_LC_13_14_6.C_ON=1'b0;
    defparam shift_srl_143_6_LC_13_14_6.SEQ_MODE=4'b1000;
    defparam shift_srl_143_6_LC_13_14_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_143_6_LC_13_14_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59737),
            .lcout(shift_srl_143Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93058),
            .ce(N__59974),
            .sr(_gnd_net_));
    defparam shift_srl_143_7_LC_13_14_7.C_ON=1'b0;
    defparam shift_srl_143_7_LC_13_14_7.SEQ_MODE=4'b1000;
    defparam shift_srl_143_7_LC_13_14_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_143_7_LC_13_14_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59731),
            .lcout(shift_srl_143Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93058),
            .ce(N__59974),
            .sr(_gnd_net_));
    defparam shift_srl_26_0_LC_13_15_0.C_ON=1'b0;
    defparam shift_srl_26_0_LC_13_15_0.SEQ_MODE=4'b1000;
    defparam shift_srl_26_0_LC_13_15_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_26_0_LC_13_15_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71543),
            .lcout(shift_srl_26Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93044),
            .ce(N__64677),
            .sr(_gnd_net_));
    defparam shift_srl_26_1_LC_13_15_1.C_ON=1'b0;
    defparam shift_srl_26_1_LC_13_15_1.SEQ_MODE=4'b1000;
    defparam shift_srl_26_1_LC_13_15_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_26_1_LC_13_15_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59725),
            .lcout(shift_srl_26Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93044),
            .ce(N__64677),
            .sr(_gnd_net_));
    defparam shift_srl_26_2_LC_13_15_2.C_ON=1'b0;
    defparam shift_srl_26_2_LC_13_15_2.SEQ_MODE=4'b1000;
    defparam shift_srl_26_2_LC_13_15_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_26_2_LC_13_15_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59719),
            .lcout(shift_srl_26Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93044),
            .ce(N__64677),
            .sr(_gnd_net_));
    defparam shift_srl_26_3_LC_13_15_3.C_ON=1'b0;
    defparam shift_srl_26_3_LC_13_15_3.SEQ_MODE=4'b1000;
    defparam shift_srl_26_3_LC_13_15_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_26_3_LC_13_15_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59815),
            .lcout(shift_srl_26Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93044),
            .ce(N__64677),
            .sr(_gnd_net_));
    defparam shift_srl_26_4_LC_13_15_4.C_ON=1'b0;
    defparam shift_srl_26_4_LC_13_15_4.SEQ_MODE=4'b1000;
    defparam shift_srl_26_4_LC_13_15_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_26_4_LC_13_15_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59809),
            .lcout(shift_srl_26Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93044),
            .ce(N__64677),
            .sr(_gnd_net_));
    defparam shift_srl_26_5_LC_13_15_5.C_ON=1'b0;
    defparam shift_srl_26_5_LC_13_15_5.SEQ_MODE=4'b1000;
    defparam shift_srl_26_5_LC_13_15_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_26_5_LC_13_15_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59803),
            .lcout(shift_srl_26Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93044),
            .ce(N__64677),
            .sr(_gnd_net_));
    defparam shift_srl_26_6_LC_13_15_6.C_ON=1'b0;
    defparam shift_srl_26_6_LC_13_15_6.SEQ_MODE=4'b1000;
    defparam shift_srl_26_6_LC_13_15_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_26_6_LC_13_15_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59797),
            .lcout(shift_srl_26Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93044),
            .ce(N__64677),
            .sr(_gnd_net_));
    defparam shift_srl_26_7_LC_13_15_7.C_ON=1'b0;
    defparam shift_srl_26_7_LC_13_15_7.SEQ_MODE=4'b1000;
    defparam shift_srl_26_7_LC_13_15_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_26_7_LC_13_15_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59791),
            .lcout(shift_srl_26Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93044),
            .ce(N__64677),
            .sr(_gnd_net_));
    defparam shift_srl_121_0_LC_13_16_0.C_ON=1'b0;
    defparam shift_srl_121_0_LC_13_16_0.SEQ_MODE=4'b1000;
    defparam shift_srl_121_0_LC_13_16_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_121_0_LC_13_16_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78473),
            .lcout(shift_srl_121Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93030),
            .ce(N__59863),
            .sr(_gnd_net_));
    defparam shift_srl_121_1_LC_13_16_1.C_ON=1'b0;
    defparam shift_srl_121_1_LC_13_16_1.SEQ_MODE=4'b1000;
    defparam shift_srl_121_1_LC_13_16_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_121_1_LC_13_16_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59785),
            .lcout(shift_srl_121Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93030),
            .ce(N__59863),
            .sr(_gnd_net_));
    defparam shift_srl_121_2_LC_13_16_2.C_ON=1'b0;
    defparam shift_srl_121_2_LC_13_16_2.SEQ_MODE=4'b1000;
    defparam shift_srl_121_2_LC_13_16_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_121_2_LC_13_16_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59779),
            .lcout(shift_srl_121Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93030),
            .ce(N__59863),
            .sr(_gnd_net_));
    defparam shift_srl_121_3_LC_13_16_3.C_ON=1'b0;
    defparam shift_srl_121_3_LC_13_16_3.SEQ_MODE=4'b1000;
    defparam shift_srl_121_3_LC_13_16_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_121_3_LC_13_16_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59773),
            .lcout(shift_srl_121Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93030),
            .ce(N__59863),
            .sr(_gnd_net_));
    defparam shift_srl_121_4_LC_13_16_4.C_ON=1'b0;
    defparam shift_srl_121_4_LC_13_16_4.SEQ_MODE=4'b1000;
    defparam shift_srl_121_4_LC_13_16_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_121_4_LC_13_16_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59899),
            .lcout(shift_srl_121Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93030),
            .ce(N__59863),
            .sr(_gnd_net_));
    defparam shift_srl_121_5_LC_13_16_5.C_ON=1'b0;
    defparam shift_srl_121_5_LC_13_16_5.SEQ_MODE=4'b1000;
    defparam shift_srl_121_5_LC_13_16_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_121_5_LC_13_16_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59893),
            .lcout(shift_srl_121Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93030),
            .ce(N__59863),
            .sr(_gnd_net_));
    defparam shift_srl_121_6_LC_13_16_6.C_ON=1'b0;
    defparam shift_srl_121_6_LC_13_16_6.SEQ_MODE=4'b1000;
    defparam shift_srl_121_6_LC_13_16_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_121_6_LC_13_16_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59887),
            .lcout(shift_srl_121Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93030),
            .ce(N__59863),
            .sr(_gnd_net_));
    defparam shift_srl_121_7_LC_13_16_7.C_ON=1'b0;
    defparam shift_srl_121_7_LC_13_16_7.SEQ_MODE=4'b1000;
    defparam shift_srl_121_7_LC_13_16_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_121_7_LC_13_16_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59881),
            .lcout(shift_srl_121Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93030),
            .ce(N__59863),
            .sr(_gnd_net_));
    defparam shift_srl_143_10_LC_13_17_0.C_ON=1'b0;
    defparam shift_srl_143_10_LC_13_17_0.SEQ_MODE=4'b1000;
    defparam shift_srl_143_10_LC_13_17_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_143_10_LC_13_17_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59950),
            .lcout(shift_srl_143Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93010),
            .ce(N__59970),
            .sr(_gnd_net_));
    defparam shift_srl_143_11_LC_13_17_1.C_ON=1'b0;
    defparam shift_srl_143_11_LC_13_17_1.SEQ_MODE=4'b1000;
    defparam shift_srl_143_11_LC_13_17_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_143_11_LC_13_17_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59839),
            .lcout(shift_srl_143Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93010),
            .ce(N__59970),
            .sr(_gnd_net_));
    defparam shift_srl_143_12_LC_13_17_2.C_ON=1'b0;
    defparam shift_srl_143_12_LC_13_17_2.SEQ_MODE=4'b1000;
    defparam shift_srl_143_12_LC_13_17_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_143_12_LC_13_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59833),
            .lcout(shift_srl_143Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93010),
            .ce(N__59970),
            .sr(_gnd_net_));
    defparam shift_srl_143_13_LC_13_17_3.C_ON=1'b0;
    defparam shift_srl_143_13_LC_13_17_3.SEQ_MODE=4'b1000;
    defparam shift_srl_143_13_LC_13_17_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_143_13_LC_13_17_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59827),
            .lcout(shift_srl_143Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93010),
            .ce(N__59970),
            .sr(_gnd_net_));
    defparam shift_srl_143_14_LC_13_17_4.C_ON=1'b0;
    defparam shift_srl_143_14_LC_13_17_4.SEQ_MODE=4'b1000;
    defparam shift_srl_143_14_LC_13_17_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_143_14_LC_13_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59821),
            .lcout(shift_srl_143Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93010),
            .ce(N__59970),
            .sr(_gnd_net_));
    defparam shift_srl_143_15_LC_13_17_5.C_ON=1'b0;
    defparam shift_srl_143_15_LC_13_17_5.SEQ_MODE=4'b1000;
    defparam shift_srl_143_15_LC_13_17_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_143_15_LC_13_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59956),
            .lcout(shift_srl_143Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93010),
            .ce(N__59970),
            .sr(_gnd_net_));
    defparam shift_srl_143_9_LC_13_17_6.C_ON=1'b0;
    defparam shift_srl_143_9_LC_13_17_6.SEQ_MODE=4'b1000;
    defparam shift_srl_143_9_LC_13_17_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_143_9_LC_13_17_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59935),
            .lcout(shift_srl_143Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93010),
            .ce(N__59970),
            .sr(_gnd_net_));
    defparam shift_srl_143_8_LC_13_17_7.C_ON=1'b0;
    defparam shift_srl_143_8_LC_13_17_7.SEQ_MODE=4'b1000;
    defparam shift_srl_143_8_LC_13_17_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_143_8_LC_13_17_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59944),
            .lcout(shift_srl_143Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93010),
            .ce(N__59970),
            .sr(_gnd_net_));
    defparam shift_srl_117_0_LC_13_18_0.C_ON=1'b0;
    defparam shift_srl_117_0_LC_13_18_0.SEQ_MODE=4'b1000;
    defparam shift_srl_117_0_LC_13_18_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_117_0_LC_13_18_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66442),
            .lcout(shift_srl_117Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93031),
            .ce(N__65064),
            .sr(_gnd_net_));
    defparam shift_srl_117_1_LC_13_18_1.C_ON=1'b0;
    defparam shift_srl_117_1_LC_13_18_1.SEQ_MODE=4'b1000;
    defparam shift_srl_117_1_LC_13_18_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_117_1_LC_13_18_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59929),
            .lcout(shift_srl_117Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93031),
            .ce(N__65064),
            .sr(_gnd_net_));
    defparam shift_srl_117_2_LC_13_18_2.C_ON=1'b0;
    defparam shift_srl_117_2_LC_13_18_2.SEQ_MODE=4'b1000;
    defparam shift_srl_117_2_LC_13_18_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_117_2_LC_13_18_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59923),
            .lcout(shift_srl_117Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93031),
            .ce(N__65064),
            .sr(_gnd_net_));
    defparam shift_srl_117_3_LC_13_18_3.C_ON=1'b0;
    defparam shift_srl_117_3_LC_13_18_3.SEQ_MODE=4'b1000;
    defparam shift_srl_117_3_LC_13_18_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_117_3_LC_13_18_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59917),
            .lcout(shift_srl_117Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93031),
            .ce(N__65064),
            .sr(_gnd_net_));
    defparam shift_srl_117_4_LC_13_18_4.C_ON=1'b0;
    defparam shift_srl_117_4_LC_13_18_4.SEQ_MODE=4'b1000;
    defparam shift_srl_117_4_LC_13_18_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_117_4_LC_13_18_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59911),
            .lcout(shift_srl_117Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93031),
            .ce(N__65064),
            .sr(_gnd_net_));
    defparam shift_srl_117_5_LC_13_18_5.C_ON=1'b0;
    defparam shift_srl_117_5_LC_13_18_5.SEQ_MODE=4'b1000;
    defparam shift_srl_117_5_LC_13_18_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_117_5_LC_13_18_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59905),
            .lcout(shift_srl_117Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93031),
            .ce(N__65064),
            .sr(_gnd_net_));
    defparam shift_srl_117_6_LC_13_18_6.C_ON=1'b0;
    defparam shift_srl_117_6_LC_13_18_6.SEQ_MODE=4'b1000;
    defparam shift_srl_117_6_LC_13_18_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_117_6_LC_13_18_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60037),
            .lcout(shift_srl_117Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93031),
            .ce(N__65064),
            .sr(_gnd_net_));
    defparam shift_srl_117_7_LC_13_18_7.C_ON=1'b0;
    defparam shift_srl_117_7_LC_13_18_7.SEQ_MODE=4'b1000;
    defparam shift_srl_117_7_LC_13_18_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_117_7_LC_13_18_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60031),
            .lcout(shift_srl_117Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93031),
            .ce(N__65064),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_143_LC_13_19_0.C_ON=1'b0;
    defparam rco_obuf_RNO_143_LC_13_19_0.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_143_LC_13_19_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 rco_obuf_RNO_143_LC_13_19_0 (
            .in0(N__91083),
            .in1(N__63762),
            .in2(N__61787),
            .in3(N__66603),
            .lcout(rco_c_143),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_142_LC_13_19_1.C_ON=1'b0;
    defparam rco_obuf_RNO_142_LC_13_19_1.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_142_LC_13_19_1.LUT_INIT=16'b1000100000000000;
    LogicCell40 rco_obuf_RNO_142_LC_13_19_1 (
            .in0(N__66602),
            .in1(N__63761),
            .in2(_gnd_net_),
            .in3(N__91082),
            .lcout(rco_c_142),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_143_RNI929B1_15_LC_13_19_2.C_ON=1'b0;
    defparam shift_srl_143_RNI929B1_15_LC_13_19_2.SEQ_MODE=4'b0000;
    defparam shift_srl_143_RNI929B1_15_LC_13_19_2.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_143_RNI929B1_15_LC_13_19_2 (
            .in0(N__61777),
            .in1(N__90350),
            .in2(N__63766),
            .in3(N__66601),
            .lcout(),
            .ltout(clk_en_0_a3_0_a2_sx_144_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_143_RNIES6841_15_LC_13_19_3.C_ON=1'b0;
    defparam shift_srl_143_RNIES6841_15_LC_13_19_3.SEQ_MODE=4'b0000;
    defparam shift_srl_143_RNIES6841_15_LC_13_19_3.LUT_INIT=16'b0000100000000000;
    LogicCell40 shift_srl_143_RNIES6841_15_LC_13_19_3 (
            .in0(N__65028),
            .in1(N__64979),
            .in2(N__59992),
            .in3(N__79335),
            .lcout(clk_en_144),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_142_RNI8HFB4_15_LC_13_19_4.C_ON=1'b0;
    defparam shift_srl_142_RNI8HFB4_15_LC_13_19_4.SEQ_MODE=4'b0000;
    defparam shift_srl_142_RNI8HFB4_15_LC_13_19_4.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_142_RNI8HFB4_15_LC_13_19_4 (
            .in0(N__64978),
            .in1(N__90349),
            .in2(N__63765),
            .in3(N__66600),
            .lcout(),
            .ltout(clk_en_0_a3_0_a2_sx_143_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_142_RNIBT1441_15_LC_13_19_5.C_ON=1'b0;
    defparam shift_srl_142_RNIBT1441_15_LC_13_19_5.SEQ_MODE=4'b0000;
    defparam shift_srl_142_RNIBT1441_15_LC_13_19_5.LUT_INIT=16'b0000110000000000;
    LogicCell40 shift_srl_142_RNIBT1441_15_LC_13_19_5 (
            .in0(_gnd_net_),
            .in1(N__65027),
            .in2(N__59977),
            .in3(N__79334),
            .lcout(clk_en_143),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_91_RNIGQ0UO_15_LC_13_19_6.C_ON=1'b0;
    defparam shift_srl_91_RNIGQ0UO_15_LC_13_19_6.SEQ_MODE=4'b0000;
    defparam shift_srl_91_RNIGQ0UO_15_LC_13_19_6.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_91_RNIGQ0UO_15_LC_13_19_6 (
            .in0(N__85160),
            .in1(N__72033),
            .in2(N__72096),
            .in3(N__75081),
            .lcout(rco_c_99),
            .ltout(rco_c_99_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_107_RNII8C2S_15_LC_13_19_7.C_ON=1'b0;
    defparam shift_srl_107_RNII8C2S_15_LC_13_19_7.SEQ_MODE=4'b0000;
    defparam shift_srl_107_RNII8C2S_15_LC_13_19_7.LUT_INIT=16'b1111000000000000;
    LogicCell40 shift_srl_107_RNII8C2S_15_LC_13_19_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__60139),
            .in3(N__64977),
            .lcout(rco_c_110),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_122_0_LC_13_20_0.C_ON=1'b0;
    defparam shift_srl_122_0_LC_13_20_0.SEQ_MODE=4'b1000;
    defparam shift_srl_122_0_LC_13_20_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_122_0_LC_13_20_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60132),
            .lcout(shift_srl_122Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93059),
            .ce(N__60052),
            .sr(_gnd_net_));
    defparam shift_srl_122_1_LC_13_20_1.C_ON=1'b0;
    defparam shift_srl_122_1_LC_13_20_1.SEQ_MODE=4'b1000;
    defparam shift_srl_122_1_LC_13_20_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_122_1_LC_13_20_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60103),
            .lcout(shift_srl_122Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93059),
            .ce(N__60052),
            .sr(_gnd_net_));
    defparam shift_srl_122_2_LC_13_20_2.C_ON=1'b0;
    defparam shift_srl_122_2_LC_13_20_2.SEQ_MODE=4'b1000;
    defparam shift_srl_122_2_LC_13_20_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_122_2_LC_13_20_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60097),
            .lcout(shift_srl_122Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93059),
            .ce(N__60052),
            .sr(_gnd_net_));
    defparam shift_srl_122_3_LC_13_20_3.C_ON=1'b0;
    defparam shift_srl_122_3_LC_13_20_3.SEQ_MODE=4'b1000;
    defparam shift_srl_122_3_LC_13_20_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_122_3_LC_13_20_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60091),
            .lcout(shift_srl_122Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93059),
            .ce(N__60052),
            .sr(_gnd_net_));
    defparam shift_srl_122_4_LC_13_20_4.C_ON=1'b0;
    defparam shift_srl_122_4_LC_13_20_4.SEQ_MODE=4'b1000;
    defparam shift_srl_122_4_LC_13_20_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_122_4_LC_13_20_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60085),
            .lcout(shift_srl_122Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93059),
            .ce(N__60052),
            .sr(_gnd_net_));
    defparam shift_srl_122_5_LC_13_20_5.C_ON=1'b0;
    defparam shift_srl_122_5_LC_13_20_5.SEQ_MODE=4'b1000;
    defparam shift_srl_122_5_LC_13_20_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_122_5_LC_13_20_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60079),
            .lcout(shift_srl_122Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93059),
            .ce(N__60052),
            .sr(_gnd_net_));
    defparam shift_srl_122_6_LC_13_20_6.C_ON=1'b0;
    defparam shift_srl_122_6_LC_13_20_6.SEQ_MODE=4'b1000;
    defparam shift_srl_122_6_LC_13_20_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_122_6_LC_13_20_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60073),
            .lcout(shift_srl_122Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93059),
            .ce(N__60052),
            .sr(_gnd_net_));
    defparam shift_srl_122_7_LC_13_20_7.C_ON=1'b0;
    defparam shift_srl_122_7_LC_13_20_7.SEQ_MODE=4'b1000;
    defparam shift_srl_122_7_LC_13_20_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_122_7_LC_13_20_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60067),
            .lcout(shift_srl_122Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93059),
            .ce(N__60052),
            .sr(_gnd_net_));
    defparam shift_srl_142_10_LC_13_21_0.C_ON=1'b0;
    defparam shift_srl_142_10_LC_13_21_0.SEQ_MODE=4'b1000;
    defparam shift_srl_142_10_LC_13_21_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_142_10_LC_13_21_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60181),
            .lcout(shift_srl_142Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93075),
            .ce(N__63655),
            .sr(_gnd_net_));
    defparam shift_srl_142_11_LC_13_21_1.C_ON=1'b0;
    defparam shift_srl_142_11_LC_13_21_1.SEQ_MODE=4'b1000;
    defparam shift_srl_142_11_LC_13_21_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_142_11_LC_13_21_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60211),
            .lcout(shift_srl_142Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93075),
            .ce(N__63655),
            .sr(_gnd_net_));
    defparam shift_srl_142_12_LC_13_21_2.C_ON=1'b0;
    defparam shift_srl_142_12_LC_13_21_2.SEQ_MODE=4'b1000;
    defparam shift_srl_142_12_LC_13_21_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_142_12_LC_13_21_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60205),
            .lcout(shift_srl_142Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93075),
            .ce(N__63655),
            .sr(_gnd_net_));
    defparam shift_srl_142_13_LC_13_21_3.C_ON=1'b0;
    defparam shift_srl_142_13_LC_13_21_3.SEQ_MODE=4'b1000;
    defparam shift_srl_142_13_LC_13_21_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_142_13_LC_13_21_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60199),
            .lcout(shift_srl_142Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93075),
            .ce(N__63655),
            .sr(_gnd_net_));
    defparam shift_srl_142_14_LC_13_21_4.C_ON=1'b0;
    defparam shift_srl_142_14_LC_13_21_4.SEQ_MODE=4'b1000;
    defparam shift_srl_142_14_LC_13_21_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_142_14_LC_13_21_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60193),
            .lcout(shift_srl_142Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93075),
            .ce(N__63655),
            .sr(_gnd_net_));
    defparam shift_srl_142_15_LC_13_21_5.C_ON=1'b0;
    defparam shift_srl_142_15_LC_13_21_5.SEQ_MODE=4'b1000;
    defparam shift_srl_142_15_LC_13_21_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_142_15_LC_13_21_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60187),
            .lcout(shift_srl_142Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93075),
            .ce(N__63655),
            .sr(_gnd_net_));
    defparam shift_srl_142_9_LC_13_21_6.C_ON=1'b0;
    defparam shift_srl_142_9_LC_13_21_6.SEQ_MODE=4'b1000;
    defparam shift_srl_142_9_LC_13_21_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_142_9_LC_13_21_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60175),
            .lcout(shift_srl_142Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93075),
            .ce(N__63655),
            .sr(_gnd_net_));
    defparam shift_srl_142_8_LC_13_21_7.C_ON=1'b0;
    defparam shift_srl_142_8_LC_13_21_7.SEQ_MODE=4'b1000;
    defparam shift_srl_142_8_LC_13_21_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_142_8_LC_13_21_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63664),
            .lcout(shift_srl_142Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93075),
            .ce(N__63655),
            .sr(_gnd_net_));
    defparam shift_srl_111_RNIBS0GS_15_LC_13_22_0.C_ON=1'b0;
    defparam shift_srl_111_RNIBS0GS_15_LC_13_22_0.SEQ_MODE=4'b0000;
    defparam shift_srl_111_RNIBS0GS_15_LC_13_22_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_111_RNIBS0GS_15_LC_13_22_0 (
            .in0(N__64947),
            .in1(N__79397),
            .in2(N__60753),
            .in3(N__90329),
            .lcout(clk_en_112),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_111_15_LC_13_22_1.C_ON=1'b0;
    defparam shift_srl_111_15_LC_13_22_1.SEQ_MODE=4'b1000;
    defparam shift_srl_111_15_LC_13_22_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_111_15_LC_13_22_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60235),
            .lcout(shift_srl_111Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93090),
            .ce(N__68114),
            .sr(_gnd_net_));
    defparam shift_srl_112_RNI6OUT_15_LC_13_22_2.C_ON=1'b0;
    defparam shift_srl_112_RNI6OUT_15_LC_13_22_2.SEQ_MODE=4'b0000;
    defparam shift_srl_112_RNI6OUT_15_LC_13_22_2.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_112_RNI6OUT_15_LC_13_22_2 (
            .in0(N__60504),
            .in1(N__66386),
            .in2(N__60333),
            .in3(N__60705),
            .lcout(rco_int_0_a3_0_a2_138_m6_0_a2_7_4_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_112_RNIFS6GS_15_LC_13_22_3.C_ON=1'b0;
    defparam shift_srl_112_RNIFS6GS_15_LC_13_22_3.SEQ_MODE=4'b0000;
    defparam shift_srl_112_RNIFS6GS_15_LC_13_22_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_112_RNIFS6GS_15_LC_13_22_3 (
            .in0(N__79398),
            .in1(N__64948),
            .in2(N__60731),
            .in3(N__60505),
            .lcout(N_91),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIDK63S_15_LC_13_22_4.C_ON=1'b0;
    defparam shift_srl_0_RNIDK63S_15_LC_13_22_4.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIDK63S_15_LC_13_22_4.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_0_RNIDK63S_15_LC_13_22_4 (
            .in0(N__64946),
            .in1(N__79396),
            .in2(_gnd_net_),
            .in3(N__90328),
            .lcout(clk_en_111),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_118_RNI6U9L3_15_LC_13_22_5.C_ON=1'b0;
    defparam shift_srl_118_RNI6U9L3_15_LC_13_22_5.SEQ_MODE=4'b0000;
    defparam shift_srl_118_RNI6U9L3_15_LC_13_22_5.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_118_RNI6U9L3_15_LC_13_22_5 (
            .in0(N__66387),
            .in1(N__64945),
            .in2(N__90474),
            .in3(N__60327),
            .lcout(clk_en_0_a3_0_a2_sx_119),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_111_14_LC_13_22_6.C_ON=1'b0;
    defparam shift_srl_111_14_LC_13_22_6.SEQ_MODE=4'b1000;
    defparam shift_srl_111_14_LC_13_22_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_111_14_LC_13_22_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60229),
            .lcout(shift_srl_111Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93090),
            .ce(N__68114),
            .sr(_gnd_net_));
    defparam shift_srl_111_13_LC_13_22_7.C_ON=1'b0;
    defparam shift_srl_111_13_LC_13_22_7.SEQ_MODE=4'b1000;
    defparam shift_srl_111_13_LC_13_22_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_111_13_LC_13_22_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67984),
            .lcout(shift_srl_111Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93090),
            .ce(N__68114),
            .sr(_gnd_net_));
    defparam shift_srl_111_0_LC_13_23_0.C_ON=1'b0;
    defparam shift_srl_111_0_LC_13_23_0.SEQ_MODE=4'b1000;
    defparam shift_srl_111_0_LC_13_23_0.LUT_INIT=16'b1100110011001100;
    LogicCell40 shift_srl_111_0_LC_13_23_0 (
            .in0(_gnd_net_),
            .in1(N__60730),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_111Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93105),
            .ce(N__68125),
            .sr(_gnd_net_));
    defparam shift_srl_111_1_LC_13_23_1.C_ON=1'b0;
    defparam shift_srl_111_1_LC_13_23_1.SEQ_MODE=4'b1000;
    defparam shift_srl_111_1_LC_13_23_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_111_1_LC_13_23_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60223),
            .lcout(shift_srl_111Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93105),
            .ce(N__68125),
            .sr(_gnd_net_));
    defparam shift_srl_111_2_LC_13_23_2.C_ON=1'b0;
    defparam shift_srl_111_2_LC_13_23_2.SEQ_MODE=4'b1000;
    defparam shift_srl_111_2_LC_13_23_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_111_2_LC_13_23_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60217),
            .lcout(shift_srl_111Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93105),
            .ce(N__68125),
            .sr(_gnd_net_));
    defparam shift_srl_111_3_LC_13_23_3.C_ON=1'b0;
    defparam shift_srl_111_3_LC_13_23_3.SEQ_MODE=4'b1000;
    defparam shift_srl_111_3_LC_13_23_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_111_3_LC_13_23_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60565),
            .lcout(shift_srl_111Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93105),
            .ce(N__68125),
            .sr(_gnd_net_));
    defparam shift_srl_111_4_LC_13_23_4.C_ON=1'b0;
    defparam shift_srl_111_4_LC_13_23_4.SEQ_MODE=4'b1000;
    defparam shift_srl_111_4_LC_13_23_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_111_4_LC_13_23_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60559),
            .lcout(shift_srl_111Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93105),
            .ce(N__68125),
            .sr(_gnd_net_));
    defparam shift_srl_111_5_LC_13_23_5.C_ON=1'b0;
    defparam shift_srl_111_5_LC_13_23_5.SEQ_MODE=4'b1000;
    defparam shift_srl_111_5_LC_13_23_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_111_5_LC_13_23_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60553),
            .lcout(shift_srl_111Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93105),
            .ce(N__68125),
            .sr(_gnd_net_));
    defparam shift_srl_111_6_LC_13_23_6.C_ON=1'b0;
    defparam shift_srl_111_6_LC_13_23_6.SEQ_MODE=4'b1000;
    defparam shift_srl_111_6_LC_13_23_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_111_6_LC_13_23_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60547),
            .lcout(shift_srl_111Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93105),
            .ce(N__68125),
            .sr(_gnd_net_));
    defparam shift_srl_111_7_LC_13_23_7.C_ON=1'b0;
    defparam shift_srl_111_7_LC_13_23_7.SEQ_MODE=4'b1000;
    defparam shift_srl_111_7_LC_13_23_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_111_7_LC_13_23_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60541),
            .lcout(shift_srl_111Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93105),
            .ce(N__68125),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIB6RUO_15_LC_13_24_0.C_ON=1'b0;
    defparam shift_srl_0_RNIB6RUO_15_LC_13_24_0.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIB6RUO_15_LC_13_24_0.LUT_INIT=16'b1100110000000000;
    LogicCell40 shift_srl_0_RNIB6RUO_15_LC_13_24_0 (
            .in0(_gnd_net_),
            .in1(N__90475),
            .in2(_gnd_net_),
            .in3(N__79464),
            .lcout(clk_en_100),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_112_RNIV16I3_15_LC_13_24_1.C_ON=1'b0;
    defparam shift_srl_112_RNIV16I3_15_LC_13_24_1.SEQ_MODE=4'b0000;
    defparam shift_srl_112_RNIV16I3_15_LC_13_24_1.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_112_RNIV16I3_15_LC_13_24_1 (
            .in0(N__64944),
            .in1(N__60530),
            .in2(_gnd_net_),
            .in3(N__60765),
            .lcout(),
            .ltout(shift_srl_112_RNIV16I3Z0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_113_RNIAO7MS_15_LC_13_24_2.C_ON=1'b0;
    defparam shift_srl_113_RNIAO7MS_15_LC_13_24_2.SEQ_MODE=4'b0000;
    defparam shift_srl_113_RNIAO7MS_15_LC_13_24_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_113_RNIAO7MS_15_LC_13_24_2 (
            .in0(N__90482),
            .in1(N__60448),
            .in2(N__60385),
            .in3(N__79465),
            .lcout(clk_en_114),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_116_RNILK5ET_15_LC_13_24_3.C_ON=1'b0;
    defparam shift_srl_116_RNILK5ET_15_LC_13_24_3.SEQ_MODE=4'b0000;
    defparam shift_srl_116_RNILK5ET_15_LC_13_24_3.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_116_RNILK5ET_15_LC_13_24_3 (
            .in0(N__79466),
            .in1(N__64951),
            .in2(_gnd_net_),
            .in3(N__65903),
            .lcout(rco_c_116),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_117_RNIK0VKT_15_LC_13_24_5.C_ON=1'b0;
    defparam shift_srl_117_RNIK0VKT_15_LC_13_24_5.SEQ_MODE=4'b0000;
    defparam shift_srl_117_RNIK0VKT_15_LC_13_24_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_117_RNIK0VKT_15_LC_13_24_5 (
            .in0(N__65904),
            .in1(N__66441),
            .in2(N__90551),
            .in3(N__61975),
            .lcout(clk_en_118),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_111_LC_13_24_6.C_ON=1'b0;
    defparam rco_obuf_RNO_111_LC_13_24_6.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_111_LC_13_24_6.LUT_INIT=16'b1010000010100000;
    LogicCell40 rco_obuf_RNO_111_LC_13_24_6 (
            .in0(N__61976),
            .in1(_gnd_net_),
            .in2(N__60776),
            .in3(_gnd_net_),
            .lcout(rco_c_111),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_116_RNI9BE15_15_LC_13_24_7.C_ON=1'b0;
    defparam shift_srl_116_RNI9BE15_15_LC_13_24_7.SEQ_MODE=4'b0000;
    defparam shift_srl_116_RNI9BE15_15_LC_13_24_7.LUT_INIT=16'b0111011111111111;
    LogicCell40 shift_srl_116_RNI9BE15_15_LC_13_24_7 (
            .in0(N__64943),
            .in1(N__65523),
            .in2(_gnd_net_),
            .in3(N__65902),
            .lcout(rco_int_0_a2_1_a2_1_120),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_199_LC_13_25_0.C_ON=1'b0;
    defparam rco_obuf_RNO_199_LC_13_25_0.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_199_LC_13_25_0.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_199_LC_13_25_0 (
            .in0(N__62506),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70452),
            .lcout(rco_c_199),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_199_0_LC_13_25_1.C_ON=1'b0;
    defparam shift_srl_199_0_LC_13_25_1.SEQ_MODE=4'b1000;
    defparam shift_srl_199_0_LC_13_25_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_199_0_LC_13_25_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62505),
            .lcout(shift_srl_199Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93142),
            .ce(N__62721),
            .sr(_gnd_net_));
    defparam shift_srl_199_1_LC_13_25_2.C_ON=1'b0;
    defparam shift_srl_199_1_LC_13_25_2.SEQ_MODE=4'b1000;
    defparam shift_srl_199_1_LC_13_25_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_199_1_LC_13_25_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60595),
            .lcout(shift_srl_199Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93142),
            .ce(N__62721),
            .sr(_gnd_net_));
    defparam shift_srl_199_2_LC_13_25_3.C_ON=1'b0;
    defparam shift_srl_199_2_LC_13_25_3.SEQ_MODE=4'b1000;
    defparam shift_srl_199_2_LC_13_25_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_199_2_LC_13_25_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60589),
            .lcout(shift_srl_199Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93142),
            .ce(N__62721),
            .sr(_gnd_net_));
    defparam shift_srl_199_3_LC_13_25_4.C_ON=1'b0;
    defparam shift_srl_199_3_LC_13_25_4.SEQ_MODE=4'b1000;
    defparam shift_srl_199_3_LC_13_25_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_199_3_LC_13_25_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60583),
            .lcout(shift_srl_199Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93142),
            .ce(N__62721),
            .sr(_gnd_net_));
    defparam shift_srl_199_4_LC_13_25_5.C_ON=1'b0;
    defparam shift_srl_199_4_LC_13_25_5.SEQ_MODE=4'b1000;
    defparam shift_srl_199_4_LC_13_25_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_199_4_LC_13_25_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60577),
            .lcout(shift_srl_199Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93142),
            .ce(N__62721),
            .sr(_gnd_net_));
    defparam shift_srl_199_5_LC_13_25_6.C_ON=1'b0;
    defparam shift_srl_199_5_LC_13_25_6.SEQ_MODE=4'b1000;
    defparam shift_srl_199_5_LC_13_25_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_199_5_LC_13_25_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60571),
            .lcout(shift_srl_199Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93142),
            .ce(N__62721),
            .sr(_gnd_net_));
    defparam shift_srl_199_6_LC_13_25_7.C_ON=1'b0;
    defparam shift_srl_199_6_LC_13_25_7.SEQ_MODE=4'b1000;
    defparam shift_srl_199_6_LC_13_25_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_199_6_LC_13_25_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60868),
            .lcout(shift_srl_199Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93142),
            .ce(N__62721),
            .sr(_gnd_net_));
    defparam shift_srl_102_10_LC_13_26_0.C_ON=1'b0;
    defparam shift_srl_102_10_LC_13_26_0.SEQ_MODE=4'b1000;
    defparam shift_srl_102_10_LC_13_26_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_102_10_LC_13_26_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62623),
            .lcout(shift_srl_102Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93160),
            .ce(N__62610),
            .sr(_gnd_net_));
    defparam shift_srl_102_11_LC_13_26_1.C_ON=1'b0;
    defparam shift_srl_102_11_LC_13_26_1.SEQ_MODE=4'b1000;
    defparam shift_srl_102_11_LC_13_26_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_102_11_LC_13_26_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60847),
            .lcout(shift_srl_102Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93160),
            .ce(N__62610),
            .sr(_gnd_net_));
    defparam shift_srl_102_12_LC_13_26_2.C_ON=1'b0;
    defparam shift_srl_102_12_LC_13_26_2.SEQ_MODE=4'b1000;
    defparam shift_srl_102_12_LC_13_26_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_102_12_LC_13_26_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60841),
            .lcout(shift_srl_102Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93160),
            .ce(N__62610),
            .sr(_gnd_net_));
    defparam shift_srl_102_13_LC_13_26_3.C_ON=1'b0;
    defparam shift_srl_102_13_LC_13_26_3.SEQ_MODE=4'b1000;
    defparam shift_srl_102_13_LC_13_26_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_102_13_LC_13_26_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60835),
            .lcout(shift_srl_102Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93160),
            .ce(N__62610),
            .sr(_gnd_net_));
    defparam shift_srl_102_14_LC_13_26_4.C_ON=1'b0;
    defparam shift_srl_102_14_LC_13_26_4.SEQ_MODE=4'b1000;
    defparam shift_srl_102_14_LC_13_26_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_102_14_LC_13_26_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60829),
            .lcout(shift_srl_102Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93160),
            .ce(N__62610),
            .sr(_gnd_net_));
    defparam shift_srl_102_15_LC_13_26_5.C_ON=1'b0;
    defparam shift_srl_102_15_LC_13_26_5.SEQ_MODE=4'b1000;
    defparam shift_srl_102_15_LC_13_26_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_102_15_LC_13_26_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60823),
            .lcout(shift_srl_102Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93160),
            .ce(N__62610),
            .sr(_gnd_net_));
    defparam shift_srl_102_7_LC_13_26_6.C_ON=1'b0;
    defparam shift_srl_102_7_LC_13_26_6.SEQ_MODE=4'b1000;
    defparam shift_srl_102_7_LC_13_26_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_102_7_LC_13_26_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62635),
            .lcout(shift_srl_102Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93160),
            .ce(N__62610),
            .sr(_gnd_net_));
    defparam shift_srl_102_8_LC_13_26_7.C_ON=1'b0;
    defparam shift_srl_102_8_LC_13_26_7.SEQ_MODE=4'b1000;
    defparam shift_srl_102_8_LC_13_26_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_102_8_LC_13_26_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60817),
            .lcout(shift_srl_102Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93160),
            .ce(N__62610),
            .sr(_gnd_net_));
    defparam shift_srl_101_RNI48LFP_15_LC_13_27_0.C_ON=1'b0;
    defparam shift_srl_101_RNI48LFP_15_LC_13_27_0.SEQ_MODE=4'b0000;
    defparam shift_srl_101_RNI48LFP_15_LC_13_27_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_101_RNI48LFP_15_LC_13_27_0 (
            .in0(N__60974),
            .in1(N__79675),
            .in2(N__90562),
            .in3(N__79541),
            .lcout(clk_en_102),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_100_15_LC_13_27_1.C_ON=1'b0;
    defparam shift_srl_100_15_LC_13_27_1.SEQ_MODE=4'b1000;
    defparam shift_srl_100_15_LC_13_27_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_100_15_LC_13_27_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60928),
            .lcout(shift_srl_100Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93179),
            .ce(N__60891),
            .sr(_gnd_net_));
    defparam shift_srl_104_RNIRO881_15_LC_13_27_2.C_ON=1'b0;
    defparam shift_srl_104_RNIRO881_15_LC_13_27_2.SEQ_MODE=4'b0000;
    defparam shift_srl_104_RNIRO881_15_LC_13_27_2.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_104_RNIRO881_15_LC_13_27_2 (
            .in0(N__60998),
            .in1(N__61089),
            .in2(_gnd_net_),
            .in3(N__79673),
            .lcout(rco_int_0_a3_0_a2_s_0_1_104),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_104_RNIOROA1_15_LC_13_27_3.C_ON=1'b0;
    defparam shift_srl_104_RNIOROA1_15_LC_13_27_3.SEQ_MODE=4'b0000;
    defparam shift_srl_104_RNIOROA1_15_LC_13_27_3.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_104_RNIOROA1_15_LC_13_27_3 (
            .in0(N__79674),
            .in1(N__60999),
            .in2(N__61096),
            .in3(N__60973),
            .lcout(rco_int_0_a3_0_a2_s_0_sx_104),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_100_14_LC_13_27_4.C_ON=1'b0;
    defparam shift_srl_100_14_LC_13_27_4.SEQ_MODE=4'b1000;
    defparam shift_srl_100_14_LC_13_27_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_100_14_LC_13_27_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60922),
            .lcout(shift_srl_100Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93179),
            .ce(N__60891),
            .sr(_gnd_net_));
    defparam shift_srl_100_13_LC_13_27_5.C_ON=1'b0;
    defparam shift_srl_100_13_LC_13_27_5.SEQ_MODE=4'b1000;
    defparam shift_srl_100_13_LC_13_27_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_100_13_LC_13_27_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60916),
            .lcout(shift_srl_100Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93179),
            .ce(N__60891),
            .sr(_gnd_net_));
    defparam shift_srl_100_12_LC_13_27_6.C_ON=1'b0;
    defparam shift_srl_100_12_LC_13_27_6.SEQ_MODE=4'b1000;
    defparam shift_srl_100_12_LC_13_27_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_100_12_LC_13_27_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60901),
            .lcout(shift_srl_100Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93179),
            .ce(N__60891),
            .sr(_gnd_net_));
    defparam shift_srl_100_11_LC_13_27_7.C_ON=1'b0;
    defparam shift_srl_100_11_LC_13_27_7.SEQ_MODE=4'b1000;
    defparam shift_srl_100_11_LC_13_27_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_100_11_LC_13_27_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60910),
            .lcout(shift_srl_100Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93179),
            .ce(N__60891),
            .sr(_gnd_net_));
    defparam shift_srl_103_10_LC_13_28_0.C_ON=1'b0;
    defparam shift_srl_103_10_LC_13_28_0.SEQ_MODE=4'b1000;
    defparam shift_srl_103_10_LC_13_28_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_103_10_LC_13_28_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61069),
            .lcout(shift_srl_103Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93201),
            .ce(N__61048),
            .sr(_gnd_net_));
    defparam shift_srl_103_11_LC_13_28_1.C_ON=1'b0;
    defparam shift_srl_103_11_LC_13_28_1.SEQ_MODE=4'b1000;
    defparam shift_srl_103_11_LC_13_28_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_103_11_LC_13_28_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61126),
            .lcout(shift_srl_103Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93201),
            .ce(N__61048),
            .sr(_gnd_net_));
    defparam shift_srl_103_12_LC_13_28_2.C_ON=1'b0;
    defparam shift_srl_103_12_LC_13_28_2.SEQ_MODE=4'b1000;
    defparam shift_srl_103_12_LC_13_28_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_103_12_LC_13_28_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61120),
            .lcout(shift_srl_103Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93201),
            .ce(N__61048),
            .sr(_gnd_net_));
    defparam shift_srl_103_13_LC_13_28_3.C_ON=1'b0;
    defparam shift_srl_103_13_LC_13_28_3.SEQ_MODE=4'b1000;
    defparam shift_srl_103_13_LC_13_28_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_103_13_LC_13_28_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61114),
            .lcout(shift_srl_103Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93201),
            .ce(N__61048),
            .sr(_gnd_net_));
    defparam shift_srl_103_14_LC_13_28_4.C_ON=1'b0;
    defparam shift_srl_103_14_LC_13_28_4.SEQ_MODE=4'b1000;
    defparam shift_srl_103_14_LC_13_28_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_103_14_LC_13_28_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61108),
            .lcout(shift_srl_103Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93201),
            .ce(N__61048),
            .sr(_gnd_net_));
    defparam shift_srl_103_15_LC_13_28_5.C_ON=1'b0;
    defparam shift_srl_103_15_LC_13_28_5.SEQ_MODE=4'b1000;
    defparam shift_srl_103_15_LC_13_28_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_103_15_LC_13_28_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61102),
            .lcout(shift_srl_103Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93201),
            .ce(N__61048),
            .sr(_gnd_net_));
    defparam shift_srl_103_9_LC_13_28_6.C_ON=1'b0;
    defparam shift_srl_103_9_LC_13_28_6.SEQ_MODE=4'b1000;
    defparam shift_srl_103_9_LC_13_28_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_103_9_LC_13_28_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61054),
            .lcout(shift_srl_103Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93201),
            .ce(N__61048),
            .sr(_gnd_net_));
    defparam shift_srl_103_8_LC_13_28_7.C_ON=1'b0;
    defparam shift_srl_103_8_LC_13_28_7.SEQ_MODE=4'b1000;
    defparam shift_srl_103_8_LC_13_28_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_103_8_LC_13_28_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61063),
            .lcout(shift_srl_103Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93201),
            .ce(N__61048),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_87_LC_14_3_2.C_ON=1'b0;
    defparam rco_obuf_RNO_87_LC_14_3_2.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_87_LC_14_3_2.LUT_INIT=16'b1000100000000000;
    LogicCell40 rco_obuf_RNO_87_LC_14_3_2 (
            .in0(N__68522),
            .in1(N__67106),
            .in2(_gnd_net_),
            .in3(N__62890),
            .lcout(rco_c_87),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_86_LC_14_4_5.C_ON=1'b0;
    defparam rco_obuf_RNO_86_LC_14_4_5.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_86_LC_14_4_5.LUT_INIT=16'b1100110000000000;
    LogicCell40 rco_obuf_RNO_86_LC_14_4_5 (
            .in0(_gnd_net_),
            .in1(N__62889),
            .in2(_gnd_net_),
            .in3(N__68505),
            .lcout(rco_c_86),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_90_0_LC_14_5_0.C_ON=1'b0;
    defparam shift_srl_90_0_LC_14_5_0.SEQ_MODE=4'b1000;
    defparam shift_srl_90_0_LC_14_5_0.LUT_INIT=16'b1100110011001100;
    LogicCell40 shift_srl_90_0_LC_14_5_0 (
            .in0(_gnd_net_),
            .in1(N__66894),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_90Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93242),
            .ce(N__61227),
            .sr(_gnd_net_));
    defparam shift_srl_90_1_LC_14_5_1.C_ON=1'b0;
    defparam shift_srl_90_1_LC_14_5_1.SEQ_MODE=4'b1000;
    defparam shift_srl_90_1_LC_14_5_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_90_1_LC_14_5_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61186),
            .lcout(shift_srl_90Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93242),
            .ce(N__61227),
            .sr(_gnd_net_));
    defparam shift_srl_90_2_LC_14_5_2.C_ON=1'b0;
    defparam shift_srl_90_2_LC_14_5_2.SEQ_MODE=4'b1000;
    defparam shift_srl_90_2_LC_14_5_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_90_2_LC_14_5_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61180),
            .lcout(shift_srl_90Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93242),
            .ce(N__61227),
            .sr(_gnd_net_));
    defparam shift_srl_90_3_LC_14_5_3.C_ON=1'b0;
    defparam shift_srl_90_3_LC_14_5_3.SEQ_MODE=4'b1000;
    defparam shift_srl_90_3_LC_14_5_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_90_3_LC_14_5_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61174),
            .lcout(shift_srl_90Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93242),
            .ce(N__61227),
            .sr(_gnd_net_));
    defparam shift_srl_90_4_LC_14_5_4.C_ON=1'b0;
    defparam shift_srl_90_4_LC_14_5_4.SEQ_MODE=4'b1000;
    defparam shift_srl_90_4_LC_14_5_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_90_4_LC_14_5_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61168),
            .lcout(shift_srl_90Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93242),
            .ce(N__61227),
            .sr(_gnd_net_));
    defparam shift_srl_90_5_LC_14_5_5.C_ON=1'b0;
    defparam shift_srl_90_5_LC_14_5_5.SEQ_MODE=4'b1000;
    defparam shift_srl_90_5_LC_14_5_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_90_5_LC_14_5_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61162),
            .lcout(shift_srl_90Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93242),
            .ce(N__61227),
            .sr(_gnd_net_));
    defparam shift_srl_90_RNITV4VM_15_LC_14_6_0.C_ON=1'b0;
    defparam shift_srl_90_RNITV4VM_15_LC_14_6_0.SEQ_MODE=4'b0000;
    defparam shift_srl_90_RNITV4VM_15_LC_14_6_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_90_RNITV4VM_15_LC_14_6_0 (
            .in0(N__68477),
            .in1(N__89458),
            .in2(N__66904),
            .in3(N__68609),
            .lcout(clk_en_91),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_90_15_LC_14_6_1.C_ON=1'b0;
    defparam shift_srl_90_15_LC_14_6_1.SEQ_MODE=4'b1000;
    defparam shift_srl_90_15_LC_14_6_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_90_15_LC_14_6_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61258),
            .lcout(shift_srl_90Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93224),
            .ce(N__61226),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNI98ETM_15_LC_14_6_3.C_ON=1'b0;
    defparam shift_srl_0_RNI98ETM_15_LC_14_6_3.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNI98ETM_15_LC_14_6_3.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_0_RNI98ETM_15_LC_14_6_3 (
            .in0(N__68608),
            .in1(N__89459),
            .in2(_gnd_net_),
            .in3(N__68478),
            .lcout(clk_en_90),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_90_14_LC_14_6_4.C_ON=1'b0;
    defparam shift_srl_90_14_LC_14_6_4.SEQ_MODE=4'b1000;
    defparam shift_srl_90_14_LC_14_6_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_90_14_LC_14_6_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61252),
            .lcout(shift_srl_90Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93224),
            .ce(N__61226),
            .sr(_gnd_net_));
    defparam shift_srl_90_13_LC_14_6_5.C_ON=1'b0;
    defparam shift_srl_90_13_LC_14_6_5.SEQ_MODE=4'b1000;
    defparam shift_srl_90_13_LC_14_6_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_90_13_LC_14_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61246),
            .lcout(shift_srl_90Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93224),
            .ce(N__61226),
            .sr(_gnd_net_));
    defparam shift_srl_90_12_LC_14_6_6.C_ON=1'b0;
    defparam shift_srl_90_12_LC_14_6_6.SEQ_MODE=4'b1000;
    defparam shift_srl_90_12_LC_14_6_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_90_12_LC_14_6_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61234),
            .lcout(shift_srl_90Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93224),
            .ce(N__61226),
            .sr(_gnd_net_));
    defparam shift_srl_90_11_LC_14_6_7.C_ON=1'b0;
    defparam shift_srl_90_11_LC_14_6_7.SEQ_MODE=4'b1000;
    defparam shift_srl_90_11_LC_14_6_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_90_11_LC_14_6_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61240),
            .lcout(shift_srl_90Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93224),
            .ce(N__61226),
            .sr(_gnd_net_));
    defparam shift_srl_87_10_LC_14_7_0.C_ON=1'b0;
    defparam shift_srl_87_10_LC_14_7_0.SEQ_MODE=4'b1000;
    defparam shift_srl_87_10_LC_14_7_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_87_10_LC_14_7_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61300),
            .lcout(shift_srl_87Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93204),
            .ce(N__64410),
            .sr(_gnd_net_));
    defparam shift_srl_87_11_LC_14_7_1.C_ON=1'b0;
    defparam shift_srl_87_11_LC_14_7_1.SEQ_MODE=4'b1000;
    defparam shift_srl_87_11_LC_14_7_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_87_11_LC_14_7_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61210),
            .lcout(shift_srl_87Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93204),
            .ce(N__64410),
            .sr(_gnd_net_));
    defparam shift_srl_87_12_LC_14_7_2.C_ON=1'b0;
    defparam shift_srl_87_12_LC_14_7_2.SEQ_MODE=4'b1000;
    defparam shift_srl_87_12_LC_14_7_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_87_12_LC_14_7_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61204),
            .lcout(shift_srl_87Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93204),
            .ce(N__64410),
            .sr(_gnd_net_));
    defparam shift_srl_87_13_LC_14_7_3.C_ON=1'b0;
    defparam shift_srl_87_13_LC_14_7_3.SEQ_MODE=4'b1000;
    defparam shift_srl_87_13_LC_14_7_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_87_13_LC_14_7_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61198),
            .lcout(shift_srl_87Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93204),
            .ce(N__64410),
            .sr(_gnd_net_));
    defparam shift_srl_87_14_LC_14_7_4.C_ON=1'b0;
    defparam shift_srl_87_14_LC_14_7_4.SEQ_MODE=4'b1000;
    defparam shift_srl_87_14_LC_14_7_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_87_14_LC_14_7_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61192),
            .lcout(shift_srl_87Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93204),
            .ce(N__64410),
            .sr(_gnd_net_));
    defparam shift_srl_87_15_LC_14_7_5.C_ON=1'b0;
    defparam shift_srl_87_15_LC_14_7_5.SEQ_MODE=4'b1000;
    defparam shift_srl_87_15_LC_14_7_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_87_15_LC_14_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61306),
            .lcout(shift_srl_87Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93204),
            .ce(N__64410),
            .sr(_gnd_net_));
    defparam shift_srl_87_9_LC_14_7_6.C_ON=1'b0;
    defparam shift_srl_87_9_LC_14_7_6.SEQ_MODE=4'b1000;
    defparam shift_srl_87_9_LC_14_7_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_87_9_LC_14_7_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61294),
            .lcout(shift_srl_87Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93204),
            .ce(N__64410),
            .sr(_gnd_net_));
    defparam shift_srl_87_8_LC_14_7_7.C_ON=1'b0;
    defparam shift_srl_87_8_LC_14_7_7.SEQ_MODE=4'b1000;
    defparam shift_srl_87_8_LC_14_7_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_87_8_LC_14_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64420),
            .lcout(shift_srl_87Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93204),
            .ce(N__64410),
            .sr(_gnd_net_));
    defparam shift_srl_86_0_LC_14_8_0.C_ON=1'b0;
    defparam shift_srl_86_0_LC_14_8_0.SEQ_MODE=4'b1000;
    defparam shift_srl_86_0_LC_14_8_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_86_0_LC_14_8_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67143),
            .lcout(shift_srl_86Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93182),
            .ce(N__67170),
            .sr(_gnd_net_));
    defparam shift_srl_86_1_LC_14_8_1.C_ON=1'b0;
    defparam shift_srl_86_1_LC_14_8_1.SEQ_MODE=4'b1000;
    defparam shift_srl_86_1_LC_14_8_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_86_1_LC_14_8_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61288),
            .lcout(shift_srl_86Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93182),
            .ce(N__67170),
            .sr(_gnd_net_));
    defparam shift_srl_86_2_LC_14_8_2.C_ON=1'b0;
    defparam shift_srl_86_2_LC_14_8_2.SEQ_MODE=4'b1000;
    defparam shift_srl_86_2_LC_14_8_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_86_2_LC_14_8_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61282),
            .lcout(shift_srl_86Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93182),
            .ce(N__67170),
            .sr(_gnd_net_));
    defparam shift_srl_86_3_LC_14_8_3.C_ON=1'b0;
    defparam shift_srl_86_3_LC_14_8_3.SEQ_MODE=4'b1000;
    defparam shift_srl_86_3_LC_14_8_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_86_3_LC_14_8_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61276),
            .lcout(shift_srl_86Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93182),
            .ce(N__67170),
            .sr(_gnd_net_));
    defparam shift_srl_86_4_LC_14_8_4.C_ON=1'b0;
    defparam shift_srl_86_4_LC_14_8_4.SEQ_MODE=4'b1000;
    defparam shift_srl_86_4_LC_14_8_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_86_4_LC_14_8_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61270),
            .lcout(shift_srl_86Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93182),
            .ce(N__67170),
            .sr(_gnd_net_));
    defparam shift_srl_86_5_LC_14_8_5.C_ON=1'b0;
    defparam shift_srl_86_5_LC_14_8_5.SEQ_MODE=4'b1000;
    defparam shift_srl_86_5_LC_14_8_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_86_5_LC_14_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61264),
            .lcout(shift_srl_86Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93182),
            .ce(N__67170),
            .sr(_gnd_net_));
    defparam shift_srl_86_12_LC_14_8_6.C_ON=1'b0;
    defparam shift_srl_86_12_LC_14_8_6.SEQ_MODE=4'b1000;
    defparam shift_srl_86_12_LC_14_8_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_86_12_LC_14_8_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61354),
            .lcout(shift_srl_86Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93182),
            .ce(N__67170),
            .sr(_gnd_net_));
    defparam shift_srl_86_11_LC_14_8_7.C_ON=1'b0;
    defparam shift_srl_86_11_LC_14_8_7.SEQ_MODE=4'b1000;
    defparam shift_srl_86_11_LC_14_8_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_86_11_LC_14_8_7 (
            .in0(N__62845),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_86Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93182),
            .ce(N__67170),
            .sr(_gnd_net_));
    defparam shift_srl_84_0_LC_14_10_0.C_ON=1'b0;
    defparam shift_srl_84_0_LC_14_10_0.SEQ_MODE=4'b1000;
    defparam shift_srl_84_0_LC_14_10_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_84_0_LC_14_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68655),
            .lcout(shift_srl_84Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93144),
            .ce(N__61456),
            .sr(_gnd_net_));
    defparam shift_srl_84_1_LC_14_10_1.C_ON=1'b0;
    defparam shift_srl_84_1_LC_14_10_1.SEQ_MODE=4'b1000;
    defparam shift_srl_84_1_LC_14_10_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_84_1_LC_14_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61348),
            .lcout(shift_srl_84Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93144),
            .ce(N__61456),
            .sr(_gnd_net_));
    defparam shift_srl_84_2_LC_14_10_2.C_ON=1'b0;
    defparam shift_srl_84_2_LC_14_10_2.SEQ_MODE=4'b1000;
    defparam shift_srl_84_2_LC_14_10_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_84_2_LC_14_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61342),
            .lcout(shift_srl_84Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93144),
            .ce(N__61456),
            .sr(_gnd_net_));
    defparam shift_srl_84_3_LC_14_10_3.C_ON=1'b0;
    defparam shift_srl_84_3_LC_14_10_3.SEQ_MODE=4'b1000;
    defparam shift_srl_84_3_LC_14_10_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_84_3_LC_14_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61336),
            .lcout(shift_srl_84Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93144),
            .ce(N__61456),
            .sr(_gnd_net_));
    defparam shift_srl_84_4_LC_14_10_4.C_ON=1'b0;
    defparam shift_srl_84_4_LC_14_10_4.SEQ_MODE=4'b1000;
    defparam shift_srl_84_4_LC_14_10_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_84_4_LC_14_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61330),
            .lcout(shift_srl_84Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93144),
            .ce(N__61456),
            .sr(_gnd_net_));
    defparam shift_srl_84_5_LC_14_10_5.C_ON=1'b0;
    defparam shift_srl_84_5_LC_14_10_5.SEQ_MODE=4'b1000;
    defparam shift_srl_84_5_LC_14_10_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_84_5_LC_14_10_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61324),
            .lcout(shift_srl_84Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93144),
            .ce(N__61456),
            .sr(_gnd_net_));
    defparam shift_srl_84_6_LC_14_10_6.C_ON=1'b0;
    defparam shift_srl_84_6_LC_14_10_6.SEQ_MODE=4'b1000;
    defparam shift_srl_84_6_LC_14_10_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_84_6_LC_14_10_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61318),
            .lcout(shift_srl_84Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93144),
            .ce(N__61456),
            .sr(_gnd_net_));
    defparam shift_srl_84_7_LC_14_10_7.C_ON=1'b0;
    defparam shift_srl_84_7_LC_14_10_7.SEQ_MODE=4'b1000;
    defparam shift_srl_84_7_LC_14_10_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_84_7_LC_14_10_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61312),
            .lcout(shift_srl_84Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93144),
            .ce(N__61456),
            .sr(_gnd_net_));
    defparam shift_srl_84_10_LC_14_11_0.C_ON=1'b0;
    defparam shift_srl_84_10_LC_14_11_0.SEQ_MODE=4'b1000;
    defparam shift_srl_84_10_LC_14_11_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_84_10_LC_14_11_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61372),
            .lcout(shift_srl_84Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93124),
            .ce(N__61455),
            .sr(_gnd_net_));
    defparam shift_srl_84_11_LC_14_11_1.C_ON=1'b0;
    defparam shift_srl_84_11_LC_14_11_1.SEQ_MODE=4'b1000;
    defparam shift_srl_84_11_LC_14_11_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_84_11_LC_14_11_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61402),
            .lcout(shift_srl_84Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93124),
            .ce(N__61455),
            .sr(_gnd_net_));
    defparam shift_srl_84_12_LC_14_11_2.C_ON=1'b0;
    defparam shift_srl_84_12_LC_14_11_2.SEQ_MODE=4'b1000;
    defparam shift_srl_84_12_LC_14_11_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_84_12_LC_14_11_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61396),
            .lcout(shift_srl_84Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93124),
            .ce(N__61455),
            .sr(_gnd_net_));
    defparam shift_srl_84_13_LC_14_11_3.C_ON=1'b0;
    defparam shift_srl_84_13_LC_14_11_3.SEQ_MODE=4'b1000;
    defparam shift_srl_84_13_LC_14_11_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_84_13_LC_14_11_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61390),
            .lcout(shift_srl_84Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93124),
            .ce(N__61455),
            .sr(_gnd_net_));
    defparam shift_srl_84_14_LC_14_11_4.C_ON=1'b0;
    defparam shift_srl_84_14_LC_14_11_4.SEQ_MODE=4'b1000;
    defparam shift_srl_84_14_LC_14_11_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_84_14_LC_14_11_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61384),
            .lcout(shift_srl_84Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93124),
            .ce(N__61455),
            .sr(_gnd_net_));
    defparam shift_srl_84_15_LC_14_11_5.C_ON=1'b0;
    defparam shift_srl_84_15_LC_14_11_5.SEQ_MODE=4'b1000;
    defparam shift_srl_84_15_LC_14_11_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_84_15_LC_14_11_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61378),
            .lcout(shift_srl_84Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93124),
            .ce(N__61455),
            .sr(_gnd_net_));
    defparam shift_srl_84_9_LC_14_11_6.C_ON=1'b0;
    defparam shift_srl_84_9_LC_14_11_6.SEQ_MODE=4'b1000;
    defparam shift_srl_84_9_LC_14_11_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_84_9_LC_14_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61360),
            .lcout(shift_srl_84Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93124),
            .ce(N__61455),
            .sr(_gnd_net_));
    defparam shift_srl_84_8_LC_14_11_7.C_ON=1'b0;
    defparam shift_srl_84_8_LC_14_11_7.SEQ_MODE=4'b1000;
    defparam shift_srl_84_8_LC_14_11_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_84_8_LC_14_11_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61366),
            .lcout(shift_srl_84Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93124),
            .ce(N__61455),
            .sr(_gnd_net_));
    defparam shift_srl_89_RNI5GFS_15_LC_14_12_0.C_ON=1'b0;
    defparam shift_srl_89_RNI5GFS_15_LC_14_12_0.SEQ_MODE=4'b0000;
    defparam shift_srl_89_RNI5GFS_15_LC_14_12_0.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_89_RNI5GFS_15_LC_14_12_0 (
            .in0(N__67104),
            .in1(N__67007),
            .in2(N__66915),
            .in3(N__66986),
            .lcout(),
            .ltout(rco_int_0_a2_0_a2_0_sx_91_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_91_RNI20EN1_15_LC_14_12_1.C_ON=1'b0;
    defparam shift_srl_91_RNI20EN1_15_LC_14_12_1.SEQ_MODE=4'b0000;
    defparam shift_srl_91_RNI20EN1_15_LC_14_12_1.LUT_INIT=16'b0000110000000000;
    LogicCell40 shift_srl_91_RNI20EN1_15_LC_14_12_1 (
            .in0(_gnd_net_),
            .in1(N__66945),
            .in2(N__61465),
            .in3(N__62858),
            .lcout(shift_srl_91_RNI20EN1Z0Z_15),
            .ltout(shift_srl_91_RNI20EN1Z0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_145_RNI4T7BG_15_LC_14_12_2.C_ON=1'b0;
    defparam shift_srl_145_RNI4T7BG_15_LC_14_12_2.SEQ_MODE=4'b0000;
    defparam shift_srl_145_RNI4T7BG_15_LC_14_12_2.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_145_RNI4T7BG_15_LC_14_12_2 (
            .in0(N__82312),
            .in1(N__71983),
            .in2(N__61462),
            .in3(N__72028),
            .lcout(rco_int_0_a2_0_a2_sx_1_153),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_83_RNIKTI68_15_LC_14_12_3.C_ON=1'b0;
    defparam shift_srl_83_RNIKTI68_15_LC_14_12_3.SEQ_MODE=4'b0000;
    defparam shift_srl_83_RNIKTI68_15_LC_14_12_3.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_83_RNIKTI68_15_LC_14_12_3 (
            .in0(N__73068),
            .in1(N__86816),
            .in2(_gnd_net_),
            .in3(N__80785),
            .lcout(),
            .ltout(shift_srl_83_RNIKTI68Z0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIGRJDL_15_LC_14_12_4.C_ON=1'b0;
    defparam shift_srl_0_RNIGRJDL_15_LC_14_12_4.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIGRJDL_15_LC_14_12_4.LUT_INIT=16'b0000000011000000;
    LogicCell40 shift_srl_0_RNIGRJDL_15_LC_14_12_4 (
            .in0(_gnd_net_),
            .in1(N__90425),
            .in2(N__61459),
            .in3(N__67354),
            .lcout(clk_en_84),
            .ltout(clk_en_84_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_88_RNIDHAGM_15_LC_14_12_5.C_ON=1'b0;
    defparam shift_srl_88_RNIDHAGM_15_LC_14_12_5.SEQ_MODE=4'b0000;
    defparam shift_srl_88_RNIDHAGM_15_LC_14_12_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_88_RNIDHAGM_15_LC_14_12_5 (
            .in0(N__66987),
            .in1(N__67105),
            .in2(N__61438),
            .in3(N__62859),
            .lcout(clk_en_89),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_86_RNI8K1L_15_LC_14_12_6.C_ON=1'b0;
    defparam shift_srl_86_RNI8K1L_15_LC_14_12_6.SEQ_MODE=4'b0000;
    defparam shift_srl_86_RNI8K1L_15_LC_14_12_6.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_86_RNI8K1L_15_LC_14_12_6 (
            .in0(N__67061),
            .in1(N__67144),
            .in2(_gnd_net_),
            .in3(N__68647),
            .lcout(shift_srl_86_RNI8K1LZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_89_15_LC_14_12_7.C_ON=1'b0;
    defparam shift_srl_89_15_LC_14_12_7.SEQ_MODE=4'b1000;
    defparam shift_srl_89_15_LC_14_12_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_89_15_LC_14_12_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61435),
            .lcout(shift_srl_89Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93106),
            .ce(N__61424),
            .sr(_gnd_net_));
    defparam shift_srl_24_7_LC_14_13_0.C_ON=1'b0;
    defparam shift_srl_24_7_LC_14_13_0.SEQ_MODE=4'b1000;
    defparam shift_srl_24_7_LC_14_13_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_24_7_LC_14_13_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61507),
            .lcout(shift_srl_24Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93091),
            .ce(N__63149),
            .sr(_gnd_net_));
    defparam shift_srl_24_5_LC_14_13_3.C_ON=1'b0;
    defparam shift_srl_24_5_LC_14_13_3.SEQ_MODE=4'b1000;
    defparam shift_srl_24_5_LC_14_13_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_24_5_LC_14_13_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61525),
            .lcout(shift_srl_24Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93091),
            .ce(N__63149),
            .sr(_gnd_net_));
    defparam shift_srl_24_4_LC_14_13_5.C_ON=1'b0;
    defparam shift_srl_24_4_LC_14_13_5.SEQ_MODE=4'b1000;
    defparam shift_srl_24_4_LC_14_13_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_24_4_LC_14_13_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61531),
            .lcout(shift_srl_24Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93091),
            .ce(N__63149),
            .sr(_gnd_net_));
    defparam shift_srl_24_8_LC_14_13_6.C_ON=1'b0;
    defparam shift_srl_24_8_LC_14_13_6.SEQ_MODE=4'b1000;
    defparam shift_srl_24_8_LC_14_13_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_24_8_LC_14_13_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61519),
            .lcout(shift_srl_24Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93091),
            .ce(N__63149),
            .sr(_gnd_net_));
    defparam shift_srl_24_6_LC_14_13_7.C_ON=1'b0;
    defparam shift_srl_24_6_LC_14_13_7.SEQ_MODE=4'b1000;
    defparam shift_srl_24_6_LC_14_13_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_24_6_LC_14_13_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61513),
            .lcout(shift_srl_24Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93091),
            .ce(N__63149),
            .sr(_gnd_net_));
    defparam shift_srl_152_10_LC_14_14_0.C_ON=1'b0;
    defparam shift_srl_152_10_LC_14_14_0.SEQ_MODE=4'b1000;
    defparam shift_srl_152_10_LC_14_14_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_152_10_LC_14_14_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61471),
            .lcout(shift_srl_152Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93076),
            .ce(N__63193),
            .sr(_gnd_net_));
    defparam shift_srl_152_11_LC_14_14_1.C_ON=1'b0;
    defparam shift_srl_152_11_LC_14_14_1.SEQ_MODE=4'b1000;
    defparam shift_srl_152_11_LC_14_14_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_152_11_LC_14_14_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61501),
            .lcout(shift_srl_152Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93076),
            .ce(N__63193),
            .sr(_gnd_net_));
    defparam shift_srl_152_12_LC_14_14_2.C_ON=1'b0;
    defparam shift_srl_152_12_LC_14_14_2.SEQ_MODE=4'b1000;
    defparam shift_srl_152_12_LC_14_14_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_152_12_LC_14_14_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61495),
            .lcout(shift_srl_152Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93076),
            .ce(N__63193),
            .sr(_gnd_net_));
    defparam shift_srl_152_13_LC_14_14_3.C_ON=1'b0;
    defparam shift_srl_152_13_LC_14_14_3.SEQ_MODE=4'b1000;
    defparam shift_srl_152_13_LC_14_14_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_152_13_LC_14_14_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61489),
            .lcout(shift_srl_152Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93076),
            .ce(N__63193),
            .sr(_gnd_net_));
    defparam shift_srl_152_14_LC_14_14_4.C_ON=1'b0;
    defparam shift_srl_152_14_LC_14_14_4.SEQ_MODE=4'b1000;
    defparam shift_srl_152_14_LC_14_14_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_152_14_LC_14_14_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61483),
            .lcout(shift_srl_152Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93076),
            .ce(N__63193),
            .sr(_gnd_net_));
    defparam shift_srl_152_15_LC_14_14_5.C_ON=1'b0;
    defparam shift_srl_152_15_LC_14_14_5.SEQ_MODE=4'b1000;
    defparam shift_srl_152_15_LC_14_14_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_152_15_LC_14_14_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61477),
            .lcout(shift_srl_152Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93076),
            .ce(N__63193),
            .sr(_gnd_net_));
    defparam shift_srl_152_9_LC_14_14_6.C_ON=1'b0;
    defparam shift_srl_152_9_LC_14_14_6.SEQ_MODE=4'b1000;
    defparam shift_srl_152_9_LC_14_14_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_152_9_LC_14_14_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61579),
            .lcout(shift_srl_152Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93076),
            .ce(N__63193),
            .sr(_gnd_net_));
    defparam shift_srl_152_8_LC_14_14_7.C_ON=1'b0;
    defparam shift_srl_152_8_LC_14_14_7.SEQ_MODE=4'b1000;
    defparam shift_srl_152_8_LC_14_14_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_152_8_LC_14_14_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63082),
            .lcout(shift_srl_152Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93076),
            .ce(N__63193),
            .sr(_gnd_net_));
    defparam shift_srl_153_10_LC_14_15_0.C_ON=1'b0;
    defparam shift_srl_153_10_LC_14_15_0.SEQ_MODE=4'b1000;
    defparam shift_srl_153_10_LC_14_15_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_153_10_LC_14_15_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61543),
            .lcout(shift_srl_153Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93060),
            .ce(N__63210),
            .sr(_gnd_net_));
    defparam shift_srl_153_11_LC_14_15_1.C_ON=1'b0;
    defparam shift_srl_153_11_LC_14_15_1.SEQ_MODE=4'b1000;
    defparam shift_srl_153_11_LC_14_15_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_153_11_LC_14_15_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61573),
            .lcout(shift_srl_153Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93060),
            .ce(N__63210),
            .sr(_gnd_net_));
    defparam shift_srl_153_12_LC_14_15_2.C_ON=1'b0;
    defparam shift_srl_153_12_LC_14_15_2.SEQ_MODE=4'b1000;
    defparam shift_srl_153_12_LC_14_15_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_153_12_LC_14_15_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61567),
            .lcout(shift_srl_153Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93060),
            .ce(N__63210),
            .sr(_gnd_net_));
    defparam shift_srl_153_13_LC_14_15_3.C_ON=1'b0;
    defparam shift_srl_153_13_LC_14_15_3.SEQ_MODE=4'b1000;
    defparam shift_srl_153_13_LC_14_15_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_153_13_LC_14_15_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61561),
            .lcout(shift_srl_153Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93060),
            .ce(N__63210),
            .sr(_gnd_net_));
    defparam shift_srl_153_14_LC_14_15_4.C_ON=1'b0;
    defparam shift_srl_153_14_LC_14_15_4.SEQ_MODE=4'b1000;
    defparam shift_srl_153_14_LC_14_15_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_153_14_LC_14_15_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61555),
            .lcout(shift_srl_153Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93060),
            .ce(N__63210),
            .sr(_gnd_net_));
    defparam shift_srl_153_15_LC_14_15_5.C_ON=1'b0;
    defparam shift_srl_153_15_LC_14_15_5.SEQ_MODE=4'b1000;
    defparam shift_srl_153_15_LC_14_15_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_153_15_LC_14_15_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61549),
            .lcout(shift_srl_153Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93060),
            .ce(N__63210),
            .sr(_gnd_net_));
    defparam shift_srl_153_9_LC_14_15_6.C_ON=1'b0;
    defparam shift_srl_153_9_LC_14_15_6.SEQ_MODE=4'b1000;
    defparam shift_srl_153_9_LC_14_15_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_153_9_LC_14_15_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61537),
            .lcout(shift_srl_153Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93060),
            .ce(N__63210),
            .sr(_gnd_net_));
    defparam shift_srl_153_8_LC_14_15_7.C_ON=1'b0;
    defparam shift_srl_153_8_LC_14_15_7.SEQ_MODE=4'b1000;
    defparam shift_srl_153_8_LC_14_15_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_153_8_LC_14_15_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61585),
            .lcout(shift_srl_153Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93060),
            .ce(N__63210),
            .sr(_gnd_net_));
    defparam shift_srl_153_0_LC_14_16_0.C_ON=1'b0;
    defparam shift_srl_153_0_LC_14_16_0.SEQ_MODE=4'b1000;
    defparam shift_srl_153_0_LC_14_16_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_153_0_LC_14_16_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61641),
            .lcout(shift_srl_153Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93045),
            .ce(N__63211),
            .sr(_gnd_net_));
    defparam shift_srl_153_1_LC_14_16_1.C_ON=1'b0;
    defparam shift_srl_153_1_LC_14_16_1.SEQ_MODE=4'b1000;
    defparam shift_srl_153_1_LC_14_16_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_153_1_LC_14_16_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61627),
            .lcout(shift_srl_153Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93045),
            .ce(N__63211),
            .sr(_gnd_net_));
    defparam shift_srl_153_2_LC_14_16_2.C_ON=1'b0;
    defparam shift_srl_153_2_LC_14_16_2.SEQ_MODE=4'b1000;
    defparam shift_srl_153_2_LC_14_16_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_153_2_LC_14_16_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61621),
            .lcout(shift_srl_153Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93045),
            .ce(N__63211),
            .sr(_gnd_net_));
    defparam shift_srl_153_3_LC_14_16_3.C_ON=1'b0;
    defparam shift_srl_153_3_LC_14_16_3.SEQ_MODE=4'b1000;
    defparam shift_srl_153_3_LC_14_16_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_153_3_LC_14_16_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61615),
            .lcout(shift_srl_153Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93045),
            .ce(N__63211),
            .sr(_gnd_net_));
    defparam shift_srl_153_4_LC_14_16_4.C_ON=1'b0;
    defparam shift_srl_153_4_LC_14_16_4.SEQ_MODE=4'b1000;
    defparam shift_srl_153_4_LC_14_16_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_153_4_LC_14_16_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61609),
            .lcout(shift_srl_153Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93045),
            .ce(N__63211),
            .sr(_gnd_net_));
    defparam shift_srl_153_5_LC_14_16_5.C_ON=1'b0;
    defparam shift_srl_153_5_LC_14_16_5.SEQ_MODE=4'b1000;
    defparam shift_srl_153_5_LC_14_16_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_153_5_LC_14_16_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61603),
            .lcout(shift_srl_153Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93045),
            .ce(N__63211),
            .sr(_gnd_net_));
    defparam shift_srl_153_6_LC_14_16_6.C_ON=1'b0;
    defparam shift_srl_153_6_LC_14_16_6.SEQ_MODE=4'b1000;
    defparam shift_srl_153_6_LC_14_16_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_153_6_LC_14_16_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61597),
            .lcout(shift_srl_153Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93045),
            .ce(N__63211),
            .sr(_gnd_net_));
    defparam shift_srl_153_7_LC_14_16_7.C_ON=1'b0;
    defparam shift_srl_153_7_LC_14_16_7.SEQ_MODE=4'b1000;
    defparam shift_srl_153_7_LC_14_16_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_153_7_LC_14_16_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61591),
            .lcout(shift_srl_153Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93045),
            .ce(N__63211),
            .sr(_gnd_net_));
    defparam shift_srl_141_10_LC_14_17_0.C_ON=1'b0;
    defparam shift_srl_141_10_LC_14_17_0.SEQ_MODE=4'b1000;
    defparam shift_srl_141_10_LC_14_17_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_141_10_LC_14_17_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61681),
            .lcout(shift_srl_141Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93023),
            .ce(N__62041),
            .sr(_gnd_net_));
    defparam shift_srl_141_11_LC_14_17_1.C_ON=1'b0;
    defparam shift_srl_141_11_LC_14_17_1.SEQ_MODE=4'b1000;
    defparam shift_srl_141_11_LC_14_17_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_141_11_LC_14_17_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61699),
            .lcout(shift_srl_141Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93023),
            .ce(N__62041),
            .sr(_gnd_net_));
    defparam shift_srl_141_12_LC_14_17_2.C_ON=1'b0;
    defparam shift_srl_141_12_LC_14_17_2.SEQ_MODE=4'b1000;
    defparam shift_srl_141_12_LC_14_17_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_141_12_LC_14_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61693),
            .lcout(shift_srl_141Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93023),
            .ce(N__62041),
            .sr(_gnd_net_));
    defparam shift_srl_141_13_LC_14_17_3.C_ON=1'b0;
    defparam shift_srl_141_13_LC_14_17_3.SEQ_MODE=4'b1000;
    defparam shift_srl_141_13_LC_14_17_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_141_13_LC_14_17_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61687),
            .lcout(shift_srl_141Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93023),
            .ce(N__62041),
            .sr(_gnd_net_));
    defparam shift_srl_141_7_LC_14_17_4.C_ON=1'b0;
    defparam shift_srl_141_7_LC_14_17_4.SEQ_MODE=4'b1000;
    defparam shift_srl_141_7_LC_14_17_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_141_7_LC_14_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61651),
            .lcout(shift_srl_141Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93023),
            .ce(N__62041),
            .sr(_gnd_net_));
    defparam shift_srl_141_9_LC_14_17_5.C_ON=1'b0;
    defparam shift_srl_141_9_LC_14_17_5.SEQ_MODE=4'b1000;
    defparam shift_srl_141_9_LC_14_17_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_141_9_LC_14_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61669),
            .lcout(shift_srl_141Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93023),
            .ce(N__62041),
            .sr(_gnd_net_));
    defparam shift_srl_141_8_LC_14_17_6.C_ON=1'b0;
    defparam shift_srl_141_8_LC_14_17_6.SEQ_MODE=4'b1000;
    defparam shift_srl_141_8_LC_14_17_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_141_8_LC_14_17_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61675),
            .lcout(shift_srl_141Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93023),
            .ce(N__62041),
            .sr(_gnd_net_));
    defparam shift_srl_141_4_LC_14_18_0.C_ON=1'b0;
    defparam shift_srl_141_4_LC_14_18_0.SEQ_MODE=4'b1000;
    defparam shift_srl_141_4_LC_14_18_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_141_4_LC_14_18_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61834),
            .lcout(shift_srl_141Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93046),
            .ce(N__62036),
            .sr(_gnd_net_));
    defparam shift_srl_141_5_LC_14_18_1.C_ON=1'b0;
    defparam shift_srl_141_5_LC_14_18_1.SEQ_MODE=4'b1000;
    defparam shift_srl_141_5_LC_14_18_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_141_5_LC_14_18_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61663),
            .lcout(shift_srl_141Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93046),
            .ce(N__62036),
            .sr(_gnd_net_));
    defparam shift_srl_141_6_LC_14_18_2.C_ON=1'b0;
    defparam shift_srl_141_6_LC_14_18_2.SEQ_MODE=4'b1000;
    defparam shift_srl_141_6_LC_14_18_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_141_6_LC_14_18_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61657),
            .lcout(shift_srl_141Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93046),
            .ce(N__62036),
            .sr(_gnd_net_));
    defparam shift_srl_141_3_LC_14_18_3.C_ON=1'b0;
    defparam shift_srl_141_3_LC_14_18_3.SEQ_MODE=4'b1000;
    defparam shift_srl_141_3_LC_14_18_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_141_3_LC_14_18_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61705),
            .lcout(shift_srl_141Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93046),
            .ce(N__62036),
            .sr(_gnd_net_));
    defparam shift_srl_141_14_LC_14_18_6.C_ON=1'b0;
    defparam shift_srl_141_14_LC_14_18_6.SEQ_MODE=4'b1000;
    defparam shift_srl_141_14_LC_14_18_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_141_14_LC_14_18_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61828),
            .lcout(shift_srl_141Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93046),
            .ce(N__62036),
            .sr(_gnd_net_));
    defparam shift_srl_141_RNIBN961_15_LC_14_19_0.C_ON=1'b0;
    defparam shift_srl_141_RNIBN961_15_LC_14_19_0.SEQ_MODE=4'b0000;
    defparam shift_srl_141_RNIBN961_15_LC_14_19_0.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_141_RNIBN961_15_LC_14_19_0 (
            .in0(N__88102),
            .in1(N__63754),
            .in2(N__61735),
            .in3(N__64877),
            .lcout(),
            .ltout(rco_int_0_a2_0_a2_0_sx_144_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_144_RNIIPPI1_15_LC_14_19_1.C_ON=1'b0;
    defparam shift_srl_144_RNIIPPI1_15_LC_14_19_1.SEQ_MODE=4'b0000;
    defparam shift_srl_144_RNIIPPI1_15_LC_14_19_1.LUT_INIT=16'b0000110000000000;
    LogicCell40 shift_srl_144_RNIIPPI1_15_LC_14_19_1 (
            .in0(_gnd_net_),
            .in1(N__61822),
            .in2(N__61795),
            .in3(N__61776),
            .lcout(shift_srl_144_RNIIPPI1Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_141_15_LC_14_19_2.C_ON=1'b0;
    defparam shift_srl_141_15_LC_14_19_2.SEQ_MODE=4'b1000;
    defparam shift_srl_141_15_LC_14_19_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_141_15_LC_14_19_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61741),
            .lcout(shift_srl_141Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93061),
            .ce(N__62037),
            .sr(_gnd_net_));
    defparam shift_srl_141_RNI9SAM_15_LC_14_19_3.C_ON=1'b0;
    defparam shift_srl_141_RNI9SAM_15_LC_14_19_3.SEQ_MODE=4'b0000;
    defparam shift_srl_141_RNI9SAM_15_LC_14_19_3.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_141_RNI9SAM_15_LC_14_19_3 (
            .in0(N__61730),
            .in1(N__88101),
            .in2(_gnd_net_),
            .in3(N__64876),
            .lcout(shift_srl_141_RNI9SAMZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_141_0_LC_14_19_4.C_ON=1'b0;
    defparam shift_srl_141_0_LC_14_19_4.SEQ_MODE=4'b1000;
    defparam shift_srl_141_0_LC_14_19_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_141_0_LC_14_19_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61731),
            .lcout(shift_srl_141Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93061),
            .ce(N__62037),
            .sr(_gnd_net_));
    defparam shift_srl_141_1_LC_14_19_5.C_ON=1'b0;
    defparam shift_srl_141_1_LC_14_19_5.SEQ_MODE=4'b1000;
    defparam shift_srl_141_1_LC_14_19_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_141_1_LC_14_19_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61717),
            .lcout(shift_srl_141Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93061),
            .ce(N__62037),
            .sr(_gnd_net_));
    defparam shift_srl_141_2_LC_14_19_6.C_ON=1'b0;
    defparam shift_srl_141_2_LC_14_19_6.SEQ_MODE=4'b1000;
    defparam shift_srl_141_2_LC_14_19_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_141_2_LC_14_19_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61711),
            .lcout(shift_srl_141Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93061),
            .ce(N__62037),
            .sr(_gnd_net_));
    defparam shift_srl_145_10_LC_14_20_0.C_ON=1'b0;
    defparam shift_srl_145_10_LC_14_20_0.SEQ_MODE=4'b1000;
    defparam shift_srl_145_10_LC_14_20_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_145_10_LC_14_20_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61849),
            .lcout(shift_srl_145Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93077),
            .ce(N__63513),
            .sr(_gnd_net_));
    defparam shift_srl_145_11_LC_14_20_1.C_ON=1'b0;
    defparam shift_srl_145_11_LC_14_20_1.SEQ_MODE=4'b1000;
    defparam shift_srl_145_11_LC_14_20_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_145_11_LC_14_20_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61879),
            .lcout(shift_srl_145Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93077),
            .ce(N__63513),
            .sr(_gnd_net_));
    defparam shift_srl_145_12_LC_14_20_2.C_ON=1'b0;
    defparam shift_srl_145_12_LC_14_20_2.SEQ_MODE=4'b1000;
    defparam shift_srl_145_12_LC_14_20_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_145_12_LC_14_20_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61873),
            .lcout(shift_srl_145Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93077),
            .ce(N__63513),
            .sr(_gnd_net_));
    defparam shift_srl_145_13_LC_14_20_3.C_ON=1'b0;
    defparam shift_srl_145_13_LC_14_20_3.SEQ_MODE=4'b1000;
    defparam shift_srl_145_13_LC_14_20_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_145_13_LC_14_20_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61867),
            .lcout(shift_srl_145Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93077),
            .ce(N__63513),
            .sr(_gnd_net_));
    defparam shift_srl_145_14_LC_14_20_4.C_ON=1'b0;
    defparam shift_srl_145_14_LC_14_20_4.SEQ_MODE=4'b1000;
    defparam shift_srl_145_14_LC_14_20_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_145_14_LC_14_20_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61861),
            .lcout(shift_srl_145Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93077),
            .ce(N__63513),
            .sr(_gnd_net_));
    defparam shift_srl_145_15_LC_14_20_5.C_ON=1'b0;
    defparam shift_srl_145_15_LC_14_20_5.SEQ_MODE=4'b1000;
    defparam shift_srl_145_15_LC_14_20_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_145_15_LC_14_20_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61855),
            .lcout(shift_srl_145Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93077),
            .ce(N__63513),
            .sr(_gnd_net_));
    defparam shift_srl_145_9_LC_14_20_6.C_ON=1'b0;
    defparam shift_srl_145_9_LC_14_20_6.SEQ_MODE=4'b1000;
    defparam shift_srl_145_9_LC_14_20_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_145_9_LC_14_20_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61843),
            .lcout(shift_srl_145Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93077),
            .ce(N__63513),
            .sr(_gnd_net_));
    defparam shift_srl_145_8_LC_14_20_7.C_ON=1'b0;
    defparam shift_srl_145_8_LC_14_20_7.SEQ_MODE=4'b1000;
    defparam shift_srl_145_8_LC_14_20_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_145_8_LC_14_20_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63520),
            .lcout(shift_srl_145Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93077),
            .ce(N__63513),
            .sr(_gnd_net_));
    defparam shift_srl_120_RNIGK6F3_15_LC_14_21_0.C_ON=1'b0;
    defparam shift_srl_120_RNIGK6F3_15_LC_14_21_0.SEQ_MODE=4'b0000;
    defparam shift_srl_120_RNIGK6F3_15_LC_14_21_0.LUT_INIT=16'b1110111000100010;
    LogicCell40 shift_srl_120_RNIGK6F3_15_LC_14_21_0 (
            .in0(_gnd_net_),
            .in1(N__65358),
            .in2(_gnd_net_),
            .in3(N__61897),
            .lcout(rco_int_0_a3_0_a2_138_m6_0_a2_7_4),
            .ltout(rco_int_0_a3_0_a2_138_m6_0_a2_7_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_138_RNIJHHQ6_15_LC_14_21_1.C_ON=1'b0;
    defparam shift_srl_138_RNIJHHQ6_15_LC_14_21_1.SEQ_MODE=4'b0000;
    defparam shift_srl_138_RNIJHHQ6_15_LC_14_21_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_138_RNIJHHQ6_15_LC_14_21_1 (
            .in0(N__65709),
            .in1(N__62182),
            .in2(N__61837),
            .in3(N__62134),
            .lcout(rco_int_0_a3_0_a2_138_m6_0_a2_7),
            .ltout(rco_int_0_a3_0_a2_138_m6_0_a2_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_139_RNI8ON031_15_LC_14_21_2.C_ON=1'b0;
    defparam shift_srl_139_RNI8ON031_15_LC_14_21_2.SEQ_MODE=4'b0000;
    defparam shift_srl_139_RNI8ON031_15_LC_14_21_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_139_RNI8ON031_15_LC_14_21_2 (
            .in0(N__90344),
            .in1(N__88112),
            .in2(N__62044),
            .in3(N__61972),
            .lcout(N_124_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNI8BA831_15_LC_14_21_3.C_ON=1'b0;
    defparam shift_srl_0_RNI8BA831_15_LC_14_21_3.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNI8BA831_15_LC_14_21_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNI8BA831_15_LC_14_21_3 (
            .in0(N__61971),
            .in1(N__90345),
            .in2(N__91155),
            .in3(N__65021),
            .lcout(N_122_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNI923K31_15_LC_14_21_4.C_ON=1'b0;
    defparam shift_srl_0_RNI923K31_15_LC_14_21_4.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNI923K31_15_LC_14_21_4.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNI923K31_15_LC_14_21_4 (
            .in0(N__65022),
            .in1(N__66611),
            .in2(N__90484),
            .in3(N__61974),
            .lcout(clk_en_142),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIIVHG41_15_LC_14_21_5.C_ON=1'b0;
    defparam shift_srl_0_RNIIVHG41_15_LC_14_21_5.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIIVHG41_15_LC_14_21_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNIIVHG41_15_LC_14_21_5 (
            .in0(N__61973),
            .in1(N__65023),
            .in2(N__90492),
            .in3(N__66536),
            .lcout(clk_en_145),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNI06OT21_15_LC_14_21_6.C_ON=1'b0;
    defparam shift_srl_0_RNI06OT21_15_LC_14_21_6.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNI06OT21_15_LC_14_21_6.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNI06OT21_15_LC_14_21_6 (
            .in0(N__65020),
            .in1(N__64975),
            .in2(N__90483),
            .in3(N__79455),
            .lcout(clk_en_139),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_120_RNIG17D2_15_LC_14_21_7.C_ON=1'b0;
    defparam shift_srl_120_RNIG17D2_15_LC_14_21_7.SEQ_MODE=4'b0000;
    defparam shift_srl_120_RNIG17D2_15_LC_14_21_7.LUT_INIT=16'b0010000000000000;
    LogicCell40 shift_srl_120_RNIG17D2_15_LC_14_21_7 (
            .in0(N__65855),
            .in1(N__61912),
            .in2(N__65603),
            .in3(N__61906),
            .lcout(shift_srl_120_RNIG17D2Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_139_0_LC_14_22_0.C_ON=1'b0;
    defparam shift_srl_139_0_LC_14_22_0.SEQ_MODE=4'b1000;
    defparam shift_srl_139_0_LC_14_22_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_139_0_LC_14_22_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88113),
            .lcout(shift_srl_139Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93107),
            .ce(N__64801),
            .sr(_gnd_net_));
    defparam shift_srl_139_1_LC_14_22_1.C_ON=1'b0;
    defparam shift_srl_139_1_LC_14_22_1.SEQ_MODE=4'b1000;
    defparam shift_srl_139_1_LC_14_22_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_139_1_LC_14_22_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61891),
            .lcout(shift_srl_139Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93107),
            .ce(N__64801),
            .sr(_gnd_net_));
    defparam shift_srl_139_2_LC_14_22_2.C_ON=1'b0;
    defparam shift_srl_139_2_LC_14_22_2.SEQ_MODE=4'b1000;
    defparam shift_srl_139_2_LC_14_22_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_139_2_LC_14_22_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61885),
            .lcout(shift_srl_139Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93107),
            .ce(N__64801),
            .sr(_gnd_net_));
    defparam shift_srl_139_3_LC_14_22_3.C_ON=1'b0;
    defparam shift_srl_139_3_LC_14_22_3.SEQ_MODE=4'b1000;
    defparam shift_srl_139_3_LC_14_22_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_139_3_LC_14_22_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62080),
            .lcout(shift_srl_139Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93107),
            .ce(N__64801),
            .sr(_gnd_net_));
    defparam shift_srl_139_4_LC_14_22_4.C_ON=1'b0;
    defparam shift_srl_139_4_LC_14_22_4.SEQ_MODE=4'b1000;
    defparam shift_srl_139_4_LC_14_22_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_139_4_LC_14_22_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62074),
            .lcout(shift_srl_139Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93107),
            .ce(N__64801),
            .sr(_gnd_net_));
    defparam shift_srl_139_5_LC_14_22_5.C_ON=1'b0;
    defparam shift_srl_139_5_LC_14_22_5.SEQ_MODE=4'b1000;
    defparam shift_srl_139_5_LC_14_22_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_139_5_LC_14_22_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62068),
            .lcout(shift_srl_139Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93107),
            .ce(N__64801),
            .sr(_gnd_net_));
    defparam shift_srl_139_6_LC_14_22_6.C_ON=1'b0;
    defparam shift_srl_139_6_LC_14_22_6.SEQ_MODE=4'b1000;
    defparam shift_srl_139_6_LC_14_22_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_139_6_LC_14_22_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62062),
            .lcout(shift_srl_139Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93107),
            .ce(N__64801),
            .sr(_gnd_net_));
    defparam shift_srl_139_7_LC_14_22_7.C_ON=1'b0;
    defparam shift_srl_139_7_LC_14_22_7.SEQ_MODE=4'b1000;
    defparam shift_srl_139_7_LC_14_22_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_139_7_LC_14_22_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62056),
            .lcout(shift_srl_139Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93107),
            .ce(N__64801),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIBCKVS_15_LC_14_23_0.C_ON=1'b0;
    defparam shift_srl_0_RNIBCKVS_15_LC_14_23_0.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIBCKVS_15_LC_14_23_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNIBCKVS_15_LC_14_23_0 (
            .in0(N__62588),
            .in1(N__64950),
            .in2(N__90552),
            .in3(N__79482),
            .lcout(clk_en_115),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_110_RNI66GS_15_LC_14_23_1.C_ON=1'b0;
    defparam shift_srl_110_RNI66GS_15_LC_14_23_1.SEQ_MODE=4'b0000;
    defparam shift_srl_110_RNI66GS_15_LC_14_23_1.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_110_RNI66GS_15_LC_14_23_1 (
            .in0(N__62423),
            .in1(N__62402),
            .in2(_gnd_net_),
            .in3(N__62302),
            .lcout(),
            .ltout(rco_int_0_a2_0_a2_s_0_1_110_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_107_RNI2EB43_15_LC_14_23_2.C_ON=1'b0;
    defparam shift_srl_107_RNI2EB43_15_LC_14_23_2.SEQ_MODE=4'b0000;
    defparam shift_srl_107_RNI2EB43_15_LC_14_23_2.LUT_INIT=16'b0000000010000000;
    LogicCell40 shift_srl_107_RNI2EB43_15_LC_14_23_2 (
            .in0(N__62370),
            .in1(N__62268),
            .in2(N__62050),
            .in3(N__62250),
            .lcout(rco_int_0_a2_0_a2_out_5),
            .ltout(rco_int_0_a2_0_a2_out_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_114_RNIG0QUS_15_LC_14_23_3.C_ON=1'b0;
    defparam shift_srl_114_RNIG0QUS_15_LC_14_23_3.SEQ_MODE=4'b0000;
    defparam shift_srl_114_RNIG0QUS_15_LC_14_23_3.LUT_INIT=16'b1010000000000000;
    LogicCell40 shift_srl_114_RNIG0QUS_15_LC_14_23_3 (
            .in0(N__79483),
            .in1(_gnd_net_),
            .in2(N__62047),
            .in3(N__62589),
            .lcout(N_162),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_110_15_LC_14_23_4.C_ON=1'b0;
    defparam shift_srl_110_15_LC_14_23_4.SEQ_MODE=4'b1000;
    defparam shift_srl_110_15_LC_14_23_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_110_15_LC_14_23_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62470),
            .lcout(shift_srl_110Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93125),
            .ce(N__62455),
            .sr(_gnd_net_));
    defparam shift_srl_110_RNI91581_15_LC_14_23_5.C_ON=1'b0;
    defparam shift_srl_110_RNI91581_15_LC_14_23_5.SEQ_MODE=4'b0000;
    defparam shift_srl_110_RNI91581_15_LC_14_23_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_110_RNI91581_15_LC_14_23_5 (
            .in0(N__62424),
            .in1(N__62403),
            .in2(N__62374),
            .in3(N__62303),
            .lcout(),
            .ltout(shift_srl_110_RNI91581Z0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_110_RNI4QDG2_15_LC_14_23_6.C_ON=1'b0;
    defparam shift_srl_110_RNI4QDG2_15_LC_14_23_6.SEQ_MODE=4'b0000;
    defparam shift_srl_110_RNI4QDG2_15_LC_14_23_6.LUT_INIT=16'b1110001011100010;
    LogicCell40 shift_srl_110_RNI4QDG2_15_LC_14_23_6 (
            .in0(_gnd_net_),
            .in1(N__62269),
            .in2(N__62254),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(shift_srl_110_RNI4QDG2Z0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_145_RNIN9307_15_LC_14_23_7.C_ON=1'b0;
    defparam shift_srl_145_RNIN9307_15_LC_14_23_7.SEQ_MODE=4'b0000;
    defparam shift_srl_145_RNIN9307_15_LC_14_23_7.LUT_INIT=16'b0100000000000000;
    LogicCell40 shift_srl_145_RNIN9307_15_LC_14_23_7 (
            .in0(N__62251),
            .in1(N__62235),
            .in2(N__62218),
            .in3(N__63590),
            .lcout(shift_srl_145_RNIN9307Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_198_RNI842R2_15_LC_14_24_0.C_ON=1'b0;
    defparam shift_srl_198_RNI842R2_15_LC_14_24_0.SEQ_MODE=4'b0000;
    defparam shift_srl_198_RNI842R2_15_LC_14_24_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_198_RNI842R2_15_LC_14_24_0 (
            .in0(N__62215),
            .in1(N__62200),
            .in2(N__70426),
            .in3(N__62181),
            .lcout(),
            .ltout(g0_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_198_RNIOVF1F_15_LC_14_24_1.C_ON=1'b0;
    defparam shift_srl_198_RNIOVF1F_15_LC_14_24_1.SEQ_MODE=4'b0000;
    defparam shift_srl_198_RNIOVF1F_15_LC_14_24_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_198_RNIOVF1F_15_LC_14_24_1 (
            .in0(N__62542),
            .in1(N__62086),
            .in2(N__62140),
            .in3(N__84244),
            .lcout(),
            .ltout(g0_16_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_183_RNIUE0UH1_15_LC_14_24_2.C_ON=1'b0;
    defparam shift_srl_183_RNIUE0UH1_15_LC_14_24_2.SEQ_MODE=4'b0000;
    defparam shift_srl_183_RNIUE0UH1_15_LC_14_24_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_183_RNIUE0UH1_15_LC_14_24_2 (
            .in0(N__70093),
            .in1(N__72216),
            .in2(N__62137),
            .in3(N__79542),
            .lcout(clk_en_199),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_144_RNISRV86_15_LC_14_24_3.C_ON=1'b0;
    defparam shift_srl_144_RNISRV86_15_LC_14_24_3.SEQ_MODE=4'b0000;
    defparam shift_srl_144_RNISRV86_15_LC_14_24_3.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_144_RNISRV86_15_LC_14_24_3 (
            .in0(N__66540),
            .in1(N__62125),
            .in2(_gnd_net_),
            .in3(N__64949),
            .lcout(g0_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_114_RNIGOM73_15_LC_14_24_4.C_ON=1'b0;
    defparam shift_srl_114_RNIGOM73_15_LC_14_24_4.SEQ_MODE=4'b0000;
    defparam shift_srl_114_RNIGOM73_15_LC_14_24_4.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_114_RNIGOM73_15_LC_14_24_4 (
            .in0(N__65739),
            .in1(N__62587),
            .in2(N__65550),
            .in3(N__65374),
            .lcout(g0_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_197_RNI3Q873_15_LC_14_24_5.C_ON=1'b0;
    defparam shift_srl_197_RNI3Q873_15_LC_14_24_5.SEQ_MODE=4'b0000;
    defparam shift_srl_197_RNI3Q873_15_LC_14_24_5.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_197_RNI3Q873_15_LC_14_24_5 (
            .in0(N__70636),
            .in1(N__72385),
            .in2(_gnd_net_),
            .in3(N__73828),
            .lcout(N_4183),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_199_10_LC_14_25_0.C_ON=1'b0;
    defparam shift_srl_199_10_LC_14_25_0.SEQ_MODE=4'b1000;
    defparam shift_srl_199_10_LC_14_25_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_199_10_LC_14_25_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62497),
            .lcout(shift_srl_199Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93161),
            .ce(N__62720),
            .sr(_gnd_net_));
    defparam shift_srl_199_11_LC_14_25_1.C_ON=1'b0;
    defparam shift_srl_199_11_LC_14_25_1.SEQ_MODE=4'b1000;
    defparam shift_srl_199_11_LC_14_25_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_199_11_LC_14_25_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62536),
            .lcout(shift_srl_199Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93161),
            .ce(N__62720),
            .sr(_gnd_net_));
    defparam shift_srl_199_12_LC_14_25_2.C_ON=1'b0;
    defparam shift_srl_199_12_LC_14_25_2.SEQ_MODE=4'b1000;
    defparam shift_srl_199_12_LC_14_25_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_199_12_LC_14_25_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62530),
            .lcout(shift_srl_199Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93161),
            .ce(N__62720),
            .sr(_gnd_net_));
    defparam shift_srl_199_13_LC_14_25_3.C_ON=1'b0;
    defparam shift_srl_199_13_LC_14_25_3.SEQ_MODE=4'b1000;
    defparam shift_srl_199_13_LC_14_25_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_199_13_LC_14_25_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62524),
            .lcout(shift_srl_199Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93161),
            .ce(N__62720),
            .sr(_gnd_net_));
    defparam shift_srl_199_14_LC_14_25_4.C_ON=1'b0;
    defparam shift_srl_199_14_LC_14_25_4.SEQ_MODE=4'b1000;
    defparam shift_srl_199_14_LC_14_25_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_199_14_LC_14_25_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62518),
            .lcout(shift_srl_199Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93161),
            .ce(N__62720),
            .sr(_gnd_net_));
    defparam shift_srl_199_15_LC_14_25_5.C_ON=1'b0;
    defparam shift_srl_199_15_LC_14_25_5.SEQ_MODE=4'b1000;
    defparam shift_srl_199_15_LC_14_25_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_199_15_LC_14_25_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62512),
            .lcout(shift_srl_199Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93161),
            .ce(N__62720),
            .sr(_gnd_net_));
    defparam shift_srl_199_9_LC_14_25_6.C_ON=1'b0;
    defparam shift_srl_199_9_LC_14_25_6.SEQ_MODE=4'b1000;
    defparam shift_srl_199_9_LC_14_25_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_199_9_LC_14_25_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62476),
            .lcout(shift_srl_199Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93161),
            .ce(N__62720),
            .sr(_gnd_net_));
    defparam shift_srl_199_8_LC_14_25_7.C_ON=1'b0;
    defparam shift_srl_199_8_LC_14_25_7.SEQ_MODE=4'b1000;
    defparam shift_srl_199_8_LC_14_25_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_199_8_LC_14_25_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62491),
            .lcout(shift_srl_199Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93161),
            .ce(N__62720),
            .sr(_gnd_net_));
    defparam shift_srl_102_0_LC_14_26_0.C_ON=1'b0;
    defparam shift_srl_102_0_LC_14_26_0.SEQ_MODE=4'b1000;
    defparam shift_srl_102_0_LC_14_26_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_102_0_LC_14_26_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62703),
            .lcout(shift_srl_102Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93181),
            .ce(N__62617),
            .sr(_gnd_net_));
    defparam shift_srl_102_1_LC_14_26_1.C_ON=1'b0;
    defparam shift_srl_102_1_LC_14_26_1.SEQ_MODE=4'b1000;
    defparam shift_srl_102_1_LC_14_26_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_102_1_LC_14_26_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62671),
            .lcout(shift_srl_102Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93181),
            .ce(N__62617),
            .sr(_gnd_net_));
    defparam shift_srl_102_2_LC_14_26_2.C_ON=1'b0;
    defparam shift_srl_102_2_LC_14_26_2.SEQ_MODE=4'b1000;
    defparam shift_srl_102_2_LC_14_26_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_102_2_LC_14_26_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62665),
            .lcout(shift_srl_102Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93181),
            .ce(N__62617),
            .sr(_gnd_net_));
    defparam shift_srl_102_3_LC_14_26_3.C_ON=1'b0;
    defparam shift_srl_102_3_LC_14_26_3.SEQ_MODE=4'b1000;
    defparam shift_srl_102_3_LC_14_26_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_102_3_LC_14_26_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62659),
            .lcout(shift_srl_102Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93181),
            .ce(N__62617),
            .sr(_gnd_net_));
    defparam shift_srl_102_4_LC_14_26_4.C_ON=1'b0;
    defparam shift_srl_102_4_LC_14_26_4.SEQ_MODE=4'b1000;
    defparam shift_srl_102_4_LC_14_26_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_102_4_LC_14_26_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62653),
            .lcout(shift_srl_102Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93181),
            .ce(N__62617),
            .sr(_gnd_net_));
    defparam shift_srl_102_5_LC_14_26_5.C_ON=1'b0;
    defparam shift_srl_102_5_LC_14_26_5.SEQ_MODE=4'b1000;
    defparam shift_srl_102_5_LC_14_26_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_102_5_LC_14_26_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62647),
            .lcout(shift_srl_102Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93181),
            .ce(N__62617),
            .sr(_gnd_net_));
    defparam shift_srl_102_6_LC_14_26_6.C_ON=1'b0;
    defparam shift_srl_102_6_LC_14_26_6.SEQ_MODE=4'b1000;
    defparam shift_srl_102_6_LC_14_26_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_102_6_LC_14_26_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62641),
            .lcout(shift_srl_102Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93181),
            .ce(N__62617),
            .sr(_gnd_net_));
    defparam shift_srl_102_9_LC_14_26_7.C_ON=1'b0;
    defparam shift_srl_102_9_LC_14_26_7.SEQ_MODE=4'b1000;
    defparam shift_srl_102_9_LC_14_26_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_102_9_LC_14_26_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62629),
            .lcout(shift_srl_102Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93181),
            .ce(N__62617),
            .sr(_gnd_net_));
    defparam shift_srl_139_9_LC_14_27_1.C_ON=1'b0;
    defparam shift_srl_139_9_LC_14_27_1.SEQ_MODE=4'b1000;
    defparam shift_srl_139_9_LC_14_27_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_139_9_LC_14_27_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62779),
            .lcout(shift_srl_139Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93203),
            .ce(N__64820),
            .sr(_gnd_net_));
    defparam shift_srl_139_8_LC_14_27_3.C_ON=1'b0;
    defparam shift_srl_139_8_LC_14_27_3.SEQ_MODE=4'b1000;
    defparam shift_srl_139_8_LC_14_27_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_139_8_LC_14_27_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62791),
            .lcout(shift_srl_139Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93203),
            .ce(N__64820),
            .sr(_gnd_net_));
    defparam shift_srl_139_11_LC_14_28_3.C_ON=1'b0;
    defparam shift_srl_139_11_LC_14_28_3.SEQ_MODE=4'b1000;
    defparam shift_srl_139_11_LC_14_28_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_139_11_LC_14_28_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62767),
            .lcout(shift_srl_139Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93223),
            .ce(N__64827),
            .sr(_gnd_net_));
    defparam shift_srl_139_10_LC_14_28_7.C_ON=1'b0;
    defparam shift_srl_139_10_LC_14_28_7.SEQ_MODE=4'b1000;
    defparam shift_srl_139_10_LC_14_28_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_139_10_LC_14_28_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62773),
            .lcout(shift_srl_139Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93223),
            .ce(N__64827),
            .sr(_gnd_net_));
    defparam shift_srl_85_10_LC_15_5_0.C_ON=1'b0;
    defparam shift_srl_85_10_LC_15_5_0.SEQ_MODE=4'b1000;
    defparam shift_srl_85_10_LC_15_5_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_85_10_LC_15_5_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62839),
            .lcout(shift_srl_85Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93264),
            .ce(N__64239),
            .sr(_gnd_net_));
    defparam shift_srl_85_11_LC_15_5_1.C_ON=1'b0;
    defparam shift_srl_85_11_LC_15_5_1.SEQ_MODE=4'b1000;
    defparam shift_srl_85_11_LC_15_5_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_85_11_LC_15_5_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62761),
            .lcout(shift_srl_85Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93264),
            .ce(N__64239),
            .sr(_gnd_net_));
    defparam shift_srl_85_12_LC_15_5_2.C_ON=1'b0;
    defparam shift_srl_85_12_LC_15_5_2.SEQ_MODE=4'b1000;
    defparam shift_srl_85_12_LC_15_5_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_85_12_LC_15_5_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62755),
            .lcout(shift_srl_85Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93264),
            .ce(N__64239),
            .sr(_gnd_net_));
    defparam shift_srl_85_13_LC_15_5_3.C_ON=1'b0;
    defparam shift_srl_85_13_LC_15_5_3.SEQ_MODE=4'b1000;
    defparam shift_srl_85_13_LC_15_5_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_85_13_LC_15_5_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62749),
            .lcout(shift_srl_85Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93264),
            .ce(N__64239),
            .sr(_gnd_net_));
    defparam shift_srl_85_14_LC_15_5_4.C_ON=1'b0;
    defparam shift_srl_85_14_LC_15_5_4.SEQ_MODE=4'b1000;
    defparam shift_srl_85_14_LC_15_5_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_85_14_LC_15_5_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62743),
            .lcout(shift_srl_85Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93264),
            .ce(N__64239),
            .sr(_gnd_net_));
    defparam shift_srl_85_15_LC_15_5_5.C_ON=1'b0;
    defparam shift_srl_85_15_LC_15_5_5.SEQ_MODE=4'b1000;
    defparam shift_srl_85_15_LC_15_5_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_85_15_LC_15_5_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62737),
            .lcout(shift_srl_85Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93264),
            .ce(N__64239),
            .sr(_gnd_net_));
    defparam shift_srl_85_9_LC_15_5_6.C_ON=1'b0;
    defparam shift_srl_85_9_LC_15_5_6.SEQ_MODE=4'b1000;
    defparam shift_srl_85_9_LC_15_5_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_85_9_LC_15_5_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62833),
            .lcout(shift_srl_85Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93264),
            .ce(N__64239),
            .sr(_gnd_net_));
    defparam shift_srl_85_8_LC_15_5_7.C_ON=1'b0;
    defparam shift_srl_85_8_LC_15_5_7.SEQ_MODE=4'b1000;
    defparam shift_srl_85_8_LC_15_5_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_85_8_LC_15_5_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64249),
            .lcout(shift_srl_85Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93264),
            .ce(N__64239),
            .sr(_gnd_net_));
    defparam shift_srl_88_10_LC_15_6_0.C_ON=1'b0;
    defparam shift_srl_88_10_LC_15_6_0.SEQ_MODE=4'b1000;
    defparam shift_srl_88_10_LC_15_6_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_88_10_LC_15_6_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62797),
            .lcout(shift_srl_88Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93244),
            .ce(N__64326),
            .sr(_gnd_net_));
    defparam shift_srl_88_11_LC_15_6_1.C_ON=1'b0;
    defparam shift_srl_88_11_LC_15_6_1.SEQ_MODE=4'b1000;
    defparam shift_srl_88_11_LC_15_6_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_88_11_LC_15_6_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62827),
            .lcout(shift_srl_88Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93244),
            .ce(N__64326),
            .sr(_gnd_net_));
    defparam shift_srl_88_12_LC_15_6_2.C_ON=1'b0;
    defparam shift_srl_88_12_LC_15_6_2.SEQ_MODE=4'b1000;
    defparam shift_srl_88_12_LC_15_6_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_88_12_LC_15_6_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62821),
            .lcout(shift_srl_88Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93244),
            .ce(N__64326),
            .sr(_gnd_net_));
    defparam shift_srl_88_13_LC_15_6_3.C_ON=1'b0;
    defparam shift_srl_88_13_LC_15_6_3.SEQ_MODE=4'b1000;
    defparam shift_srl_88_13_LC_15_6_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_88_13_LC_15_6_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62815),
            .lcout(shift_srl_88Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93244),
            .ce(N__64326),
            .sr(_gnd_net_));
    defparam shift_srl_88_14_LC_15_6_4.C_ON=1'b0;
    defparam shift_srl_88_14_LC_15_6_4.SEQ_MODE=4'b1000;
    defparam shift_srl_88_14_LC_15_6_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_88_14_LC_15_6_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62809),
            .lcout(shift_srl_88Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93244),
            .ce(N__64326),
            .sr(_gnd_net_));
    defparam shift_srl_88_15_LC_15_6_5.C_ON=1'b0;
    defparam shift_srl_88_15_LC_15_6_5.SEQ_MODE=4'b1000;
    defparam shift_srl_88_15_LC_15_6_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_88_15_LC_15_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62803),
            .lcout(shift_srl_88Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93244),
            .ce(N__64326),
            .sr(_gnd_net_));
    defparam shift_srl_88_9_LC_15_6_6.C_ON=1'b0;
    defparam shift_srl_88_9_LC_15_6_6.SEQ_MODE=4'b1000;
    defparam shift_srl_88_9_LC_15_6_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_88_9_LC_15_6_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62914),
            .lcout(shift_srl_88Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93244),
            .ce(N__64326),
            .sr(_gnd_net_));
    defparam shift_srl_88_8_LC_15_6_7.C_ON=1'b0;
    defparam shift_srl_88_8_LC_15_6_7.SEQ_MODE=4'b1000;
    defparam shift_srl_88_8_LC_15_6_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_88_8_LC_15_6_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64333),
            .lcout(shift_srl_88Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93244),
            .ce(N__64326),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_88_LC_15_7_0.C_ON=1'b0;
    defparam rco_obuf_RNO_88_LC_15_7_0.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_88_LC_15_7_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 rco_obuf_RNO_88_LC_15_7_0 (
            .in0(N__62881),
            .in1(N__66985),
            .in2(N__68509),
            .in3(N__67100),
            .lcout(rco_c_88),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_59_RNILFPCL_15_LC_15_7_3.C_ON=1'b0;
    defparam shift_srl_59_RNILFPCL_15_LC_15_7_3.SEQ_MODE=4'b0000;
    defparam shift_srl_59_RNILFPCL_15_LC_15_7_3.LUT_INIT=16'b0100000000000000;
    LogicCell40 shift_srl_59_RNILFPCL_15_LC_15_7_3 (
            .in0(N__67353),
            .in1(N__86821),
            .in2(N__73072),
            .in3(N__80774),
            .lcout(rco_c_83),
            .ltout(rco_c_83_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_84_RNI7UOLL_15_LC_15_7_4.C_ON=1'b0;
    defparam shift_srl_84_RNI7UOLL_15_LC_15_7_4.SEQ_MODE=4'b0000;
    defparam shift_srl_84_RNI7UOLL_15_LC_15_7_4.LUT_INIT=16'b1100000000000000;
    LogicCell40 shift_srl_84_RNI7UOLL_15_LC_15_7_4 (
            .in0(_gnd_net_),
            .in1(N__89973),
            .in2(N__62893),
            .in3(N__68682),
            .lcout(clk_en_85),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIOFL2M_15_LC_15_7_5.C_ON=1'b0;
    defparam shift_srl_0_RNIOFL2M_15_LC_15_7_5.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIOFL2M_15_LC_15_7_5.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_0_RNIOFL2M_15_LC_15_7_5 (
            .in0(N__89978),
            .in1(N__62877),
            .in2(_gnd_net_),
            .in3(N__68481),
            .lcout(clk_en_87),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_87_RNIIUC7M_15_LC_15_7_6.C_ON=1'b0;
    defparam shift_srl_87_RNIIUC7M_15_LC_15_7_6.SEQ_MODE=4'b0000;
    defparam shift_srl_87_RNIIUC7M_15_LC_15_7_6.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_87_RNIIUC7M_15_LC_15_7_6 (
            .in0(N__68479),
            .in1(N__89974),
            .in2(N__62888),
            .in3(N__67099),
            .lcout(clk_en_88),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_85_RNIV442M_15_LC_15_7_7.C_ON=1'b0;
    defparam shift_srl_85_RNIV442M_15_LC_15_7_7.SEQ_MODE=4'b0000;
    defparam shift_srl_85_RNIV442M_15_LC_15_7_7.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_85_RNIV442M_15_LC_15_7_7 (
            .in0(N__68681),
            .in1(N__67057),
            .in2(N__90244),
            .in3(N__68480),
            .lcout(clk_en_86),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_86_10_LC_15_8_0.C_ON=1'b0;
    defparam shift_srl_86_10_LC_15_8_0.SEQ_MODE=4'b1000;
    defparam shift_srl_86_10_LC_15_8_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_86_10_LC_15_8_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62950),
            .lcout(shift_srl_86Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93205),
            .ce(N__67169),
            .sr(_gnd_net_));
    defparam shift_srl_86_7_LC_15_8_1.C_ON=1'b0;
    defparam shift_srl_86_7_LC_15_8_1.SEQ_MODE=4'b1000;
    defparam shift_srl_86_7_LC_15_8_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_86_7_LC_15_8_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62968),
            .lcout(shift_srl_86Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93205),
            .ce(N__67169),
            .sr(_gnd_net_));
    defparam shift_srl_86_6_LC_15_8_2.C_ON=1'b0;
    defparam shift_srl_86_6_LC_15_8_2.SEQ_MODE=4'b1000;
    defparam shift_srl_86_6_LC_15_8_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_86_6_LC_15_8_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62974),
            .lcout(shift_srl_86Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93205),
            .ce(N__67169),
            .sr(_gnd_net_));
    defparam shift_srl_86_13_LC_15_8_3.C_ON=1'b0;
    defparam shift_srl_86_13_LC_15_8_3.SEQ_MODE=4'b1000;
    defparam shift_srl_86_13_LC_15_8_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_86_13_LC_15_8_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62962),
            .lcout(shift_srl_86Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93205),
            .ce(N__67169),
            .sr(_gnd_net_));
    defparam shift_srl_86_14_LC_15_8_4.C_ON=1'b0;
    defparam shift_srl_86_14_LC_15_8_4.SEQ_MODE=4'b1000;
    defparam shift_srl_86_14_LC_15_8_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_86_14_LC_15_8_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62956),
            .lcout(shift_srl_86Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93205),
            .ce(N__67169),
            .sr(_gnd_net_));
    defparam shift_srl_86_9_LC_15_8_5.C_ON=1'b0;
    defparam shift_srl_86_9_LC_15_8_5.SEQ_MODE=4'b1000;
    defparam shift_srl_86_9_LC_15_8_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_86_9_LC_15_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62938),
            .lcout(shift_srl_86Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93205),
            .ce(N__67169),
            .sr(_gnd_net_));
    defparam shift_srl_86_8_LC_15_8_6.C_ON=1'b0;
    defparam shift_srl_86_8_LC_15_8_6.SEQ_MODE=4'b1000;
    defparam shift_srl_86_8_LC_15_8_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_86_8_LC_15_8_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62944),
            .lcout(shift_srl_86Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93205),
            .ce(N__67169),
            .sr(_gnd_net_));
    defparam shift_srl_43_12_LC_15_9_3.C_ON=1'b0;
    defparam shift_srl_43_12_LC_15_9_3.SEQ_MODE=4'b1000;
    defparam shift_srl_43_12_LC_15_9_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_43_12_LC_15_9_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62932),
            .lcout(shift_srl_43Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93184),
            .ce(N__68998),
            .sr(_gnd_net_));
    defparam shift_srl_43_6_LC_15_10_0.C_ON=1'b0;
    defparam shift_srl_43_6_LC_15_10_0.SEQ_MODE=4'b1000;
    defparam shift_srl_43_6_LC_15_10_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_43_6_LC_15_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62980),
            .lcout(shift_srl_43Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93162),
            .ce(N__68997),
            .sr(_gnd_net_));
    defparam shift_srl_43_11_LC_15_10_1.C_ON=1'b0;
    defparam shift_srl_43_11_LC_15_10_1.SEQ_MODE=4'b1000;
    defparam shift_srl_43_11_LC_15_10_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_43_11_LC_15_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62926),
            .lcout(shift_srl_43Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93162),
            .ce(N__68997),
            .sr(_gnd_net_));
    defparam shift_srl_43_10_LC_15_10_2.C_ON=1'b0;
    defparam shift_srl_43_10_LC_15_10_2.SEQ_MODE=4'b1000;
    defparam shift_srl_43_10_LC_15_10_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_43_10_LC_15_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63010),
            .lcout(shift_srl_43Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93162),
            .ce(N__68997),
            .sr(_gnd_net_));
    defparam shift_srl_43_13_LC_15_10_3.C_ON=1'b0;
    defparam shift_srl_43_13_LC_15_10_3.SEQ_MODE=4'b1000;
    defparam shift_srl_43_13_LC_15_10_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_43_13_LC_15_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62920),
            .lcout(shift_srl_43Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93162),
            .ce(N__68997),
            .sr(_gnd_net_));
    defparam shift_srl_43_14_LC_15_10_4.C_ON=1'b0;
    defparam shift_srl_43_14_LC_15_10_4.SEQ_MODE=4'b1000;
    defparam shift_srl_43_14_LC_15_10_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_43_14_LC_15_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63022),
            .lcout(shift_srl_43Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93162),
            .ce(N__68997),
            .sr(_gnd_net_));
    defparam shift_srl_43_15_LC_15_10_5.C_ON=1'b0;
    defparam shift_srl_43_15_LC_15_10_5.SEQ_MODE=4'b1000;
    defparam shift_srl_43_15_LC_15_10_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_43_15_LC_15_10_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63016),
            .lcout(shift_srl_43Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93162),
            .ce(N__68997),
            .sr(_gnd_net_));
    defparam shift_srl_43_9_LC_15_10_6.C_ON=1'b0;
    defparam shift_srl_43_9_LC_15_10_6.SEQ_MODE=4'b1000;
    defparam shift_srl_43_9_LC_15_10_6.LUT_INIT=16'b1100110011001100;
    LogicCell40 shift_srl_43_9_LC_15_10_6 (
            .in0(_gnd_net_),
            .in1(N__63004),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_43Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93162),
            .ce(N__68997),
            .sr(_gnd_net_));
    defparam shift_srl_43_0_LC_15_11_0.C_ON=1'b0;
    defparam shift_srl_43_0_LC_15_11_0.SEQ_MODE=4'b1000;
    defparam shift_srl_43_0_LC_15_11_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_43_0_LC_15_11_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73261),
            .lcout(shift_srl_43Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93145),
            .ce(N__68990),
            .sr(_gnd_net_));
    defparam shift_srl_43_8_LC_15_11_1.C_ON=1'b0;
    defparam shift_srl_43_8_LC_15_11_1.SEQ_MODE=4'b1000;
    defparam shift_srl_43_8_LC_15_11_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_43_8_LC_15_11_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63058),
            .lcout(shift_srl_43Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93145),
            .ce(N__68990),
            .sr(_gnd_net_));
    defparam shift_srl_43_2_LC_15_11_2.C_ON=1'b0;
    defparam shift_srl_43_2_LC_15_11_2.SEQ_MODE=4'b1000;
    defparam shift_srl_43_2_LC_15_11_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_43_2_LC_15_11_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63070),
            .lcout(shift_srl_43Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93145),
            .ce(N__68990),
            .sr(_gnd_net_));
    defparam shift_srl_43_3_LC_15_11_3.C_ON=1'b0;
    defparam shift_srl_43_3_LC_15_11_3.SEQ_MODE=4'b1000;
    defparam shift_srl_43_3_LC_15_11_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_43_3_LC_15_11_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62998),
            .lcout(shift_srl_43Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93145),
            .ce(N__68990),
            .sr(_gnd_net_));
    defparam shift_srl_43_4_LC_15_11_4.C_ON=1'b0;
    defparam shift_srl_43_4_LC_15_11_4.SEQ_MODE=4'b1000;
    defparam shift_srl_43_4_LC_15_11_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_43_4_LC_15_11_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62992),
            .lcout(shift_srl_43Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93145),
            .ce(N__68990),
            .sr(_gnd_net_));
    defparam shift_srl_43_5_LC_15_11_5.C_ON=1'b0;
    defparam shift_srl_43_5_LC_15_11_5.SEQ_MODE=4'b1000;
    defparam shift_srl_43_5_LC_15_11_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_43_5_LC_15_11_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62986),
            .lcout(shift_srl_43Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93145),
            .ce(N__68990),
            .sr(_gnd_net_));
    defparam shift_srl_43_1_LC_15_11_6.C_ON=1'b0;
    defparam shift_srl_43_1_LC_15_11_6.SEQ_MODE=4'b1000;
    defparam shift_srl_43_1_LC_15_11_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_43_1_LC_15_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63076),
            .lcout(shift_srl_43Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93145),
            .ce(N__68990),
            .sr(_gnd_net_));
    defparam shift_srl_43_7_LC_15_11_7.C_ON=1'b0;
    defparam shift_srl_43_7_LC_15_11_7.SEQ_MODE=4'b1000;
    defparam shift_srl_43_7_LC_15_11_7.LUT_INIT=16'b1100110011001100;
    LogicCell40 shift_srl_43_7_LC_15_11_7 (
            .in0(_gnd_net_),
            .in1(N__63064),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_43Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93145),
            .ce(N__68990),
            .sr(_gnd_net_));
    defparam shift_srl_99_6_LC_15_12_0.C_ON=1'b0;
    defparam shift_srl_99_6_LC_15_12_0.SEQ_MODE=4'b1000;
    defparam shift_srl_99_6_LC_15_12_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_99_6_LC_15_12_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67663),
            .lcout(shift_srl_99Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93126),
            .ce(N__67650),
            .sr(_gnd_net_));
    defparam shift_srl_24_10_LC_15_13_0.C_ON=1'b0;
    defparam shift_srl_24_10_LC_15_13_0.SEQ_MODE=4'b1000;
    defparam shift_srl_24_10_LC_15_13_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_24_10_LC_15_13_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63160),
            .lcout(shift_srl_24Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93108),
            .ce(N__63154),
            .sr(_gnd_net_));
    defparam shift_srl_24_11_LC_15_13_1.C_ON=1'b0;
    defparam shift_srl_24_11_LC_15_13_1.SEQ_MODE=4'b1000;
    defparam shift_srl_24_11_LC_15_13_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_24_11_LC_15_13_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63052),
            .lcout(shift_srl_24Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93108),
            .ce(N__63154),
            .sr(_gnd_net_));
    defparam shift_srl_24_12_LC_15_13_2.C_ON=1'b0;
    defparam shift_srl_24_12_LC_15_13_2.SEQ_MODE=4'b1000;
    defparam shift_srl_24_12_LC_15_13_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_24_12_LC_15_13_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63046),
            .lcout(shift_srl_24Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93108),
            .ce(N__63154),
            .sr(_gnd_net_));
    defparam shift_srl_24_13_LC_15_13_3.C_ON=1'b0;
    defparam shift_srl_24_13_LC_15_13_3.SEQ_MODE=4'b1000;
    defparam shift_srl_24_13_LC_15_13_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_24_13_LC_15_13_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63040),
            .lcout(shift_srl_24Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93108),
            .ce(N__63154),
            .sr(_gnd_net_));
    defparam shift_srl_24_14_LC_15_13_4.C_ON=1'b0;
    defparam shift_srl_24_14_LC_15_13_4.SEQ_MODE=4'b1000;
    defparam shift_srl_24_14_LC_15_13_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_24_14_LC_15_13_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63034),
            .lcout(shift_srl_24Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93108),
            .ce(N__63154),
            .sr(_gnd_net_));
    defparam shift_srl_24_15_LC_15_13_5.C_ON=1'b0;
    defparam shift_srl_24_15_LC_15_13_5.SEQ_MODE=4'b1000;
    defparam shift_srl_24_15_LC_15_13_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_24_15_LC_15_13_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63028),
            .lcout(shift_srl_24Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93108),
            .ce(N__63154),
            .sr(_gnd_net_));
    defparam shift_srl_24_9_LC_15_13_6.C_ON=1'b0;
    defparam shift_srl_24_9_LC_15_13_6.SEQ_MODE=4'b1000;
    defparam shift_srl_24_9_LC_15_13_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_24_9_LC_15_13_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63166),
            .lcout(shift_srl_24Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93108),
            .ce(N__63154),
            .sr(_gnd_net_));
    defparam shift_srl_152_0_LC_15_14_0.C_ON=1'b0;
    defparam shift_srl_152_0_LC_15_14_0.SEQ_MODE=4'b1000;
    defparam shift_srl_152_0_LC_15_14_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_152_0_LC_15_14_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63241),
            .lcout(shift_srl_152Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93092),
            .ce(N__63192),
            .sr(_gnd_net_));
    defparam shift_srl_152_1_LC_15_14_1.C_ON=1'b0;
    defparam shift_srl_152_1_LC_15_14_1.SEQ_MODE=4'b1000;
    defparam shift_srl_152_1_LC_15_14_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_152_1_LC_15_14_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63124),
            .lcout(shift_srl_152Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93092),
            .ce(N__63192),
            .sr(_gnd_net_));
    defparam shift_srl_152_2_LC_15_14_2.C_ON=1'b0;
    defparam shift_srl_152_2_LC_15_14_2.SEQ_MODE=4'b1000;
    defparam shift_srl_152_2_LC_15_14_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_152_2_LC_15_14_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63118),
            .lcout(shift_srl_152Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93092),
            .ce(N__63192),
            .sr(_gnd_net_));
    defparam shift_srl_152_3_LC_15_14_3.C_ON=1'b0;
    defparam shift_srl_152_3_LC_15_14_3.SEQ_MODE=4'b1000;
    defparam shift_srl_152_3_LC_15_14_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_152_3_LC_15_14_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63112),
            .lcout(shift_srl_152Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93092),
            .ce(N__63192),
            .sr(_gnd_net_));
    defparam shift_srl_152_4_LC_15_14_4.C_ON=1'b0;
    defparam shift_srl_152_4_LC_15_14_4.SEQ_MODE=4'b1000;
    defparam shift_srl_152_4_LC_15_14_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_152_4_LC_15_14_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63106),
            .lcout(shift_srl_152Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93092),
            .ce(N__63192),
            .sr(_gnd_net_));
    defparam shift_srl_152_5_LC_15_14_5.C_ON=1'b0;
    defparam shift_srl_152_5_LC_15_14_5.SEQ_MODE=4'b1000;
    defparam shift_srl_152_5_LC_15_14_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_152_5_LC_15_14_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63100),
            .lcout(shift_srl_152Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93092),
            .ce(N__63192),
            .sr(_gnd_net_));
    defparam shift_srl_152_6_LC_15_14_6.C_ON=1'b0;
    defparam shift_srl_152_6_LC_15_14_6.SEQ_MODE=4'b1000;
    defparam shift_srl_152_6_LC_15_14_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_152_6_LC_15_14_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63094),
            .lcout(shift_srl_152Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93092),
            .ce(N__63192),
            .sr(_gnd_net_));
    defparam shift_srl_152_7_LC_15_14_7.C_ON=1'b0;
    defparam shift_srl_152_7_LC_15_14_7.SEQ_MODE=4'b1000;
    defparam shift_srl_152_7_LC_15_14_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_152_7_LC_15_14_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63088),
            .lcout(shift_srl_152Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93092),
            .ce(N__63192),
            .sr(_gnd_net_));
    defparam shift_srl_152_RNIV45F1_15_LC_15_15_2.C_ON=1'b0;
    defparam shift_srl_152_RNIV45F1_15_LC_15_15_2.SEQ_MODE=4'b0000;
    defparam shift_srl_152_RNIV45F1_15_LC_15_15_2.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_152_RNIV45F1_15_LC_15_15_2 (
            .in0(N__66800),
            .in1(N__90423),
            .in2(N__63248),
            .in3(N__63407),
            .lcout(),
            .ltout(clk_en_0_a3_0_a2_sx_153_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_152_RNIRVDB61_15_LC_15_15_3.C_ON=1'b0;
    defparam shift_srl_152_RNIRVDB61_15_LC_15_15_3.SEQ_MODE=4'b0000;
    defparam shift_srl_152_RNIRVDB61_15_LC_15_15_3.LUT_INIT=16'b0000110000000000;
    LogicCell40 shift_srl_152_RNIRVDB61_15_LC_15_15_3 (
            .in0(_gnd_net_),
            .in1(N__77816),
            .in2(N__63214),
            .in3(N__79555),
            .lcout(clk_en_153),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIM32R51_15_LC_15_15_4.C_ON=1'b0;
    defparam shift_srl_0_RNIM32R51_15_LC_15_15_4.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIM32R51_15_LC_15_15_4.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNIM32R51_15_LC_15_15_4 (
            .in0(N__79556),
            .in1(N__90422),
            .in2(N__66808),
            .in3(N__77820),
            .lcout(clk_en_151),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_91_RNIUH4HP_15_LC_15_15_5.C_ON=1'b0;
    defparam shift_srl_91_RNIUH4HP_15_LC_15_15_5.SEQ_MODE=4'b0000;
    defparam shift_srl_91_RNIUH4HP_15_LC_15_15_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_91_RNIUH4HP_15_LC_15_15_5 (
            .in0(N__85090),
            .in1(N__72029),
            .in2(N__72097),
            .in3(N__77815),
            .lcout(),
            .ltout(shift_srl_91_RNIUH4HPZ0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_91_RNISQ8S41_15_LC_15_15_6.C_ON=1'b0;
    defparam shift_srl_91_RNISQ8S41_15_LC_15_15_6.SEQ_MODE=4'b0000;
    defparam shift_srl_91_RNISQ8S41_15_LC_15_15_6.LUT_INIT=16'b1111000010101010;
    LogicCell40 shift_srl_91_RNISQ8S41_15_LC_15_15_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__63199),
            .in3(N__75053),
            .lcout(rco_c_145),
            .ltout(rco_c_145_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_151_RNIOV4161_15_LC_15_15_7.C_ON=1'b0;
    defparam shift_srl_151_RNIOV4161_15_LC_15_15_7.SEQ_MODE=4'b0000;
    defparam shift_srl_151_RNIOV4161_15_LC_15_15_7.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_151_RNIOV4161_15_LC_15_15_7 (
            .in0(N__63408),
            .in1(N__66804),
            .in2(N__63196),
            .in3(N__90424),
            .lcout(clk_en_152),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_151_0_LC_15_16_0.C_ON=1'b0;
    defparam shift_srl_151_0_LC_15_16_0.SEQ_MODE=4'b1000;
    defparam shift_srl_151_0_LC_15_16_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_151_0_LC_15_16_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63405),
            .lcout(shift_srl_151Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93062),
            .ce(N__63358),
            .sr(_gnd_net_));
    defparam shift_srl_151_1_LC_15_16_1.C_ON=1'b0;
    defparam shift_srl_151_1_LC_15_16_1.SEQ_MODE=4'b1000;
    defparam shift_srl_151_1_LC_15_16_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_151_1_LC_15_16_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63178),
            .lcout(shift_srl_151Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93062),
            .ce(N__63358),
            .sr(_gnd_net_));
    defparam shift_srl_151_2_LC_15_16_2.C_ON=1'b0;
    defparam shift_srl_151_2_LC_15_16_2.SEQ_MODE=4'b1000;
    defparam shift_srl_151_2_LC_15_16_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_151_2_LC_15_16_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63172),
            .lcout(shift_srl_151Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93062),
            .ce(N__63358),
            .sr(_gnd_net_));
    defparam shift_srl_151_3_LC_15_16_3.C_ON=1'b0;
    defparam shift_srl_151_3_LC_15_16_3.SEQ_MODE=4'b1000;
    defparam shift_srl_151_3_LC_15_16_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_151_3_LC_15_16_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63307),
            .lcout(shift_srl_151Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93062),
            .ce(N__63358),
            .sr(_gnd_net_));
    defparam shift_srl_151_4_LC_15_16_4.C_ON=1'b0;
    defparam shift_srl_151_4_LC_15_16_4.SEQ_MODE=4'b1000;
    defparam shift_srl_151_4_LC_15_16_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_151_4_LC_15_16_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63301),
            .lcout(shift_srl_151Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93062),
            .ce(N__63358),
            .sr(_gnd_net_));
    defparam shift_srl_151_5_LC_15_16_5.C_ON=1'b0;
    defparam shift_srl_151_5_LC_15_16_5.SEQ_MODE=4'b1000;
    defparam shift_srl_151_5_LC_15_16_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_151_5_LC_15_16_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63295),
            .lcout(shift_srl_151Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93062),
            .ce(N__63358),
            .sr(_gnd_net_));
    defparam shift_srl_151_6_LC_15_16_6.C_ON=1'b0;
    defparam shift_srl_151_6_LC_15_16_6.SEQ_MODE=4'b1000;
    defparam shift_srl_151_6_LC_15_16_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_151_6_LC_15_16_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63289),
            .lcout(shift_srl_151Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93062),
            .ce(N__63358),
            .sr(_gnd_net_));
    defparam shift_srl_151_7_LC_15_16_7.C_ON=1'b0;
    defparam shift_srl_151_7_LC_15_16_7.SEQ_MODE=4'b1000;
    defparam shift_srl_151_7_LC_15_16_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_151_7_LC_15_16_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63283),
            .lcout(shift_srl_151Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93062),
            .ce(N__63358),
            .sr(_gnd_net_));
    defparam shift_srl_151_10_LC_15_17_0.C_ON=1'b0;
    defparam shift_srl_151_10_LC_15_17_0.SEQ_MODE=4'b1000;
    defparam shift_srl_151_10_LC_15_17_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_151_10_LC_15_17_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63376),
            .lcout(shift_srl_151Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93038),
            .ce(N__63357),
            .sr(_gnd_net_));
    defparam shift_srl_151_11_LC_15_17_1.C_ON=1'b0;
    defparam shift_srl_151_11_LC_15_17_1.SEQ_MODE=4'b1000;
    defparam shift_srl_151_11_LC_15_17_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_151_11_LC_15_17_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63277),
            .lcout(shift_srl_151Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93038),
            .ce(N__63357),
            .sr(_gnd_net_));
    defparam shift_srl_151_12_LC_15_17_2.C_ON=1'b0;
    defparam shift_srl_151_12_LC_15_17_2.SEQ_MODE=4'b1000;
    defparam shift_srl_151_12_LC_15_17_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_151_12_LC_15_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63271),
            .lcout(shift_srl_151Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93038),
            .ce(N__63357),
            .sr(_gnd_net_));
    defparam shift_srl_151_13_LC_15_17_3.C_ON=1'b0;
    defparam shift_srl_151_13_LC_15_17_3.SEQ_MODE=4'b1000;
    defparam shift_srl_151_13_LC_15_17_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_151_13_LC_15_17_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63265),
            .lcout(shift_srl_151Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93038),
            .ce(N__63357),
            .sr(_gnd_net_));
    defparam shift_srl_151_14_LC_15_17_4.C_ON=1'b0;
    defparam shift_srl_151_14_LC_15_17_4.SEQ_MODE=4'b1000;
    defparam shift_srl_151_14_LC_15_17_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_151_14_LC_15_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63439),
            .lcout(shift_srl_151Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93038),
            .ce(N__63357),
            .sr(_gnd_net_));
    defparam shift_srl_151_15_LC_15_17_5.C_ON=1'b0;
    defparam shift_srl_151_15_LC_15_17_5.SEQ_MODE=4'b1000;
    defparam shift_srl_151_15_LC_15_17_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_151_15_LC_15_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63433),
            .lcout(shift_srl_151Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93038),
            .ce(N__63357),
            .sr(_gnd_net_));
    defparam shift_srl_151_9_LC_15_17_6.C_ON=1'b0;
    defparam shift_srl_151_9_LC_15_17_6.SEQ_MODE=4'b1000;
    defparam shift_srl_151_9_LC_15_17_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_151_9_LC_15_17_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63364),
            .lcout(shift_srl_151Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93038),
            .ce(N__63357),
            .sr(_gnd_net_));
    defparam shift_srl_151_8_LC_15_17_7.C_ON=1'b0;
    defparam shift_srl_151_8_LC_15_17_7.SEQ_MODE=4'b1000;
    defparam shift_srl_151_8_LC_15_17_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_151_8_LC_15_17_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63370),
            .lcout(shift_srl_151Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93038),
            .ce(N__63357),
            .sr(_gnd_net_));
    defparam shift_srl_140_10_LC_15_18_0.C_ON=1'b0;
    defparam shift_srl_140_10_LC_15_18_0.SEQ_MODE=4'b1000;
    defparam shift_srl_140_10_LC_15_18_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_140_10_LC_15_18_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63487),
            .lcout(shift_srl_140Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93063),
            .ce(N__63622),
            .sr(_gnd_net_));
    defparam shift_srl_140_11_LC_15_18_1.C_ON=1'b0;
    defparam shift_srl_140_11_LC_15_18_1.SEQ_MODE=4'b1000;
    defparam shift_srl_140_11_LC_15_18_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_140_11_LC_15_18_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63331),
            .lcout(shift_srl_140Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93063),
            .ce(N__63622),
            .sr(_gnd_net_));
    defparam shift_srl_140_12_LC_15_18_2.C_ON=1'b0;
    defparam shift_srl_140_12_LC_15_18_2.SEQ_MODE=4'b1000;
    defparam shift_srl_140_12_LC_15_18_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_140_12_LC_15_18_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63325),
            .lcout(shift_srl_140Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93063),
            .ce(N__63622),
            .sr(_gnd_net_));
    defparam shift_srl_140_13_LC_15_18_3.C_ON=1'b0;
    defparam shift_srl_140_13_LC_15_18_3.SEQ_MODE=4'b1000;
    defparam shift_srl_140_13_LC_15_18_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_140_13_LC_15_18_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63319),
            .lcout(shift_srl_140Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93063),
            .ce(N__63622),
            .sr(_gnd_net_));
    defparam shift_srl_140_14_LC_15_18_4.C_ON=1'b0;
    defparam shift_srl_140_14_LC_15_18_4.SEQ_MODE=4'b1000;
    defparam shift_srl_140_14_LC_15_18_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_140_14_LC_15_18_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63313),
            .lcout(shift_srl_140Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93063),
            .ce(N__63622),
            .sr(_gnd_net_));
    defparam shift_srl_140_15_LC_15_18_5.C_ON=1'b0;
    defparam shift_srl_140_15_LC_15_18_5.SEQ_MODE=4'b1000;
    defparam shift_srl_140_15_LC_15_18_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_140_15_LC_15_18_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63493),
            .lcout(shift_srl_140Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93063),
            .ce(N__63622),
            .sr(_gnd_net_));
    defparam shift_srl_140_9_LC_15_18_6.C_ON=1'b0;
    defparam shift_srl_140_9_LC_15_18_6.SEQ_MODE=4'b1000;
    defparam shift_srl_140_9_LC_15_18_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_140_9_LC_15_18_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63481),
            .lcout(shift_srl_140Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93063),
            .ce(N__63622),
            .sr(_gnd_net_));
    defparam shift_srl_140_8_LC_15_18_7.C_ON=1'b0;
    defparam shift_srl_140_8_LC_15_18_7.SEQ_MODE=4'b1000;
    defparam shift_srl_140_8_LC_15_18_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_140_8_LC_15_18_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63628),
            .lcout(shift_srl_140Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93063),
            .ce(N__63622),
            .sr(_gnd_net_));
    defparam shift_srl_140_0_LC_15_19_0.C_ON=1'b0;
    defparam shift_srl_140_0_LC_15_19_0.SEQ_MODE=4'b1000;
    defparam shift_srl_140_0_LC_15_19_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_140_0_LC_15_19_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64879),
            .lcout(shift_srl_140Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93078),
            .ce(N__63621),
            .sr(_gnd_net_));
    defparam shift_srl_140_1_LC_15_19_1.C_ON=1'b0;
    defparam shift_srl_140_1_LC_15_19_1.SEQ_MODE=4'b1000;
    defparam shift_srl_140_1_LC_15_19_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_140_1_LC_15_19_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63475),
            .lcout(shift_srl_140Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93078),
            .ce(N__63621),
            .sr(_gnd_net_));
    defparam shift_srl_140_2_LC_15_19_2.C_ON=1'b0;
    defparam shift_srl_140_2_LC_15_19_2.SEQ_MODE=4'b1000;
    defparam shift_srl_140_2_LC_15_19_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_140_2_LC_15_19_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63469),
            .lcout(shift_srl_140Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93078),
            .ce(N__63621),
            .sr(_gnd_net_));
    defparam shift_srl_140_3_LC_15_19_3.C_ON=1'b0;
    defparam shift_srl_140_3_LC_15_19_3.SEQ_MODE=4'b1000;
    defparam shift_srl_140_3_LC_15_19_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_140_3_LC_15_19_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63463),
            .lcout(shift_srl_140Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93078),
            .ce(N__63621),
            .sr(_gnd_net_));
    defparam shift_srl_140_4_LC_15_19_4.C_ON=1'b0;
    defparam shift_srl_140_4_LC_15_19_4.SEQ_MODE=4'b1000;
    defparam shift_srl_140_4_LC_15_19_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_140_4_LC_15_19_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63457),
            .lcout(shift_srl_140Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93078),
            .ce(N__63621),
            .sr(_gnd_net_));
    defparam shift_srl_140_5_LC_15_19_5.C_ON=1'b0;
    defparam shift_srl_140_5_LC_15_19_5.SEQ_MODE=4'b1000;
    defparam shift_srl_140_5_LC_15_19_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_140_5_LC_15_19_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63451),
            .lcout(shift_srl_140Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93078),
            .ce(N__63621),
            .sr(_gnd_net_));
    defparam shift_srl_140_6_LC_15_19_6.C_ON=1'b0;
    defparam shift_srl_140_6_LC_15_19_6.SEQ_MODE=4'b1000;
    defparam shift_srl_140_6_LC_15_19_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_140_6_LC_15_19_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63445),
            .lcout(shift_srl_140Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93078),
            .ce(N__63621),
            .sr(_gnd_net_));
    defparam shift_srl_140_7_LC_15_19_7.C_ON=1'b0;
    defparam shift_srl_140_7_LC_15_19_7.SEQ_MODE=4'b1000;
    defparam shift_srl_140_7_LC_15_19_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_140_7_LC_15_19_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63634),
            .lcout(shift_srl_140Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93078),
            .ce(N__63621),
            .sr(_gnd_net_));
    defparam shift_srl_145_0_LC_15_20_0.C_ON=1'b0;
    defparam shift_srl_145_0_LC_15_20_0.SEQ_MODE=4'b1000;
    defparam shift_srl_145_0_LC_15_20_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_145_0_LC_15_20_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63583),
            .lcout(shift_srl_145Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93093),
            .ce(N__63514),
            .sr(_gnd_net_));
    defparam shift_srl_145_1_LC_15_20_1.C_ON=1'b0;
    defparam shift_srl_145_1_LC_15_20_1.SEQ_MODE=4'b1000;
    defparam shift_srl_145_1_LC_15_20_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_145_1_LC_15_20_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63562),
            .lcout(shift_srl_145Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93093),
            .ce(N__63514),
            .sr(_gnd_net_));
    defparam shift_srl_145_2_LC_15_20_2.C_ON=1'b0;
    defparam shift_srl_145_2_LC_15_20_2.SEQ_MODE=4'b1000;
    defparam shift_srl_145_2_LC_15_20_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_145_2_LC_15_20_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63556),
            .lcout(shift_srl_145Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93093),
            .ce(N__63514),
            .sr(_gnd_net_));
    defparam shift_srl_145_3_LC_15_20_3.C_ON=1'b0;
    defparam shift_srl_145_3_LC_15_20_3.SEQ_MODE=4'b1000;
    defparam shift_srl_145_3_LC_15_20_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_145_3_LC_15_20_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63550),
            .lcout(shift_srl_145Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93093),
            .ce(N__63514),
            .sr(_gnd_net_));
    defparam shift_srl_145_4_LC_15_20_4.C_ON=1'b0;
    defparam shift_srl_145_4_LC_15_20_4.SEQ_MODE=4'b1000;
    defparam shift_srl_145_4_LC_15_20_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_145_4_LC_15_20_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63544),
            .lcout(shift_srl_145Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93093),
            .ce(N__63514),
            .sr(_gnd_net_));
    defparam shift_srl_145_5_LC_15_20_5.C_ON=1'b0;
    defparam shift_srl_145_5_LC_15_20_5.SEQ_MODE=4'b1000;
    defparam shift_srl_145_5_LC_15_20_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_145_5_LC_15_20_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63538),
            .lcout(shift_srl_145Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93093),
            .ce(N__63514),
            .sr(_gnd_net_));
    defparam shift_srl_145_6_LC_15_20_6.C_ON=1'b0;
    defparam shift_srl_145_6_LC_15_20_6.SEQ_MODE=4'b1000;
    defparam shift_srl_145_6_LC_15_20_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_145_6_LC_15_20_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63532),
            .lcout(shift_srl_145Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93093),
            .ce(N__63514),
            .sr(_gnd_net_));
    defparam shift_srl_145_7_LC_15_20_7.C_ON=1'b0;
    defparam shift_srl_145_7_LC_15_20_7.SEQ_MODE=4'b1000;
    defparam shift_srl_145_7_LC_15_20_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_145_7_LC_15_20_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63526),
            .lcout(shift_srl_145Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93093),
            .ce(N__63514),
            .sr(_gnd_net_));
    defparam shift_srl_142_0_LC_15_21_0.C_ON=1'b0;
    defparam shift_srl_142_0_LC_15_21_0.SEQ_MODE=4'b1000;
    defparam shift_srl_142_0_LC_15_21_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_142_0_LC_15_21_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63748),
            .lcout(shift_srl_142Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93109),
            .ce(N__63654),
            .sr(_gnd_net_));
    defparam shift_srl_142_1_LC_15_21_1.C_ON=1'b0;
    defparam shift_srl_142_1_LC_15_21_1.SEQ_MODE=4'b1000;
    defparam shift_srl_142_1_LC_15_21_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_142_1_LC_15_21_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63706),
            .lcout(shift_srl_142Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93109),
            .ce(N__63654),
            .sr(_gnd_net_));
    defparam shift_srl_142_2_LC_15_21_2.C_ON=1'b0;
    defparam shift_srl_142_2_LC_15_21_2.SEQ_MODE=4'b1000;
    defparam shift_srl_142_2_LC_15_21_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_142_2_LC_15_21_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63700),
            .lcout(shift_srl_142Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93109),
            .ce(N__63654),
            .sr(_gnd_net_));
    defparam shift_srl_142_3_LC_15_21_3.C_ON=1'b0;
    defparam shift_srl_142_3_LC_15_21_3.SEQ_MODE=4'b1000;
    defparam shift_srl_142_3_LC_15_21_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_142_3_LC_15_21_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63694),
            .lcout(shift_srl_142Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93109),
            .ce(N__63654),
            .sr(_gnd_net_));
    defparam shift_srl_142_4_LC_15_21_4.C_ON=1'b0;
    defparam shift_srl_142_4_LC_15_21_4.SEQ_MODE=4'b1000;
    defparam shift_srl_142_4_LC_15_21_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_142_4_LC_15_21_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63688),
            .lcout(shift_srl_142Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93109),
            .ce(N__63654),
            .sr(_gnd_net_));
    defparam shift_srl_142_5_LC_15_21_5.C_ON=1'b0;
    defparam shift_srl_142_5_LC_15_21_5.SEQ_MODE=4'b1000;
    defparam shift_srl_142_5_LC_15_21_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_142_5_LC_15_21_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63682),
            .lcout(shift_srl_142Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93109),
            .ce(N__63654),
            .sr(_gnd_net_));
    defparam shift_srl_142_6_LC_15_21_6.C_ON=1'b0;
    defparam shift_srl_142_6_LC_15_21_6.SEQ_MODE=4'b1000;
    defparam shift_srl_142_6_LC_15_21_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_142_6_LC_15_21_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63676),
            .lcout(shift_srl_142Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93109),
            .ce(N__63654),
            .sr(_gnd_net_));
    defparam shift_srl_142_7_LC_15_21_7.C_ON=1'b0;
    defparam shift_srl_142_7_LC_15_21_7.SEQ_MODE=4'b1000;
    defparam shift_srl_142_7_LC_15_21_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_142_7_LC_15_21_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63670),
            .lcout(shift_srl_142Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93109),
            .ce(N__63654),
            .sr(_gnd_net_));
    defparam shift_srl_120_10_LC_15_22_0.C_ON=1'b0;
    defparam shift_srl_120_10_LC_15_22_0.SEQ_MODE=4'b1000;
    defparam shift_srl_120_10_LC_15_22_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_120_10_LC_15_22_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63892),
            .lcout(shift_srl_120Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93127),
            .ce(N__65191),
            .sr(_gnd_net_));
    defparam shift_srl_120_11_LC_15_22_1.C_ON=1'b0;
    defparam shift_srl_120_11_LC_15_22_1.SEQ_MODE=4'b1000;
    defparam shift_srl_120_11_LC_15_22_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_120_11_LC_15_22_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63922),
            .lcout(shift_srl_120Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93127),
            .ce(N__65191),
            .sr(_gnd_net_));
    defparam shift_srl_120_12_LC_15_22_2.C_ON=1'b0;
    defparam shift_srl_120_12_LC_15_22_2.SEQ_MODE=4'b1000;
    defparam shift_srl_120_12_LC_15_22_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_120_12_LC_15_22_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63916),
            .lcout(shift_srl_120Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93127),
            .ce(N__65191),
            .sr(_gnd_net_));
    defparam shift_srl_120_13_LC_15_22_3.C_ON=1'b0;
    defparam shift_srl_120_13_LC_15_22_3.SEQ_MODE=4'b1000;
    defparam shift_srl_120_13_LC_15_22_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_120_13_LC_15_22_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63910),
            .lcout(shift_srl_120Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93127),
            .ce(N__65191),
            .sr(_gnd_net_));
    defparam shift_srl_120_14_LC_15_22_4.C_ON=1'b0;
    defparam shift_srl_120_14_LC_15_22_4.SEQ_MODE=4'b1000;
    defparam shift_srl_120_14_LC_15_22_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_120_14_LC_15_22_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63904),
            .lcout(shift_srl_120Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93127),
            .ce(N__65191),
            .sr(_gnd_net_));
    defparam shift_srl_120_15_LC_15_22_5.C_ON=1'b0;
    defparam shift_srl_120_15_LC_15_22_5.SEQ_MODE=4'b1000;
    defparam shift_srl_120_15_LC_15_22_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_120_15_LC_15_22_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63898),
            .lcout(shift_srl_120Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93127),
            .ce(N__65191),
            .sr(_gnd_net_));
    defparam shift_srl_120_9_LC_15_22_6.C_ON=1'b0;
    defparam shift_srl_120_9_LC_15_22_6.SEQ_MODE=4'b1000;
    defparam shift_srl_120_9_LC_15_22_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_120_9_LC_15_22_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63886),
            .lcout(shift_srl_120Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93127),
            .ce(N__65191),
            .sr(_gnd_net_));
    defparam shift_srl_120_8_LC_15_22_7.C_ON=1'b0;
    defparam shift_srl_120_8_LC_15_22_7.SEQ_MODE=4'b1000;
    defparam shift_srl_120_8_LC_15_22_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_120_8_LC_15_22_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65113),
            .lcout(shift_srl_120Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93127),
            .ce(N__65191),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_115_LC_15_23_0.C_ON=1'b0;
    defparam rco_obuf_RNO_115_LC_15_23_0.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_115_LC_15_23_0.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_115_LC_15_23_0 (
            .in0(N__63835),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63873),
            .lcout(rco_c_115),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_115_0_LC_15_23_1.C_ON=1'b0;
    defparam shift_srl_115_0_LC_15_23_1.SEQ_MODE=4'b1000;
    defparam shift_srl_115_0_LC_15_23_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_115_0_LC_15_23_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63834),
            .lcout(shift_srl_115Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93146),
            .ce(N__64073),
            .sr(_gnd_net_));
    defparam shift_srl_115_1_LC_15_23_2.C_ON=1'b0;
    defparam shift_srl_115_1_LC_15_23_2.SEQ_MODE=4'b1000;
    defparam shift_srl_115_1_LC_15_23_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_115_1_LC_15_23_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63970),
            .lcout(shift_srl_115Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93146),
            .ce(N__64073),
            .sr(_gnd_net_));
    defparam shift_srl_115_2_LC_15_23_3.C_ON=1'b0;
    defparam shift_srl_115_2_LC_15_23_3.SEQ_MODE=4'b1000;
    defparam shift_srl_115_2_LC_15_23_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_115_2_LC_15_23_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63964),
            .lcout(shift_srl_115Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93146),
            .ce(N__64073),
            .sr(_gnd_net_));
    defparam shift_srl_115_3_LC_15_23_4.C_ON=1'b0;
    defparam shift_srl_115_3_LC_15_23_4.SEQ_MODE=4'b1000;
    defparam shift_srl_115_3_LC_15_23_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_115_3_LC_15_23_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63958),
            .lcout(shift_srl_115Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93146),
            .ce(N__64073),
            .sr(_gnd_net_));
    defparam shift_srl_115_4_LC_15_23_5.C_ON=1'b0;
    defparam shift_srl_115_4_LC_15_23_5.SEQ_MODE=4'b1000;
    defparam shift_srl_115_4_LC_15_23_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_115_4_LC_15_23_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63952),
            .lcout(shift_srl_115Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93146),
            .ce(N__64073),
            .sr(_gnd_net_));
    defparam shift_srl_115_5_LC_15_23_6.C_ON=1'b0;
    defparam shift_srl_115_5_LC_15_23_6.SEQ_MODE=4'b1000;
    defparam shift_srl_115_5_LC_15_23_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_115_5_LC_15_23_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63946),
            .lcout(shift_srl_115Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93146),
            .ce(N__64073),
            .sr(_gnd_net_));
    defparam shift_srl_115_6_LC_15_23_7.C_ON=1'b0;
    defparam shift_srl_115_6_LC_15_23_7.SEQ_MODE=4'b1000;
    defparam shift_srl_115_6_LC_15_23_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_115_6_LC_15_23_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63940),
            .lcout(shift_srl_115Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93146),
            .ce(N__64073),
            .sr(_gnd_net_));
    defparam shift_srl_115_10_LC_15_24_0.C_ON=1'b0;
    defparam shift_srl_115_10_LC_15_24_0.SEQ_MODE=4'b1000;
    defparam shift_srl_115_10_LC_15_24_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_115_10_LC_15_24_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64108),
            .lcout(shift_srl_115Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93163),
            .ce(N__64080),
            .sr(_gnd_net_));
    defparam shift_srl_115_11_LC_15_24_1.C_ON=1'b0;
    defparam shift_srl_115_11_LC_15_24_1.SEQ_MODE=4'b1000;
    defparam shift_srl_115_11_LC_15_24_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_115_11_LC_15_24_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63934),
            .lcout(shift_srl_115Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93163),
            .ce(N__64080),
            .sr(_gnd_net_));
    defparam shift_srl_115_12_LC_15_24_2.C_ON=1'b0;
    defparam shift_srl_115_12_LC_15_24_2.SEQ_MODE=4'b1000;
    defparam shift_srl_115_12_LC_15_24_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_115_12_LC_15_24_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63928),
            .lcout(shift_srl_115Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93163),
            .ce(N__64080),
            .sr(_gnd_net_));
    defparam shift_srl_115_13_LC_15_24_3.C_ON=1'b0;
    defparam shift_srl_115_13_LC_15_24_3.SEQ_MODE=4'b1000;
    defparam shift_srl_115_13_LC_15_24_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_115_13_LC_15_24_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64135),
            .lcout(shift_srl_115Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93163),
            .ce(N__64080),
            .sr(_gnd_net_));
    defparam shift_srl_115_14_LC_15_24_4.C_ON=1'b0;
    defparam shift_srl_115_14_LC_15_24_4.SEQ_MODE=4'b1000;
    defparam shift_srl_115_14_LC_15_24_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_115_14_LC_15_24_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64129),
            .lcout(shift_srl_115Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93163),
            .ce(N__64080),
            .sr(_gnd_net_));
    defparam shift_srl_115_9_LC_15_24_5.C_ON=1'b0;
    defparam shift_srl_115_9_LC_15_24_5.SEQ_MODE=4'b1000;
    defparam shift_srl_115_9_LC_15_24_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_115_9_LC_15_24_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64102),
            .lcout(shift_srl_115Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93163),
            .ce(N__64080),
            .sr(_gnd_net_));
    defparam shift_srl_115_8_LC_15_24_6.C_ON=1'b0;
    defparam shift_srl_115_8_LC_15_24_6.SEQ_MODE=4'b1000;
    defparam shift_srl_115_8_LC_15_24_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_115_8_LC_15_24_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64090),
            .lcout(shift_srl_115Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93163),
            .ce(N__64080),
            .sr(_gnd_net_));
    defparam shift_srl_115_7_LC_15_24_7.C_ON=1'b0;
    defparam shift_srl_115_7_LC_15_24_7.SEQ_MODE=4'b1000;
    defparam shift_srl_115_7_LC_15_24_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_115_7_LC_15_24_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64096),
            .lcout(shift_srl_115Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93163),
            .ce(N__64080),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_194_LC_15_25_0.C_ON=1'b0;
    defparam rco_obuf_RNO_194_LC_15_25_0.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_194_LC_15_25_0.LUT_INIT=16'b1000100000000000;
    LogicCell40 rco_obuf_RNO_194_LC_15_25_0 (
            .in0(N__73864),
            .in1(N__91531),
            .in2(_gnd_net_),
            .in3(N__73903),
            .lcout(rco_c_194),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_193_LC_15_25_1.C_ON=1'b0;
    defparam rco_obuf_RNO_193_LC_15_25_1.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_193_LC_15_25_1.LUT_INIT=16'b1000100010001000;
    LogicCell40 rco_obuf_RNO_193_LC_15_25_1 (
            .in0(N__91530),
            .in1(N__73863),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(rco_c_193),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_184_LC_15_25_2.C_ON=1'b0;
    defparam rco_obuf_RNO_184_LC_15_25_2.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_184_LC_15_25_2.LUT_INIT=16'b1100110000000000;
    LogicCell40 rco_obuf_RNO_184_LC_15_25_2 (
            .in0(_gnd_net_),
            .in1(N__91528),
            .in2(_gnd_net_),
            .in3(N__91691),
            .lcout(rco_c_184),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_187_LC_15_25_3.C_ON=1'b0;
    defparam rco_obuf_RNO_187_LC_15_25_3.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_187_LC_15_25_3.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_187_LC_15_25_3 (
            .in0(N__80359),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__91532),
            .lcout(rco_c_187),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_191_LC_15_25_4.C_ON=1'b0;
    defparam rco_obuf_RNO_191_LC_15_25_4.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_191_LC_15_25_4.LUT_INIT=16'b1100110000000000;
    LogicCell40 rco_obuf_RNO_191_LC_15_25_4 (
            .in0(_gnd_net_),
            .in1(N__91529),
            .in2(_gnd_net_),
            .in3(N__74260),
            .lcout(rco_c_191),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_195_LC_15_25_5.C_ON=1'b0;
    defparam rco_obuf_RNO_195_LC_15_25_5.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_195_LC_15_25_5.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_195_LC_15_25_5 (
            .in0(N__73834),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__91533),
            .lcout(rco_c_195),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_194_0_LC_15_25_6.C_ON=1'b0;
    defparam shift_srl_194_0_LC_15_25_6.SEQ_MODE=4'b1000;
    defparam shift_srl_194_0_LC_15_25_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_194_0_LC_15_25_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73902),
            .lcout(shift_srl_194Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93183),
            .ce(N__72265),
            .sr(_gnd_net_));
    defparam shift_srl_194_1_LC_15_25_7.C_ON=1'b0;
    defparam shift_srl_194_1_LC_15_25_7.SEQ_MODE=4'b1000;
    defparam shift_srl_194_1_LC_15_25_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_194_1_LC_15_25_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64174),
            .lcout(shift_srl_194Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93183),
            .ce(N__72265),
            .sr(_gnd_net_));
    defparam shift_srl_139_12_LC_15_28_2.C_ON=1'b0;
    defparam shift_srl_139_12_LC_15_28_2.SEQ_MODE=4'b1000;
    defparam shift_srl_139_12_LC_15_28_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_139_12_LC_15_28_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64168),
            .lcout(shift_srl_139Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93243),
            .ce(N__64828),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_90_LC_16_3_1.C_ON=1'b0;
    defparam rco_obuf_RNO_90_LC_16_3_1.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_90_LC_16_3_1.LUT_INIT=16'b1000100000000000;
    LogicCell40 rco_obuf_RNO_90_LC_16_3_1 (
            .in0(N__66914),
            .in1(N__68611),
            .in2(_gnd_net_),
            .in3(N__68519),
            .lcout(rco_c_90),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_91_LC_16_3_7.C_ON=1'b0;
    defparam rco_obuf_RNO_91_LC_16_3_7.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_91_LC_16_3_7.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_91_LC_16_3_7 (
            .in0(N__72111),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68520),
            .lcout(rco_c_91),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_94_8_LC_16_4_2.C_ON=1'b0;
    defparam shift_srl_94_8_LC_16_4_2.SEQ_MODE=4'b1000;
    defparam shift_srl_94_8_LC_16_4_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_94_8_LC_16_4_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66643),
            .lcout(shift_srl_94Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93300),
            .ce(N__72650),
            .sr(_gnd_net_));
    defparam shift_srl_85_0_LC_16_5_0.C_ON=1'b0;
    defparam shift_srl_85_0_LC_16_5_0.SEQ_MODE=4'b1000;
    defparam shift_srl_85_0_LC_16_5_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_85_0_LC_16_5_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67047),
            .lcout(shift_srl_85Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93284),
            .ce(N__64243),
            .sr(_gnd_net_));
    defparam shift_srl_85_1_LC_16_5_1.C_ON=1'b0;
    defparam shift_srl_85_1_LC_16_5_1.SEQ_MODE=4'b1000;
    defparam shift_srl_85_1_LC_16_5_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_85_1_LC_16_5_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64291),
            .lcout(shift_srl_85Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93284),
            .ce(N__64243),
            .sr(_gnd_net_));
    defparam shift_srl_85_2_LC_16_5_2.C_ON=1'b0;
    defparam shift_srl_85_2_LC_16_5_2.SEQ_MODE=4'b1000;
    defparam shift_srl_85_2_LC_16_5_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_85_2_LC_16_5_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64285),
            .lcout(shift_srl_85Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93284),
            .ce(N__64243),
            .sr(_gnd_net_));
    defparam shift_srl_85_3_LC_16_5_3.C_ON=1'b0;
    defparam shift_srl_85_3_LC_16_5_3.SEQ_MODE=4'b1000;
    defparam shift_srl_85_3_LC_16_5_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_85_3_LC_16_5_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64279),
            .lcout(shift_srl_85Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93284),
            .ce(N__64243),
            .sr(_gnd_net_));
    defparam shift_srl_85_4_LC_16_5_4.C_ON=1'b0;
    defparam shift_srl_85_4_LC_16_5_4.SEQ_MODE=4'b1000;
    defparam shift_srl_85_4_LC_16_5_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_85_4_LC_16_5_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64273),
            .lcout(shift_srl_85Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93284),
            .ce(N__64243),
            .sr(_gnd_net_));
    defparam shift_srl_85_5_LC_16_5_5.C_ON=1'b0;
    defparam shift_srl_85_5_LC_16_5_5.SEQ_MODE=4'b1000;
    defparam shift_srl_85_5_LC_16_5_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_85_5_LC_16_5_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64267),
            .lcout(shift_srl_85Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93284),
            .ce(N__64243),
            .sr(_gnd_net_));
    defparam shift_srl_85_6_LC_16_5_6.C_ON=1'b0;
    defparam shift_srl_85_6_LC_16_5_6.SEQ_MODE=4'b1000;
    defparam shift_srl_85_6_LC_16_5_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_85_6_LC_16_5_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64261),
            .lcout(shift_srl_85Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93284),
            .ce(N__64243),
            .sr(_gnd_net_));
    defparam shift_srl_85_7_LC_16_5_7.C_ON=1'b0;
    defparam shift_srl_85_7_LC_16_5_7.SEQ_MODE=4'b1000;
    defparam shift_srl_85_7_LC_16_5_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_85_7_LC_16_5_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64255),
            .lcout(shift_srl_85Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93284),
            .ce(N__64243),
            .sr(_gnd_net_));
    defparam shift_srl_88_0_LC_16_6_0.C_ON=1'b0;
    defparam shift_srl_88_0_LC_16_6_0.SEQ_MODE=4'b1000;
    defparam shift_srl_88_0_LC_16_6_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_88_0_LC_16_6_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66973),
            .lcout(shift_srl_88Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93265),
            .ce(N__64327),
            .sr(_gnd_net_));
    defparam shift_srl_88_1_LC_16_6_1.C_ON=1'b0;
    defparam shift_srl_88_1_LC_16_6_1.SEQ_MODE=4'b1000;
    defparam shift_srl_88_1_LC_16_6_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_88_1_LC_16_6_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64222),
            .lcout(shift_srl_88Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93265),
            .ce(N__64327),
            .sr(_gnd_net_));
    defparam shift_srl_88_2_LC_16_6_2.C_ON=1'b0;
    defparam shift_srl_88_2_LC_16_6_2.SEQ_MODE=4'b1000;
    defparam shift_srl_88_2_LC_16_6_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_88_2_LC_16_6_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64369),
            .lcout(shift_srl_88Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93265),
            .ce(N__64327),
            .sr(_gnd_net_));
    defparam shift_srl_88_3_LC_16_6_3.C_ON=1'b0;
    defparam shift_srl_88_3_LC_16_6_3.SEQ_MODE=4'b1000;
    defparam shift_srl_88_3_LC_16_6_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_88_3_LC_16_6_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64363),
            .lcout(shift_srl_88Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93265),
            .ce(N__64327),
            .sr(_gnd_net_));
    defparam shift_srl_88_4_LC_16_6_4.C_ON=1'b0;
    defparam shift_srl_88_4_LC_16_6_4.SEQ_MODE=4'b1000;
    defparam shift_srl_88_4_LC_16_6_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_88_4_LC_16_6_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64357),
            .lcout(shift_srl_88Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93265),
            .ce(N__64327),
            .sr(_gnd_net_));
    defparam shift_srl_88_5_LC_16_6_5.C_ON=1'b0;
    defparam shift_srl_88_5_LC_16_6_5.SEQ_MODE=4'b1000;
    defparam shift_srl_88_5_LC_16_6_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_88_5_LC_16_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64351),
            .lcout(shift_srl_88Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93265),
            .ce(N__64327),
            .sr(_gnd_net_));
    defparam shift_srl_88_6_LC_16_6_6.C_ON=1'b0;
    defparam shift_srl_88_6_LC_16_6_6.SEQ_MODE=4'b1000;
    defparam shift_srl_88_6_LC_16_6_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_88_6_LC_16_6_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64345),
            .lcout(shift_srl_88Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93265),
            .ce(N__64327),
            .sr(_gnd_net_));
    defparam shift_srl_88_7_LC_16_6_7.C_ON=1'b0;
    defparam shift_srl_88_7_LC_16_6_7.SEQ_MODE=4'b1000;
    defparam shift_srl_88_7_LC_16_6_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_88_7_LC_16_6_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64339),
            .lcout(shift_srl_88Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93265),
            .ce(N__64327),
            .sr(_gnd_net_));
    defparam shift_srl_87_0_LC_16_7_0.C_ON=1'b0;
    defparam shift_srl_87_0_LC_16_7_0.SEQ_MODE=4'b1000;
    defparam shift_srl_87_0_LC_16_7_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_87_0_LC_16_7_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67110),
            .lcout(shift_srl_87Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93246),
            .ce(N__64411),
            .sr(_gnd_net_));
    defparam shift_srl_87_1_LC_16_7_1.C_ON=1'b0;
    defparam shift_srl_87_1_LC_16_7_1.SEQ_MODE=4'b1000;
    defparam shift_srl_87_1_LC_16_7_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_87_1_LC_16_7_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64303),
            .lcout(shift_srl_87Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93246),
            .ce(N__64411),
            .sr(_gnd_net_));
    defparam shift_srl_87_2_LC_16_7_2.C_ON=1'b0;
    defparam shift_srl_87_2_LC_16_7_2.SEQ_MODE=4'b1000;
    defparam shift_srl_87_2_LC_16_7_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_87_2_LC_16_7_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64297),
            .lcout(shift_srl_87Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93246),
            .ce(N__64411),
            .sr(_gnd_net_));
    defparam shift_srl_87_3_LC_16_7_3.C_ON=1'b0;
    defparam shift_srl_87_3_LC_16_7_3.SEQ_MODE=4'b1000;
    defparam shift_srl_87_3_LC_16_7_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_87_3_LC_16_7_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64450),
            .lcout(shift_srl_87Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93246),
            .ce(N__64411),
            .sr(_gnd_net_));
    defparam shift_srl_87_4_LC_16_7_4.C_ON=1'b0;
    defparam shift_srl_87_4_LC_16_7_4.SEQ_MODE=4'b1000;
    defparam shift_srl_87_4_LC_16_7_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_87_4_LC_16_7_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64444),
            .lcout(shift_srl_87Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93246),
            .ce(N__64411),
            .sr(_gnd_net_));
    defparam shift_srl_87_5_LC_16_7_5.C_ON=1'b0;
    defparam shift_srl_87_5_LC_16_7_5.SEQ_MODE=4'b1000;
    defparam shift_srl_87_5_LC_16_7_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_87_5_LC_16_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64438),
            .lcout(shift_srl_87Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93246),
            .ce(N__64411),
            .sr(_gnd_net_));
    defparam shift_srl_87_6_LC_16_7_6.C_ON=1'b0;
    defparam shift_srl_87_6_LC_16_7_6.SEQ_MODE=4'b1000;
    defparam shift_srl_87_6_LC_16_7_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_87_6_LC_16_7_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64432),
            .lcout(shift_srl_87Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93246),
            .ce(N__64411),
            .sr(_gnd_net_));
    defparam shift_srl_87_7_LC_16_7_7.C_ON=1'b0;
    defparam shift_srl_87_7_LC_16_7_7.SEQ_MODE=4'b1000;
    defparam shift_srl_87_7_LC_16_7_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_87_7_LC_16_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64426),
            .lcout(shift_srl_87Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93246),
            .ce(N__64411),
            .sr(_gnd_net_));
    defparam shift_srl_99_10_LC_16_8_0.C_ON=1'b0;
    defparam shift_srl_99_10_LC_16_8_0.SEQ_MODE=4'b1000;
    defparam shift_srl_99_10_LC_16_8_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_99_10_LC_16_8_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64504),
            .lcout(shift_srl_99Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93226),
            .ce(N__67640),
            .sr(_gnd_net_));
    defparam shift_srl_99_11_LC_16_8_1.C_ON=1'b0;
    defparam shift_srl_99_11_LC_16_8_1.SEQ_MODE=4'b1000;
    defparam shift_srl_99_11_LC_16_8_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_99_11_LC_16_8_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64393),
            .lcout(shift_srl_99Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93226),
            .ce(N__67640),
            .sr(_gnd_net_));
    defparam shift_srl_99_12_LC_16_8_2.C_ON=1'b0;
    defparam shift_srl_99_12_LC_16_8_2.SEQ_MODE=4'b1000;
    defparam shift_srl_99_12_LC_16_8_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_99_12_LC_16_8_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64387),
            .lcout(shift_srl_99Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93226),
            .ce(N__67640),
            .sr(_gnd_net_));
    defparam shift_srl_99_13_LC_16_8_3.C_ON=1'b0;
    defparam shift_srl_99_13_LC_16_8_3.SEQ_MODE=4'b1000;
    defparam shift_srl_99_13_LC_16_8_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_99_13_LC_16_8_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64381),
            .lcout(shift_srl_99Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93226),
            .ce(N__67640),
            .sr(_gnd_net_));
    defparam shift_srl_99_14_LC_16_8_4.C_ON=1'b0;
    defparam shift_srl_99_14_LC_16_8_4.SEQ_MODE=4'b1000;
    defparam shift_srl_99_14_LC_16_8_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_99_14_LC_16_8_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64375),
            .lcout(shift_srl_99Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93226),
            .ce(N__67640),
            .sr(_gnd_net_));
    defparam shift_srl_99_9_LC_16_8_5.C_ON=1'b0;
    defparam shift_srl_99_9_LC_16_8_5.SEQ_MODE=4'b1000;
    defparam shift_srl_99_9_LC_16_8_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_99_9_LC_16_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64498),
            .lcout(shift_srl_99Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93226),
            .ce(N__67640),
            .sr(_gnd_net_));
    defparam shift_srl_99_8_LC_16_8_6.C_ON=1'b0;
    defparam shift_srl_99_8_LC_16_8_6.SEQ_MODE=4'b1000;
    defparam shift_srl_99_8_LC_16_8_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_99_8_LC_16_8_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64480),
            .lcout(shift_srl_99Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93226),
            .ce(N__67640),
            .sr(_gnd_net_));
    defparam shift_srl_99_7_LC_16_8_7.C_ON=1'b0;
    defparam shift_srl_99_7_LC_16_8_7.SEQ_MODE=4'b1000;
    defparam shift_srl_99_7_LC_16_8_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_99_7_LC_16_8_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64492),
            .lcout(shift_srl_99Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93226),
            .ce(N__67640),
            .sr(_gnd_net_));
    defparam shift_srl_42_6_LC_16_9_0.C_ON=1'b0;
    defparam shift_srl_42_6_LC_16_9_0.SEQ_MODE=4'b1000;
    defparam shift_srl_42_6_LC_16_9_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_42_6_LC_16_9_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64468),
            .lcout(shift_srl_42Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93207),
            .ce(N__67295),
            .sr(_gnd_net_));
    defparam shift_srl_42_7_LC_16_9_1.C_ON=1'b0;
    defparam shift_srl_42_7_LC_16_9_1.SEQ_MODE=4'b1000;
    defparam shift_srl_42_7_LC_16_9_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_42_7_LC_16_9_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64474),
            .lcout(shift_srl_42Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93207),
            .ce(N__67295),
            .sr(_gnd_net_));
    defparam shift_srl_42_5_LC_16_9_7.C_ON=1'b0;
    defparam shift_srl_42_5_LC_16_9_7.SEQ_MODE=4'b1000;
    defparam shift_srl_42_5_LC_16_9_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_42_5_LC_16_9_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64618),
            .lcout(shift_srl_42Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93207),
            .ce(N__67295),
            .sr(_gnd_net_));
    defparam shift_srl_42_10_LC_16_10_0.C_ON=1'b0;
    defparam shift_srl_42_10_LC_16_10_0.SEQ_MODE=4'b1000;
    defparam shift_srl_42_10_LC_16_10_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_42_10_LC_16_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64567),
            .lcout(shift_srl_42Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93185),
            .ce(N__67302),
            .sr(_gnd_net_));
    defparam shift_srl_42_11_LC_16_10_1.C_ON=1'b0;
    defparam shift_srl_42_11_LC_16_10_1.SEQ_MODE=4'b1000;
    defparam shift_srl_42_11_LC_16_10_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_42_11_LC_16_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64462),
            .lcout(shift_srl_42Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93185),
            .ce(N__67302),
            .sr(_gnd_net_));
    defparam shift_srl_42_12_LC_16_10_2.C_ON=1'b0;
    defparam shift_srl_42_12_LC_16_10_2.SEQ_MODE=4'b1000;
    defparam shift_srl_42_12_LC_16_10_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_42_12_LC_16_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64456),
            .lcout(shift_srl_42Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93185),
            .ce(N__67302),
            .sr(_gnd_net_));
    defparam shift_srl_42_13_LC_16_10_3.C_ON=1'b0;
    defparam shift_srl_42_13_LC_16_10_3.SEQ_MODE=4'b1000;
    defparam shift_srl_42_13_LC_16_10_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_42_13_LC_16_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64585),
            .lcout(shift_srl_42Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93185),
            .ce(N__67302),
            .sr(_gnd_net_));
    defparam shift_srl_42_14_LC_16_10_4.C_ON=1'b0;
    defparam shift_srl_42_14_LC_16_10_4.SEQ_MODE=4'b1000;
    defparam shift_srl_42_14_LC_16_10_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_42_14_LC_16_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64579),
            .lcout(shift_srl_42Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93185),
            .ce(N__67302),
            .sr(_gnd_net_));
    defparam shift_srl_42_15_LC_16_10_5.C_ON=1'b0;
    defparam shift_srl_42_15_LC_16_10_5.SEQ_MODE=4'b1000;
    defparam shift_srl_42_15_LC_16_10_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_42_15_LC_16_10_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64573),
            .lcout(shift_srl_42Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93185),
            .ce(N__67302),
            .sr(_gnd_net_));
    defparam shift_srl_42_9_LC_16_10_6.C_ON=1'b0;
    defparam shift_srl_42_9_LC_16_10_6.SEQ_MODE=4'b1000;
    defparam shift_srl_42_9_LC_16_10_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_42_9_LC_16_10_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64555),
            .lcout(shift_srl_42Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93185),
            .ce(N__67302),
            .sr(_gnd_net_));
    defparam shift_srl_42_8_LC_16_10_7.C_ON=1'b0;
    defparam shift_srl_42_8_LC_16_10_7.SEQ_MODE=4'b1000;
    defparam shift_srl_42_8_LC_16_10_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_42_8_LC_16_10_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64561),
            .lcout(shift_srl_42Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93185),
            .ce(N__67302),
            .sr(_gnd_net_));
    defparam shift_srl_59_8_LC_16_11_0.C_ON=1'b0;
    defparam shift_srl_59_8_LC_16_11_0.SEQ_MODE=4'b1000;
    defparam shift_srl_59_8_LC_16_11_0.LUT_INIT=16'b1100110011001100;
    LogicCell40 shift_srl_59_8_LC_16_11_0 (
            .in0(_gnd_net_),
            .in1(N__71269),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_59Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93164),
            .ce(N__73108),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_43_LC_16_12_0.C_ON=1'b0;
    defparam rco_obuf_RNO_43_LC_16_12_0.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_43_LC_16_12_0.LUT_INIT=16'b1000100000000000;
    LogicCell40 rco_obuf_RNO_43_LC_16_12_0 (
            .in0(N__73232),
            .in1(N__69120),
            .in2(_gnd_net_),
            .in3(N__73271),
            .lcout(rco_c_43),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_42_LC_16_12_1.C_ON=1'b0;
    defparam rco_obuf_RNO_42_LC_16_12_1.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_42_LC_16_12_1.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_42_LC_16_12_1 (
            .in0(N__69119),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73231),
            .lcout(rco_c_42),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_42_0_LC_16_12_2.C_ON=1'b0;
    defparam shift_srl_42_0_LC_16_12_2.SEQ_MODE=4'b1000;
    defparam shift_srl_42_0_LC_16_12_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_42_0_LC_16_12_2 (
            .in0(N__73230),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_42Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93147),
            .ce(N__67303),
            .sr(_gnd_net_));
    defparam shift_srl_42_1_LC_16_12_3.C_ON=1'b0;
    defparam shift_srl_42_1_LC_16_12_3.SEQ_MODE=4'b1000;
    defparam shift_srl_42_1_LC_16_12_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_42_1_LC_16_12_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64642),
            .lcout(shift_srl_42Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93147),
            .ce(N__67303),
            .sr(_gnd_net_));
    defparam shift_srl_42_2_LC_16_12_4.C_ON=1'b0;
    defparam shift_srl_42_2_LC_16_12_4.SEQ_MODE=4'b1000;
    defparam shift_srl_42_2_LC_16_12_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_42_2_LC_16_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64636),
            .lcout(shift_srl_42Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93147),
            .ce(N__67303),
            .sr(_gnd_net_));
    defparam shift_srl_42_3_LC_16_12_5.C_ON=1'b0;
    defparam shift_srl_42_3_LC_16_12_5.SEQ_MODE=4'b1000;
    defparam shift_srl_42_3_LC_16_12_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_42_3_LC_16_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64630),
            .lcout(shift_srl_42Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93147),
            .ce(N__67303),
            .sr(_gnd_net_));
    defparam shift_srl_42_4_LC_16_12_6.C_ON=1'b0;
    defparam shift_srl_42_4_LC_16_12_6.SEQ_MODE=4'b1000;
    defparam shift_srl_42_4_LC_16_12_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_42_4_LC_16_12_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64624),
            .lcout(shift_srl_42Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93147),
            .ce(N__67303),
            .sr(_gnd_net_));
    defparam shift_srl_26_10_LC_16_15_0.C_ON=1'b0;
    defparam shift_srl_26_10_LC_16_15_0.SEQ_MODE=4'b1000;
    defparam shift_srl_26_10_LC_16_15_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_26_10_LC_16_15_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64702),
            .lcout(shift_srl_26Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93094),
            .ce(N__64681),
            .sr(_gnd_net_));
    defparam shift_srl_26_11_LC_16_15_1.C_ON=1'b0;
    defparam shift_srl_26_11_LC_16_15_1.SEQ_MODE=4'b1000;
    defparam shift_srl_26_11_LC_16_15_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_26_11_LC_16_15_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64609),
            .lcout(shift_srl_26Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93094),
            .ce(N__64681),
            .sr(_gnd_net_));
    defparam shift_srl_26_12_LC_16_15_2.C_ON=1'b0;
    defparam shift_srl_26_12_LC_16_15_2.SEQ_MODE=4'b1000;
    defparam shift_srl_26_12_LC_16_15_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_26_12_LC_16_15_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64603),
            .lcout(shift_srl_26Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93094),
            .ce(N__64681),
            .sr(_gnd_net_));
    defparam shift_srl_26_13_LC_16_15_3.C_ON=1'b0;
    defparam shift_srl_26_13_LC_16_15_3.SEQ_MODE=4'b1000;
    defparam shift_srl_26_13_LC_16_15_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_26_13_LC_16_15_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64597),
            .lcout(shift_srl_26Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93094),
            .ce(N__64681),
            .sr(_gnd_net_));
    defparam shift_srl_26_14_LC_16_15_4.C_ON=1'b0;
    defparam shift_srl_26_14_LC_16_15_4.SEQ_MODE=4'b1000;
    defparam shift_srl_26_14_LC_16_15_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_26_14_LC_16_15_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64591),
            .lcout(shift_srl_26Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93094),
            .ce(N__64681),
            .sr(_gnd_net_));
    defparam shift_srl_26_15_LC_16_15_5.C_ON=1'b0;
    defparam shift_srl_26_15_LC_16_15_5.SEQ_MODE=4'b1000;
    defparam shift_srl_26_15_LC_16_15_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_26_15_LC_16_15_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64708),
            .lcout(shift_srl_26Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93094),
            .ce(N__64681),
            .sr(_gnd_net_));
    defparam shift_srl_26_9_LC_16_15_6.C_ON=1'b0;
    defparam shift_srl_26_9_LC_16_15_6.SEQ_MODE=4'b1000;
    defparam shift_srl_26_9_LC_16_15_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_26_9_LC_16_15_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64687),
            .lcout(shift_srl_26Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93094),
            .ce(N__64681),
            .sr(_gnd_net_));
    defparam shift_srl_26_8_LC_16_15_7.C_ON=1'b0;
    defparam shift_srl_26_8_LC_16_15_7.SEQ_MODE=4'b1000;
    defparam shift_srl_26_8_LC_16_15_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_26_8_LC_16_15_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64696),
            .lcout(shift_srl_26Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93094),
            .ce(N__64681),
            .sr(_gnd_net_));
    defparam shift_srl_28_10_LC_16_16_0.C_ON=1'b0;
    defparam shift_srl_28_10_LC_16_16_0.SEQ_MODE=4'b1000;
    defparam shift_srl_28_10_LC_16_16_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_28_10_LC_16_16_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64648),
            .lcout(shift_srl_28Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93079),
            .ce(N__67716),
            .sr(_gnd_net_));
    defparam shift_srl_28_0_LC_16_16_1.C_ON=1'b0;
    defparam shift_srl_28_0_LC_16_16_1.SEQ_MODE=4'b1000;
    defparam shift_srl_28_0_LC_16_16_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_28_0_LC_16_16_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83839),
            .lcout(shift_srl_28Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93079),
            .ce(N__67716),
            .sr(_gnd_net_));
    defparam shift_srl_28_1_LC_16_16_2.C_ON=1'b0;
    defparam shift_srl_28_1_LC_16_16_2.SEQ_MODE=4'b1000;
    defparam shift_srl_28_1_LC_16_16_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_28_1_LC_16_16_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64660),
            .lcout(shift_srl_28Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93079),
            .ce(N__67716),
            .sr(_gnd_net_));
    defparam shift_srl_28_11_LC_16_16_3.C_ON=1'b0;
    defparam shift_srl_28_11_LC_16_16_3.SEQ_MODE=4'b1000;
    defparam shift_srl_28_11_LC_16_16_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_28_11_LC_16_16_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64654),
            .lcout(shift_srl_28Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93079),
            .ce(N__67716),
            .sr(_gnd_net_));
    defparam shift_srl_28_3_LC_16_16_4.C_ON=1'b0;
    defparam shift_srl_28_3_LC_16_16_4.SEQ_MODE=4'b1000;
    defparam shift_srl_28_3_LC_16_16_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_28_3_LC_16_16_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64768),
            .lcout(shift_srl_28Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93079),
            .ce(N__67716),
            .sr(_gnd_net_));
    defparam shift_srl_28_15_LC_16_16_5.C_ON=1'b0;
    defparam shift_srl_28_15_LC_16_16_5.SEQ_MODE=4'b1000;
    defparam shift_srl_28_15_LC_16_16_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_28_15_LC_16_16_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64732),
            .lcout(shift_srl_28Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93079),
            .ce(N__67716),
            .sr(_gnd_net_));
    defparam shift_srl_28_9_LC_16_16_6.C_ON=1'b0;
    defparam shift_srl_28_9_LC_16_16_6.SEQ_MODE=4'b1000;
    defparam shift_srl_28_9_LC_16_16_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_28_9_LC_16_16_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64750),
            .lcout(shift_srl_28Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93079),
            .ce(N__67716),
            .sr(_gnd_net_));
    defparam shift_srl_28_2_LC_16_16_7.C_ON=1'b0;
    defparam shift_srl_28_2_LC_16_16_7.SEQ_MODE=4'b1000;
    defparam shift_srl_28_2_LC_16_16_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_28_2_LC_16_16_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64774),
            .lcout(shift_srl_28Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93079),
            .ce(N__67716),
            .sr(_gnd_net_));
    defparam shift_srl_28_4_LC_16_17_0.C_ON=1'b0;
    defparam shift_srl_28_4_LC_16_17_0.SEQ_MODE=4'b1000;
    defparam shift_srl_28_4_LC_16_17_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_28_4_LC_16_17_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64762),
            .lcout(shift_srl_28Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93053),
            .ce(N__67717),
            .sr(_gnd_net_));
    defparam shift_srl_28_12_LC_16_17_1.C_ON=1'b0;
    defparam shift_srl_28_12_LC_16_17_1.SEQ_MODE=4'b1000;
    defparam shift_srl_28_12_LC_16_17_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_28_12_LC_16_17_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64756),
            .lcout(shift_srl_28Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93053),
            .ce(N__67717),
            .sr(_gnd_net_));
    defparam shift_srl_28_8_LC_16_17_2.C_ON=1'b0;
    defparam shift_srl_28_8_LC_16_17_2.SEQ_MODE=4'b1000;
    defparam shift_srl_28_8_LC_16_17_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_28_8_LC_16_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65107),
            .lcout(shift_srl_28Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93053),
            .ce(N__67717),
            .sr(_gnd_net_));
    defparam shift_srl_28_13_LC_16_17_3.C_ON=1'b0;
    defparam shift_srl_28_13_LC_16_17_3.SEQ_MODE=4'b1000;
    defparam shift_srl_28_13_LC_16_17_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_28_13_LC_16_17_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64744),
            .lcout(shift_srl_28Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93053),
            .ce(N__67717),
            .sr(_gnd_net_));
    defparam shift_srl_28_14_LC_16_17_4.C_ON=1'b0;
    defparam shift_srl_28_14_LC_16_17_4.SEQ_MODE=4'b1000;
    defparam shift_srl_28_14_LC_16_17_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_28_14_LC_16_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64738),
            .lcout(shift_srl_28Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93053),
            .ce(N__67717),
            .sr(_gnd_net_));
    defparam shift_srl_28_5_LC_16_17_5.C_ON=1'b0;
    defparam shift_srl_28_5_LC_16_17_5.SEQ_MODE=4'b1000;
    defparam shift_srl_28_5_LC_16_17_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_28_5_LC_16_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64726),
            .lcout(shift_srl_28Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93053),
            .ce(N__67717),
            .sr(_gnd_net_));
    defparam shift_srl_28_6_LC_16_17_6.C_ON=1'b0;
    defparam shift_srl_28_6_LC_16_17_6.SEQ_MODE=4'b1000;
    defparam shift_srl_28_6_LC_16_17_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_28_6_LC_16_17_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64720),
            .lcout(shift_srl_28Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93053),
            .ce(N__67717),
            .sr(_gnd_net_));
    defparam shift_srl_28_7_LC_16_17_7.C_ON=1'b0;
    defparam shift_srl_28_7_LC_16_17_7.SEQ_MODE=4'b1000;
    defparam shift_srl_28_7_LC_16_17_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_28_7_LC_16_17_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64714),
            .lcout(shift_srl_28Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93053),
            .ce(N__67717),
            .sr(_gnd_net_));
    defparam shift_srl_117_8_LC_16_18_0.C_ON=1'b0;
    defparam shift_srl_117_8_LC_16_18_0.SEQ_MODE=4'b1000;
    defparam shift_srl_117_8_LC_16_18_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_117_8_LC_16_18_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65101),
            .lcout(shift_srl_117Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93080),
            .ce(N__65068),
            .sr(_gnd_net_));
    defparam shift_srl_117_9_LC_16_18_1.C_ON=1'b0;
    defparam shift_srl_117_9_LC_16_18_1.SEQ_MODE=4'b1000;
    defparam shift_srl_117_9_LC_16_18_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_117_9_LC_16_18_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65089),
            .lcout(shift_srl_117Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93080),
            .ce(N__65068),
            .sr(_gnd_net_));
    defparam shift_srl_107_RNI5QTS21_15_LC_16_19_0.C_ON=1'b0;
    defparam shift_srl_107_RNI5QTS21_15_LC_16_19_0.SEQ_MODE=4'b0000;
    defparam shift_srl_107_RNI5QTS21_15_LC_16_19_0.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_107_RNI5QTS21_15_LC_16_19_0 (
            .in0(N__79392),
            .in1(N__65032),
            .in2(_gnd_net_),
            .in3(N__64983),
            .lcout(rco_c_138),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_140_RNI85IA_15_LC_16_19_1.C_ON=1'b0;
    defparam shift_srl_140_RNI85IA_15_LC_16_19_1.SEQ_MODE=4'b0000;
    defparam shift_srl_140_RNI85IA_15_LC_16_19_1.LUT_INIT=16'b1100110000000000;
    LogicCell40 shift_srl_140_RNI85IA_15_LC_16_19_1 (
            .in0(_gnd_net_),
            .in1(N__64878),
            .in2(_gnd_net_),
            .in3(N__88097),
            .lcout(shift_srl_140_RNI85IAZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_139_15_LC_16_19_4.C_ON=1'b0;
    defparam shift_srl_139_15_LC_16_19_4.SEQ_MODE=4'b1000;
    defparam shift_srl_139_15_LC_16_19_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_139_15_LC_16_19_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64855),
            .lcout(shift_srl_139Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93095),
            .ce(N__64811),
            .sr(_gnd_net_));
    defparam shift_srl_139_14_LC_16_19_5.C_ON=1'b0;
    defparam shift_srl_139_14_LC_16_19_5.SEQ_MODE=4'b1000;
    defparam shift_srl_139_14_LC_16_19_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_139_14_LC_16_19_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64834),
            .lcout(shift_srl_139Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93095),
            .ce(N__64811),
            .sr(_gnd_net_));
    defparam shift_srl_139_13_LC_16_19_6.C_ON=1'b0;
    defparam shift_srl_139_13_LC_16_19_6.SEQ_MODE=4'b1000;
    defparam shift_srl_139_13_LC_16_19_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_139_13_LC_16_19_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64849),
            .lcout(shift_srl_139Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93095),
            .ce(N__64811),
            .sr(_gnd_net_));
    defparam shift_srl_162_10_LC_16_20_0.C_ON=1'b0;
    defparam shift_srl_162_10_LC_16_20_0.SEQ_MODE=4'b1000;
    defparam shift_srl_162_10_LC_16_20_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_162_10_LC_16_20_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65137),
            .lcout(shift_srl_162Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93110),
            .ce(N__69889),
            .sr(_gnd_net_));
    defparam shift_srl_162_11_LC_16_20_1.C_ON=1'b0;
    defparam shift_srl_162_11_LC_16_20_1.SEQ_MODE=4'b1000;
    defparam shift_srl_162_11_LC_16_20_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_162_11_LC_16_20_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65155),
            .lcout(shift_srl_162Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93110),
            .ce(N__69889),
            .sr(_gnd_net_));
    defparam shift_srl_162_6_LC_16_20_2.C_ON=1'b0;
    defparam shift_srl_162_6_LC_16_20_2.SEQ_MODE=4'b1000;
    defparam shift_srl_162_6_LC_16_20_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_162_6_LC_16_20_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67894),
            .lcout(shift_srl_162Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93110),
            .ce(N__69889),
            .sr(_gnd_net_));
    defparam shift_srl_162_7_LC_16_20_3.C_ON=1'b0;
    defparam shift_srl_162_7_LC_16_20_3.SEQ_MODE=4'b1000;
    defparam shift_srl_162_7_LC_16_20_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_162_7_LC_16_20_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65149),
            .lcout(shift_srl_162Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93110),
            .ce(N__69889),
            .sr(_gnd_net_));
    defparam shift_srl_162_14_LC_16_20_4.C_ON=1'b0;
    defparam shift_srl_162_14_LC_16_20_4.SEQ_MODE=4'b1000;
    defparam shift_srl_162_14_LC_16_20_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_162_14_LC_16_20_4 (
            .in0(N__67876),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_162Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93110),
            .ce(N__69889),
            .sr(_gnd_net_));
    defparam shift_srl_162_15_LC_16_20_5.C_ON=1'b0;
    defparam shift_srl_162_15_LC_16_20_5.SEQ_MODE=4'b1000;
    defparam shift_srl_162_15_LC_16_20_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_162_15_LC_16_20_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65143),
            .lcout(shift_srl_162Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93110),
            .ce(N__69889),
            .sr(_gnd_net_));
    defparam shift_srl_162_9_LC_16_20_6.C_ON=1'b0;
    defparam shift_srl_162_9_LC_16_20_6.SEQ_MODE=4'b1000;
    defparam shift_srl_162_9_LC_16_20_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_162_9_LC_16_20_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65125),
            .lcout(shift_srl_162Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93110),
            .ce(N__69889),
            .sr(_gnd_net_));
    defparam shift_srl_162_8_LC_16_20_7.C_ON=1'b0;
    defparam shift_srl_162_8_LC_16_20_7.SEQ_MODE=4'b1000;
    defparam shift_srl_162_8_LC_16_20_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_162_8_LC_16_20_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65131),
            .lcout(shift_srl_162Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93110),
            .ce(N__69889),
            .sr(_gnd_net_));
    defparam shift_srl_120_6_LC_16_21_0.C_ON=1'b0;
    defparam shift_srl_120_6_LC_16_21_0.SEQ_MODE=4'b1000;
    defparam shift_srl_120_6_LC_16_21_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_120_6_LC_16_21_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65245),
            .lcout(shift_srl_120Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93128),
            .ce(N__65190),
            .sr(_gnd_net_));
    defparam shift_srl_120_7_LC_16_21_1.C_ON=1'b0;
    defparam shift_srl_120_7_LC_16_21_1.SEQ_MODE=4'b1000;
    defparam shift_srl_120_7_LC_16_21_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_120_7_LC_16_21_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65119),
            .lcout(shift_srl_120Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93128),
            .ce(N__65190),
            .sr(_gnd_net_));
    defparam shift_srl_120_3_LC_16_21_4.C_ON=1'b0;
    defparam shift_srl_120_3_LC_16_21_4.SEQ_MODE=4'b1000;
    defparam shift_srl_120_3_LC_16_21_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_120_3_LC_16_21_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65197),
            .lcout(shift_srl_120Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93128),
            .ce(N__65190),
            .sr(_gnd_net_));
    defparam shift_srl_120_5_LC_16_21_5.C_ON=1'b0;
    defparam shift_srl_120_5_LC_16_21_5.SEQ_MODE=4'b1000;
    defparam shift_srl_120_5_LC_16_21_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_120_5_LC_16_21_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65233),
            .lcout(shift_srl_120Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93128),
            .ce(N__65190),
            .sr(_gnd_net_));
    defparam shift_srl_120_4_LC_16_21_7.C_ON=1'b0;
    defparam shift_srl_120_4_LC_16_21_7.SEQ_MODE=4'b1000;
    defparam shift_srl_120_4_LC_16_21_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_120_4_LC_16_21_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65239),
            .lcout(shift_srl_120Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93128),
            .ce(N__65190),
            .sr(_gnd_net_));
    defparam shift_srl_119_RNIVCFDU_15_LC_16_22_0.C_ON=1'b0;
    defparam shift_srl_119_RNIVCFDU_15_LC_16_22_0.SEQ_MODE=4'b0000;
    defparam shift_srl_119_RNIVCFDU_15_LC_16_22_0.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_119_RNIVCFDU_15_LC_16_22_0 (
            .in0(N__90485),
            .in1(N__65851),
            .in2(_gnd_net_),
            .in3(N__65970),
            .lcout(clk_en_120),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_119_LC_16_22_1.C_ON=1'b0;
    defparam rco_obuf_RNO_119_LC_16_22_1.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_119_LC_16_22_1.LUT_INIT=16'b1010000010100000;
    LogicCell40 rco_obuf_RNO_119_LC_16_22_1 (
            .in0(N__65971),
            .in1(_gnd_net_),
            .in2(N__65859),
            .in3(_gnd_net_),
            .lcout(rco_c_119),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_120_0_LC_16_22_2.C_ON=1'b0;
    defparam shift_srl_120_0_LC_16_22_2.SEQ_MODE=4'b1000;
    defparam shift_srl_120_0_LC_16_22_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_120_0_LC_16_22_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65602),
            .lcout(shift_srl_120Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93148),
            .ce(N__65186),
            .sr(_gnd_net_));
    defparam shift_srl_120_1_LC_16_22_3.C_ON=1'b0;
    defparam shift_srl_120_1_LC_16_22_3.SEQ_MODE=4'b1000;
    defparam shift_srl_120_1_LC_16_22_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_120_1_LC_16_22_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65209),
            .lcout(shift_srl_120Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93148),
            .ce(N__65186),
            .sr(_gnd_net_));
    defparam shift_srl_120_2_LC_16_22_4.C_ON=1'b0;
    defparam shift_srl_120_2_LC_16_22_4.SEQ_MODE=4'b1000;
    defparam shift_srl_120_2_LC_16_22_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_120_2_LC_16_22_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65203),
            .lcout(shift_srl_120Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93148),
            .ce(N__65186),
            .sr(_gnd_net_));
    defparam shift_srl_127_10_LC_16_23_0.C_ON=1'b0;
    defparam shift_srl_127_10_LC_16_23_0.SEQ_MODE=4'b1000;
    defparam shift_srl_127_10_LC_16_23_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_127_10_LC_16_23_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65767),
            .lcout(shift_srl_127Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93165),
            .ce(N__68214),
            .sr(_gnd_net_));
    defparam shift_srl_127_11_LC_16_23_1.C_ON=1'b0;
    defparam shift_srl_127_11_LC_16_23_1.SEQ_MODE=4'b1000;
    defparam shift_srl_127_11_LC_16_23_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_127_11_LC_16_23_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65161),
            .lcout(shift_srl_127Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93165),
            .ce(N__68214),
            .sr(_gnd_net_));
    defparam shift_srl_127_12_LC_16_23_2.C_ON=1'b0;
    defparam shift_srl_127_12_LC_16_23_2.SEQ_MODE=4'b1000;
    defparam shift_srl_127_12_LC_16_23_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_127_12_LC_16_23_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65791),
            .lcout(shift_srl_127Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93165),
            .ce(N__68214),
            .sr(_gnd_net_));
    defparam shift_srl_127_13_LC_16_23_3.C_ON=1'b0;
    defparam shift_srl_127_13_LC_16_23_3.SEQ_MODE=4'b1000;
    defparam shift_srl_127_13_LC_16_23_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_127_13_LC_16_23_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65785),
            .lcout(shift_srl_127Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93165),
            .ce(N__68214),
            .sr(_gnd_net_));
    defparam shift_srl_127_14_LC_16_23_4.C_ON=1'b0;
    defparam shift_srl_127_14_LC_16_23_4.SEQ_MODE=4'b1000;
    defparam shift_srl_127_14_LC_16_23_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_127_14_LC_16_23_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65779),
            .lcout(shift_srl_127Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93165),
            .ce(N__68214),
            .sr(_gnd_net_));
    defparam shift_srl_127_15_LC_16_23_5.C_ON=1'b0;
    defparam shift_srl_127_15_LC_16_23_5.SEQ_MODE=4'b1000;
    defparam shift_srl_127_15_LC_16_23_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_127_15_LC_16_23_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65773),
            .lcout(shift_srl_127Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93165),
            .ce(N__68214),
            .sr(_gnd_net_));
    defparam shift_srl_127_9_LC_16_23_6.C_ON=1'b0;
    defparam shift_srl_127_9_LC_16_23_6.SEQ_MODE=4'b1000;
    defparam shift_srl_127_9_LC_16_23_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_127_9_LC_16_23_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65761),
            .lcout(shift_srl_127Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93165),
            .ce(N__68214),
            .sr(_gnd_net_));
    defparam shift_srl_127_8_LC_16_23_7.C_ON=1'b0;
    defparam shift_srl_127_8_LC_16_23_7.SEQ_MODE=4'b1000;
    defparam shift_srl_127_8_LC_16_23_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_127_8_LC_16_23_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68221),
            .lcout(shift_srl_127Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93165),
            .ce(N__68214),
            .sr(_gnd_net_));
    defparam shift_srl_118_RNIGPI901_15_LC_16_24_0.C_ON=1'b0;
    defparam shift_srl_118_RNIGPI901_15_LC_16_24_0.SEQ_MODE=4'b0000;
    defparam shift_srl_118_RNIGPI901_15_LC_16_24_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_118_RNIGPI901_15_LC_16_24_0 (
            .in0(N__65514),
            .in1(N__65716),
            .in2(N__65380),
            .in3(N__65973),
            .lcout(rco_c_127),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_120_RNI4H9H_15_LC_16_24_2.C_ON=1'b0;
    defparam shift_srl_120_RNI4H9H_15_LC_16_24_2.SEQ_MODE=4'b0000;
    defparam shift_srl_120_RNI4H9H_15_LC_16_24_2.LUT_INIT=16'b1010101000000000;
    LogicCell40 shift_srl_120_RNI4H9H_15_LC_16_24_2 (
            .in0(N__65604),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65843),
            .lcout(rco_int_0_a2_1_a2_0_120),
            .ltout(rco_int_0_a2_1_a2_0_120_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_124_RNI19QN1_15_LC_16_24_3.C_ON=1'b0;
    defparam shift_srl_124_RNI19QN1_15_LC_16_24_3.SEQ_MODE=4'b0000;
    defparam shift_srl_124_RNI19QN1_15_LC_16_24_3.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_124_RNI19QN1_15_LC_16_24_3 (
            .in0(N__90449),
            .in1(N__65453),
            .in2(N__65383),
            .in3(N__65375),
            .lcout(),
            .ltout(clk_en_0_a3_0_a2_1_127_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_126_RNI604A01_15_LC_16_24_4.C_ON=1'b0;
    defparam shift_srl_126_RNI604A01_15_LC_16_24_4.SEQ_MODE=4'b0000;
    defparam shift_srl_126_RNI604A01_15_LC_16_24_4.LUT_INIT=16'b0000100000000000;
    LogicCell40 shift_srl_126_RNI604A01_15_LC_16_24_4 (
            .in0(N__66073),
            .in1(N__66036),
            .in2(N__65980),
            .in3(N__65972),
            .lcout(clk_en_127),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_119_15_LC_16_24_6.C_ON=1'b0;
    defparam shift_srl_119_15_LC_16_24_6.SEQ_MODE=4'b1000;
    defparam shift_srl_119_15_LC_16_24_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_119_15_LC_16_24_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65929),
            .lcout(shift_srl_119Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93186),
            .ce(N__68302),
            .sr(_gnd_net_));
    defparam shift_srl_119_14_LC_16_24_7.C_ON=1'b0;
    defparam shift_srl_119_14_LC_16_24_7.SEQ_MODE=4'b1000;
    defparam shift_srl_119_14_LC_16_24_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_119_14_LC_16_24_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66112),
            .lcout(shift_srl_119Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93186),
            .ce(N__68302),
            .sr(_gnd_net_));
    defparam shift_srl_118_RNIP44VT_15_LC_16_25_0.C_ON=1'b0;
    defparam shift_srl_118_RNIP44VT_15_LC_16_25_0.SEQ_MODE=4'b0000;
    defparam shift_srl_118_RNIP44VT_15_LC_16_25_0.LUT_INIT=16'b0100010000000000;
    LogicCell40 shift_srl_118_RNIP44VT_15_LC_16_25_0 (
            .in0(N__65923),
            .in1(N__65911),
            .in2(_gnd_net_),
            .in3(N__79531),
            .lcout(clk_en_119),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_119_0_LC_16_25_1.C_ON=1'b0;
    defparam shift_srl_119_0_LC_16_25_1.SEQ_MODE=4'b1000;
    defparam shift_srl_119_0_LC_16_25_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_119_0_LC_16_25_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65844),
            .lcout(shift_srl_119Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93206),
            .ce(N__68285),
            .sr(_gnd_net_));
    defparam shift_srl_119_1_LC_16_25_2.C_ON=1'b0;
    defparam shift_srl_119_1_LC_16_25_2.SEQ_MODE=4'b1000;
    defparam shift_srl_119_1_LC_16_25_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_119_1_LC_16_25_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65815),
            .lcout(shift_srl_119Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93206),
            .ce(N__68285),
            .sr(_gnd_net_));
    defparam shift_srl_119_2_LC_16_25_3.C_ON=1'b0;
    defparam shift_srl_119_2_LC_16_25_3.SEQ_MODE=4'b1000;
    defparam shift_srl_119_2_LC_16_25_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_119_2_LC_16_25_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65809),
            .lcout(shift_srl_119Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93206),
            .ce(N__68285),
            .sr(_gnd_net_));
    defparam shift_srl_119_3_LC_16_25_4.C_ON=1'b0;
    defparam shift_srl_119_3_LC_16_25_4.SEQ_MODE=4'b1000;
    defparam shift_srl_119_3_LC_16_25_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_119_3_LC_16_25_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65803),
            .lcout(shift_srl_119Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93206),
            .ce(N__68285),
            .sr(_gnd_net_));
    defparam shift_srl_119_4_LC_16_25_5.C_ON=1'b0;
    defparam shift_srl_119_4_LC_16_25_5.SEQ_MODE=4'b1000;
    defparam shift_srl_119_4_LC_16_25_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_119_4_LC_16_25_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65797),
            .lcout(shift_srl_119Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93206),
            .ce(N__68285),
            .sr(_gnd_net_));
    defparam shift_srl_119_10_LC_16_26_0.C_ON=1'b0;
    defparam shift_srl_119_10_LC_16_26_0.SEQ_MODE=4'b1000;
    defparam shift_srl_119_10_LC_16_26_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_119_10_LC_16_26_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66103),
            .lcout(shift_srl_119Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93225),
            .ce(N__68301),
            .sr(_gnd_net_));
    defparam shift_srl_119_11_LC_16_26_1.C_ON=1'b0;
    defparam shift_srl_119_11_LC_16_26_1.SEQ_MODE=4'b1000;
    defparam shift_srl_119_11_LC_16_26_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_119_11_LC_16_26_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66118),
            .lcout(shift_srl_119Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93225),
            .ce(N__68301),
            .sr(_gnd_net_));
    defparam shift_srl_119_13_LC_16_26_3.C_ON=1'b0;
    defparam shift_srl_119_13_LC_16_26_3.SEQ_MODE=4'b1000;
    defparam shift_srl_119_13_LC_16_26_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_119_13_LC_16_26_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68308),
            .lcout(shift_srl_119Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93225),
            .ce(N__68301),
            .sr(_gnd_net_));
    defparam shift_srl_119_9_LC_16_26_4.C_ON=1'b0;
    defparam shift_srl_119_9_LC_16_26_4.SEQ_MODE=4'b1000;
    defparam shift_srl_119_9_LC_16_26_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_119_9_LC_16_26_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66097),
            .lcout(shift_srl_119Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93225),
            .ce(N__68301),
            .sr(_gnd_net_));
    defparam shift_srl_119_8_LC_16_26_5.C_ON=1'b0;
    defparam shift_srl_119_8_LC_16_26_5.SEQ_MODE=4'b1000;
    defparam shift_srl_119_8_LC_16_26_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_119_8_LC_16_26_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68155),
            .lcout(shift_srl_119Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93225),
            .ce(N__68301),
            .sr(_gnd_net_));
    defparam shift_srl_119_5_LC_16_26_6.C_ON=1'b0;
    defparam shift_srl_119_5_LC_16_26_6.SEQ_MODE=4'b1000;
    defparam shift_srl_119_5_LC_16_26_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_119_5_LC_16_26_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66091),
            .lcout(shift_srl_119Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93225),
            .ce(N__68301),
            .sr(_gnd_net_));
    defparam shift_srl_40_9_LC_16_27_1.C_ON=1'b0;
    defparam shift_srl_40_9_LC_16_27_1.SEQ_MODE=4'b1000;
    defparam shift_srl_40_9_LC_16_27_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_40_9_LC_16_27_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66085),
            .lcout(shift_srl_40Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93245),
            .ce(N__69672),
            .sr(_gnd_net_));
    defparam shift_srl_40_8_LC_16_27_4.C_ON=1'b0;
    defparam shift_srl_40_8_LC_16_27_4.SEQ_MODE=4'b1000;
    defparam shift_srl_40_8_LC_16_27_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_40_8_LC_16_27_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66079),
            .lcout(shift_srl_40Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93245),
            .ce(N__69672),
            .sr(_gnd_net_));
    defparam shift_srl_40_7_LC_16_27_7.C_ON=1'b0;
    defparam shift_srl_40_7_LC_16_27_7.SEQ_MODE=4'b1000;
    defparam shift_srl_40_7_LC_16_27_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_40_7_LC_16_27_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68386),
            .lcout(shift_srl_40Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93245),
            .ce(N__69672),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_117_LC_16_29_2.C_ON=1'b0;
    defparam rco_obuf_RNO_117_LC_16_29_2.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_117_LC_16_29_2.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_117_LC_16_29_2 (
            .in0(N__66495),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66466),
            .lcout(rco_c_117),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_133_LC_16_30_6.C_ON=1'b0;
    defparam rco_obuf_RNO_133_LC_16_30_6.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_133_LC_16_30_6.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_133_LC_16_30_6 (
            .in0(N__66309),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66258),
            .lcout(rco_c_133),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_58_LC_16_32_6.C_ON=1'b0;
    defparam rco_obuf_RNO_58_LC_16_32_6.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_58_LC_16_32_6.LUT_INIT=16'b1000100010001000;
    LogicCell40 rco_obuf_RNO_58_LC_16_32_6 (
            .in0(N__77082),
            .in1(N__81490),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(rco_c_58),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_85_LC_17_2_1.C_ON=1'b0;
    defparam rco_obuf_RNO_85_LC_17_2_1.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_85_LC_17_2_1.LUT_INIT=16'b1000100000000000;
    LogicCell40 rco_obuf_RNO_85_LC_17_2_1 (
            .in0(N__68529),
            .in1(N__67063),
            .in2(_gnd_net_),
            .in3(N__68680),
            .lcout(rco_c_85),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_92_10_LC_17_3_0.C_ON=1'b0;
    defparam shift_srl_92_10_LC_17_3_0.SEQ_MODE=4'b1000;
    defparam shift_srl_92_10_LC_17_3_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_92_10_LC_17_3_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66661),
            .lcout(shift_srl_92Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93343),
            .ce(N__70758),
            .sr(_gnd_net_));
    defparam shift_srl_92_11_LC_17_3_1.C_ON=1'b0;
    defparam shift_srl_92_11_LC_17_3_1.SEQ_MODE=4'b1000;
    defparam shift_srl_92_11_LC_17_3_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_92_11_LC_17_3_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66142),
            .lcout(shift_srl_92Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93343),
            .ce(N__70758),
            .sr(_gnd_net_));
    defparam shift_srl_92_12_LC_17_3_2.C_ON=1'b0;
    defparam shift_srl_92_12_LC_17_3_2.SEQ_MODE=4'b1000;
    defparam shift_srl_92_12_LC_17_3_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_92_12_LC_17_3_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66136),
            .lcout(shift_srl_92Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93343),
            .ce(N__70758),
            .sr(_gnd_net_));
    defparam shift_srl_92_13_LC_17_3_3.C_ON=1'b0;
    defparam shift_srl_92_13_LC_17_3_3.SEQ_MODE=4'b1000;
    defparam shift_srl_92_13_LC_17_3_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_92_13_LC_17_3_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66130),
            .lcout(shift_srl_92Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93343),
            .ce(N__70758),
            .sr(_gnd_net_));
    defparam shift_srl_92_14_LC_17_3_4.C_ON=1'b0;
    defparam shift_srl_92_14_LC_17_3_4.SEQ_MODE=4'b1000;
    defparam shift_srl_92_14_LC_17_3_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_92_14_LC_17_3_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66124),
            .lcout(shift_srl_92Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93343),
            .ce(N__70758),
            .sr(_gnd_net_));
    defparam shift_srl_92_15_LC_17_3_5.C_ON=1'b0;
    defparam shift_srl_92_15_LC_17_3_5.SEQ_MODE=4'b1000;
    defparam shift_srl_92_15_LC_17_3_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_92_15_LC_17_3_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66667),
            .lcout(shift_srl_92Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93343),
            .ce(N__70758),
            .sr(_gnd_net_));
    defparam shift_srl_92_9_LC_17_3_6.C_ON=1'b0;
    defparam shift_srl_92_9_LC_17_3_6.SEQ_MODE=4'b1000;
    defparam shift_srl_92_9_LC_17_3_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_92_9_LC_17_3_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70771),
            .lcout(shift_srl_92Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93343),
            .ce(N__70758),
            .sr(_gnd_net_));
    defparam shift_srl_94_10_LC_17_4_0.C_ON=1'b0;
    defparam shift_srl_94_10_LC_17_4_0.SEQ_MODE=4'b1000;
    defparam shift_srl_94_10_LC_17_4_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_94_10_LC_17_4_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66649),
            .lcout(shift_srl_94Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93321),
            .ce(N__72654),
            .sr(_gnd_net_));
    defparam shift_srl_94_9_LC_17_4_1.C_ON=1'b0;
    defparam shift_srl_94_9_LC_17_4_1.SEQ_MODE=4'b1000;
    defparam shift_srl_94_9_LC_17_4_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_94_9_LC_17_4_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66655),
            .lcout(shift_srl_94Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93321),
            .ce(N__72654),
            .sr(_gnd_net_));
    defparam shift_srl_94_7_LC_17_4_3.C_ON=1'b0;
    defparam shift_srl_94_7_LC_17_4_3.SEQ_MODE=4'b1000;
    defparam shift_srl_94_7_LC_17_4_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_94_7_LC_17_4_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66637),
            .lcout(shift_srl_94Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93321),
            .ce(N__72654),
            .sr(_gnd_net_));
    defparam shift_srl_94_6_LC_17_4_4.C_ON=1'b0;
    defparam shift_srl_94_6_LC_17_4_4.SEQ_MODE=4'b1000;
    defparam shift_srl_94_6_LC_17_4_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_94_6_LC_17_4_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66631),
            .lcout(shift_srl_94Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93321),
            .ce(N__72654),
            .sr(_gnd_net_));
    defparam shift_srl_94_5_LC_17_4_5.C_ON=1'b0;
    defparam shift_srl_94_5_LC_17_4_5.SEQ_MODE=4'b1000;
    defparam shift_srl_94_5_LC_17_4_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_94_5_LC_17_4_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72664),
            .lcout(shift_srl_94Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93321),
            .ce(N__72654),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_141_LC_17_5_0.C_ON=1'b0;
    defparam rco_obuf_RNO_141_LC_17_5_0.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_141_LC_17_5_0.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_141_LC_17_5_0 (
            .in0(N__91110),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66625),
            .lcout(rco_c_141),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_144_LC_17_5_1.C_ON=1'b0;
    defparam rco_obuf_RNO_144_LC_17_5_1.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_144_LC_17_5_1.LUT_INIT=16'b1100110000000000;
    LogicCell40 rco_obuf_RNO_144_LC_17_5_1 (
            .in0(_gnd_net_),
            .in1(N__91111),
            .in2(_gnd_net_),
            .in3(N__66547),
            .lcout(rco_c_144),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_150_LC_17_5_3.C_ON=1'b0;
    defparam rco_obuf_RNO_150_LC_17_5_3.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_150_LC_17_5_3.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_150_LC_17_5_3 (
            .in0(N__82175),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66807),
            .lcout(rco_c_150),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_173_LC_17_5_4.C_ON=1'b0;
    defparam rco_obuf_RNO_173_LC_17_5_4.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_173_LC_17_5_4.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_173_LC_17_5_4 (
            .in0(N__85989),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75976),
            .lcout(rco_c_173),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_176_LC_17_5_5.C_ON=1'b0;
    defparam rco_obuf_RNO_176_LC_17_5_5.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_176_LC_17_5_5.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_176_LC_17_5_5 (
            .in0(N__80548),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85990),
            .lcout(rco_c_176),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_179_LC_17_5_6.C_ON=1'b0;
    defparam rco_obuf_RNO_179_LC_17_5_6.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_179_LC_17_5_6.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_179_LC_17_5_6 (
            .in0(N__85991),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78172),
            .lcout(rco_c_179),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_182_LC_17_5_7.C_ON=1'b0;
    defparam rco_obuf_RNO_182_LC_17_5_7.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_182_LC_17_5_7.LUT_INIT=16'b1100110000000000;
    LogicCell40 rco_obuf_RNO_182_LC_17_5_7 (
            .in0(_gnd_net_),
            .in1(N__75850),
            .in2(_gnd_net_),
            .in3(N__85992),
            .lcout(rco_c_182),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_95_10_LC_17_6_0.C_ON=1'b0;
    defparam shift_srl_95_10_LC_17_6_0.SEQ_MODE=4'b1000;
    defparam shift_srl_95_10_LC_17_6_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_95_10_LC_17_6_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66856),
            .lcout(shift_srl_95Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93285),
            .ce(N__69548),
            .sr(_gnd_net_));
    defparam shift_srl_95_11_LC_17_6_1.C_ON=1'b0;
    defparam shift_srl_95_11_LC_17_6_1.SEQ_MODE=4'b1000;
    defparam shift_srl_95_11_LC_17_6_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_95_11_LC_17_6_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66685),
            .lcout(shift_srl_95Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93285),
            .ce(N__69548),
            .sr(_gnd_net_));
    defparam shift_srl_95_12_LC_17_6_2.C_ON=1'b0;
    defparam shift_srl_95_12_LC_17_6_2.SEQ_MODE=4'b1000;
    defparam shift_srl_95_12_LC_17_6_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_95_12_LC_17_6_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66679),
            .lcout(shift_srl_95Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93285),
            .ce(N__69548),
            .sr(_gnd_net_));
    defparam shift_srl_95_13_LC_17_6_3.C_ON=1'b0;
    defparam shift_srl_95_13_LC_17_6_3.SEQ_MODE=4'b1000;
    defparam shift_srl_95_13_LC_17_6_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_95_13_LC_17_6_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66673),
            .lcout(shift_srl_95Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93285),
            .ce(N__69548),
            .sr(_gnd_net_));
    defparam shift_srl_95_9_LC_17_6_4.C_ON=1'b0;
    defparam shift_srl_95_9_LC_17_6_4.SEQ_MODE=4'b1000;
    defparam shift_srl_95_9_LC_17_6_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_95_9_LC_17_6_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66850),
            .lcout(shift_srl_95Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93285),
            .ce(N__69548),
            .sr(_gnd_net_));
    defparam shift_srl_95_8_LC_17_6_5.C_ON=1'b0;
    defparam shift_srl_95_8_LC_17_6_5.SEQ_MODE=4'b1000;
    defparam shift_srl_95_8_LC_17_6_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_95_8_LC_17_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67189),
            .lcout(shift_srl_95Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93285),
            .ce(N__69548),
            .sr(_gnd_net_));
    defparam shift_srl_95_0_LC_17_7_0.C_ON=1'b0;
    defparam shift_srl_95_0_LC_17_7_0.SEQ_MODE=4'b1000;
    defparam shift_srl_95_0_LC_17_7_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_95_0_LC_17_7_0 (
            .in0(N__69382),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_95Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93267),
            .ce(N__69552),
            .sr(_gnd_net_));
    defparam shift_srl_95_1_LC_17_7_1.C_ON=1'b0;
    defparam shift_srl_95_1_LC_17_7_1.SEQ_MODE=4'b1000;
    defparam shift_srl_95_1_LC_17_7_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_95_1_LC_17_7_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66844),
            .lcout(shift_srl_95Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93267),
            .ce(N__69552),
            .sr(_gnd_net_));
    defparam shift_srl_95_2_LC_17_7_2.C_ON=1'b0;
    defparam shift_srl_95_2_LC_17_7_2.SEQ_MODE=4'b1000;
    defparam shift_srl_95_2_LC_17_7_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_95_2_LC_17_7_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66838),
            .lcout(shift_srl_95Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93267),
            .ce(N__69552),
            .sr(_gnd_net_));
    defparam shift_srl_95_3_LC_17_7_3.C_ON=1'b0;
    defparam shift_srl_95_3_LC_17_7_3.SEQ_MODE=4'b1000;
    defparam shift_srl_95_3_LC_17_7_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_95_3_LC_17_7_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66832),
            .lcout(shift_srl_95Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93267),
            .ce(N__69552),
            .sr(_gnd_net_));
    defparam shift_srl_95_4_LC_17_7_4.C_ON=1'b0;
    defparam shift_srl_95_4_LC_17_7_4.SEQ_MODE=4'b1000;
    defparam shift_srl_95_4_LC_17_7_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_95_4_LC_17_7_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66826),
            .lcout(shift_srl_95Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93267),
            .ce(N__69552),
            .sr(_gnd_net_));
    defparam shift_srl_95_5_LC_17_7_5.C_ON=1'b0;
    defparam shift_srl_95_5_LC_17_7_5.SEQ_MODE=4'b1000;
    defparam shift_srl_95_5_LC_17_7_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_95_5_LC_17_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66820),
            .lcout(shift_srl_95Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93267),
            .ce(N__69552),
            .sr(_gnd_net_));
    defparam shift_srl_95_6_LC_17_7_6.C_ON=1'b0;
    defparam shift_srl_95_6_LC_17_7_6.SEQ_MODE=4'b1000;
    defparam shift_srl_95_6_LC_17_7_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_95_6_LC_17_7_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66814),
            .lcout(shift_srl_95Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93267),
            .ce(N__69552),
            .sr(_gnd_net_));
    defparam shift_srl_95_7_LC_17_7_7.C_ON=1'b0;
    defparam shift_srl_95_7_LC_17_7_7.SEQ_MODE=4'b1000;
    defparam shift_srl_95_7_LC_17_7_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_95_7_LC_17_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67195),
            .lcout(shift_srl_95Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93267),
            .ce(N__69552),
            .sr(_gnd_net_));
    defparam shift_srl_86_15_LC_17_8_0.C_ON=1'b0;
    defparam shift_srl_86_15_LC_17_8_0.SEQ_MODE=4'b1000;
    defparam shift_srl_86_15_LC_17_8_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_86_15_LC_17_8_0 (
            .in0(N__67183),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_86Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93248),
            .ce(N__67174),
            .sr(_gnd_net_));
    defparam shift_srl_94_RNI43JJN_15_LC_17_8_1.C_ON=1'b0;
    defparam shift_srl_94_RNI43JJN_15_LC_17_8_1.SEQ_MODE=4'b0000;
    defparam shift_srl_94_RNI43JJN_15_LC_17_8_1.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_94_RNI43JJN_15_LC_17_8_1 (
            .in0(N__72713),
            .in1(N__89944),
            .in2(_gnd_net_),
            .in3(N__72763),
            .lcout(clk_en_95),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_86_RNI23PP_15_LC_17_8_2.C_ON=1'b0;
    defparam shift_srl_86_RNI23PP_15_LC_17_8_2.SEQ_MODE=4'b0000;
    defparam shift_srl_86_RNI23PP_15_LC_17_8_2.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_86_RNI23PP_15_LC_17_8_2 (
            .in0(N__68671),
            .in1(N__67136),
            .in2(N__67117),
            .in3(N__67062),
            .lcout(),
            .ltout(rco_int_0_a2_0_a2_0_sx_89_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_89_RNIPCQF1_15_LC_17_8_3.C_ON=1'b0;
    defparam shift_srl_89_RNIPCQF1_15_LC_17_8_3.SEQ_MODE=4'b0000;
    defparam shift_srl_89_RNIPCQF1_15_LC_17_8_3.LUT_INIT=16'b0000110000000000;
    LogicCell40 shift_srl_89_RNIPCQF1_15_LC_17_8_3 (
            .in0(_gnd_net_),
            .in1(N__67018),
            .in2(N__66991),
            .in3(N__66988),
            .lcout(shift_srl_89_RNIPCQF1Z0Z_15),
            .ltout(shift_srl_89_RNIPCQF1Z0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_91_RNIOVG12_15_LC_17_8_4.C_ON=1'b0;
    defparam shift_srl_91_RNIOVG12_15_LC_17_8_4.SEQ_MODE=4'b0000;
    defparam shift_srl_91_RNIOVG12_15_LC_17_8_4.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_91_RNIOVG12_15_LC_17_8_4 (
            .in0(N__66946),
            .in1(N__66916),
            .in2(N__66865),
            .in3(N__68419),
            .lcout(shift_srl_91_RNIOVG12Z0Z_15),
            .ltout(shift_srl_91_RNIOVG12Z0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_91_RNIHF9GN_15_LC_17_8_5.C_ON=1'b0;
    defparam shift_srl_91_RNIHF9GN_15_LC_17_8_5.SEQ_MODE=4'b0000;
    defparam shift_srl_91_RNIHF9GN_15_LC_17_8_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_91_RNIHF9GN_15_LC_17_8_5 (
            .in0(N__74767),
            .in1(N__81331),
            .in2(N__66862),
            .in3(N__75078),
            .lcout(rco_c_93),
            .ltout(rco_c_93_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIEADNO_15_LC_17_8_6.C_ON=1'b0;
    defparam shift_srl_0_RNIEADNO_15_LC_17_8_6.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIEADNO_15_LC_17_8_6.LUT_INIT=16'b1000000010000000;
    LogicCell40 shift_srl_0_RNIEADNO_15_LC_17_8_6 (
            .in0(N__89943),
            .in1(N__72819),
            .in2(N__66859),
            .in3(_gnd_net_),
            .lcout(clk_en_99),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNITE8QN_15_LC_17_8_7.C_ON=1'b0;
    defparam shift_srl_0_RNITE8QN_15_LC_17_8_7.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNITE8QN_15_LC_17_8_7.LUT_INIT=16'b1100000000000000;
    LogicCell40 shift_srl_0_RNITE8QN_15_LC_17_8_7 (
            .in0(_gnd_net_),
            .in1(N__89945),
            .in2(N__72877),
            .in3(N__72764),
            .lcout(clk_en_96),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_40_LC_17_9_0.C_ON=1'b0;
    defparam rco_obuf_RNO_40_LC_17_9_0.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_40_LC_17_9_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 rco_obuf_RNO_40_LC_17_9_0 (
            .in0(N__74756),
            .in1(N__74705),
            .in2(N__85230),
            .in3(N__74498),
            .lcout(rco_c_40),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_41_RNILJSKA_15_LC_17_9_1.C_ON=1'b0;
    defparam shift_srl_41_RNILJSKA_15_LC_17_9_1.SEQ_MODE=4'b0000;
    defparam shift_srl_41_RNILJSKA_15_LC_17_9_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_41_RNILJSKA_15_LC_17_9_1 (
            .in0(N__74704),
            .in1(N__67236),
            .in2(N__90228),
            .in3(N__78798),
            .lcout(clk_en_42),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_39_RNIR6K3A_15_LC_17_9_2.C_ON=1'b0;
    defparam shift_srl_39_RNIR6K3A_15_LC_17_9_2.SEQ_MODE=4'b0000;
    defparam shift_srl_39_RNIR6K3A_15_LC_17_9_2.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_39_RNIR6K3A_15_LC_17_9_2 (
            .in0(N__74755),
            .in1(N__74497),
            .in2(_gnd_net_),
            .in3(N__85216),
            .lcout(rco_c_39),
            .ltout(rco_c_39_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNICR3HN_15_LC_17_9_3.C_ON=1'b0;
    defparam shift_srl_0_RNICR3HN_15_LC_17_9_3.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNICR3HN_15_LC_17_9_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNICR3HN_15_LC_17_9_3 (
            .in0(N__89931),
            .in1(N__68549),
            .in2(N__67270),
            .in3(N__75080),
            .lcout(clk_en_94),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIMIE4A_15_LC_17_9_4.C_ON=1'b0;
    defparam shift_srl_0_RNIMIE4A_15_LC_17_9_4.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIMIE4A_15_LC_17_9_4.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNIMIE4A_15_LC_17_9_4 (
            .in0(N__74754),
            .in1(N__74496),
            .in2(N__90212),
            .in3(N__85217),
            .lcout(clk_en_40),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_97_RNI13S31_15_LC_17_9_5.C_ON=1'b0;
    defparam shift_srl_97_RNI13S31_15_LC_17_9_5.SEQ_MODE=4'b0000;
    defparam shift_srl_97_RNI13S31_15_LC_17_9_5.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_97_RNI13S31_15_LC_17_9_5 (
            .in0(N__89930),
            .in1(N__70847),
            .in2(N__72883),
            .in3(N__69446),
            .lcout(),
            .ltout(clk_en_0_a3_0_a2_sx_98_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_97_RNIII5KO_15_LC_17_9_6.C_ON=1'b0;
    defparam shift_srl_97_RNIII5KO_15_LC_17_9_6.SEQ_MODE=4'b0000;
    defparam shift_srl_97_RNIII5KO_15_LC_17_9_6.LUT_INIT=16'b0000100000000000;
    LogicCell40 shift_srl_97_RNIII5KO_15_LC_17_9_6 (
            .in0(N__75079),
            .in1(N__67235),
            .in2(N__67219),
            .in3(N__68550),
            .lcout(clk_en_98),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_97_LC_17_9_7.C_ON=1'b0;
    defparam rco_obuf_RNO_97_LC_17_9_7.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_97_LC_17_9_7.LUT_INIT=16'b1000000000000000;
    LogicCell40 rco_obuf_RNO_97_LC_17_9_7 (
            .in0(N__72881),
            .in1(N__69447),
            .in2(N__72776),
            .in3(N__70848),
            .lcout(rco_c_97),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_45_0_LC_17_10_0.C_ON=1'b0;
    defparam shift_srl_45_0_LC_17_10_0.SEQ_MODE=4'b1000;
    defparam shift_srl_45_0_LC_17_10_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_45_0_LC_17_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76190),
            .lcout(shift_srl_45Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93208),
            .ce(N__69073),
            .sr(_gnd_net_));
    defparam shift_srl_45_1_LC_17_10_1.C_ON=1'b0;
    defparam shift_srl_45_1_LC_17_10_1.SEQ_MODE=4'b1000;
    defparam shift_srl_45_1_LC_17_10_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_45_1_LC_17_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67396),
            .lcout(shift_srl_45Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93208),
            .ce(N__69073),
            .sr(_gnd_net_));
    defparam shift_srl_45_2_LC_17_10_2.C_ON=1'b0;
    defparam shift_srl_45_2_LC_17_10_2.SEQ_MODE=4'b1000;
    defparam shift_srl_45_2_LC_17_10_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_45_2_LC_17_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67390),
            .lcout(shift_srl_45Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93208),
            .ce(N__69073),
            .sr(_gnd_net_));
    defparam shift_srl_45_3_LC_17_10_3.C_ON=1'b0;
    defparam shift_srl_45_3_LC_17_10_3.SEQ_MODE=4'b1000;
    defparam shift_srl_45_3_LC_17_10_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_45_3_LC_17_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67384),
            .lcout(shift_srl_45Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93208),
            .ce(N__69073),
            .sr(_gnd_net_));
    defparam shift_srl_45_4_LC_17_10_4.C_ON=1'b0;
    defparam shift_srl_45_4_LC_17_10_4.SEQ_MODE=4'b1000;
    defparam shift_srl_45_4_LC_17_10_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_45_4_LC_17_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67378),
            .lcout(shift_srl_45Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93208),
            .ce(N__69073),
            .sr(_gnd_net_));
    defparam shift_srl_45_5_LC_17_10_5.C_ON=1'b0;
    defparam shift_srl_45_5_LC_17_10_5.SEQ_MODE=4'b1000;
    defparam shift_srl_45_5_LC_17_10_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_45_5_LC_17_10_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67372),
            .lcout(shift_srl_45Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93208),
            .ce(N__69073),
            .sr(_gnd_net_));
    defparam shift_srl_45_6_LC_17_10_6.C_ON=1'b0;
    defparam shift_srl_45_6_LC_17_10_6.SEQ_MODE=4'b1000;
    defparam shift_srl_45_6_LC_17_10_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_45_6_LC_17_10_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67366),
            .lcout(shift_srl_45Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93208),
            .ce(N__69073),
            .sr(_gnd_net_));
    defparam shift_srl_45_7_LC_17_10_7.C_ON=1'b0;
    defparam shift_srl_45_7_LC_17_10_7.SEQ_MODE=4'b1000;
    defparam shift_srl_45_7_LC_17_10_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_45_7_LC_17_10_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67360),
            .lcout(shift_srl_45Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93208),
            .ce(N__69073),
            .sr(_gnd_net_));
    defparam shift_srl_59_RNI1I66D_15_LC_17_11_0.C_ON=1'b0;
    defparam shift_srl_59_RNI1I66D_15_LC_17_11_0.SEQ_MODE=4'b0000;
    defparam shift_srl_59_RNI1I66D_15_LC_17_11_0.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_59_RNI1I66D_15_LC_17_11_0 (
            .in0(N__81288),
            .in1(N__85003),
            .in2(N__81587),
            .in3(N__81479),
            .lcout(rco_int_0_a2_0_a2_83_m6_0_a2_sx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_59_15_LC_17_11_1.C_ON=1'b0;
    defparam shift_srl_59_15_LC_17_11_1.SEQ_MODE=4'b1000;
    defparam shift_srl_59_15_LC_17_11_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_59_15_LC_17_11_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67330),
            .lcout(shift_srl_59Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93187),
            .ce(N__73101),
            .sr(_gnd_net_));
    defparam shift_srl_59_14_LC_17_11_2.C_ON=1'b0;
    defparam shift_srl_59_14_LC_17_11_2.SEQ_MODE=4'b1000;
    defparam shift_srl_59_14_LC_17_11_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_59_14_LC_17_11_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67450),
            .lcout(shift_srl_59Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93187),
            .ce(N__73101),
            .sr(_gnd_net_));
    defparam shift_srl_59_13_LC_17_11_3.C_ON=1'b0;
    defparam shift_srl_59_13_LC_17_11_3.SEQ_MODE=4'b1000;
    defparam shift_srl_59_13_LC_17_11_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_59_13_LC_17_11_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67444),
            .lcout(shift_srl_59Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93187),
            .ce(N__73101),
            .sr(_gnd_net_));
    defparam shift_srl_59_12_LC_17_11_4.C_ON=1'b0;
    defparam shift_srl_59_12_LC_17_11_4.SEQ_MODE=4'b1000;
    defparam shift_srl_59_12_LC_17_11_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_59_12_LC_17_11_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67438),
            .lcout(shift_srl_59Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93187),
            .ce(N__73101),
            .sr(_gnd_net_));
    defparam shift_srl_59_11_LC_17_11_5.C_ON=1'b0;
    defparam shift_srl_59_11_LC_17_11_5.SEQ_MODE=4'b1000;
    defparam shift_srl_59_11_LC_17_11_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_59_11_LC_17_11_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67432),
            .lcout(shift_srl_59Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93187),
            .ce(N__73101),
            .sr(_gnd_net_));
    defparam shift_srl_59_10_LC_17_11_6.C_ON=1'b0;
    defparam shift_srl_59_10_LC_17_11_6.SEQ_MODE=4'b1000;
    defparam shift_srl_59_10_LC_17_11_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_59_10_LC_17_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67420),
            .lcout(shift_srl_59Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93187),
            .ce(N__73101),
            .sr(_gnd_net_));
    defparam shift_srl_59_9_LC_17_11_7.C_ON=1'b0;
    defparam shift_srl_59_9_LC_17_11_7.SEQ_MODE=4'b1000;
    defparam shift_srl_59_9_LC_17_11_7.LUT_INIT=16'b1100110011001100;
    LogicCell40 shift_srl_59_9_LC_17_11_7 (
            .in0(_gnd_net_),
            .in1(N__67426),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_59Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93187),
            .ce(N__73101),
            .sr(_gnd_net_));
    defparam shift_srl_98_0_LC_17_12_0.C_ON=1'b0;
    defparam shift_srl_98_0_LC_17_12_0.SEQ_MODE=4'b1000;
    defparam shift_srl_98_0_LC_17_12_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_98_0_LC_17_12_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69417),
            .lcout(shift_srl_98Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93166),
            .ce(N__67554),
            .sr(_gnd_net_));
    defparam shift_srl_98_1_LC_17_12_1.C_ON=1'b0;
    defparam shift_srl_98_1_LC_17_12_1.SEQ_MODE=4'b1000;
    defparam shift_srl_98_1_LC_17_12_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_98_1_LC_17_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67414),
            .lcout(shift_srl_98Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93166),
            .ce(N__67554),
            .sr(_gnd_net_));
    defparam shift_srl_98_2_LC_17_12_2.C_ON=1'b0;
    defparam shift_srl_98_2_LC_17_12_2.SEQ_MODE=4'b1000;
    defparam shift_srl_98_2_LC_17_12_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_98_2_LC_17_12_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67408),
            .lcout(shift_srl_98Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93166),
            .ce(N__67554),
            .sr(_gnd_net_));
    defparam shift_srl_98_3_LC_17_12_3.C_ON=1'b0;
    defparam shift_srl_98_3_LC_17_12_3.SEQ_MODE=4'b1000;
    defparam shift_srl_98_3_LC_17_12_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_98_3_LC_17_12_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67402),
            .lcout(shift_srl_98Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93166),
            .ce(N__67554),
            .sr(_gnd_net_));
    defparam shift_srl_98_4_LC_17_12_4.C_ON=1'b0;
    defparam shift_srl_98_4_LC_17_12_4.SEQ_MODE=4'b1000;
    defparam shift_srl_98_4_LC_17_12_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_98_4_LC_17_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67498),
            .lcout(shift_srl_98Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93166),
            .ce(N__67554),
            .sr(_gnd_net_));
    defparam shift_srl_98_5_LC_17_12_5.C_ON=1'b0;
    defparam shift_srl_98_5_LC_17_12_5.SEQ_MODE=4'b1000;
    defparam shift_srl_98_5_LC_17_12_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_98_5_LC_17_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67492),
            .lcout(shift_srl_98Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93166),
            .ce(N__67554),
            .sr(_gnd_net_));
    defparam shift_srl_98_6_LC_17_12_6.C_ON=1'b0;
    defparam shift_srl_98_6_LC_17_12_6.SEQ_MODE=4'b1000;
    defparam shift_srl_98_6_LC_17_12_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_98_6_LC_17_12_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67486),
            .lcout(shift_srl_98Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93166),
            .ce(N__67554),
            .sr(_gnd_net_));
    defparam shift_srl_98_7_LC_17_12_7.C_ON=1'b0;
    defparam shift_srl_98_7_LC_17_12_7.SEQ_MODE=4'b1000;
    defparam shift_srl_98_7_LC_17_12_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_98_7_LC_17_12_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67480),
            .lcout(shift_srl_98Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93166),
            .ce(N__67554),
            .sr(_gnd_net_));
    defparam shift_srl_98_10_LC_17_13_0.C_ON=1'b0;
    defparam shift_srl_98_10_LC_17_13_0.SEQ_MODE=4'b1000;
    defparam shift_srl_98_10_LC_17_13_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_98_10_LC_17_13_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67579),
            .lcout(shift_srl_98Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93149),
            .ce(N__67561),
            .sr(_gnd_net_));
    defparam shift_srl_98_11_LC_17_13_1.C_ON=1'b0;
    defparam shift_srl_98_11_LC_17_13_1.SEQ_MODE=4'b1000;
    defparam shift_srl_98_11_LC_17_13_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_98_11_LC_17_13_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67474),
            .lcout(shift_srl_98Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93149),
            .ce(N__67561),
            .sr(_gnd_net_));
    defparam shift_srl_98_12_LC_17_13_2.C_ON=1'b0;
    defparam shift_srl_98_12_LC_17_13_2.SEQ_MODE=4'b1000;
    defparam shift_srl_98_12_LC_17_13_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_98_12_LC_17_13_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67468),
            .lcout(shift_srl_98Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93149),
            .ce(N__67561),
            .sr(_gnd_net_));
    defparam shift_srl_98_13_LC_17_13_3.C_ON=1'b0;
    defparam shift_srl_98_13_LC_17_13_3.SEQ_MODE=4'b1000;
    defparam shift_srl_98_13_LC_17_13_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_98_13_LC_17_13_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67462),
            .lcout(shift_srl_98Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93149),
            .ce(N__67561),
            .sr(_gnd_net_));
    defparam shift_srl_98_14_LC_17_13_4.C_ON=1'b0;
    defparam shift_srl_98_14_LC_17_13_4.SEQ_MODE=4'b1000;
    defparam shift_srl_98_14_LC_17_13_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_98_14_LC_17_13_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67456),
            .lcout(shift_srl_98Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93149),
            .ce(N__67561),
            .sr(_gnd_net_));
    defparam shift_srl_98_15_LC_17_13_5.C_ON=1'b0;
    defparam shift_srl_98_15_LC_17_13_5.SEQ_MODE=4'b1000;
    defparam shift_srl_98_15_LC_17_13_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_98_15_LC_17_13_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67585),
            .lcout(shift_srl_98Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93149),
            .ce(N__67561),
            .sr(_gnd_net_));
    defparam shift_srl_98_9_LC_17_13_6.C_ON=1'b0;
    defparam shift_srl_98_9_LC_17_13_6.SEQ_MODE=4'b1000;
    defparam shift_srl_98_9_LC_17_13_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_98_9_LC_17_13_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67567),
            .lcout(shift_srl_98Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93149),
            .ce(N__67561),
            .sr(_gnd_net_));
    defparam shift_srl_98_8_LC_17_13_7.C_ON=1'b0;
    defparam shift_srl_98_8_LC_17_13_7.SEQ_MODE=4'b1000;
    defparam shift_srl_98_8_LC_17_13_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_98_8_LC_17_13_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67573),
            .lcout(shift_srl_98Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93149),
            .ce(N__67561),
            .sr(_gnd_net_));
    defparam shift_srl_99_RNI699Q_15_LC_17_14_0.C_ON=1'b0;
    defparam shift_srl_99_RNI699Q_15_LC_17_14_0.SEQ_MODE=4'b0000;
    defparam shift_srl_99_RNI699Q_15_LC_17_14_0.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_99_RNI699Q_15_LC_17_14_0 (
            .in0(N__67524),
            .in1(N__68418),
            .in2(_gnd_net_),
            .in3(N__81903),
            .lcout(rco_int_0_a2_0_a2_99_m6_0_a2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_99_15_LC_17_14_1.C_ON=1'b0;
    defparam shift_srl_99_15_LC_17_14_1.SEQ_MODE=4'b1000;
    defparam shift_srl_99_15_LC_17_14_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_99_15_LC_17_14_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67537),
            .lcout(shift_srl_99Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93129),
            .ce(N__67651),
            .sr(_gnd_net_));
    defparam shift_srl_99_0_LC_17_14_2.C_ON=1'b0;
    defparam shift_srl_99_0_LC_17_14_2.SEQ_MODE=4'b1000;
    defparam shift_srl_99_0_LC_17_14_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_99_0_LC_17_14_2 (
            .in0(N__67525),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_99Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93129),
            .ce(N__67651),
            .sr(_gnd_net_));
    defparam shift_srl_99_1_LC_17_14_3.C_ON=1'b0;
    defparam shift_srl_99_1_LC_17_14_3.SEQ_MODE=4'b1000;
    defparam shift_srl_99_1_LC_17_14_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_99_1_LC_17_14_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67516),
            .lcout(shift_srl_99Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93129),
            .ce(N__67651),
            .sr(_gnd_net_));
    defparam shift_srl_99_2_LC_17_14_4.C_ON=1'b0;
    defparam shift_srl_99_2_LC_17_14_4.SEQ_MODE=4'b1000;
    defparam shift_srl_99_2_LC_17_14_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_99_2_LC_17_14_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67510),
            .lcout(shift_srl_99Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93129),
            .ce(N__67651),
            .sr(_gnd_net_));
    defparam shift_srl_99_3_LC_17_14_5.C_ON=1'b0;
    defparam shift_srl_99_3_LC_17_14_5.SEQ_MODE=4'b1000;
    defparam shift_srl_99_3_LC_17_14_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_99_3_LC_17_14_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67504),
            .lcout(shift_srl_99Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93129),
            .ce(N__67651),
            .sr(_gnd_net_));
    defparam shift_srl_99_4_LC_17_14_6.C_ON=1'b0;
    defparam shift_srl_99_4_LC_17_14_6.SEQ_MODE=4'b1000;
    defparam shift_srl_99_4_LC_17_14_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_99_4_LC_17_14_6 (
            .in0(N__67675),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_99Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93129),
            .ce(N__67651),
            .sr(_gnd_net_));
    defparam shift_srl_99_5_LC_17_14_7.C_ON=1'b0;
    defparam shift_srl_99_5_LC_17_14_7.SEQ_MODE=4'b1000;
    defparam shift_srl_99_5_LC_17_14_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_99_5_LC_17_14_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67669),
            .lcout(shift_srl_99Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93129),
            .ce(N__67651),
            .sr(_gnd_net_));
    defparam shift_srl_29_9_LC_17_15_0.C_ON=1'b0;
    defparam shift_srl_29_9_LC_17_15_0.SEQ_MODE=4'b1000;
    defparam shift_srl_29_9_LC_17_15_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_29_9_LC_17_15_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67738),
            .lcout(shift_srl_29Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93111),
            .ce(N__67761),
            .sr(_gnd_net_));
    defparam shift_srl_29_2_LC_17_15_1.C_ON=1'b0;
    defparam shift_srl_29_2_LC_17_15_1.SEQ_MODE=4'b1000;
    defparam shift_srl_29_2_LC_17_15_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_29_2_LC_17_15_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67795),
            .lcout(shift_srl_29Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93111),
            .ce(N__67761),
            .sr(_gnd_net_));
    defparam shift_srl_29_3_LC_17_15_2.C_ON=1'b0;
    defparam shift_srl_29_3_LC_17_15_2.SEQ_MODE=4'b1000;
    defparam shift_srl_29_3_LC_17_15_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_29_3_LC_17_15_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67615),
            .lcout(shift_srl_29Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93111),
            .ce(N__67761),
            .sr(_gnd_net_));
    defparam shift_srl_29_7_LC_17_15_3.C_ON=1'b0;
    defparam shift_srl_29_7_LC_17_15_3.SEQ_MODE=4'b1000;
    defparam shift_srl_29_7_LC_17_15_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_29_7_LC_17_15_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67591),
            .lcout(shift_srl_29Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93111),
            .ce(N__67761),
            .sr(_gnd_net_));
    defparam shift_srl_29_4_LC_17_15_4.C_ON=1'b0;
    defparam shift_srl_29_4_LC_17_15_4.SEQ_MODE=4'b1000;
    defparam shift_srl_29_4_LC_17_15_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_29_4_LC_17_15_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67609),
            .lcout(shift_srl_29Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93111),
            .ce(N__67761),
            .sr(_gnd_net_));
    defparam shift_srl_29_5_LC_17_15_5.C_ON=1'b0;
    defparam shift_srl_29_5_LC_17_15_5.SEQ_MODE=4'b1000;
    defparam shift_srl_29_5_LC_17_15_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_29_5_LC_17_15_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67603),
            .lcout(shift_srl_29Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93111),
            .ce(N__67761),
            .sr(_gnd_net_));
    defparam shift_srl_29_6_LC_17_15_6.C_ON=1'b0;
    defparam shift_srl_29_6_LC_17_15_6.SEQ_MODE=4'b1000;
    defparam shift_srl_29_6_LC_17_15_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_29_6_LC_17_15_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67597),
            .lcout(shift_srl_29Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93111),
            .ce(N__67761),
            .sr(_gnd_net_));
    defparam shift_srl_29_8_LC_17_15_7.C_ON=1'b0;
    defparam shift_srl_29_8_LC_17_15_7.SEQ_MODE=4'b1000;
    defparam shift_srl_29_8_LC_17_15_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_29_8_LC_17_15_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67744),
            .lcout(shift_srl_29Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93111),
            .ce(N__67761),
            .sr(_gnd_net_));
    defparam shift_srl_27_RNIAA521_15_LC_17_16_0.C_ON=1'b0;
    defparam shift_srl_27_RNIAA521_15_LC_17_16_0.SEQ_MODE=4'b0000;
    defparam shift_srl_27_RNIAA521_15_LC_17_16_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_27_RNIAA521_15_LC_17_16_0 (
            .in0(N__71527),
            .in1(N__71501),
            .in2(N__71431),
            .in3(N__83794),
            .lcout(rco_int_0_a2_0_a2_out_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_27_RNIN5N67_15_LC_17_16_1.C_ON=1'b0;
    defparam shift_srl_27_RNIN5N67_15_LC_17_16_1.SEQ_MODE=4'b0000;
    defparam shift_srl_27_RNIN5N67_15_LC_17_16_1.LUT_INIT=16'b1010101000000000;
    LogicCell40 shift_srl_27_RNIN5N67_15_LC_17_16_1 (
            .in0(N__85178),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67704),
            .lcout(rco_c_27),
            .ltout(rco_c_27_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIIHH77_15_LC_17_16_2.C_ON=1'b0;
    defparam shift_srl_0_RNIIHH77_15_LC_17_16_2.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIIHH77_15_LC_17_16_2.LUT_INIT=16'b1111000000000000;
    LogicCell40 shift_srl_0_RNIIHH77_15_LC_17_16_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__67720),
            .in3(N__90430),
            .lcout(clk_en_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_28_RNICQNH7_15_LC_17_16_3.C_ON=1'b0;
    defparam shift_srl_28_RNICQNH7_15_LC_17_16_3.SEQ_MODE=4'b0000;
    defparam shift_srl_28_RNICQNH7_15_LC_17_16_3.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_28_RNICQNH7_15_LC_17_16_3 (
            .in0(N__85177),
            .in1(N__67705),
            .in2(_gnd_net_),
            .in3(N__83838),
            .lcout(rco_c_28),
            .ltout(rco_c_28_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNI76II7_15_LC_17_16_4.C_ON=1'b0;
    defparam shift_srl_0_RNI76II7_15_LC_17_16_4.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNI76II7_15_LC_17_16_4.LUT_INIT=16'b1111000000000000;
    LogicCell40 shift_srl_0_RNI76II7_15_LC_17_16_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__67684),
            .in3(N__90429),
            .lcout(clk_en_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_27_RNIP5TN_15_LC_17_16_5.C_ON=1'b0;
    defparam shift_srl_27_RNIP5TN_15_LC_17_16_5.SEQ_MODE=4'b0000;
    defparam shift_srl_27_RNIP5TN_15_LC_17_16_5.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_27_RNIP5TN_15_LC_17_16_5 (
            .in0(N__71426),
            .in1(N__71500),
            .in2(_gnd_net_),
            .in3(N__71526),
            .lcout(shift_srl_27_RNIP5TNZ0Z_15),
            .ltout(shift_srl_27_RNIP5TNZ0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_29_RNILNCS1_15_LC_17_16_6.C_ON=1'b0;
    defparam shift_srl_29_RNILNCS1_15_LC_17_16_6.SEQ_MODE=4'b0000;
    defparam shift_srl_29_RNILNCS1_15_LC_17_16_6.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_29_RNILNCS1_15_LC_17_16_6 (
            .in0(N__83888),
            .in1(N__83837),
            .in2(N__67681),
            .in3(N__83795),
            .lcout(rco_int_0_a2_0_a2_out_2),
            .ltout(rco_int_0_a2_0_a2_out_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_29_RNI2JU08_15_LC_17_16_7.C_ON=1'b0;
    defparam shift_srl_29_RNI2JU08_15_LC_17_16_7.SEQ_MODE=4'b0000;
    defparam shift_srl_29_RNI2JU08_15_LC_17_16_7.LUT_INIT=16'b1010000010100000;
    LogicCell40 shift_srl_29_RNI2JU08_15_LC_17_16_7 (
            .in0(N__85176),
            .in1(_gnd_net_),
            .in2(N__67678),
            .in3(_gnd_net_),
            .lcout(rco_c_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_29_10_LC_17_17_0.C_ON=1'b0;
    defparam shift_srl_29_10_LC_17_17_0.SEQ_MODE=4'b1000;
    defparam shift_srl_29_10_LC_17_17_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_29_10_LC_17_17_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67822),
            .lcout(shift_srl_29Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93069),
            .ce(N__67768),
            .sr(_gnd_net_));
    defparam shift_srl_29_11_LC_17_17_1.C_ON=1'b0;
    defparam shift_srl_29_11_LC_17_17_1.SEQ_MODE=4'b1000;
    defparam shift_srl_29_11_LC_17_17_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_29_11_LC_17_17_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67813),
            .lcout(shift_srl_29Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93069),
            .ce(N__67768),
            .sr(_gnd_net_));
    defparam shift_srl_29_12_LC_17_17_2.C_ON=1'b0;
    defparam shift_srl_29_12_LC_17_17_2.SEQ_MODE=4'b1000;
    defparam shift_srl_29_12_LC_17_17_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_29_12_LC_17_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67807),
            .lcout(shift_srl_29Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93069),
            .ce(N__67768),
            .sr(_gnd_net_));
    defparam shift_srl_29_13_LC_17_17_3.C_ON=1'b0;
    defparam shift_srl_29_13_LC_17_17_3.SEQ_MODE=4'b1000;
    defparam shift_srl_29_13_LC_17_17_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_29_13_LC_17_17_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67801),
            .lcout(shift_srl_29Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93069),
            .ce(N__67768),
            .sr(_gnd_net_));
    defparam shift_srl_29_1_LC_17_17_4.C_ON=1'b0;
    defparam shift_srl_29_1_LC_17_17_4.SEQ_MODE=4'b1000;
    defparam shift_srl_29_1_LC_17_17_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_29_1_LC_17_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67786),
            .lcout(shift_srl_29Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93069),
            .ce(N__67768),
            .sr(_gnd_net_));
    defparam shift_srl_29_15_LC_17_17_5.C_ON=1'b0;
    defparam shift_srl_29_15_LC_17_17_5.SEQ_MODE=4'b1000;
    defparam shift_srl_29_15_LC_17_17_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_29_15_LC_17_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67774),
            .lcout(shift_srl_29Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93069),
            .ce(N__67768),
            .sr(_gnd_net_));
    defparam shift_srl_29_0_LC_17_17_6.C_ON=1'b0;
    defparam shift_srl_29_0_LC_17_17_6.SEQ_MODE=4'b1000;
    defparam shift_srl_29_0_LC_17_17_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_29_0_LC_17_17_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83883),
            .lcout(shift_srl_29Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93069),
            .ce(N__67768),
            .sr(_gnd_net_));
    defparam shift_srl_29_14_LC_17_17_7.C_ON=1'b0;
    defparam shift_srl_29_14_LC_17_17_7.SEQ_MODE=4'b1000;
    defparam shift_srl_29_14_LC_17_17_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_29_14_LC_17_17_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67780),
            .lcout(shift_srl_29Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93069),
            .ce(N__67768),
            .sr(_gnd_net_));
    defparam shift_srl_38_7_LC_17_18_0.C_ON=1'b0;
    defparam shift_srl_38_7_LC_17_18_0.SEQ_MODE=4'b1000;
    defparam shift_srl_38_7_LC_17_18_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_38_7_LC_17_18_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69700),
            .lcout(shift_srl_38Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93096),
            .ce(N__69784),
            .sr(_gnd_net_));
    defparam shift_srl_38_14_LC_17_18_1.C_ON=1'b0;
    defparam shift_srl_38_14_LC_17_18_1.SEQ_MODE=4'b1000;
    defparam shift_srl_38_14_LC_17_18_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_38_14_LC_17_18_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67870),
            .lcout(shift_srl_38Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93096),
            .ce(N__69784),
            .sr(_gnd_net_));
    defparam shift_srl_38_13_LC_17_18_2.C_ON=1'b0;
    defparam shift_srl_38_13_LC_17_18_2.SEQ_MODE=4'b1000;
    defparam shift_srl_38_13_LC_17_18_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_38_13_LC_17_18_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69814),
            .lcout(shift_srl_38Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93096),
            .ce(N__69784),
            .sr(_gnd_net_));
    defparam shift_srl_158_0_LC_17_19_0.C_ON=1'b0;
    defparam shift_srl_158_0_LC_17_19_0.SEQ_MODE=4'b1000;
    defparam shift_srl_158_0_LC_17_19_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_158_0_LC_17_19_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77277),
            .lcout(shift_srl_158Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93112),
            .ce(N__70045),
            .sr(_gnd_net_));
    defparam shift_srl_158_1_LC_17_19_1.C_ON=1'b0;
    defparam shift_srl_158_1_LC_17_19_1.SEQ_MODE=4'b1000;
    defparam shift_srl_158_1_LC_17_19_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_158_1_LC_17_19_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67864),
            .lcout(shift_srl_158Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93112),
            .ce(N__70045),
            .sr(_gnd_net_));
    defparam shift_srl_158_2_LC_17_19_2.C_ON=1'b0;
    defparam shift_srl_158_2_LC_17_19_2.SEQ_MODE=4'b1000;
    defparam shift_srl_158_2_LC_17_19_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_158_2_LC_17_19_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67858),
            .lcout(shift_srl_158Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93112),
            .ce(N__70045),
            .sr(_gnd_net_));
    defparam shift_srl_158_3_LC_17_19_3.C_ON=1'b0;
    defparam shift_srl_158_3_LC_17_19_3.SEQ_MODE=4'b1000;
    defparam shift_srl_158_3_LC_17_19_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_158_3_LC_17_19_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67852),
            .lcout(shift_srl_158Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93112),
            .ce(N__70045),
            .sr(_gnd_net_));
    defparam shift_srl_158_4_LC_17_19_4.C_ON=1'b0;
    defparam shift_srl_158_4_LC_17_19_4.SEQ_MODE=4'b1000;
    defparam shift_srl_158_4_LC_17_19_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_158_4_LC_17_19_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67846),
            .lcout(shift_srl_158Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93112),
            .ce(N__70045),
            .sr(_gnd_net_));
    defparam shift_srl_158_5_LC_17_19_5.C_ON=1'b0;
    defparam shift_srl_158_5_LC_17_19_5.SEQ_MODE=4'b1000;
    defparam shift_srl_158_5_LC_17_19_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_158_5_LC_17_19_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67840),
            .lcout(shift_srl_158Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93112),
            .ce(N__70045),
            .sr(_gnd_net_));
    defparam shift_srl_158_6_LC_17_19_6.C_ON=1'b0;
    defparam shift_srl_158_6_LC_17_19_6.SEQ_MODE=4'b1000;
    defparam shift_srl_158_6_LC_17_19_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_158_6_LC_17_19_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67834),
            .lcout(shift_srl_158Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93112),
            .ce(N__70045),
            .sr(_gnd_net_));
    defparam shift_srl_158_7_LC_17_19_7.C_ON=1'b0;
    defparam shift_srl_158_7_LC_17_19_7.SEQ_MODE=4'b1000;
    defparam shift_srl_158_7_LC_17_19_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_158_7_LC_17_19_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67828),
            .lcout(shift_srl_158Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93112),
            .ce(N__70045),
            .sr(_gnd_net_));
    defparam shift_srl_162_0_LC_17_20_0.C_ON=1'b0;
    defparam shift_srl_162_0_LC_17_20_0.SEQ_MODE=4'b1000;
    defparam shift_srl_162_0_LC_17_20_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_162_0_LC_17_20_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77391),
            .lcout(shift_srl_162Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93130),
            .ce(N__69888),
            .sr(_gnd_net_));
    defparam shift_srl_162_1_LC_17_20_1.C_ON=1'b0;
    defparam shift_srl_162_1_LC_17_20_1.SEQ_MODE=4'b1000;
    defparam shift_srl_162_1_LC_17_20_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_162_1_LC_17_20_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67924),
            .lcout(shift_srl_162Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93130),
            .ce(N__69888),
            .sr(_gnd_net_));
    defparam shift_srl_162_2_LC_17_20_2.C_ON=1'b0;
    defparam shift_srl_162_2_LC_17_20_2.SEQ_MODE=4'b1000;
    defparam shift_srl_162_2_LC_17_20_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_162_2_LC_17_20_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67918),
            .lcout(shift_srl_162Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93130),
            .ce(N__69888),
            .sr(_gnd_net_));
    defparam shift_srl_162_3_LC_17_20_3.C_ON=1'b0;
    defparam shift_srl_162_3_LC_17_20_3.SEQ_MODE=4'b1000;
    defparam shift_srl_162_3_LC_17_20_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_162_3_LC_17_20_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67912),
            .lcout(shift_srl_162Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93130),
            .ce(N__69888),
            .sr(_gnd_net_));
    defparam shift_srl_162_4_LC_17_20_4.C_ON=1'b0;
    defparam shift_srl_162_4_LC_17_20_4.SEQ_MODE=4'b1000;
    defparam shift_srl_162_4_LC_17_20_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_162_4_LC_17_20_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67906),
            .lcout(shift_srl_162Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93130),
            .ce(N__69888),
            .sr(_gnd_net_));
    defparam shift_srl_162_5_LC_17_20_5.C_ON=1'b0;
    defparam shift_srl_162_5_LC_17_20_5.SEQ_MODE=4'b1000;
    defparam shift_srl_162_5_LC_17_20_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_162_5_LC_17_20_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67900),
            .lcout(shift_srl_162Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93130),
            .ce(N__69888),
            .sr(_gnd_net_));
    defparam shift_srl_162_12_LC_17_20_6.C_ON=1'b0;
    defparam shift_srl_162_12_LC_17_20_6.SEQ_MODE=4'b1000;
    defparam shift_srl_162_12_LC_17_20_6.LUT_INIT=16'b1100110011001100;
    LogicCell40 shift_srl_162_12_LC_17_20_6 (
            .in0(_gnd_net_),
            .in1(N__67888),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_162Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93130),
            .ce(N__69888),
            .sr(_gnd_net_));
    defparam shift_srl_162_13_LC_17_20_7.C_ON=1'b0;
    defparam shift_srl_162_13_LC_17_20_7.SEQ_MODE=4'b1000;
    defparam shift_srl_162_13_LC_17_20_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_162_13_LC_17_20_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67882),
            .lcout(shift_srl_162Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93130),
            .ce(N__69888),
            .sr(_gnd_net_));
    defparam shift_srl_156_0_LC_17_21_0.C_ON=1'b0;
    defparam shift_srl_156_0_LC_17_21_0.SEQ_MODE=4'b1000;
    defparam shift_srl_156_0_LC_17_21_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_156_0_LC_17_21_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77670),
            .lcout(shift_srl_156Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93150),
            .ce(N__70108),
            .sr(_gnd_net_));
    defparam shift_srl_156_1_LC_17_21_1.C_ON=1'b0;
    defparam shift_srl_156_1_LC_17_21_1.SEQ_MODE=4'b1000;
    defparam shift_srl_156_1_LC_17_21_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_156_1_LC_17_21_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67972),
            .lcout(shift_srl_156Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93150),
            .ce(N__70108),
            .sr(_gnd_net_));
    defparam shift_srl_156_2_LC_17_21_2.C_ON=1'b0;
    defparam shift_srl_156_2_LC_17_21_2.SEQ_MODE=4'b1000;
    defparam shift_srl_156_2_LC_17_21_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_156_2_LC_17_21_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67966),
            .lcout(shift_srl_156Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93150),
            .ce(N__70108),
            .sr(_gnd_net_));
    defparam shift_srl_156_3_LC_17_21_3.C_ON=1'b0;
    defparam shift_srl_156_3_LC_17_21_3.SEQ_MODE=4'b1000;
    defparam shift_srl_156_3_LC_17_21_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_156_3_LC_17_21_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67960),
            .lcout(shift_srl_156Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93150),
            .ce(N__70108),
            .sr(_gnd_net_));
    defparam shift_srl_156_4_LC_17_21_4.C_ON=1'b0;
    defparam shift_srl_156_4_LC_17_21_4.SEQ_MODE=4'b1000;
    defparam shift_srl_156_4_LC_17_21_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_156_4_LC_17_21_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67954),
            .lcout(shift_srl_156Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93150),
            .ce(N__70108),
            .sr(_gnd_net_));
    defparam shift_srl_156_5_LC_17_21_5.C_ON=1'b0;
    defparam shift_srl_156_5_LC_17_21_5.SEQ_MODE=4'b1000;
    defparam shift_srl_156_5_LC_17_21_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_156_5_LC_17_21_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67948),
            .lcout(shift_srl_156Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93150),
            .ce(N__70108),
            .sr(_gnd_net_));
    defparam shift_srl_156_6_LC_17_21_6.C_ON=1'b0;
    defparam shift_srl_156_6_LC_17_21_6.SEQ_MODE=4'b1000;
    defparam shift_srl_156_6_LC_17_21_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_156_6_LC_17_21_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67942),
            .lcout(shift_srl_156Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93150),
            .ce(N__70108),
            .sr(_gnd_net_));
    defparam shift_srl_156_7_LC_17_21_7.C_ON=1'b0;
    defparam shift_srl_156_7_LC_17_21_7.SEQ_MODE=4'b1000;
    defparam shift_srl_156_7_LC_17_21_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_156_7_LC_17_21_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67936),
            .lcout(shift_srl_156Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93150),
            .ce(N__70108),
            .sr(_gnd_net_));
    defparam shift_srl_187_0_LC_17_22_0.C_ON=1'b0;
    defparam shift_srl_187_0_LC_17_22_0.SEQ_MODE=4'b1000;
    defparam shift_srl_187_0_LC_17_22_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_187_0_LC_17_22_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86162),
            .lcout(shift_srl_187Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93167),
            .ce(N__70149),
            .sr(_gnd_net_));
    defparam shift_srl_187_1_LC_17_22_1.C_ON=1'b0;
    defparam shift_srl_187_1_LC_17_22_1.SEQ_MODE=4'b1000;
    defparam shift_srl_187_1_LC_17_22_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_187_1_LC_17_22_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67930),
            .lcout(shift_srl_187Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93167),
            .ce(N__70149),
            .sr(_gnd_net_));
    defparam shift_srl_187_2_LC_17_22_2.C_ON=1'b0;
    defparam shift_srl_187_2_LC_17_22_2.SEQ_MODE=4'b1000;
    defparam shift_srl_187_2_LC_17_22_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_187_2_LC_17_22_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68032),
            .lcout(shift_srl_187Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93167),
            .ce(N__70149),
            .sr(_gnd_net_));
    defparam shift_srl_187_3_LC_17_22_3.C_ON=1'b0;
    defparam shift_srl_187_3_LC_17_22_3.SEQ_MODE=4'b1000;
    defparam shift_srl_187_3_LC_17_22_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_187_3_LC_17_22_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68026),
            .lcout(shift_srl_187Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93167),
            .ce(N__70149),
            .sr(_gnd_net_));
    defparam shift_srl_187_4_LC_17_22_4.C_ON=1'b0;
    defparam shift_srl_187_4_LC_17_22_4.SEQ_MODE=4'b1000;
    defparam shift_srl_187_4_LC_17_22_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_187_4_LC_17_22_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68020),
            .lcout(shift_srl_187Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93167),
            .ce(N__70149),
            .sr(_gnd_net_));
    defparam shift_srl_187_5_LC_17_22_5.C_ON=1'b0;
    defparam shift_srl_187_5_LC_17_22_5.SEQ_MODE=4'b1000;
    defparam shift_srl_187_5_LC_17_22_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_187_5_LC_17_22_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68014),
            .lcout(shift_srl_187Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93167),
            .ce(N__70149),
            .sr(_gnd_net_));
    defparam shift_srl_187_6_LC_17_22_6.C_ON=1'b0;
    defparam shift_srl_187_6_LC_17_22_6.SEQ_MODE=4'b1000;
    defparam shift_srl_187_6_LC_17_22_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_187_6_LC_17_22_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68008),
            .lcout(shift_srl_187Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93167),
            .ce(N__70149),
            .sr(_gnd_net_));
    defparam shift_srl_187_7_LC_17_22_7.C_ON=1'b0;
    defparam shift_srl_187_7_LC_17_22_7.SEQ_MODE=4'b1000;
    defparam shift_srl_187_7_LC_17_22_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_187_7_LC_17_22_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68002),
            .lcout(shift_srl_187Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93167),
            .ce(N__70149),
            .sr(_gnd_net_));
    defparam shift_srl_111_10_LC_17_23_0.C_ON=1'b0;
    defparam shift_srl_111_10_LC_17_23_0.SEQ_MODE=4'b1000;
    defparam shift_srl_111_10_LC_17_23_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_111_10_LC_17_23_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68149),
            .lcout(shift_srl_111Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93188),
            .ce(N__68124),
            .sr(_gnd_net_));
    defparam shift_srl_111_11_LC_17_23_1.C_ON=1'b0;
    defparam shift_srl_111_11_LC_17_23_1.SEQ_MODE=4'b1000;
    defparam shift_srl_111_11_LC_17_23_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_111_11_LC_17_23_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67996),
            .lcout(shift_srl_111Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93188),
            .ce(N__68124),
            .sr(_gnd_net_));
    defparam shift_srl_111_12_LC_17_23_2.C_ON=1'b0;
    defparam shift_srl_111_12_LC_17_23_2.SEQ_MODE=4'b1000;
    defparam shift_srl_111_12_LC_17_23_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_111_12_LC_17_23_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67990),
            .lcout(shift_srl_111Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93188),
            .ce(N__68124),
            .sr(_gnd_net_));
    defparam shift_srl_111_9_LC_17_23_3.C_ON=1'b0;
    defparam shift_srl_111_9_LC_17_23_3.SEQ_MODE=4'b1000;
    defparam shift_srl_111_9_LC_17_23_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_111_9_LC_17_23_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68131),
            .lcout(shift_srl_111Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93188),
            .ce(N__68124),
            .sr(_gnd_net_));
    defparam shift_srl_111_8_LC_17_23_4.C_ON=1'b0;
    defparam shift_srl_111_8_LC_17_23_4.SEQ_MODE=4'b1000;
    defparam shift_srl_111_8_LC_17_23_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_111_8_LC_17_23_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68143),
            .lcout(shift_srl_111Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93188),
            .ce(N__68124),
            .sr(_gnd_net_));
    defparam shift_srl_127_0_LC_17_24_0.C_ON=1'b0;
    defparam shift_srl_127_0_LC_17_24_0.SEQ_MODE=4'b1000;
    defparam shift_srl_127_0_LC_17_24_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_127_0_LC_17_24_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68082),
            .lcout(shift_srl_127Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93209),
            .ce(N__68215),
            .sr(_gnd_net_));
    defparam shift_srl_127_1_LC_17_24_1.C_ON=1'b0;
    defparam shift_srl_127_1_LC_17_24_1.SEQ_MODE=4'b1000;
    defparam shift_srl_127_1_LC_17_24_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_127_1_LC_17_24_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68068),
            .lcout(shift_srl_127Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93209),
            .ce(N__68215),
            .sr(_gnd_net_));
    defparam shift_srl_127_2_LC_17_24_2.C_ON=1'b0;
    defparam shift_srl_127_2_LC_17_24_2.SEQ_MODE=4'b1000;
    defparam shift_srl_127_2_LC_17_24_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_127_2_LC_17_24_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68062),
            .lcout(shift_srl_127Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93209),
            .ce(N__68215),
            .sr(_gnd_net_));
    defparam shift_srl_127_3_LC_17_24_3.C_ON=1'b0;
    defparam shift_srl_127_3_LC_17_24_3.SEQ_MODE=4'b1000;
    defparam shift_srl_127_3_LC_17_24_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_127_3_LC_17_24_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68056),
            .lcout(shift_srl_127Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93209),
            .ce(N__68215),
            .sr(_gnd_net_));
    defparam shift_srl_127_4_LC_17_24_4.C_ON=1'b0;
    defparam shift_srl_127_4_LC_17_24_4.SEQ_MODE=4'b1000;
    defparam shift_srl_127_4_LC_17_24_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_127_4_LC_17_24_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68050),
            .lcout(shift_srl_127Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93209),
            .ce(N__68215),
            .sr(_gnd_net_));
    defparam shift_srl_127_5_LC_17_24_5.C_ON=1'b0;
    defparam shift_srl_127_5_LC_17_24_5.SEQ_MODE=4'b1000;
    defparam shift_srl_127_5_LC_17_24_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_127_5_LC_17_24_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68044),
            .lcout(shift_srl_127Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93209),
            .ce(N__68215),
            .sr(_gnd_net_));
    defparam shift_srl_127_6_LC_17_24_6.C_ON=1'b0;
    defparam shift_srl_127_6_LC_17_24_6.SEQ_MODE=4'b1000;
    defparam shift_srl_127_6_LC_17_24_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_127_6_LC_17_24_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68038),
            .lcout(shift_srl_127Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93209),
            .ce(N__68215),
            .sr(_gnd_net_));
    defparam shift_srl_127_7_LC_17_24_7.C_ON=1'b0;
    defparam shift_srl_127_7_LC_17_24_7.SEQ_MODE=4'b1000;
    defparam shift_srl_127_7_LC_17_24_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_127_7_LC_17_24_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68227),
            .lcout(shift_srl_127Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93209),
            .ce(N__68215),
            .sr(_gnd_net_));
    defparam shift_srl_173_0_LC_17_25_0.C_ON=1'b0;
    defparam shift_srl_173_0_LC_17_25_0.SEQ_MODE=4'b1000;
    defparam shift_srl_173_0_LC_17_25_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_173_0_LC_17_25_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75965),
            .lcout(shift_srl_173Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93227),
            .ce(N__80579),
            .sr(_gnd_net_));
    defparam shift_srl_173_1_LC_17_25_1.C_ON=1'b0;
    defparam shift_srl_173_1_LC_17_25_1.SEQ_MODE=4'b1000;
    defparam shift_srl_173_1_LC_17_25_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_173_1_LC_17_25_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68197),
            .lcout(shift_srl_173Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93227),
            .ce(N__80579),
            .sr(_gnd_net_));
    defparam shift_srl_173_2_LC_17_25_2.C_ON=1'b0;
    defparam shift_srl_173_2_LC_17_25_2.SEQ_MODE=4'b1000;
    defparam shift_srl_173_2_LC_17_25_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_173_2_LC_17_25_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68191),
            .lcout(shift_srl_173Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93227),
            .ce(N__80579),
            .sr(_gnd_net_));
    defparam shift_srl_173_3_LC_17_25_3.C_ON=1'b0;
    defparam shift_srl_173_3_LC_17_25_3.SEQ_MODE=4'b1000;
    defparam shift_srl_173_3_LC_17_25_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_173_3_LC_17_25_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68185),
            .lcout(shift_srl_173Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93227),
            .ce(N__80579),
            .sr(_gnd_net_));
    defparam shift_srl_173_4_LC_17_25_4.C_ON=1'b0;
    defparam shift_srl_173_4_LC_17_25_4.SEQ_MODE=4'b1000;
    defparam shift_srl_173_4_LC_17_25_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_173_4_LC_17_25_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68179),
            .lcout(shift_srl_173Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93227),
            .ce(N__80579),
            .sr(_gnd_net_));
    defparam shift_srl_173_5_LC_17_25_5.C_ON=1'b0;
    defparam shift_srl_173_5_LC_17_25_5.SEQ_MODE=4'b1000;
    defparam shift_srl_173_5_LC_17_25_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_173_5_LC_17_25_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68173),
            .lcout(shift_srl_173Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93227),
            .ce(N__80579),
            .sr(_gnd_net_));
    defparam shift_srl_173_6_LC_17_25_6.C_ON=1'b0;
    defparam shift_srl_173_6_LC_17_25_6.SEQ_MODE=4'b1000;
    defparam shift_srl_173_6_LC_17_25_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_173_6_LC_17_25_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68167),
            .lcout(shift_srl_173Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93227),
            .ce(N__80579),
            .sr(_gnd_net_));
    defparam shift_srl_173_7_LC_17_25_7.C_ON=1'b0;
    defparam shift_srl_173_7_LC_17_25_7.SEQ_MODE=4'b1000;
    defparam shift_srl_173_7_LC_17_25_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_173_7_LC_17_25_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68161),
            .lcout(shift_srl_173Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93227),
            .ce(N__80579),
            .sr(_gnd_net_));
    defparam shift_srl_119_7_LC_17_26_1.C_ON=1'b0;
    defparam shift_srl_119_7_LC_17_26_1.SEQ_MODE=4'b1000;
    defparam shift_srl_119_7_LC_17_26_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_119_7_LC_17_26_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68320),
            .lcout(shift_srl_119Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93247),
            .ce(N__68294),
            .sr(_gnd_net_));
    defparam shift_srl_119_6_LC_17_26_4.C_ON=1'b0;
    defparam shift_srl_119_6_LC_17_26_4.SEQ_MODE=4'b1000;
    defparam shift_srl_119_6_LC_17_26_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_119_6_LC_17_26_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68326),
            .lcout(shift_srl_119Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93247),
            .ce(N__68294),
            .sr(_gnd_net_));
    defparam shift_srl_119_12_LC_17_26_6.C_ON=1'b0;
    defparam shift_srl_119_12_LC_17_26_6.SEQ_MODE=4'b1000;
    defparam shift_srl_119_12_LC_17_26_6.LUT_INIT=16'b1100110011001100;
    LogicCell40 shift_srl_119_12_LC_17_26_6 (
            .in0(_gnd_net_),
            .in1(N__68314),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_119Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93247),
            .ce(N__68294),
            .sr(_gnd_net_));
    defparam shift_srl_40_0_LC_17_27_0.C_ON=1'b0;
    defparam shift_srl_40_0_LC_17_27_0.SEQ_MODE=4'b1000;
    defparam shift_srl_40_0_LC_17_27_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_40_0_LC_17_27_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74714),
            .lcout(shift_srl_40Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93266),
            .ce(N__69671),
            .sr(_gnd_net_));
    defparam shift_srl_40_1_LC_17_27_1.C_ON=1'b0;
    defparam shift_srl_40_1_LC_17_27_1.SEQ_MODE=4'b1000;
    defparam shift_srl_40_1_LC_17_27_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_40_1_LC_17_27_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68263),
            .lcout(shift_srl_40Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93266),
            .ce(N__69671),
            .sr(_gnd_net_));
    defparam shift_srl_40_2_LC_17_27_2.C_ON=1'b0;
    defparam shift_srl_40_2_LC_17_27_2.SEQ_MODE=4'b1000;
    defparam shift_srl_40_2_LC_17_27_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_40_2_LC_17_27_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68257),
            .lcout(shift_srl_40Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93266),
            .ce(N__69671),
            .sr(_gnd_net_));
    defparam shift_srl_40_3_LC_17_27_3.C_ON=1'b0;
    defparam shift_srl_40_3_LC_17_27_3.SEQ_MODE=4'b1000;
    defparam shift_srl_40_3_LC_17_27_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_40_3_LC_17_27_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68251),
            .lcout(shift_srl_40Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93266),
            .ce(N__69671),
            .sr(_gnd_net_));
    defparam shift_srl_40_4_LC_17_27_4.C_ON=1'b0;
    defparam shift_srl_40_4_LC_17_27_4.SEQ_MODE=4'b1000;
    defparam shift_srl_40_4_LC_17_27_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_40_4_LC_17_27_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68245),
            .lcout(shift_srl_40Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93266),
            .ce(N__69671),
            .sr(_gnd_net_));
    defparam shift_srl_40_5_LC_17_27_5.C_ON=1'b0;
    defparam shift_srl_40_5_LC_17_27_5.SEQ_MODE=4'b1000;
    defparam shift_srl_40_5_LC_17_27_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_40_5_LC_17_27_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68239),
            .lcout(shift_srl_40Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93266),
            .ce(N__69671),
            .sr(_gnd_net_));
    defparam shift_srl_40_6_LC_17_27_6.C_ON=1'b0;
    defparam shift_srl_40_6_LC_17_27_6.SEQ_MODE=4'b1000;
    defparam shift_srl_40_6_LC_17_27_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_40_6_LC_17_27_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68233),
            .lcout(shift_srl_40Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93266),
            .ce(N__69671),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_54_LC_17_29_3.C_ON=1'b0;
    defparam rco_obuf_RNO_54_LC_17_29_3.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_54_LC_17_29_3.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_54_LC_17_29_3 (
            .in0(N__77069),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77023),
            .lcout(rco_c_54),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_198_6_LC_17_30_0.C_ON=1'b0;
    defparam shift_srl_198_6_LC_17_30_0.SEQ_MODE=4'b1000;
    defparam shift_srl_198_6_LC_17_30_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_198_6_LC_17_30_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70369),
            .lcout(shift_srl_198Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93320),
            .ce(N__72205),
            .sr(_gnd_net_));
    defparam shift_srl_198_7_LC_17_30_1.C_ON=1'b0;
    defparam shift_srl_198_7_LC_17_30_1.SEQ_MODE=4'b1000;
    defparam shift_srl_198_7_LC_17_30_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_198_7_LC_17_30_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68362),
            .lcout(shift_srl_198Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93320),
            .ce(N__72205),
            .sr(_gnd_net_));
    defparam shift_srl_93_0_LC_18_2_0.C_ON=1'b0;
    defparam shift_srl_93_0_LC_18_2_0.SEQ_MODE=4'b1000;
    defparam shift_srl_93_0_LC_18_2_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_93_0_LC_18_2_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69519),
            .lcout(shift_srl_93Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93380),
            .ce(N__70571),
            .sr(_gnd_net_));
    defparam shift_srl_93_1_LC_18_2_1.C_ON=1'b0;
    defparam shift_srl_93_1_LC_18_2_1.SEQ_MODE=4'b1000;
    defparam shift_srl_93_1_LC_18_2_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_93_1_LC_18_2_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68356),
            .lcout(shift_srl_93Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93380),
            .ce(N__70571),
            .sr(_gnd_net_));
    defparam shift_srl_93_2_LC_18_2_2.C_ON=1'b0;
    defparam shift_srl_93_2_LC_18_2_2.SEQ_MODE=4'b1000;
    defparam shift_srl_93_2_LC_18_2_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_93_2_LC_18_2_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68350),
            .lcout(shift_srl_93Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93380),
            .ce(N__70571),
            .sr(_gnd_net_));
    defparam shift_srl_93_3_LC_18_2_3.C_ON=1'b0;
    defparam shift_srl_93_3_LC_18_2_3.SEQ_MODE=4'b1000;
    defparam shift_srl_93_3_LC_18_2_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_93_3_LC_18_2_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68344),
            .lcout(shift_srl_93Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93380),
            .ce(N__70571),
            .sr(_gnd_net_));
    defparam shift_srl_93_4_LC_18_2_4.C_ON=1'b0;
    defparam shift_srl_93_4_LC_18_2_4.SEQ_MODE=4'b1000;
    defparam shift_srl_93_4_LC_18_2_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_93_4_LC_18_2_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68338),
            .lcout(shift_srl_93Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93380),
            .ce(N__70571),
            .sr(_gnd_net_));
    defparam shift_srl_93_5_LC_18_2_5.C_ON=1'b0;
    defparam shift_srl_93_5_LC_18_2_5.SEQ_MODE=4'b1000;
    defparam shift_srl_93_5_LC_18_2_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_93_5_LC_18_2_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68332),
            .lcout(shift_srl_93Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93380),
            .ce(N__70571),
            .sr(_gnd_net_));
    defparam shift_srl_93_6_LC_18_2_6.C_ON=1'b0;
    defparam shift_srl_93_6_LC_18_2_6.SEQ_MODE=4'b1000;
    defparam shift_srl_93_6_LC_18_2_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_93_6_LC_18_2_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68692),
            .lcout(shift_srl_93Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93380),
            .ce(N__70571),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_84_LC_18_3_1.C_ON=1'b0;
    defparam rco_obuf_RNO_84_LC_18_3_1.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_84_LC_18_3_1.LUT_INIT=16'b1100110000000000;
    LogicCell40 rco_obuf_RNO_84_LC_18_3_1 (
            .in0(_gnd_net_),
            .in1(N__68686),
            .in2(_gnd_net_),
            .in3(N__68517),
            .lcout(rco_c_84),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_89_LC_18_3_2.C_ON=1'b0;
    defparam rco_obuf_RNO_89_LC_18_3_2.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_89_LC_18_3_2.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_89_LC_18_3_2 (
            .in0(N__68518),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68610),
            .lcout(rco_c_89),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIIR15N_15_LC_18_3_4.C_ON=1'b0;
    defparam shift_srl_0_RNIIR15N_15_LC_18_3_4.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIIR15N_15_LC_18_3_4.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_0_RNIIR15N_15_LC_18_3_4 (
            .in0(N__68515),
            .in1(N__90230),
            .in2(_gnd_net_),
            .in3(N__72110),
            .lcout(clk_en_92),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNI8R4FN_15_LC_18_3_5.C_ON=1'b0;
    defparam shift_srl_0_RNI8R4FN_15_LC_18_3_5.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNI8R4FN_15_LC_18_3_5.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_0_RNI8R4FN_15_LC_18_3_5 (
            .in0(N__90229),
            .in1(N__68559),
            .in2(_gnd_net_),
            .in3(N__68516),
            .lcout(clk_en_93),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_92_LC_18_3_6.C_ON=1'b0;
    defparam rco_obuf_RNO_92_LC_18_3_6.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_92_LC_18_3_6.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_92_LC_18_3_6 (
            .in0(N__68560),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68521),
            .lcout(rco_c_92),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_92_0_LC_18_3_7.C_ON=1'b0;
    defparam shift_srl_92_0_LC_18_3_7.SEQ_MODE=4'b1000;
    defparam shift_srl_92_0_LC_18_3_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_92_0_LC_18_3_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68411),
            .lcout(shift_srl_92Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93363),
            .ce(N__70757),
            .sr(_gnd_net_));
    defparam shift_srl_93_10_LC_18_4_0.C_ON=1'b0;
    defparam shift_srl_93_10_LC_18_4_0.SEQ_MODE=4'b1000;
    defparam shift_srl_93_10_LC_18_4_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_93_10_LC_18_4_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68704),
            .lcout(shift_srl_93Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93345),
            .ce(N__70576),
            .sr(_gnd_net_));
    defparam shift_srl_93_11_LC_18_4_1.C_ON=1'b0;
    defparam shift_srl_93_11_LC_18_4_1.SEQ_MODE=4'b1000;
    defparam shift_srl_93_11_LC_18_4_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_93_11_LC_18_4_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68392),
            .lcout(shift_srl_93Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93345),
            .ce(N__70576),
            .sr(_gnd_net_));
    defparam shift_srl_93_12_LC_18_4_2.C_ON=1'b0;
    defparam shift_srl_93_12_LC_18_4_2.SEQ_MODE=4'b1000;
    defparam shift_srl_93_12_LC_18_4_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_93_12_LC_18_4_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68728),
            .lcout(shift_srl_93Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93345),
            .ce(N__70576),
            .sr(_gnd_net_));
    defparam shift_srl_93_13_LC_18_4_3.C_ON=1'b0;
    defparam shift_srl_93_13_LC_18_4_3.SEQ_MODE=4'b1000;
    defparam shift_srl_93_13_LC_18_4_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_93_13_LC_18_4_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68722),
            .lcout(shift_srl_93Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93345),
            .ce(N__70576),
            .sr(_gnd_net_));
    defparam shift_srl_93_14_LC_18_4_4.C_ON=1'b0;
    defparam shift_srl_93_14_LC_18_4_4.SEQ_MODE=4'b1000;
    defparam shift_srl_93_14_LC_18_4_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_93_14_LC_18_4_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68716),
            .lcout(shift_srl_93Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93345),
            .ce(N__70576),
            .sr(_gnd_net_));
    defparam shift_srl_93_15_LC_18_4_5.C_ON=1'b0;
    defparam shift_srl_93_15_LC_18_4_5.SEQ_MODE=4'b1000;
    defparam shift_srl_93_15_LC_18_4_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_93_15_LC_18_4_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68710),
            .lcout(shift_srl_93Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93345),
            .ce(N__70576),
            .sr(_gnd_net_));
    defparam shift_srl_93_9_LC_18_4_6.C_ON=1'b0;
    defparam shift_srl_93_9_LC_18_4_6.SEQ_MODE=4'b1000;
    defparam shift_srl_93_9_LC_18_4_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_93_9_LC_18_4_6 (
            .in0(N__70597),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_93Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93345),
            .ce(N__70576),
            .sr(_gnd_net_));
    defparam shift_srl_46_0_LC_18_5_0.C_ON=1'b0;
    defparam shift_srl_46_0_LC_18_5_0.SEQ_MODE=4'b1000;
    defparam shift_srl_46_0_LC_18_5_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_46_0_LC_18_5_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74369),
            .lcout(shift_srl_46Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93323),
            .ce(N__70872),
            .sr(_gnd_net_));
    defparam shift_srl_46_1_LC_18_5_1.C_ON=1'b0;
    defparam shift_srl_46_1_LC_18_5_1.SEQ_MODE=4'b1000;
    defparam shift_srl_46_1_LC_18_5_1.LUT_INIT=16'b1100110011001100;
    LogicCell40 shift_srl_46_1_LC_18_5_1 (
            .in0(_gnd_net_),
            .in1(N__68698),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_46Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93323),
            .ce(N__70872),
            .sr(_gnd_net_));
    defparam shift_srl_46_10_LC_18_5_2.C_ON=1'b0;
    defparam shift_srl_46_10_LC_18_5_2.SEQ_MODE=4'b1000;
    defparam shift_srl_46_10_LC_18_5_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_46_10_LC_18_5_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68770),
            .lcout(shift_srl_46Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93323),
            .ce(N__70872),
            .sr(_gnd_net_));
    defparam shift_srl_46_3_LC_18_5_3.C_ON=1'b0;
    defparam shift_srl_46_3_LC_18_5_3.SEQ_MODE=4'b1000;
    defparam shift_srl_46_3_LC_18_5_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_46_3_LC_18_5_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68758),
            .lcout(shift_srl_46Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93323),
            .ce(N__70872),
            .sr(_gnd_net_));
    defparam shift_srl_46_4_LC_18_5_4.C_ON=1'b0;
    defparam shift_srl_46_4_LC_18_5_4.SEQ_MODE=4'b1000;
    defparam shift_srl_46_4_LC_18_5_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_46_4_LC_18_5_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68782),
            .lcout(shift_srl_46Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93323),
            .ce(N__70872),
            .sr(_gnd_net_));
    defparam shift_srl_46_8_LC_18_5_5.C_ON=1'b0;
    defparam shift_srl_46_8_LC_18_5_5.SEQ_MODE=4'b1000;
    defparam shift_srl_46_8_LC_18_5_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_46_8_LC_18_5_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70927),
            .lcout(shift_srl_46Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93323),
            .ce(N__70872),
            .sr(_gnd_net_));
    defparam shift_srl_46_9_LC_18_5_6.C_ON=1'b0;
    defparam shift_srl_46_9_LC_18_5_6.SEQ_MODE=4'b1000;
    defparam shift_srl_46_9_LC_18_5_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_46_9_LC_18_5_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68776),
            .lcout(shift_srl_46Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93323),
            .ce(N__70872),
            .sr(_gnd_net_));
    defparam shift_srl_46_2_LC_18_5_7.C_ON=1'b0;
    defparam shift_srl_46_2_LC_18_5_7.SEQ_MODE=4'b1000;
    defparam shift_srl_46_2_LC_18_5_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_46_2_LC_18_5_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68764),
            .lcout(shift_srl_46Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93323),
            .ce(N__70872),
            .sr(_gnd_net_));
    defparam shift_srl_97_10_LC_18_6_0.C_ON=1'b0;
    defparam shift_srl_97_10_LC_18_6_0.SEQ_MODE=4'b1000;
    defparam shift_srl_97_10_LC_18_6_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_97_10_LC_18_6_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68830),
            .lcout(shift_srl_97Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93302),
            .ce(N__70944),
            .sr(_gnd_net_));
    defparam shift_srl_97_11_LC_18_6_1.C_ON=1'b0;
    defparam shift_srl_97_11_LC_18_6_1.SEQ_MODE=4'b1000;
    defparam shift_srl_97_11_LC_18_6_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_97_11_LC_18_6_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68752),
            .lcout(shift_srl_97Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93302),
            .ce(N__70944),
            .sr(_gnd_net_));
    defparam shift_srl_97_12_LC_18_6_2.C_ON=1'b0;
    defparam shift_srl_97_12_LC_18_6_2.SEQ_MODE=4'b1000;
    defparam shift_srl_97_12_LC_18_6_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_97_12_LC_18_6_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68746),
            .lcout(shift_srl_97Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93302),
            .ce(N__70944),
            .sr(_gnd_net_));
    defparam shift_srl_97_13_LC_18_6_3.C_ON=1'b0;
    defparam shift_srl_97_13_LC_18_6_3.SEQ_MODE=4'b1000;
    defparam shift_srl_97_13_LC_18_6_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_97_13_LC_18_6_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68740),
            .lcout(shift_srl_97Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93302),
            .ce(N__70944),
            .sr(_gnd_net_));
    defparam shift_srl_97_14_LC_18_6_4.C_ON=1'b0;
    defparam shift_srl_97_14_LC_18_6_4.SEQ_MODE=4'b1000;
    defparam shift_srl_97_14_LC_18_6_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_97_14_LC_18_6_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68734),
            .lcout(shift_srl_97Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93302),
            .ce(N__70944),
            .sr(_gnd_net_));
    defparam shift_srl_97_15_LC_18_6_5.C_ON=1'b0;
    defparam shift_srl_97_15_LC_18_6_5.SEQ_MODE=4'b1000;
    defparam shift_srl_97_15_LC_18_6_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_97_15_LC_18_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68836),
            .lcout(shift_srl_97Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93302),
            .ce(N__70944),
            .sr(_gnd_net_));
    defparam shift_srl_97_9_LC_18_6_6.C_ON=1'b0;
    defparam shift_srl_97_9_LC_18_6_6.SEQ_MODE=4'b1000;
    defparam shift_srl_97_9_LC_18_6_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_97_9_LC_18_6_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68824),
            .lcout(shift_srl_97Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93302),
            .ce(N__70944),
            .sr(_gnd_net_));
    defparam shift_srl_97_8_LC_18_6_7.C_ON=1'b0;
    defparam shift_srl_97_8_LC_18_6_7.SEQ_MODE=4'b1000;
    defparam shift_srl_97_8_LC_18_6_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_97_8_LC_18_6_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70951),
            .lcout(shift_srl_97Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93302),
            .ce(N__70944),
            .sr(_gnd_net_));
    defparam shift_srl_94_15_LC_18_7_0.C_ON=1'b0;
    defparam shift_srl_94_15_LC_18_7_0.SEQ_MODE=4'b1000;
    defparam shift_srl_94_15_LC_18_7_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_94_15_LC_18_7_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68800),
            .lcout(shift_srl_94Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93287),
            .ce(N__72646),
            .sr(_gnd_net_));
    defparam shift_srl_95_RNIHJ49_15_LC_18_7_1.C_ON=1'b0;
    defparam shift_srl_95_RNIHJ49_15_LC_18_7_1.SEQ_MODE=4'b0000;
    defparam shift_srl_95_RNIHJ49_15_LC_18_7_1.LUT_INIT=16'b1100110000000000;
    LogicCell40 shift_srl_95_RNIHJ49_15_LC_18_7_1 (
            .in0(_gnd_net_),
            .in1(N__72712),
            .in2(_gnd_net_),
            .in3(N__69381),
            .lcout(shift_srl_95_RNIHJ49Z0Z_15),
            .ltout(shift_srl_95_RNIHJ49Z0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_96_RNINU35O_15_LC_18_7_2.C_ON=1'b0;
    defparam shift_srl_96_RNINU35O_15_LC_18_7_2.SEQ_MODE=4'b0000;
    defparam shift_srl_96_RNINU35O_15_LC_18_7_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_96_RNINU35O_15_LC_18_7_2 (
            .in0(N__89916),
            .in1(N__72765),
            .in2(N__68818),
            .in3(N__69450),
            .lcout(clk_en_97),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_96_LC_18_7_3.C_ON=1'b0;
    defparam rco_obuf_RNO_96_LC_18_7_3.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_96_LC_18_7_3.LUT_INIT=16'b1010000000000000;
    LogicCell40 rco_obuf_RNO_96_LC_18_7_3 (
            .in0(N__72766),
            .in1(_gnd_net_),
            .in2(N__69454),
            .in3(N__72873),
            .lcout(rco_c_96),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_94_14_LC_18_7_4.C_ON=1'b0;
    defparam shift_srl_94_14_LC_18_7_4.SEQ_MODE=4'b1000;
    defparam shift_srl_94_14_LC_18_7_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_94_14_LC_18_7_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68794),
            .lcout(shift_srl_94Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93287),
            .ce(N__72646),
            .sr(_gnd_net_));
    defparam shift_srl_94_13_LC_18_7_5.C_ON=1'b0;
    defparam shift_srl_94_13_LC_18_7_5.SEQ_MODE=4'b1000;
    defparam shift_srl_94_13_LC_18_7_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_94_13_LC_18_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68788),
            .lcout(shift_srl_94Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93287),
            .ce(N__72646),
            .sr(_gnd_net_));
    defparam shift_srl_94_12_LC_18_7_6.C_ON=1'b0;
    defparam shift_srl_94_12_LC_18_7_6.SEQ_MODE=4'b1000;
    defparam shift_srl_94_12_LC_18_7_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_94_12_LC_18_7_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68878),
            .lcout(shift_srl_94Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93287),
            .ce(N__72646),
            .sr(_gnd_net_));
    defparam shift_srl_94_11_LC_18_7_7.C_ON=1'b0;
    defparam shift_srl_94_11_LC_18_7_7.SEQ_MODE=4'b1000;
    defparam shift_srl_94_11_LC_18_7_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_94_11_LC_18_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68890),
            .lcout(shift_srl_94Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93287),
            .ce(N__72646),
            .sr(_gnd_net_));
    defparam shift_srl_96_12_LC_18_8_0.C_ON=1'b0;
    defparam shift_srl_96_12_LC_18_8_0.SEQ_MODE=4'b1000;
    defparam shift_srl_96_12_LC_18_8_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_96_12_LC_18_8_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68842),
            .lcout(shift_srl_96Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93269),
            .ce(N__68907),
            .sr(_gnd_net_));
    defparam shift_srl_96_1_LC_18_8_1.C_ON=1'b0;
    defparam shift_srl_96_1_LC_18_8_1.SEQ_MODE=4'b1000;
    defparam shift_srl_96_1_LC_18_8_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_96_1_LC_18_8_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68854),
            .lcout(shift_srl_96Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93269),
            .ce(N__68907),
            .sr(_gnd_net_));
    defparam shift_srl_96_2_LC_18_8_2.C_ON=1'b0;
    defparam shift_srl_96_2_LC_18_8_2.SEQ_MODE=4'b1000;
    defparam shift_srl_96_2_LC_18_8_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_96_2_LC_18_8_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68872),
            .lcout(shift_srl_96Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93269),
            .ce(N__68907),
            .sr(_gnd_net_));
    defparam shift_srl_96_3_LC_18_8_3.C_ON=1'b0;
    defparam shift_srl_96_3_LC_18_8_3.SEQ_MODE=4'b1000;
    defparam shift_srl_96_3_LC_18_8_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_96_3_LC_18_8_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68866),
            .lcout(shift_srl_96Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93269),
            .ce(N__68907),
            .sr(_gnd_net_));
    defparam shift_srl_96_4_LC_18_8_4.C_ON=1'b0;
    defparam shift_srl_96_4_LC_18_8_4.SEQ_MODE=4'b1000;
    defparam shift_srl_96_4_LC_18_8_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_96_4_LC_18_8_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68860),
            .lcout(shift_srl_96Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93269),
            .ce(N__68907),
            .sr(_gnd_net_));
    defparam shift_srl_96_0_LC_18_8_5.C_ON=1'b0;
    defparam shift_srl_96_0_LC_18_8_5.SEQ_MODE=4'b1000;
    defparam shift_srl_96_0_LC_18_8_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_96_0_LC_18_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69448),
            .lcout(shift_srl_96Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93269),
            .ce(N__68907),
            .sr(_gnd_net_));
    defparam shift_srl_96_10_LC_18_8_6.C_ON=1'b0;
    defparam shift_srl_96_10_LC_18_8_6.SEQ_MODE=4'b1000;
    defparam shift_srl_96_10_LC_18_8_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_96_10_LC_18_8_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68926),
            .lcout(shift_srl_96Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93269),
            .ce(N__68907),
            .sr(_gnd_net_));
    defparam shift_srl_96_11_LC_18_8_7.C_ON=1'b0;
    defparam shift_srl_96_11_LC_18_8_7.SEQ_MODE=4'b1000;
    defparam shift_srl_96_11_LC_18_8_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_96_11_LC_18_8_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68848),
            .lcout(shift_srl_96Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93269),
            .ce(N__68907),
            .sr(_gnd_net_));
    defparam shift_srl_96_6_LC_18_9_0.C_ON=1'b0;
    defparam shift_srl_96_6_LC_18_9_0.SEQ_MODE=4'b1000;
    defparam shift_srl_96_6_LC_18_9_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_96_6_LC_18_9_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68950),
            .lcout(shift_srl_96Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93250),
            .ce(N__68908),
            .sr(_gnd_net_));
    defparam shift_srl_96_7_LC_18_9_1.C_ON=1'b0;
    defparam shift_srl_96_7_LC_18_9_1.SEQ_MODE=4'b1000;
    defparam shift_srl_96_7_LC_18_9_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_96_7_LC_18_9_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68962),
            .lcout(shift_srl_96Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93250),
            .ce(N__68908),
            .sr(_gnd_net_));
    defparam shift_srl_96_5_LC_18_9_2.C_ON=1'b0;
    defparam shift_srl_96_5_LC_18_9_2.SEQ_MODE=4'b1000;
    defparam shift_srl_96_5_LC_18_9_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_96_5_LC_18_9_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68956),
            .lcout(shift_srl_96Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93250),
            .ce(N__68908),
            .sr(_gnd_net_));
    defparam shift_srl_96_13_LC_18_9_3.C_ON=1'b0;
    defparam shift_srl_96_13_LC_18_9_3.SEQ_MODE=4'b1000;
    defparam shift_srl_96_13_LC_18_9_3.LUT_INIT=16'b1100110011001100;
    LogicCell40 shift_srl_96_13_LC_18_9_3 (
            .in0(_gnd_net_),
            .in1(N__68944),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_96Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93250),
            .ce(N__68908),
            .sr(_gnd_net_));
    defparam shift_srl_96_14_LC_18_9_4.C_ON=1'b0;
    defparam shift_srl_96_14_LC_18_9_4.SEQ_MODE=4'b1000;
    defparam shift_srl_96_14_LC_18_9_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_96_14_LC_18_9_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68938),
            .lcout(shift_srl_96Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93250),
            .ce(N__68908),
            .sr(_gnd_net_));
    defparam shift_srl_96_15_LC_18_9_5.C_ON=1'b0;
    defparam shift_srl_96_15_LC_18_9_5.SEQ_MODE=4'b1000;
    defparam shift_srl_96_15_LC_18_9_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_96_15_LC_18_9_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68932),
            .lcout(shift_srl_96Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93250),
            .ce(N__68908),
            .sr(_gnd_net_));
    defparam shift_srl_96_9_LC_18_9_6.C_ON=1'b0;
    defparam shift_srl_96_9_LC_18_9_6.SEQ_MODE=4'b1000;
    defparam shift_srl_96_9_LC_18_9_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_96_9_LC_18_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68914),
            .lcout(shift_srl_96Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93250),
            .ce(N__68908),
            .sr(_gnd_net_));
    defparam shift_srl_96_8_LC_18_9_7.C_ON=1'b0;
    defparam shift_srl_96_8_LC_18_9_7.SEQ_MODE=4'b1000;
    defparam shift_srl_96_8_LC_18_9_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_96_8_LC_18_9_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68920),
            .lcout(shift_srl_96Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93250),
            .ce(N__68908),
            .sr(_gnd_net_));
    defparam shift_srl_45_10_LC_18_10_0.C_ON=1'b0;
    defparam shift_srl_45_10_LC_18_10_0.SEQ_MODE=4'b1000;
    defparam shift_srl_45_10_LC_18_10_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_45_10_LC_18_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69016),
            .lcout(shift_srl_45Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93228),
            .ce(N__69072),
            .sr(_gnd_net_));
    defparam shift_srl_45_11_LC_18_10_1.C_ON=1'b0;
    defparam shift_srl_45_11_LC_18_10_1.SEQ_MODE=4'b1000;
    defparam shift_srl_45_11_LC_18_10_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_45_11_LC_18_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69046),
            .lcout(shift_srl_45Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93228),
            .ce(N__69072),
            .sr(_gnd_net_));
    defparam shift_srl_45_12_LC_18_10_2.C_ON=1'b0;
    defparam shift_srl_45_12_LC_18_10_2.SEQ_MODE=4'b1000;
    defparam shift_srl_45_12_LC_18_10_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_45_12_LC_18_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69040),
            .lcout(shift_srl_45Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93228),
            .ce(N__69072),
            .sr(_gnd_net_));
    defparam shift_srl_45_13_LC_18_10_3.C_ON=1'b0;
    defparam shift_srl_45_13_LC_18_10_3.SEQ_MODE=4'b1000;
    defparam shift_srl_45_13_LC_18_10_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_45_13_LC_18_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69034),
            .lcout(shift_srl_45Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93228),
            .ce(N__69072),
            .sr(_gnd_net_));
    defparam shift_srl_45_14_LC_18_10_4.C_ON=1'b0;
    defparam shift_srl_45_14_LC_18_10_4.SEQ_MODE=4'b1000;
    defparam shift_srl_45_14_LC_18_10_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_45_14_LC_18_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69028),
            .lcout(shift_srl_45Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93228),
            .ce(N__69072),
            .sr(_gnd_net_));
    defparam shift_srl_45_15_LC_18_10_5.C_ON=1'b0;
    defparam shift_srl_45_15_LC_18_10_5.SEQ_MODE=4'b1000;
    defparam shift_srl_45_15_LC_18_10_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_45_15_LC_18_10_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69022),
            .lcout(shift_srl_45Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93228),
            .ce(N__69072),
            .sr(_gnd_net_));
    defparam shift_srl_45_9_LC_18_10_6.C_ON=1'b0;
    defparam shift_srl_45_9_LC_18_10_6.SEQ_MODE=4'b1000;
    defparam shift_srl_45_9_LC_18_10_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_45_9_LC_18_10_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69004),
            .lcout(shift_srl_45Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93228),
            .ce(N__69072),
            .sr(_gnd_net_));
    defparam shift_srl_45_8_LC_18_10_7.C_ON=1'b0;
    defparam shift_srl_45_8_LC_18_10_7.SEQ_MODE=4'b1000;
    defparam shift_srl_45_8_LC_18_10_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_45_8_LC_18_10_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69010),
            .lcout(shift_srl_45Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93228),
            .ce(N__69072),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIANPAC_15_LC_18_11_0.C_ON=1'b0;
    defparam shift_srl_0_RNIANPAC_15_LC_18_11_0.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIANPAC_15_LC_18_11_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNIANPAC_15_LC_18_11_0 (
            .in0(N__75148),
            .in1(N__90025),
            .in2(N__69110),
            .in3(N__76861),
            .lcout(clk_en_48),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_42_RNI6QCRA_15_LC_18_11_1.C_ON=1'b0;
    defparam shift_srl_42_RNI6QCRA_15_LC_18_11_1.SEQ_MODE=4'b0000;
    defparam shift_srl_42_RNI6QCRA_15_LC_18_11_1.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_42_RNI6QCRA_15_LC_18_11_1 (
            .in0(N__90022),
            .in1(N__69095),
            .in2(_gnd_net_),
            .in3(N__73239),
            .lcout(clk_en_43),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_23_RNI0DK37_15_LC_18_11_2.C_ON=1'b0;
    defparam shift_srl_23_RNI0DK37_15_LC_18_11_2.SEQ_MODE=4'b0000;
    defparam shift_srl_23_RNI0DK37_15_LC_18_11_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_23_RNI0DK37_15_LC_18_11_2 (
            .in0(N__69304),
            .in1(N__74479),
            .in2(N__69277),
            .in3(N__69238),
            .lcout(),
            .ltout(shift_srl_23_RNI0DK37Z0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_7_RNIEFOK9_15_LC_18_11_3.C_ON=1'b0;
    defparam shift_srl_7_RNIEFOK9_15_LC_18_11_3.SEQ_MODE=4'b0000;
    defparam shift_srl_7_RNIEFOK9_15_LC_18_11_3.LUT_INIT=16'b1111000010101010;
    LogicCell40 shift_srl_7_RNIEFOK9_15_LC_18_11_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__69196),
            .in3(N__69192),
            .lcout(rco_c_37),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_43_RNIO436B_15_LC_18_11_4.C_ON=1'b0;
    defparam shift_srl_43_RNIO436B_15_LC_18_11_4.SEQ_MODE=4'b0000;
    defparam shift_srl_43_RNIO436B_15_LC_18_11_4.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_43_RNIO436B_15_LC_18_11_4 (
            .in0(N__73240),
            .in1(N__73279),
            .in2(N__69109),
            .in3(N__90024),
            .lcout(clk_en_44),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_41_RNIQ72KA_15_LC_18_11_5.C_ON=1'b0;
    defparam shift_srl_41_RNIQ72KA_15_LC_18_11_5.SEQ_MODE=4'b0000;
    defparam shift_srl_41_RNIQ72KA_15_LC_18_11_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_41_RNIQ72KA_15_LC_18_11_5 (
            .in0(N__74763),
            .in1(N__81289),
            .in2(N__74700),
            .in3(N__78786),
            .lcout(rco_c_41),
            .ltout(rco_c_41_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_45_RNIV52OB_15_LC_18_11_6.C_ON=1'b0;
    defparam shift_srl_45_RNIV52OB_15_LC_18_11_6.SEQ_MODE=4'b0000;
    defparam shift_srl_45_RNIV52OB_15_LC_18_11_6.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_45_RNIV52OB_15_LC_18_11_6 (
            .in0(N__75147),
            .in1(N__90023),
            .in2(N__69133),
            .in3(N__76189),
            .lcout(clk_en_46),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIBJVKB_15_LC_18_11_7.C_ON=1'b0;
    defparam shift_srl_0_RNIBJVKB_15_LC_18_11_7.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIBJVKB_15_LC_18_11_7.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_0_RNIBJVKB_15_LC_18_11_7 (
            .in0(N__90026),
            .in1(N__69102),
            .in2(_gnd_net_),
            .in3(N__75146),
            .lcout(clk_en_45),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_44_0_LC_18_12_0.C_ON=1'b0;
    defparam shift_srl_44_0_LC_18_12_0.SEQ_MODE=4'b1000;
    defparam shift_srl_44_0_LC_18_12_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_44_0_LC_18_12_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73291),
            .lcout(shift_srl_44Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93189),
            .ce(N__71211),
            .sr(_gnd_net_));
    defparam shift_srl_44_1_LC_18_12_1.C_ON=1'b0;
    defparam shift_srl_44_1_LC_18_12_1.SEQ_MODE=4'b1000;
    defparam shift_srl_44_1_LC_18_12_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_44_1_LC_18_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69058),
            .lcout(shift_srl_44Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93189),
            .ce(N__71211),
            .sr(_gnd_net_));
    defparam shift_srl_44_2_LC_18_12_2.C_ON=1'b0;
    defparam shift_srl_44_2_LC_18_12_2.SEQ_MODE=4'b1000;
    defparam shift_srl_44_2_LC_18_12_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_44_2_LC_18_12_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69052),
            .lcout(shift_srl_44Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93189),
            .ce(N__71211),
            .sr(_gnd_net_));
    defparam shift_srl_44_3_LC_18_12_3.C_ON=1'b0;
    defparam shift_srl_44_3_LC_18_12_3.SEQ_MODE=4'b1000;
    defparam shift_srl_44_3_LC_18_12_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_44_3_LC_18_12_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69358),
            .lcout(shift_srl_44Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93189),
            .ce(N__71211),
            .sr(_gnd_net_));
    defparam shift_srl_44_4_LC_18_12_4.C_ON=1'b0;
    defparam shift_srl_44_4_LC_18_12_4.SEQ_MODE=4'b1000;
    defparam shift_srl_44_4_LC_18_12_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_44_4_LC_18_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69352),
            .lcout(shift_srl_44Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93189),
            .ce(N__71211),
            .sr(_gnd_net_));
    defparam shift_srl_44_5_LC_18_12_5.C_ON=1'b0;
    defparam shift_srl_44_5_LC_18_12_5.SEQ_MODE=4'b1000;
    defparam shift_srl_44_5_LC_18_12_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_44_5_LC_18_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69346),
            .lcout(shift_srl_44Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93189),
            .ce(N__71211),
            .sr(_gnd_net_));
    defparam shift_srl_44_6_LC_18_12_6.C_ON=1'b0;
    defparam shift_srl_44_6_LC_18_12_6.SEQ_MODE=4'b1000;
    defparam shift_srl_44_6_LC_18_12_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_44_6_LC_18_12_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69340),
            .lcout(shift_srl_44Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93189),
            .ce(N__71211),
            .sr(_gnd_net_));
    defparam shift_srl_44_7_LC_18_12_7.C_ON=1'b0;
    defparam shift_srl_44_7_LC_18_12_7.SEQ_MODE=4'b1000;
    defparam shift_srl_44_7_LC_18_12_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_44_7_LC_18_12_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69334),
            .lcout(shift_srl_44Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93189),
            .ce(N__71211),
            .sr(_gnd_net_));
    defparam shift_srl_48_0_LC_18_13_0.C_ON=1'b0;
    defparam shift_srl_48_0_LC_18_13_0.SEQ_MODE=4'b1000;
    defparam shift_srl_48_0_LC_18_13_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_48_0_LC_18_13_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76612),
            .lcout(shift_srl_48Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93168),
            .ce(N__73379),
            .sr(_gnd_net_));
    defparam shift_srl_48_1_LC_18_13_1.C_ON=1'b0;
    defparam shift_srl_48_1_LC_18_13_1.SEQ_MODE=4'b1000;
    defparam shift_srl_48_1_LC_18_13_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_48_1_LC_18_13_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69328),
            .lcout(shift_srl_48Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93168),
            .ce(N__73379),
            .sr(_gnd_net_));
    defparam shift_srl_48_2_LC_18_13_2.C_ON=1'b0;
    defparam shift_srl_48_2_LC_18_13_2.SEQ_MODE=4'b1000;
    defparam shift_srl_48_2_LC_18_13_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_48_2_LC_18_13_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69322),
            .lcout(shift_srl_48Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93168),
            .ce(N__73379),
            .sr(_gnd_net_));
    defparam shift_srl_48_3_LC_18_13_3.C_ON=1'b0;
    defparam shift_srl_48_3_LC_18_13_3.SEQ_MODE=4'b1000;
    defparam shift_srl_48_3_LC_18_13_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_48_3_LC_18_13_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69316),
            .lcout(shift_srl_48Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93168),
            .ce(N__73379),
            .sr(_gnd_net_));
    defparam shift_srl_48_4_LC_18_13_4.C_ON=1'b0;
    defparam shift_srl_48_4_LC_18_13_4.SEQ_MODE=4'b1000;
    defparam shift_srl_48_4_LC_18_13_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_48_4_LC_18_13_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69310),
            .lcout(shift_srl_48Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93168),
            .ce(N__73379),
            .sr(_gnd_net_));
    defparam shift_srl_48_5_LC_18_13_5.C_ON=1'b0;
    defparam shift_srl_48_5_LC_18_13_5.SEQ_MODE=4'b1000;
    defparam shift_srl_48_5_LC_18_13_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_48_5_LC_18_13_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69469),
            .lcout(shift_srl_48Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93168),
            .ce(N__73379),
            .sr(_gnd_net_));
    defparam shift_srl_48_6_LC_18_13_6.C_ON=1'b0;
    defparam shift_srl_48_6_LC_18_13_6.SEQ_MODE=4'b1000;
    defparam shift_srl_48_6_LC_18_13_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_48_6_LC_18_13_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69463),
            .lcout(shift_srl_48Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93168),
            .ce(N__73379),
            .sr(_gnd_net_));
    defparam shift_srl_48_10_LC_18_13_7.C_ON=1'b0;
    defparam shift_srl_48_10_LC_18_13_7.SEQ_MODE=4'b1000;
    defparam shift_srl_48_10_LC_18_13_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_48_10_LC_18_13_7 (
            .in0(N__71329),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_48Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93168),
            .ce(N__73379),
            .sr(_gnd_net_));
    defparam shift_srl_94_RNI2F961_15_LC_18_14_0.C_ON=1'b0;
    defparam shift_srl_94_RNI2F961_15_LC_18_14_0.SEQ_MODE=4'b0000;
    defparam shift_srl_94_RNI2F961_15_LC_18_14_0.LUT_INIT=16'b1110111000100010;
    LogicCell40 shift_srl_94_RNI2F961_15_LC_18_14_0 (
            .in0(_gnd_net_),
            .in1(N__72717),
            .in2(_gnd_net_),
            .in3(N__69403),
            .lcout(shift_srl_94_RNI2F961Z0Z_15),
            .ltout(shift_srl_94_RNI2F961Z0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_33_RNILVDN1_15_LC_18_14_1.C_ON=1'b0;
    defparam shift_srl_33_RNILVDN1_15_LC_18_14_1.SEQ_MODE=4'b0000;
    defparam shift_srl_33_RNILVDN1_15_LC_18_14_1.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_33_RNILVDN1_15_LC_18_14_1 (
            .in0(N__87323),
            .in1(N__83349),
            .in2(N__69457),
            .in3(N__85575),
            .lcout(rco_int_0_a2_0_a2_99_m6_0_a2_9_sx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_98_RNIA7Q31_15_LC_18_14_2.C_ON=1'b0;
    defparam shift_srl_98_RNIA7Q31_15_LC_18_14_2.SEQ_MODE=4'b0000;
    defparam shift_srl_98_RNIA7Q31_15_LC_18_14_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_98_RNIA7Q31_15_LC_18_14_2 (
            .in0(N__69449),
            .in1(N__69418),
            .in2(N__70852),
            .in3(N__69369),
            .lcout(shift_srl_98_RNIA7Q31Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_37_RNI094V1_15_LC_18_14_3.C_ON=1'b0;
    defparam shift_srl_37_RNI094V1_15_LC_18_14_3.SEQ_MODE=4'b0000;
    defparam shift_srl_37_RNI094V1_15_LC_18_14_3.LUT_INIT=16'b1111111101010101;
    LogicCell40 shift_srl_37_RNI094V1_15_LC_18_14_3 (
            .in0(N__71554),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71305),
            .lcout(),
            .ltout(rco_int_0_a2_0_a2_99_m6_0_a2_9_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_33_RNI3MSM5_15_LC_18_14_4.C_ON=1'b0;
    defparam shift_srl_33_RNI3MSM5_15_LC_18_14_4.SEQ_MODE=4'b0000;
    defparam shift_srl_33_RNI3MSM5_15_LC_18_14_4.LUT_INIT=16'b0000000000001000;
    LogicCell40 shift_srl_33_RNI3MSM5_15_LC_18_14_4 (
            .in0(N__71389),
            .in1(N__69397),
            .in2(N__69391),
            .in3(N__69388),
            .lcout(rco_int_0_a2_0_a2_99_m6_0_a2_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_95_15_LC_18_14_5.C_ON=1'b0;
    defparam shift_srl_95_15_LC_18_14_5.SEQ_MODE=4'b1000;
    defparam shift_srl_95_15_LC_18_14_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_95_15_LC_18_14_5 (
            .in0(N__69559),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_95Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93151),
            .ce(N__69553),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_34_LC_18_14_6.C_ON=1'b0;
    defparam rco_obuf_RNO_34_LC_18_14_6.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_34_LC_18_14_6.LUT_INIT=16'b1000000000000000;
    LogicCell40 rco_obuf_RNO_34_LC_18_14_6 (
            .in0(N__83350),
            .in1(N__87363),
            .in2(N__85579),
            .in3(N__87324),
            .lcout(rco_c_34),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_95_14_LC_18_14_7.C_ON=1'b0;
    defparam shift_srl_95_14_LC_18_14_7.SEQ_MODE=4'b1000;
    defparam shift_srl_95_14_LC_18_14_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_95_14_LC_18_14_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69574),
            .lcout(shift_srl_95Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93151),
            .ce(N__69553),
            .sr(_gnd_net_));
    defparam shift_srl_40_fast_RNI31DI_15_LC_18_15_0.C_ON=1'b0;
    defparam shift_srl_40_fast_RNI31DI_15_LC_18_15_0.SEQ_MODE=4'b0000;
    defparam shift_srl_40_fast_RNI31DI_15_LC_18_15_0.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_40_fast_RNI31DI_15_LC_18_15_0 (
            .in0(N__69520),
            .in1(N__78797),
            .in2(_gnd_net_),
            .in3(N__69502),
            .lcout(rco_int_0_a2_0_a2_93_m6_0_a2_4_7_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_40_fast_15_LC_18_15_1.C_ON=1'b0;
    defparam shift_srl_40_fast_15_LC_18_15_1.SEQ_MODE=4'b1000;
    defparam shift_srl_40_fast_15_LC_18_15_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_40_fast_15_LC_18_15_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69496),
            .lcout(shift_srl_40_fastZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93131),
            .ce(N__69673),
            .sr(_gnd_net_));
    defparam shift_srl_40_14_LC_18_15_2.C_ON=1'b0;
    defparam shift_srl_40_14_LC_18_15_2.SEQ_MODE=4'b1000;
    defparam shift_srl_40_14_LC_18_15_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_40_14_LC_18_15_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69487),
            .lcout(shift_srl_40Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93131),
            .ce(N__69673),
            .sr(_gnd_net_));
    defparam shift_srl_40_15_LC_18_15_3.C_ON=1'b0;
    defparam shift_srl_40_15_LC_18_15_3.SEQ_MODE=4'b1000;
    defparam shift_srl_40_15_LC_18_15_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_40_15_LC_18_15_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69495),
            .lcout(shift_srl_40Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93131),
            .ce(N__69673),
            .sr(_gnd_net_));
    defparam shift_srl_40_13_LC_18_15_4.C_ON=1'b0;
    defparam shift_srl_40_13_LC_18_15_4.SEQ_MODE=4'b1000;
    defparam shift_srl_40_13_LC_18_15_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_40_13_LC_18_15_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69481),
            .lcout(shift_srl_40Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93131),
            .ce(N__69673),
            .sr(_gnd_net_));
    defparam shift_srl_40_12_LC_18_15_5.C_ON=1'b0;
    defparam shift_srl_40_12_LC_18_15_5.SEQ_MODE=4'b1000;
    defparam shift_srl_40_12_LC_18_15_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_40_12_LC_18_15_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69475),
            .lcout(shift_srl_40Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93131),
            .ce(N__69673),
            .sr(_gnd_net_));
    defparam shift_srl_40_11_LC_18_15_6.C_ON=1'b0;
    defparam shift_srl_40_11_LC_18_15_6.SEQ_MODE=4'b1000;
    defparam shift_srl_40_11_LC_18_15_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_40_11_LC_18_15_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69679),
            .lcout(shift_srl_40Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93131),
            .ce(N__69673),
            .sr(_gnd_net_));
    defparam shift_srl_40_10_LC_18_15_7.C_ON=1'b0;
    defparam shift_srl_40_10_LC_18_15_7.SEQ_MODE=4'b1000;
    defparam shift_srl_40_10_LC_18_15_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_40_10_LC_18_15_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69694),
            .lcout(shift_srl_40Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93131),
            .ce(N__69673),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_30_LC_18_16_0.C_ON=1'b0;
    defparam rco_obuf_RNO_30_LC_18_16_0.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_30_LC_18_16_0.LUT_INIT=16'b1000100000000000;
    LogicCell40 rco_obuf_RNO_30_LC_18_16_0 (
            .in0(N__69658),
            .in1(N__83722),
            .in2(_gnd_net_),
            .in3(N__85179),
            .lcout(rco_c_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_30_0_LC_18_16_1.C_ON=1'b0;
    defparam shift_srl_30_0_LC_18_16_1.SEQ_MODE=4'b1000;
    defparam shift_srl_30_0_LC_18_16_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_30_0_LC_18_16_1 (
            .in0(N__83721),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_30Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93113),
            .ce(N__79834),
            .sr(_gnd_net_));
    defparam shift_srl_30_1_LC_18_16_2.C_ON=1'b0;
    defparam shift_srl_30_1_LC_18_16_2.SEQ_MODE=4'b1000;
    defparam shift_srl_30_1_LC_18_16_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_30_1_LC_18_16_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69631),
            .lcout(shift_srl_30Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93113),
            .ce(N__79834),
            .sr(_gnd_net_));
    defparam shift_srl_30_2_LC_18_16_3.C_ON=1'b0;
    defparam shift_srl_30_2_LC_18_16_3.SEQ_MODE=4'b1000;
    defparam shift_srl_30_2_LC_18_16_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_30_2_LC_18_16_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69625),
            .lcout(shift_srl_30Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93113),
            .ce(N__79834),
            .sr(_gnd_net_));
    defparam shift_srl_30_3_LC_18_16_4.C_ON=1'b0;
    defparam shift_srl_30_3_LC_18_16_4.SEQ_MODE=4'b1000;
    defparam shift_srl_30_3_LC_18_16_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_30_3_LC_18_16_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69619),
            .lcout(shift_srl_30Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93113),
            .ce(N__79834),
            .sr(_gnd_net_));
    defparam shift_srl_30_4_LC_18_16_5.C_ON=1'b0;
    defparam shift_srl_30_4_LC_18_16_5.SEQ_MODE=4'b1000;
    defparam shift_srl_30_4_LC_18_16_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_30_4_LC_18_16_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69613),
            .lcout(shift_srl_30Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93113),
            .ce(N__79834),
            .sr(_gnd_net_));
    defparam shift_srl_30_5_LC_18_16_6.C_ON=1'b0;
    defparam shift_srl_30_5_LC_18_16_6.SEQ_MODE=4'b1000;
    defparam shift_srl_30_5_LC_18_16_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_30_5_LC_18_16_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69607),
            .lcout(shift_srl_30Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93113),
            .ce(N__79834),
            .sr(_gnd_net_));
    defparam shift_srl_30_6_LC_18_16_7.C_ON=1'b0;
    defparam shift_srl_30_6_LC_18_16_7.SEQ_MODE=4'b1000;
    defparam shift_srl_30_6_LC_18_16_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_30_6_LC_18_16_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69601),
            .lcout(shift_srl_30Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93113),
            .ce(N__79834),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNI9RIL9_15_LC_18_17_0.C_ON=1'b0;
    defparam shift_srl_0_RNI9RIL9_15_LC_18_17_0.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNI9RIL9_15_LC_18_17_0.LUT_INIT=16'b1100110000000000;
    LogicCell40 shift_srl_0_RNI9RIL9_15_LC_18_17_0 (
            .in0(_gnd_net_),
            .in1(N__90431),
            .in2(_gnd_net_),
            .in3(N__81322),
            .lcout(clk_en_38),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_38_0_LC_18_17_1.C_ON=1'b0;
    defparam shift_srl_38_0_LC_18_17_1.SEQ_MODE=4'b1000;
    defparam shift_srl_38_0_LC_18_17_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_38_0_LC_18_17_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79744),
            .lcout(shift_srl_38Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93084),
            .ce(N__69773),
            .sr(_gnd_net_));
    defparam shift_srl_38_1_LC_18_17_2.C_ON=1'b0;
    defparam shift_srl_38_1_LC_18_17_2.SEQ_MODE=4'b1000;
    defparam shift_srl_38_1_LC_18_17_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_38_1_LC_18_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69736),
            .lcout(shift_srl_38Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93084),
            .ce(N__69773),
            .sr(_gnd_net_));
    defparam shift_srl_38_2_LC_18_17_3.C_ON=1'b0;
    defparam shift_srl_38_2_LC_18_17_3.SEQ_MODE=4'b1000;
    defparam shift_srl_38_2_LC_18_17_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_38_2_LC_18_17_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69730),
            .lcout(shift_srl_38Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93084),
            .ce(N__69773),
            .sr(_gnd_net_));
    defparam shift_srl_38_3_LC_18_17_4.C_ON=1'b0;
    defparam shift_srl_38_3_LC_18_17_4.SEQ_MODE=4'b1000;
    defparam shift_srl_38_3_LC_18_17_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_38_3_LC_18_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69724),
            .lcout(shift_srl_38Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93084),
            .ce(N__69773),
            .sr(_gnd_net_));
    defparam shift_srl_38_4_LC_18_17_5.C_ON=1'b0;
    defparam shift_srl_38_4_LC_18_17_5.SEQ_MODE=4'b1000;
    defparam shift_srl_38_4_LC_18_17_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_38_4_LC_18_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69718),
            .lcout(shift_srl_38Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93084),
            .ce(N__69773),
            .sr(_gnd_net_));
    defparam shift_srl_38_5_LC_18_17_6.C_ON=1'b0;
    defparam shift_srl_38_5_LC_18_17_6.SEQ_MODE=4'b1000;
    defparam shift_srl_38_5_LC_18_17_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_38_5_LC_18_17_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69712),
            .lcout(shift_srl_38Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93084),
            .ce(N__69773),
            .sr(_gnd_net_));
    defparam shift_srl_38_6_LC_18_17_7.C_ON=1'b0;
    defparam shift_srl_38_6_LC_18_17_7.SEQ_MODE=4'b1000;
    defparam shift_srl_38_6_LC_18_17_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_38_6_LC_18_17_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69706),
            .lcout(shift_srl_38Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93084),
            .ce(N__69773),
            .sr(_gnd_net_));
    defparam shift_srl_38_10_LC_18_18_0.C_ON=1'b0;
    defparam shift_srl_38_10_LC_18_18_0.SEQ_MODE=4'b1000;
    defparam shift_srl_38_10_LC_18_18_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_38_10_LC_18_18_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69802),
            .lcout(shift_srl_38Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93114),
            .ce(N__69780),
            .sr(_gnd_net_));
    defparam shift_srl_38_11_LC_18_18_1.C_ON=1'b0;
    defparam shift_srl_38_11_LC_18_18_1.SEQ_MODE=4'b1000;
    defparam shift_srl_38_11_LC_18_18_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_38_11_LC_18_18_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69826),
            .lcout(shift_srl_38Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93114),
            .ce(N__69780),
            .sr(_gnd_net_));
    defparam shift_srl_38_12_LC_18_18_2.C_ON=1'b0;
    defparam shift_srl_38_12_LC_18_18_2.SEQ_MODE=4'b1000;
    defparam shift_srl_38_12_LC_18_18_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_38_12_LC_18_18_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69820),
            .lcout(shift_srl_38Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93114),
            .ce(N__69780),
            .sr(_gnd_net_));
    defparam shift_srl_38_15_LC_18_18_5.C_ON=1'b0;
    defparam shift_srl_38_15_LC_18_18_5.SEQ_MODE=4'b1000;
    defparam shift_srl_38_15_LC_18_18_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_38_15_LC_18_18_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69808),
            .lcout(shift_srl_38Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93114),
            .ce(N__69780),
            .sr(_gnd_net_));
    defparam shift_srl_38_9_LC_18_18_6.C_ON=1'b0;
    defparam shift_srl_38_9_LC_18_18_6.SEQ_MODE=4'b1000;
    defparam shift_srl_38_9_LC_18_18_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_38_9_LC_18_18_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69790),
            .lcout(shift_srl_38Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93114),
            .ce(N__69780),
            .sr(_gnd_net_));
    defparam shift_srl_38_8_LC_18_18_7.C_ON=1'b0;
    defparam shift_srl_38_8_LC_18_18_7.SEQ_MODE=4'b1000;
    defparam shift_srl_38_8_LC_18_18_7.LUT_INIT=16'b1100110011001100;
    LogicCell40 shift_srl_38_8_LC_18_18_7 (
            .in0(_gnd_net_),
            .in1(N__69796),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_38Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93114),
            .ce(N__69780),
            .sr(_gnd_net_));
    defparam shift_srl_158_10_LC_18_19_0.C_ON=1'b0;
    defparam shift_srl_158_10_LC_18_19_0.SEQ_MODE=4'b1000;
    defparam shift_srl_158_10_LC_18_19_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_158_10_LC_18_19_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69973),
            .lcout(shift_srl_158Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93132),
            .ce(N__70044),
            .sr(_gnd_net_));
    defparam shift_srl_158_11_LC_18_19_1.C_ON=1'b0;
    defparam shift_srl_158_11_LC_18_19_1.SEQ_MODE=4'b1000;
    defparam shift_srl_158_11_LC_18_19_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_158_11_LC_18_19_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69754),
            .lcout(shift_srl_158Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93132),
            .ce(N__70044),
            .sr(_gnd_net_));
    defparam shift_srl_158_12_LC_18_19_2.C_ON=1'b0;
    defparam shift_srl_158_12_LC_18_19_2.SEQ_MODE=4'b1000;
    defparam shift_srl_158_12_LC_18_19_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_158_12_LC_18_19_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69748),
            .lcout(shift_srl_158Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93132),
            .ce(N__70044),
            .sr(_gnd_net_));
    defparam shift_srl_158_13_LC_18_19_3.C_ON=1'b0;
    defparam shift_srl_158_13_LC_18_19_3.SEQ_MODE=4'b1000;
    defparam shift_srl_158_13_LC_18_19_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_158_13_LC_18_19_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69742),
            .lcout(shift_srl_158Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93132),
            .ce(N__70044),
            .sr(_gnd_net_));
    defparam shift_srl_158_14_LC_18_19_4.C_ON=1'b0;
    defparam shift_srl_158_14_LC_18_19_4.SEQ_MODE=4'b1000;
    defparam shift_srl_158_14_LC_18_19_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_158_14_LC_18_19_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69985),
            .lcout(shift_srl_158Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93132),
            .ce(N__70044),
            .sr(_gnd_net_));
    defparam shift_srl_158_15_LC_18_19_5.C_ON=1'b0;
    defparam shift_srl_158_15_LC_18_19_5.SEQ_MODE=4'b1000;
    defparam shift_srl_158_15_LC_18_19_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_158_15_LC_18_19_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69979),
            .lcout(shift_srl_158Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93132),
            .ce(N__70044),
            .sr(_gnd_net_));
    defparam shift_srl_158_9_LC_18_19_6.C_ON=1'b0;
    defparam shift_srl_158_9_LC_18_19_6.SEQ_MODE=4'b1000;
    defparam shift_srl_158_9_LC_18_19_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_158_9_LC_18_19_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69961),
            .lcout(shift_srl_158Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93132),
            .ce(N__70044),
            .sr(_gnd_net_));
    defparam shift_srl_158_8_LC_18_19_7.C_ON=1'b0;
    defparam shift_srl_158_8_LC_18_19_7.SEQ_MODE=4'b1000;
    defparam shift_srl_158_8_LC_18_19_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_158_8_LC_18_19_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69967),
            .lcout(shift_srl_158Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93132),
            .ce(N__70044),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_158_LC_18_20_0.C_ON=1'b0;
    defparam rco_obuf_RNO_158_LC_18_20_0.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_158_LC_18_20_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 rco_obuf_RNO_158_LC_18_20_0 (
            .in0(N__77278),
            .in1(N__77903),
            .in2(N__87869),
            .in3(N__77551),
            .lcout(rco_c_158),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_157_LC_18_20_1.C_ON=1'b0;
    defparam rco_obuf_RNO_157_LC_18_20_1.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_157_LC_18_20_1.LUT_INIT=16'b1100000000000000;
    LogicCell40 rco_obuf_RNO_157_LC_18_20_1 (
            .in0(_gnd_net_),
            .in1(N__77902),
            .in2(N__77556),
            .in3(N__87844),
            .lcout(rco_c_157),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_145_RNI4O2P61_15_LC_18_20_3.C_ON=1'b0;
    defparam shift_srl_145_RNI4O2P61_15_LC_18_20_3.SEQ_MODE=4'b0000;
    defparam shift_srl_145_RNI4O2P61_15_LC_18_20_3.LUT_INIT=16'b0000010000000000;
    LogicCell40 shift_srl_145_RNI4O2P61_15_LC_18_20_3 (
            .in0(N__69910),
            .in1(N__85172),
            .in2(N__71956),
            .in3(N__75077),
            .lcout(rco_c_153),
            .ltout(rco_c_153_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_161_RNIHFCL81_15_LC_18_20_4.C_ON=1'b0;
    defparam shift_srl_161_RNIHFCL81_15_LC_18_20_4.SEQ_MODE=4'b0000;
    defparam shift_srl_161_RNIHFCL81_15_LC_18_20_4.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_161_RNIHFCL81_15_LC_18_20_4 (
            .in0(N__77377),
            .in1(N__90488),
            .in2(N__69892),
            .in3(N__69842),
            .lcout(clk_en_162),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_160_RNIFA2R1_15_LC_18_20_5.C_ON=1'b0;
    defparam shift_srl_160_RNIFA2R1_15_LC_18_20_5.SEQ_MODE=4'b0000;
    defparam shift_srl_160_RNIFA2R1_15_LC_18_20_5.LUT_INIT=16'b1100110000000000;
    LogicCell40 shift_srl_160_RNIFA2R1_15_LC_18_20_5 (
            .in0(_gnd_net_),
            .in1(N__71634),
            .in2(_gnd_net_),
            .in3(N__77430),
            .lcout(shift_srl_160_RNIFA2R1Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_157_RNIPSMT71_15_LC_18_20_6.C_ON=1'b0;
    defparam shift_srl_157_RNIPSMT71_15_LC_18_20_6.SEQ_MODE=4'b0000;
    defparam shift_srl_157_RNIPSMT71_15_LC_18_20_6.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_157_RNIPSMT71_15_LC_18_20_6 (
            .in0(N__87842),
            .in1(N__90487),
            .in2(N__77907),
            .in3(N__77547),
            .lcout(clk_en_158),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_155_RNIAOD371_15_LC_18_20_7.C_ON=1'b0;
    defparam shift_srl_155_RNIAOD371_15_LC_18_20_7.SEQ_MODE=4'b0000;
    defparam shift_srl_155_RNIAOD371_15_LC_18_20_7.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_155_RNIAOD371_15_LC_18_20_7 (
            .in0(N__77652),
            .in1(N__77611),
            .in2(N__90553),
            .in3(N__87843),
            .lcout(clk_en_156),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_156_10_LC_18_21_0.C_ON=1'b0;
    defparam shift_srl_156_10_LC_18_21_0.SEQ_MODE=4'b1000;
    defparam shift_srl_156_10_LC_18_21_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_156_10_LC_18_21_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69991),
            .lcout(shift_srl_156Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93169),
            .ce(N__70107),
            .sr(_gnd_net_));
    defparam shift_srl_156_11_LC_18_21_1.C_ON=1'b0;
    defparam shift_srl_156_11_LC_18_21_1.SEQ_MODE=4'b1000;
    defparam shift_srl_156_11_LC_18_21_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_156_11_LC_18_21_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70021),
            .lcout(shift_srl_156Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93169),
            .ce(N__70107),
            .sr(_gnd_net_));
    defparam shift_srl_156_12_LC_18_21_2.C_ON=1'b0;
    defparam shift_srl_156_12_LC_18_21_2.SEQ_MODE=4'b1000;
    defparam shift_srl_156_12_LC_18_21_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_156_12_LC_18_21_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70015),
            .lcout(shift_srl_156Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93169),
            .ce(N__70107),
            .sr(_gnd_net_));
    defparam shift_srl_156_13_LC_18_21_3.C_ON=1'b0;
    defparam shift_srl_156_13_LC_18_21_3.SEQ_MODE=4'b1000;
    defparam shift_srl_156_13_LC_18_21_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_156_13_LC_18_21_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70009),
            .lcout(shift_srl_156Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93169),
            .ce(N__70107),
            .sr(_gnd_net_));
    defparam shift_srl_156_14_LC_18_21_4.C_ON=1'b0;
    defparam shift_srl_156_14_LC_18_21_4.SEQ_MODE=4'b1000;
    defparam shift_srl_156_14_LC_18_21_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_156_14_LC_18_21_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70003),
            .lcout(shift_srl_156Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93169),
            .ce(N__70107),
            .sr(_gnd_net_));
    defparam shift_srl_156_15_LC_18_21_5.C_ON=1'b0;
    defparam shift_srl_156_15_LC_18_21_5.SEQ_MODE=4'b1000;
    defparam shift_srl_156_15_LC_18_21_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_156_15_LC_18_21_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69997),
            .lcout(shift_srl_156Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93169),
            .ce(N__70107),
            .sr(_gnd_net_));
    defparam shift_srl_156_9_LC_18_21_6.C_ON=1'b0;
    defparam shift_srl_156_9_LC_18_21_6.SEQ_MODE=4'b1000;
    defparam shift_srl_156_9_LC_18_21_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_156_9_LC_18_21_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70114),
            .lcout(shift_srl_156Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93169),
            .ce(N__70107),
            .sr(_gnd_net_));
    defparam shift_srl_156_8_LC_18_21_7.C_ON=1'b0;
    defparam shift_srl_156_8_LC_18_21_7.SEQ_MODE=4'b1000;
    defparam shift_srl_156_8_LC_18_21_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_156_8_LC_18_21_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70120),
            .lcout(shift_srl_156Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93169),
            .ce(N__70107),
            .sr(_gnd_net_));
    defparam shift_srl_183_RNIJQ6N6_15_LC_18_22_0.C_ON=1'b0;
    defparam shift_srl_183_RNIJQ6N6_15_LC_18_22_0.SEQ_MODE=4'b0000;
    defparam shift_srl_183_RNIJQ6N6_15_LC_18_22_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_183_RNIJQ6N6_15_LC_18_22_0 (
            .in0(N__82334),
            .in1(N__75830),
            .in2(N__70069),
            .in3(N__87988),
            .lcout(g0_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_183_15_LC_18_22_1.C_ON=1'b0;
    defparam shift_srl_183_15_LC_18_22_1.SEQ_MODE=4'b1000;
    defparam shift_srl_183_15_LC_18_22_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_183_15_LC_18_22_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71764),
            .lcout(shift_srl_183Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93190),
            .ce(N__71869),
            .sr(_gnd_net_));
    defparam shift_srl_183_RNILCAQ2_15_LC_18_22_2.C_ON=1'b0;
    defparam shift_srl_183_RNILCAQ2_15_LC_18_22_2.SEQ_MODE=4'b0000;
    defparam shift_srl_183_RNILCAQ2_15_LC_18_22_2.LUT_INIT=16'b1100110000000000;
    LogicCell40 shift_srl_183_RNILCAQ2_15_LC_18_22_2 (
            .in0(_gnd_net_),
            .in1(N__70064),
            .in2(_gnd_net_),
            .in3(N__75829),
            .lcout(rco_int_0_a3_0_a2_0_183),
            .ltout(rco_int_0_a3_0_a2_0_183_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_184_RNISMFI5_15_LC_18_22_3.C_ON=1'b0;
    defparam shift_srl_184_RNISMFI5_15_LC_18_22_3.SEQ_MODE=4'b0000;
    defparam shift_srl_184_RNISMFI5_15_LC_18_22_3.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_184_RNISMFI5_15_LC_18_22_3 (
            .in0(N__91688),
            .in1(N__90486),
            .in2(N__70081),
            .in3(N__84236),
            .lcout(),
            .ltout(clk_en_0_a2_0_a2_1_187_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_184_RNI9QERE1_15_LC_18_22_4.C_ON=1'b0;
    defparam shift_srl_184_RNI9QERE1_15_LC_18_22_4.SEQ_MODE=4'b0000;
    defparam shift_srl_184_RNI9QERE1_15_LC_18_22_4.LUT_INIT=16'b0000010000000000;
    LogicCell40 shift_srl_184_RNI9QERE1_15_LC_18_22_4 (
            .in0(N__70075),
            .in1(N__77823),
            .in2(N__70078),
            .in3(N__79532),
            .lcout(clk_en_187),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_186_RNIH8MC4_15_LC_18_22_5.C_ON=1'b0;
    defparam shift_srl_186_RNIH8MC4_15_LC_18_22_5.SEQ_MODE=4'b0000;
    defparam shift_srl_186_RNIH8MC4_15_LC_18_22_5.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_186_RNIH8MC4_15_LC_18_22_5 (
            .in0(N__91814),
            .in1(N__91762),
            .in2(N__88005),
            .in3(N__82335),
            .lcout(clk_en_0_a2_0_a2_sx_187),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_183_0_LC_18_22_6.C_ON=1'b0;
    defparam shift_srl_183_0_LC_18_22_6.SEQ_MODE=4'b1000;
    defparam shift_srl_183_0_LC_18_22_6.LUT_INIT=16'b1100110011001100;
    LogicCell40 shift_srl_183_0_LC_18_22_6 (
            .in0(_gnd_net_),
            .in1(N__70065),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_183Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93190),
            .ce(N__71869),
            .sr(_gnd_net_));
    defparam shift_srl_183_1_LC_18_22_7.C_ON=1'b0;
    defparam shift_srl_183_1_LC_18_22_7.SEQ_MODE=4'b1000;
    defparam shift_srl_183_1_LC_18_22_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_183_1_LC_18_22_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70051),
            .lcout(shift_srl_183Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93190),
            .ce(N__71869),
            .sr(_gnd_net_));
    defparam shift_srl_187_10_LC_18_23_0.C_ON=1'b0;
    defparam shift_srl_187_10_LC_18_23_0.SEQ_MODE=4'b1000;
    defparam shift_srl_187_10_LC_18_23_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_187_10_LC_18_23_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70171),
            .lcout(shift_srl_187Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93210),
            .ce(N__70153),
            .sr(_gnd_net_));
    defparam shift_srl_187_11_LC_18_23_1.C_ON=1'b0;
    defparam shift_srl_187_11_LC_18_23_1.SEQ_MODE=4'b1000;
    defparam shift_srl_187_11_LC_18_23_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_187_11_LC_18_23_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70201),
            .lcout(shift_srl_187Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93210),
            .ce(N__70153),
            .sr(_gnd_net_));
    defparam shift_srl_187_12_LC_18_23_2.C_ON=1'b0;
    defparam shift_srl_187_12_LC_18_23_2.SEQ_MODE=4'b1000;
    defparam shift_srl_187_12_LC_18_23_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_187_12_LC_18_23_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70195),
            .lcout(shift_srl_187Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93210),
            .ce(N__70153),
            .sr(_gnd_net_));
    defparam shift_srl_187_13_LC_18_23_3.C_ON=1'b0;
    defparam shift_srl_187_13_LC_18_23_3.SEQ_MODE=4'b1000;
    defparam shift_srl_187_13_LC_18_23_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_187_13_LC_18_23_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70189),
            .lcout(shift_srl_187Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93210),
            .ce(N__70153),
            .sr(_gnd_net_));
    defparam shift_srl_187_14_LC_18_23_4.C_ON=1'b0;
    defparam shift_srl_187_14_LC_18_23_4.SEQ_MODE=4'b1000;
    defparam shift_srl_187_14_LC_18_23_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_187_14_LC_18_23_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70183),
            .lcout(shift_srl_187Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93210),
            .ce(N__70153),
            .sr(_gnd_net_));
    defparam shift_srl_187_15_LC_18_23_5.C_ON=1'b0;
    defparam shift_srl_187_15_LC_18_23_5.SEQ_MODE=4'b1000;
    defparam shift_srl_187_15_LC_18_23_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_187_15_LC_18_23_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70177),
            .lcout(shift_srl_187Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93210),
            .ce(N__70153),
            .sr(_gnd_net_));
    defparam shift_srl_187_9_LC_18_23_6.C_ON=1'b0;
    defparam shift_srl_187_9_LC_18_23_6.SEQ_MODE=4'b1000;
    defparam shift_srl_187_9_LC_18_23_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_187_9_LC_18_23_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70159),
            .lcout(shift_srl_187Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93210),
            .ce(N__70153),
            .sr(_gnd_net_));
    defparam shift_srl_187_8_LC_18_23_7.C_ON=1'b0;
    defparam shift_srl_187_8_LC_18_23_7.SEQ_MODE=4'b1000;
    defparam shift_srl_187_8_LC_18_23_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_187_8_LC_18_23_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70165),
            .lcout(shift_srl_187Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93210),
            .ce(N__70153),
            .sr(_gnd_net_));
    defparam shift_srl_194_10_LC_18_24_0.C_ON=1'b0;
    defparam shift_srl_194_10_LC_18_24_0.SEQ_MODE=4'b1000;
    defparam shift_srl_194_10_LC_18_24_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_194_10_LC_18_24_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70234),
            .lcout(shift_srl_194Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93229),
            .ce(N__72261),
            .sr(_gnd_net_));
    defparam shift_srl_194_11_LC_18_24_1.C_ON=1'b0;
    defparam shift_srl_194_11_LC_18_24_1.SEQ_MODE=4'b1000;
    defparam shift_srl_194_11_LC_18_24_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_194_11_LC_18_24_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70126),
            .lcout(shift_srl_194Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93229),
            .ce(N__72261),
            .sr(_gnd_net_));
    defparam shift_srl_194_12_LC_18_24_2.C_ON=1'b0;
    defparam shift_srl_194_12_LC_18_24_2.SEQ_MODE=4'b1000;
    defparam shift_srl_194_12_LC_18_24_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_194_12_LC_18_24_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70258),
            .lcout(shift_srl_194Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93229),
            .ce(N__72261),
            .sr(_gnd_net_));
    defparam shift_srl_194_13_LC_18_24_3.C_ON=1'b0;
    defparam shift_srl_194_13_LC_18_24_3.SEQ_MODE=4'b1000;
    defparam shift_srl_194_13_LC_18_24_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_194_13_LC_18_24_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70252),
            .lcout(shift_srl_194Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93229),
            .ce(N__72261),
            .sr(_gnd_net_));
    defparam shift_srl_194_14_LC_18_24_4.C_ON=1'b0;
    defparam shift_srl_194_14_LC_18_24_4.SEQ_MODE=4'b1000;
    defparam shift_srl_194_14_LC_18_24_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_194_14_LC_18_24_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70246),
            .lcout(shift_srl_194Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93229),
            .ce(N__72261),
            .sr(_gnd_net_));
    defparam shift_srl_194_15_LC_18_24_5.C_ON=1'b0;
    defparam shift_srl_194_15_LC_18_24_5.SEQ_MODE=4'b1000;
    defparam shift_srl_194_15_LC_18_24_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_194_15_LC_18_24_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70240),
            .lcout(shift_srl_194Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93229),
            .ce(N__72261),
            .sr(_gnd_net_));
    defparam shift_srl_194_9_LC_18_24_6.C_ON=1'b0;
    defparam shift_srl_194_9_LC_18_24_6.SEQ_MODE=4'b1000;
    defparam shift_srl_194_9_LC_18_24_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_194_9_LC_18_24_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70294),
            .lcout(shift_srl_194Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93229),
            .ce(N__72261),
            .sr(_gnd_net_));
    defparam shift_srl_194_2_LC_18_25_0.C_ON=1'b0;
    defparam shift_srl_194_2_LC_18_25_0.SEQ_MODE=4'b1000;
    defparam shift_srl_194_2_LC_18_25_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_194_2_LC_18_25_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70228),
            .lcout(shift_srl_194Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93249),
            .ce(N__72254),
            .sr(_gnd_net_));
    defparam shift_srl_194_3_LC_18_25_1.C_ON=1'b0;
    defparam shift_srl_194_3_LC_18_25_1.SEQ_MODE=4'b1000;
    defparam shift_srl_194_3_LC_18_25_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_194_3_LC_18_25_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70219),
            .lcout(shift_srl_194Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93249),
            .ce(N__72254),
            .sr(_gnd_net_));
    defparam shift_srl_194_4_LC_18_25_2.C_ON=1'b0;
    defparam shift_srl_194_4_LC_18_25_2.SEQ_MODE=4'b1000;
    defparam shift_srl_194_4_LC_18_25_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_194_4_LC_18_25_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70213),
            .lcout(shift_srl_194Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93249),
            .ce(N__72254),
            .sr(_gnd_net_));
    defparam shift_srl_194_5_LC_18_25_3.C_ON=1'b0;
    defparam shift_srl_194_5_LC_18_25_3.SEQ_MODE=4'b1000;
    defparam shift_srl_194_5_LC_18_25_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_194_5_LC_18_25_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70207),
            .lcout(shift_srl_194Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93249),
            .ce(N__72254),
            .sr(_gnd_net_));
    defparam shift_srl_194_6_LC_18_25_4.C_ON=1'b0;
    defparam shift_srl_194_6_LC_18_25_4.SEQ_MODE=4'b1000;
    defparam shift_srl_194_6_LC_18_25_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_194_6_LC_18_25_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70312),
            .lcout(shift_srl_194Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93249),
            .ce(N__72254),
            .sr(_gnd_net_));
    defparam shift_srl_194_7_LC_18_25_5.C_ON=1'b0;
    defparam shift_srl_194_7_LC_18_25_5.SEQ_MODE=4'b1000;
    defparam shift_srl_194_7_LC_18_25_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_194_7_LC_18_25_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70306),
            .lcout(shift_srl_194Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93249),
            .ce(N__72254),
            .sr(_gnd_net_));
    defparam shift_srl_194_8_LC_18_25_7.C_ON=1'b0;
    defparam shift_srl_194_8_LC_18_25_7.SEQ_MODE=4'b1000;
    defparam shift_srl_194_8_LC_18_25_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_194_8_LC_18_25_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70300),
            .lcout(shift_srl_194Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93249),
            .ce(N__72254),
            .sr(_gnd_net_));
    defparam shift_srl_175_0_LC_18_26_0.C_ON=1'b0;
    defparam shift_srl_175_0_LC_18_26_0.SEQ_MODE=4'b1000;
    defparam shift_srl_175_0_LC_18_26_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_175_0_LC_18_26_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76051),
            .lcout(shift_srl_175Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93268),
            .ce(N__74124),
            .sr(_gnd_net_));
    defparam shift_srl_175_1_LC_18_26_1.C_ON=1'b0;
    defparam shift_srl_175_1_LC_18_26_1.SEQ_MODE=4'b1000;
    defparam shift_srl_175_1_LC_18_26_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_175_1_LC_18_26_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70288),
            .lcout(shift_srl_175Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93268),
            .ce(N__74124),
            .sr(_gnd_net_));
    defparam shift_srl_175_2_LC_18_26_2.C_ON=1'b0;
    defparam shift_srl_175_2_LC_18_26_2.SEQ_MODE=4'b1000;
    defparam shift_srl_175_2_LC_18_26_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_175_2_LC_18_26_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70282),
            .lcout(shift_srl_175Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93268),
            .ce(N__74124),
            .sr(_gnd_net_));
    defparam shift_srl_175_3_LC_18_26_3.C_ON=1'b0;
    defparam shift_srl_175_3_LC_18_26_3.SEQ_MODE=4'b1000;
    defparam shift_srl_175_3_LC_18_26_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_175_3_LC_18_26_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70276),
            .lcout(shift_srl_175Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93268),
            .ce(N__74124),
            .sr(_gnd_net_));
    defparam shift_srl_175_4_LC_18_26_4.C_ON=1'b0;
    defparam shift_srl_175_4_LC_18_26_4.SEQ_MODE=4'b1000;
    defparam shift_srl_175_4_LC_18_26_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_175_4_LC_18_26_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70270),
            .lcout(shift_srl_175Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93268),
            .ce(N__74124),
            .sr(_gnd_net_));
    defparam shift_srl_175_5_LC_18_26_5.C_ON=1'b0;
    defparam shift_srl_175_5_LC_18_26_5.SEQ_MODE=4'b1000;
    defparam shift_srl_175_5_LC_18_26_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_175_5_LC_18_26_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70264),
            .lcout(shift_srl_175Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93268),
            .ce(N__74124),
            .sr(_gnd_net_));
    defparam shift_srl_175_6_LC_18_26_6.C_ON=1'b0;
    defparam shift_srl_175_6_LC_18_26_6.SEQ_MODE=4'b1000;
    defparam shift_srl_175_6_LC_18_26_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_175_6_LC_18_26_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70360),
            .lcout(shift_srl_175Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93268),
            .ce(N__74124),
            .sr(_gnd_net_));
    defparam shift_srl_175_7_LC_18_26_7.C_ON=1'b0;
    defparam shift_srl_175_7_LC_18_26_7.SEQ_MODE=4'b1000;
    defparam shift_srl_175_7_LC_18_26_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_175_7_LC_18_26_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70354),
            .lcout(shift_srl_175Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93268),
            .ce(N__74124),
            .sr(_gnd_net_));
    defparam shift_srl_198_10_LC_18_27_0.C_ON=1'b0;
    defparam shift_srl_198_10_LC_18_27_0.SEQ_MODE=4'b1000;
    defparam shift_srl_198_10_LC_18_27_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_198_10_LC_18_27_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70318),
            .lcout(shift_srl_198Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93286),
            .ce(N__72204),
            .sr(_gnd_net_));
    defparam shift_srl_198_11_LC_18_27_1.C_ON=1'b0;
    defparam shift_srl_198_11_LC_18_27_1.SEQ_MODE=4'b1000;
    defparam shift_srl_198_11_LC_18_27_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_198_11_LC_18_27_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70348),
            .lcout(shift_srl_198Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93286),
            .ce(N__72204),
            .sr(_gnd_net_));
    defparam shift_srl_198_12_LC_18_27_2.C_ON=1'b0;
    defparam shift_srl_198_12_LC_18_27_2.SEQ_MODE=4'b1000;
    defparam shift_srl_198_12_LC_18_27_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_198_12_LC_18_27_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70342),
            .lcout(shift_srl_198Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93286),
            .ce(N__72204),
            .sr(_gnd_net_));
    defparam shift_srl_198_13_LC_18_27_3.C_ON=1'b0;
    defparam shift_srl_198_13_LC_18_27_3.SEQ_MODE=4'b1000;
    defparam shift_srl_198_13_LC_18_27_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_198_13_LC_18_27_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70336),
            .lcout(shift_srl_198Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93286),
            .ce(N__72204),
            .sr(_gnd_net_));
    defparam shift_srl_198_14_LC_18_27_4.C_ON=1'b0;
    defparam shift_srl_198_14_LC_18_27_4.SEQ_MODE=4'b1000;
    defparam shift_srl_198_14_LC_18_27_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_198_14_LC_18_27_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70330),
            .lcout(shift_srl_198Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93286),
            .ce(N__72204),
            .sr(_gnd_net_));
    defparam shift_srl_198_15_LC_18_27_5.C_ON=1'b0;
    defparam shift_srl_198_15_LC_18_27_5.SEQ_MODE=4'b1000;
    defparam shift_srl_198_15_LC_18_27_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_198_15_LC_18_27_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70324),
            .lcout(shift_srl_198Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93286),
            .ce(N__72204),
            .sr(_gnd_net_));
    defparam shift_srl_198_9_LC_18_27_6.C_ON=1'b0;
    defparam shift_srl_198_9_LC_18_27_6.SEQ_MODE=4'b1000;
    defparam shift_srl_198_9_LC_18_27_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_198_9_LC_18_27_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70489),
            .lcout(shift_srl_198Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93286),
            .ce(N__72204),
            .sr(_gnd_net_));
    defparam shift_srl_198_8_LC_18_27_7.C_ON=1'b0;
    defparam shift_srl_198_8_LC_18_27_7.SEQ_MODE=4'b1000;
    defparam shift_srl_198_8_LC_18_27_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_198_8_LC_18_27_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70498),
            .lcout(shift_srl_198Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93286),
            .ce(N__72204),
            .sr(_gnd_net_));
    defparam shift_srl_197_RNIMMFGH1_15_LC_18_28_0.C_ON=1'b0;
    defparam shift_srl_197_RNIMMFGH1_15_LC_18_28_0.SEQ_MODE=4'b0000;
    defparam shift_srl_197_RNIMMFGH1_15_LC_18_28_0.LUT_INIT=16'b1100110000000000;
    LogicCell40 shift_srl_197_RNIMMFGH1_15_LC_18_28_0 (
            .in0(_gnd_net_),
            .in1(N__72235),
            .in2(_gnd_net_),
            .in3(N__91516),
            .lcout(rco_c_197),
            .ltout(rco_c_197_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_198_RNI336TH1_15_LC_18_28_1.C_ON=1'b0;
    defparam shift_srl_198_RNI336TH1_15_LC_18_28_1.SEQ_MODE=4'b0000;
    defparam shift_srl_198_RNI336TH1_15_LC_18_28_1.LUT_INIT=16'b1010000010100000;
    LogicCell40 shift_srl_198_RNI336TH1_15_LC_18_28_1 (
            .in0(N__70416),
            .in1(_gnd_net_),
            .in2(N__70462),
            .in3(_gnd_net_),
            .lcout(rco_c_198),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_198_0_LC_18_28_2.C_ON=1'b0;
    defparam shift_srl_198_0_LC_18_28_2.SEQ_MODE=4'b1000;
    defparam shift_srl_198_0_LC_18_28_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_198_0_LC_18_28_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70415),
            .lcout(shift_srl_198Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93301),
            .ce(N__72200),
            .sr(_gnd_net_));
    defparam shift_srl_198_1_LC_18_28_3.C_ON=1'b0;
    defparam shift_srl_198_1_LC_18_28_3.SEQ_MODE=4'b1000;
    defparam shift_srl_198_1_LC_18_28_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_198_1_LC_18_28_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70399),
            .lcout(shift_srl_198Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93301),
            .ce(N__72200),
            .sr(_gnd_net_));
    defparam shift_srl_198_2_LC_18_28_4.C_ON=1'b0;
    defparam shift_srl_198_2_LC_18_28_4.SEQ_MODE=4'b1000;
    defparam shift_srl_198_2_LC_18_28_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_198_2_LC_18_28_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70393),
            .lcout(shift_srl_198Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93301),
            .ce(N__72200),
            .sr(_gnd_net_));
    defparam shift_srl_198_3_LC_18_28_5.C_ON=1'b0;
    defparam shift_srl_198_3_LC_18_28_5.SEQ_MODE=4'b1000;
    defparam shift_srl_198_3_LC_18_28_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_198_3_LC_18_28_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70387),
            .lcout(shift_srl_198Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93301),
            .ce(N__72200),
            .sr(_gnd_net_));
    defparam shift_srl_198_4_LC_18_28_6.C_ON=1'b0;
    defparam shift_srl_198_4_LC_18_28_6.SEQ_MODE=4'b1000;
    defparam shift_srl_198_4_LC_18_28_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_198_4_LC_18_28_6 (
            .in0(N__70381),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_198Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93301),
            .ce(N__72200),
            .sr(_gnd_net_));
    defparam shift_srl_198_5_LC_18_28_7.C_ON=1'b0;
    defparam shift_srl_198_5_LC_18_28_7.SEQ_MODE=4'b1000;
    defparam shift_srl_198_5_LC_18_28_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_198_5_LC_18_28_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70375),
            .lcout(shift_srl_198Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93301),
            .ce(N__72200),
            .sr(_gnd_net_));
    defparam shift_srl_197_0_LC_18_29_0.C_ON=1'b0;
    defparam shift_srl_197_0_LC_18_29_0.SEQ_MODE=4'b1000;
    defparam shift_srl_197_0_LC_18_29_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_197_0_LC_18_29_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70629),
            .lcout(shift_srl_197Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93322),
            .ce(N__72405),
            .sr(_gnd_net_));
    defparam shift_srl_197_7_LC_18_29_1.C_ON=1'b0;
    defparam shift_srl_197_7_LC_18_29_1.SEQ_MODE=4'b1000;
    defparam shift_srl_197_7_LC_18_29_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_197_7_LC_18_29_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70522),
            .lcout(shift_srl_197Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93322),
            .ce(N__72405),
            .sr(_gnd_net_));
    defparam shift_srl_197_2_LC_18_29_2.C_ON=1'b0;
    defparam shift_srl_197_2_LC_18_29_2.SEQ_MODE=4'b1000;
    defparam shift_srl_197_2_LC_18_29_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_197_2_LC_18_29_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70510),
            .lcout(shift_srl_197Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93322),
            .ce(N__72405),
            .sr(_gnd_net_));
    defparam shift_srl_197_3_LC_18_29_3.C_ON=1'b0;
    defparam shift_srl_197_3_LC_18_29_3.SEQ_MODE=4'b1000;
    defparam shift_srl_197_3_LC_18_29_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_197_3_LC_18_29_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70546),
            .lcout(shift_srl_197Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93322),
            .ce(N__72405),
            .sr(_gnd_net_));
    defparam shift_srl_197_4_LC_18_29_4.C_ON=1'b0;
    defparam shift_srl_197_4_LC_18_29_4.SEQ_MODE=4'b1000;
    defparam shift_srl_197_4_LC_18_29_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_197_4_LC_18_29_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70540),
            .lcout(shift_srl_197Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93322),
            .ce(N__72405),
            .sr(_gnd_net_));
    defparam shift_srl_197_5_LC_18_29_5.C_ON=1'b0;
    defparam shift_srl_197_5_LC_18_29_5.SEQ_MODE=4'b1000;
    defparam shift_srl_197_5_LC_18_29_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_197_5_LC_18_29_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70534),
            .lcout(shift_srl_197Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93322),
            .ce(N__72405),
            .sr(_gnd_net_));
    defparam shift_srl_197_6_LC_18_29_6.C_ON=1'b0;
    defparam shift_srl_197_6_LC_18_29_6.SEQ_MODE=4'b1000;
    defparam shift_srl_197_6_LC_18_29_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_197_6_LC_18_29_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70528),
            .lcout(shift_srl_197Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93322),
            .ce(N__72405),
            .sr(_gnd_net_));
    defparam shift_srl_197_1_LC_18_29_7.C_ON=1'b0;
    defparam shift_srl_197_1_LC_18_29_7.SEQ_MODE=4'b1000;
    defparam shift_srl_197_1_LC_18_29_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_197_1_LC_18_29_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70516),
            .lcout(shift_srl_197Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93322),
            .ce(N__72405),
            .sr(_gnd_net_));
    defparam shift_srl_197_10_LC_18_30_0.C_ON=1'b0;
    defparam shift_srl_197_10_LC_18_30_0.SEQ_MODE=4'b1000;
    defparam shift_srl_197_10_LC_18_30_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_197_10_LC_18_30_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70615),
            .lcout(shift_srl_197Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93344),
            .ce(N__72409),
            .sr(_gnd_net_));
    defparam shift_srl_197_11_LC_18_30_1.C_ON=1'b0;
    defparam shift_srl_197_11_LC_18_30_1.SEQ_MODE=4'b1000;
    defparam shift_srl_197_11_LC_18_30_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_197_11_LC_18_30_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70504),
            .lcout(shift_srl_197Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93344),
            .ce(N__72409),
            .sr(_gnd_net_));
    defparam shift_srl_197_12_LC_18_30_2.C_ON=1'b0;
    defparam shift_srl_197_12_LC_18_30_2.SEQ_MODE=4'b1000;
    defparam shift_srl_197_12_LC_18_30_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_197_12_LC_18_30_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70660),
            .lcout(shift_srl_197Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93344),
            .ce(N__72409),
            .sr(_gnd_net_));
    defparam shift_srl_197_13_LC_18_30_3.C_ON=1'b0;
    defparam shift_srl_197_13_LC_18_30_3.SEQ_MODE=4'b1000;
    defparam shift_srl_197_13_LC_18_30_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_197_13_LC_18_30_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70654),
            .lcout(shift_srl_197Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93344),
            .ce(N__72409),
            .sr(_gnd_net_));
    defparam shift_srl_197_14_LC_18_30_4.C_ON=1'b0;
    defparam shift_srl_197_14_LC_18_30_4.SEQ_MODE=4'b1000;
    defparam shift_srl_197_14_LC_18_30_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_197_14_LC_18_30_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70648),
            .lcout(shift_srl_197Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93344),
            .ce(N__72409),
            .sr(_gnd_net_));
    defparam shift_srl_197_15_LC_18_30_5.C_ON=1'b0;
    defparam shift_srl_197_15_LC_18_30_5.SEQ_MODE=4'b1000;
    defparam shift_srl_197_15_LC_18_30_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_197_15_LC_18_30_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70642),
            .lcout(shift_srl_197Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93344),
            .ce(N__72409),
            .sr(_gnd_net_));
    defparam shift_srl_197_9_LC_18_30_6.C_ON=1'b0;
    defparam shift_srl_197_9_LC_18_30_6.SEQ_MODE=4'b1000;
    defparam shift_srl_197_9_LC_18_30_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_197_9_LC_18_30_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70603),
            .lcout(shift_srl_197Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93344),
            .ce(N__72409),
            .sr(_gnd_net_));
    defparam shift_srl_197_8_LC_18_30_7.C_ON=1'b0;
    defparam shift_srl_197_8_LC_18_30_7.SEQ_MODE=4'b1000;
    defparam shift_srl_197_8_LC_18_30_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_197_8_LC_18_30_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70609),
            .lcout(shift_srl_197Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93344),
            .ce(N__72409),
            .sr(_gnd_net_));
    defparam shift_srl_93_8_LC_19_2_2.C_ON=1'b0;
    defparam shift_srl_93_8_LC_19_2_2.SEQ_MODE=4'b1000;
    defparam shift_srl_93_8_LC_19_2_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_93_8_LC_19_2_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70582),
            .lcout(shift_srl_93Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93395),
            .ce(N__70575),
            .sr(_gnd_net_));
    defparam shift_srl_93_7_LC_19_2_4.C_ON=1'b0;
    defparam shift_srl_93_7_LC_19_2_4.SEQ_MODE=4'b1000;
    defparam shift_srl_93_7_LC_19_2_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_93_7_LC_19_2_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70588),
            .lcout(shift_srl_93Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93395),
            .ce(N__70575),
            .sr(_gnd_net_));
    defparam shift_srl_92_1_LC_19_3_0.C_ON=1'b0;
    defparam shift_srl_92_1_LC_19_3_0.SEQ_MODE=4'b1000;
    defparam shift_srl_92_1_LC_19_3_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_92_1_LC_19_3_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70819),
            .lcout(shift_srl_92Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93382),
            .ce(N__70762),
            .sr(_gnd_net_));
    defparam shift_srl_92_2_LC_19_3_1.C_ON=1'b0;
    defparam shift_srl_92_2_LC_19_3_1.SEQ_MODE=4'b1000;
    defparam shift_srl_92_2_LC_19_3_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_92_2_LC_19_3_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70813),
            .lcout(shift_srl_92Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93382),
            .ce(N__70762),
            .sr(_gnd_net_));
    defparam shift_srl_92_3_LC_19_3_2.C_ON=1'b0;
    defparam shift_srl_92_3_LC_19_3_2.SEQ_MODE=4'b1000;
    defparam shift_srl_92_3_LC_19_3_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_92_3_LC_19_3_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70807),
            .lcout(shift_srl_92Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93382),
            .ce(N__70762),
            .sr(_gnd_net_));
    defparam shift_srl_92_4_LC_19_3_3.C_ON=1'b0;
    defparam shift_srl_92_4_LC_19_3_3.SEQ_MODE=4'b1000;
    defparam shift_srl_92_4_LC_19_3_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_92_4_LC_19_3_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70801),
            .lcout(shift_srl_92Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93382),
            .ce(N__70762),
            .sr(_gnd_net_));
    defparam shift_srl_92_5_LC_19_3_4.C_ON=1'b0;
    defparam shift_srl_92_5_LC_19_3_4.SEQ_MODE=4'b1000;
    defparam shift_srl_92_5_LC_19_3_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_92_5_LC_19_3_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70795),
            .lcout(shift_srl_92Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93382),
            .ce(N__70762),
            .sr(_gnd_net_));
    defparam shift_srl_92_6_LC_19_3_5.C_ON=1'b0;
    defparam shift_srl_92_6_LC_19_3_5.SEQ_MODE=4'b1000;
    defparam shift_srl_92_6_LC_19_3_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_92_6_LC_19_3_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70789),
            .lcout(shift_srl_92Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93382),
            .ce(N__70762),
            .sr(_gnd_net_));
    defparam shift_srl_92_7_LC_19_3_6.C_ON=1'b0;
    defparam shift_srl_92_7_LC_19_3_6.SEQ_MODE=4'b1000;
    defparam shift_srl_92_7_LC_19_3_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_92_7_LC_19_3_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70783),
            .lcout(shift_srl_92Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93382),
            .ce(N__70762),
            .sr(_gnd_net_));
    defparam shift_srl_92_8_LC_19_3_7.C_ON=1'b0;
    defparam shift_srl_92_8_LC_19_3_7.SEQ_MODE=4'b1000;
    defparam shift_srl_92_8_LC_19_3_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_92_8_LC_19_3_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70777),
            .lcout(shift_srl_92Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93382),
            .ce(N__70762),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_146_LC_19_4_5.C_ON=1'b0;
    defparam rco_obuf_RNO_146_LC_19_4_5.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_146_LC_19_4_5.LUT_INIT=16'b1100110000000000;
    LogicCell40 rco_obuf_RNO_146_LC_19_4_5 (
            .in0(_gnd_net_),
            .in1(N__70729),
            .in2(_gnd_net_),
            .in3(N__82220),
            .lcout(rco_c_146),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_46_7_LC_19_5_0.C_ON=1'b0;
    defparam shift_srl_46_7_LC_19_5_0.SEQ_MODE=4'b1000;
    defparam shift_srl_46_7_LC_19_5_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_46_7_LC_19_5_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70891),
            .lcout(shift_srl_46Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93347),
            .ce(N__70873),
            .sr(_gnd_net_));
    defparam shift_srl_46_11_LC_19_5_1.C_ON=1'b0;
    defparam shift_srl_46_11_LC_19_5_1.SEQ_MODE=4'b1000;
    defparam shift_srl_46_11_LC_19_5_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_46_11_LC_19_5_1 (
            .in0(N__70921),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_46Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93347),
            .ce(N__70873),
            .sr(_gnd_net_));
    defparam shift_srl_46_12_LC_19_5_2.C_ON=1'b0;
    defparam shift_srl_46_12_LC_19_5_2.SEQ_MODE=4'b1000;
    defparam shift_srl_46_12_LC_19_5_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_46_12_LC_19_5_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70915),
            .lcout(shift_srl_46Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93347),
            .ce(N__70873),
            .sr(_gnd_net_));
    defparam shift_srl_46_13_LC_19_5_3.C_ON=1'b0;
    defparam shift_srl_46_13_LC_19_5_3.SEQ_MODE=4'b1000;
    defparam shift_srl_46_13_LC_19_5_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_46_13_LC_19_5_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70909),
            .lcout(shift_srl_46Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93347),
            .ce(N__70873),
            .sr(_gnd_net_));
    defparam shift_srl_46_14_LC_19_5_4.C_ON=1'b0;
    defparam shift_srl_46_14_LC_19_5_4.SEQ_MODE=4'b1000;
    defparam shift_srl_46_14_LC_19_5_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_46_14_LC_19_5_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70903),
            .lcout(shift_srl_46Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93347),
            .ce(N__70873),
            .sr(_gnd_net_));
    defparam shift_srl_46_15_LC_19_5_5.C_ON=1'b0;
    defparam shift_srl_46_15_LC_19_5_5.SEQ_MODE=4'b1000;
    defparam shift_srl_46_15_LC_19_5_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_46_15_LC_19_5_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70897),
            .lcout(shift_srl_46Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93347),
            .ce(N__70873),
            .sr(_gnd_net_));
    defparam shift_srl_46_6_LC_19_5_6.C_ON=1'b0;
    defparam shift_srl_46_6_LC_19_5_6.SEQ_MODE=4'b1000;
    defparam shift_srl_46_6_LC_19_5_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_46_6_LC_19_5_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70879),
            .lcout(shift_srl_46Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93347),
            .ce(N__70873),
            .sr(_gnd_net_));
    defparam shift_srl_46_5_LC_19_5_7.C_ON=1'b0;
    defparam shift_srl_46_5_LC_19_5_7.SEQ_MODE=4'b1000;
    defparam shift_srl_46_5_LC_19_5_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_46_5_LC_19_5_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70885),
            .lcout(shift_srl_46Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93347),
            .ce(N__70873),
            .sr(_gnd_net_));
    defparam shift_srl_97_0_LC_19_6_0.C_ON=1'b0;
    defparam shift_srl_97_0_LC_19_6_0.SEQ_MODE=4'b1000;
    defparam shift_srl_97_0_LC_19_6_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_97_0_LC_19_6_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70843),
            .lcout(shift_srl_97Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93325),
            .ce(N__70945),
            .sr(_gnd_net_));
    defparam shift_srl_97_1_LC_19_6_1.C_ON=1'b0;
    defparam shift_srl_97_1_LC_19_6_1.SEQ_MODE=4'b1000;
    defparam shift_srl_97_1_LC_19_6_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_97_1_LC_19_6_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70993),
            .lcout(shift_srl_97Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93325),
            .ce(N__70945),
            .sr(_gnd_net_));
    defparam shift_srl_97_2_LC_19_6_2.C_ON=1'b0;
    defparam shift_srl_97_2_LC_19_6_2.SEQ_MODE=4'b1000;
    defparam shift_srl_97_2_LC_19_6_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_97_2_LC_19_6_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70987),
            .lcout(shift_srl_97Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93325),
            .ce(N__70945),
            .sr(_gnd_net_));
    defparam shift_srl_97_3_LC_19_6_3.C_ON=1'b0;
    defparam shift_srl_97_3_LC_19_6_3.SEQ_MODE=4'b1000;
    defparam shift_srl_97_3_LC_19_6_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_97_3_LC_19_6_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70981),
            .lcout(shift_srl_97Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93325),
            .ce(N__70945),
            .sr(_gnd_net_));
    defparam shift_srl_97_4_LC_19_6_4.C_ON=1'b0;
    defparam shift_srl_97_4_LC_19_6_4.SEQ_MODE=4'b1000;
    defparam shift_srl_97_4_LC_19_6_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_97_4_LC_19_6_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70975),
            .lcout(shift_srl_97Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93325),
            .ce(N__70945),
            .sr(_gnd_net_));
    defparam shift_srl_97_5_LC_19_6_5.C_ON=1'b0;
    defparam shift_srl_97_5_LC_19_6_5.SEQ_MODE=4'b1000;
    defparam shift_srl_97_5_LC_19_6_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_97_5_LC_19_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70969),
            .lcout(shift_srl_97Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93325),
            .ce(N__70945),
            .sr(_gnd_net_));
    defparam shift_srl_97_6_LC_19_6_6.C_ON=1'b0;
    defparam shift_srl_97_6_LC_19_6_6.SEQ_MODE=4'b1000;
    defparam shift_srl_97_6_LC_19_6_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_97_6_LC_19_6_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70963),
            .lcout(shift_srl_97Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93325),
            .ce(N__70945),
            .sr(_gnd_net_));
    defparam shift_srl_97_7_LC_19_6_7.C_ON=1'b0;
    defparam shift_srl_97_7_LC_19_6_7.SEQ_MODE=4'b1000;
    defparam shift_srl_97_7_LC_19_6_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_97_7_LC_19_6_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70957),
            .lcout(shift_srl_97Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93325),
            .ce(N__70945),
            .sr(_gnd_net_));
    defparam shift_srl_51_10_LC_19_7_0.C_ON=1'b0;
    defparam shift_srl_51_10_LC_19_7_0.SEQ_MODE=4'b1000;
    defparam shift_srl_51_10_LC_19_7_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_51_10_LC_19_7_0 (
            .in0(N__73015),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_51Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93304),
            .ce(N__72982),
            .sr(_gnd_net_));
    defparam shift_srl_51_11_LC_19_7_1.C_ON=1'b0;
    defparam shift_srl_51_11_LC_19_7_1.SEQ_MODE=4'b1000;
    defparam shift_srl_51_11_LC_19_7_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_51_11_LC_19_7_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70933),
            .lcout(shift_srl_51Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93304),
            .ce(N__72982),
            .sr(_gnd_net_));
    defparam shift_srl_51_12_LC_19_7_2.C_ON=1'b0;
    defparam shift_srl_51_12_LC_19_7_2.SEQ_MODE=4'b1000;
    defparam shift_srl_51_12_LC_19_7_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_51_12_LC_19_7_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71041),
            .lcout(shift_srl_51Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93304),
            .ce(N__72982),
            .sr(_gnd_net_));
    defparam shift_srl_51_13_LC_19_7_3.C_ON=1'b0;
    defparam shift_srl_51_13_LC_19_7_3.SEQ_MODE=4'b1000;
    defparam shift_srl_51_13_LC_19_7_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_51_13_LC_19_7_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71035),
            .lcout(shift_srl_51Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93304),
            .ce(N__72982),
            .sr(_gnd_net_));
    defparam shift_srl_51_14_LC_19_7_4.C_ON=1'b0;
    defparam shift_srl_51_14_LC_19_7_4.SEQ_MODE=4'b1000;
    defparam shift_srl_51_14_LC_19_7_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_51_14_LC_19_7_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71029),
            .lcout(shift_srl_51Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93304),
            .ce(N__72982),
            .sr(_gnd_net_));
    defparam shift_srl_51_15_LC_19_7_5.C_ON=1'b0;
    defparam shift_srl_51_15_LC_19_7_5.SEQ_MODE=4'b1000;
    defparam shift_srl_51_15_LC_19_7_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_51_15_LC_19_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71023),
            .lcout(shift_srl_51Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93304),
            .ce(N__72982),
            .sr(_gnd_net_));
    defparam shift_srl_51_7_LC_19_7_6.C_ON=1'b0;
    defparam shift_srl_51_7_LC_19_7_6.SEQ_MODE=4'b1000;
    defparam shift_srl_51_7_LC_19_7_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_51_7_LC_19_7_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71017),
            .lcout(shift_srl_51Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93304),
            .ce(N__72982),
            .sr(_gnd_net_));
    defparam shift_srl_51_6_LC_19_7_7.C_ON=1'b0;
    defparam shift_srl_51_6_LC_19_7_7.SEQ_MODE=4'b1000;
    defparam shift_srl_51_6_LC_19_7_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_51_6_LC_19_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72895),
            .lcout(shift_srl_51Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93304),
            .ce(N__72982),
            .sr(_gnd_net_));
    defparam shift_srl_53_0_LC_19_8_0.C_ON=1'b0;
    defparam shift_srl_53_0_LC_19_8_0.SEQ_MODE=4'b1000;
    defparam shift_srl_53_0_LC_19_8_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_53_0_LC_19_8_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73042),
            .lcout(shift_srl_53Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93288),
            .ce(N__73008),
            .sr(_gnd_net_));
    defparam shift_srl_53_1_LC_19_8_1.C_ON=1'b0;
    defparam shift_srl_53_1_LC_19_8_1.SEQ_MODE=4'b1000;
    defparam shift_srl_53_1_LC_19_8_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_53_1_LC_19_8_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71011),
            .lcout(shift_srl_53Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93288),
            .ce(N__73008),
            .sr(_gnd_net_));
    defparam shift_srl_53_2_LC_19_8_2.C_ON=1'b0;
    defparam shift_srl_53_2_LC_19_8_2.SEQ_MODE=4'b1000;
    defparam shift_srl_53_2_LC_19_8_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_53_2_LC_19_8_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71005),
            .lcout(shift_srl_53Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93288),
            .ce(N__73008),
            .sr(_gnd_net_));
    defparam shift_srl_53_3_LC_19_8_3.C_ON=1'b0;
    defparam shift_srl_53_3_LC_19_8_3.SEQ_MODE=4'b1000;
    defparam shift_srl_53_3_LC_19_8_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_53_3_LC_19_8_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70999),
            .lcout(shift_srl_53Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93288),
            .ce(N__73008),
            .sr(_gnd_net_));
    defparam shift_srl_53_4_LC_19_8_4.C_ON=1'b0;
    defparam shift_srl_53_4_LC_19_8_4.SEQ_MODE=4'b1000;
    defparam shift_srl_53_4_LC_19_8_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_53_4_LC_19_8_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71089),
            .lcout(shift_srl_53Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93288),
            .ce(N__73008),
            .sr(_gnd_net_));
    defparam shift_srl_53_5_LC_19_8_5.C_ON=1'b0;
    defparam shift_srl_53_5_LC_19_8_5.SEQ_MODE=4'b1000;
    defparam shift_srl_53_5_LC_19_8_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_53_5_LC_19_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71083),
            .lcout(shift_srl_53Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93288),
            .ce(N__73008),
            .sr(_gnd_net_));
    defparam shift_srl_53_6_LC_19_8_6.C_ON=1'b0;
    defparam shift_srl_53_6_LC_19_8_6.SEQ_MODE=4'b1000;
    defparam shift_srl_53_6_LC_19_8_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_53_6_LC_19_8_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71077),
            .lcout(shift_srl_53Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93288),
            .ce(N__73008),
            .sr(_gnd_net_));
    defparam shift_srl_53_7_LC_19_8_7.C_ON=1'b0;
    defparam shift_srl_53_7_LC_19_8_7.SEQ_MODE=4'b1000;
    defparam shift_srl_53_7_LC_19_8_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_53_7_LC_19_8_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71071),
            .lcout(shift_srl_53Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93288),
            .ce(N__73008),
            .sr(_gnd_net_));
    defparam shift_srl_53_10_LC_19_9_0.C_ON=1'b0;
    defparam shift_srl_53_10_LC_19_9_0.SEQ_MODE=4'b1000;
    defparam shift_srl_53_10_LC_19_9_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_53_10_LC_19_9_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71137),
            .lcout(shift_srl_53Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93271),
            .ce(N__73009),
            .sr(_gnd_net_));
    defparam shift_srl_53_11_LC_19_9_1.C_ON=1'b0;
    defparam shift_srl_53_11_LC_19_9_1.SEQ_MODE=4'b1000;
    defparam shift_srl_53_11_LC_19_9_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_53_11_LC_19_9_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71065),
            .lcout(shift_srl_53Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93271),
            .ce(N__73009),
            .sr(_gnd_net_));
    defparam shift_srl_53_12_LC_19_9_2.C_ON=1'b0;
    defparam shift_srl_53_12_LC_19_9_2.SEQ_MODE=4'b1000;
    defparam shift_srl_53_12_LC_19_9_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_53_12_LC_19_9_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71059),
            .lcout(shift_srl_53Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93271),
            .ce(N__73009),
            .sr(_gnd_net_));
    defparam shift_srl_53_13_LC_19_9_3.C_ON=1'b0;
    defparam shift_srl_53_13_LC_19_9_3.SEQ_MODE=4'b1000;
    defparam shift_srl_53_13_LC_19_9_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_53_13_LC_19_9_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71053),
            .lcout(shift_srl_53Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93271),
            .ce(N__73009),
            .sr(_gnd_net_));
    defparam shift_srl_53_14_LC_19_9_4.C_ON=1'b0;
    defparam shift_srl_53_14_LC_19_9_4.SEQ_MODE=4'b1000;
    defparam shift_srl_53_14_LC_19_9_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_53_14_LC_19_9_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71047),
            .lcout(shift_srl_53Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93271),
            .ce(N__73009),
            .sr(_gnd_net_));
    defparam shift_srl_53_15_LC_19_9_5.C_ON=1'b0;
    defparam shift_srl_53_15_LC_19_9_5.SEQ_MODE=4'b1000;
    defparam shift_srl_53_15_LC_19_9_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_53_15_LC_19_9_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71143),
            .lcout(shift_srl_53Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93271),
            .ce(N__73009),
            .sr(_gnd_net_));
    defparam shift_srl_53_9_LC_19_9_6.C_ON=1'b0;
    defparam shift_srl_53_9_LC_19_9_6.SEQ_MODE=4'b1000;
    defparam shift_srl_53_9_LC_19_9_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_53_9_LC_19_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71125),
            .lcout(shift_srl_53Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93271),
            .ce(N__73009),
            .sr(_gnd_net_));
    defparam shift_srl_53_8_LC_19_9_7.C_ON=1'b0;
    defparam shift_srl_53_8_LC_19_9_7.SEQ_MODE=4'b1000;
    defparam shift_srl_53_8_LC_19_9_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_53_8_LC_19_9_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71131),
            .lcout(shift_srl_53Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93271),
            .ce(N__73009),
            .sr(_gnd_net_));
    defparam shift_srl_41_10_LC_19_10_0.C_ON=1'b0;
    defparam shift_srl_41_10_LC_19_10_0.SEQ_MODE=4'b1000;
    defparam shift_srl_41_10_LC_19_10_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_41_10_LC_19_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71191),
            .lcout(shift_srl_41Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93251),
            .ce(N__78687),
            .sr(_gnd_net_));
    defparam shift_srl_41_11_LC_19_10_1.C_ON=1'b0;
    defparam shift_srl_41_11_LC_19_10_1.SEQ_MODE=4'b1000;
    defparam shift_srl_41_11_LC_19_10_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_41_11_LC_19_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71119),
            .lcout(shift_srl_41Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93251),
            .ce(N__78687),
            .sr(_gnd_net_));
    defparam shift_srl_41_12_LC_19_10_2.C_ON=1'b0;
    defparam shift_srl_41_12_LC_19_10_2.SEQ_MODE=4'b1000;
    defparam shift_srl_41_12_LC_19_10_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_41_12_LC_19_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71113),
            .lcout(shift_srl_41Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93251),
            .ce(N__78687),
            .sr(_gnd_net_));
    defparam shift_srl_41_13_LC_19_10_3.C_ON=1'b0;
    defparam shift_srl_41_13_LC_19_10_3.SEQ_MODE=4'b1000;
    defparam shift_srl_41_13_LC_19_10_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_41_13_LC_19_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71107),
            .lcout(shift_srl_41Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93251),
            .ce(N__78687),
            .sr(_gnd_net_));
    defparam shift_srl_41_14_LC_19_10_4.C_ON=1'b0;
    defparam shift_srl_41_14_LC_19_10_4.SEQ_MODE=4'b1000;
    defparam shift_srl_41_14_LC_19_10_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_41_14_LC_19_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71101),
            .lcout(shift_srl_41Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93251),
            .ce(N__78687),
            .sr(_gnd_net_));
    defparam shift_srl_41_15_LC_19_10_5.C_ON=1'b0;
    defparam shift_srl_41_15_LC_19_10_5.SEQ_MODE=4'b1000;
    defparam shift_srl_41_15_LC_19_10_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_41_15_LC_19_10_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71095),
            .lcout(shift_srl_41Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93251),
            .ce(N__78687),
            .sr(_gnd_net_));
    defparam shift_srl_41_9_LC_19_10_6.C_ON=1'b0;
    defparam shift_srl_41_9_LC_19_10_6.SEQ_MODE=4'b1000;
    defparam shift_srl_41_9_LC_19_10_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_41_9_LC_19_10_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71185),
            .lcout(shift_srl_41Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93251),
            .ce(N__78687),
            .sr(_gnd_net_));
    defparam shift_srl_41_8_LC_19_10_7.C_ON=1'b0;
    defparam shift_srl_41_8_LC_19_10_7.SEQ_MODE=4'b1000;
    defparam shift_srl_41_8_LC_19_10_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_41_8_LC_19_10_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78703),
            .lcout(shift_srl_41Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93251),
            .ce(N__78687),
            .sr(_gnd_net_));
    defparam shift_srl_59_0_LC_19_11_0.C_ON=1'b0;
    defparam shift_srl_59_0_LC_19_11_0.SEQ_MODE=4'b1000;
    defparam shift_srl_59_0_LC_19_11_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_59_0_LC_19_11_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81586),
            .lcout(shift_srl_59Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93230),
            .ce(N__73089),
            .sr(_gnd_net_));
    defparam shift_srl_59_1_LC_19_11_1.C_ON=1'b0;
    defparam shift_srl_59_1_LC_19_11_1.SEQ_MODE=4'b1000;
    defparam shift_srl_59_1_LC_19_11_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_59_1_LC_19_11_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71179),
            .lcout(shift_srl_59Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93230),
            .ce(N__73089),
            .sr(_gnd_net_));
    defparam shift_srl_59_2_LC_19_11_2.C_ON=1'b0;
    defparam shift_srl_59_2_LC_19_11_2.SEQ_MODE=4'b1000;
    defparam shift_srl_59_2_LC_19_11_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_59_2_LC_19_11_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71173),
            .lcout(shift_srl_59Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93230),
            .ce(N__73089),
            .sr(_gnd_net_));
    defparam shift_srl_59_3_LC_19_11_3.C_ON=1'b0;
    defparam shift_srl_59_3_LC_19_11_3.SEQ_MODE=4'b1000;
    defparam shift_srl_59_3_LC_19_11_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_59_3_LC_19_11_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71167),
            .lcout(shift_srl_59Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93230),
            .ce(N__73089),
            .sr(_gnd_net_));
    defparam shift_srl_59_4_LC_19_11_4.C_ON=1'b0;
    defparam shift_srl_59_4_LC_19_11_4.SEQ_MODE=4'b1000;
    defparam shift_srl_59_4_LC_19_11_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_59_4_LC_19_11_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71161),
            .lcout(shift_srl_59Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93230),
            .ce(N__73089),
            .sr(_gnd_net_));
    defparam shift_srl_59_5_LC_19_11_5.C_ON=1'b0;
    defparam shift_srl_59_5_LC_19_11_5.SEQ_MODE=4'b1000;
    defparam shift_srl_59_5_LC_19_11_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_59_5_LC_19_11_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71155),
            .lcout(shift_srl_59Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93230),
            .ce(N__73089),
            .sr(_gnd_net_));
    defparam shift_srl_59_6_LC_19_11_6.C_ON=1'b0;
    defparam shift_srl_59_6_LC_19_11_6.SEQ_MODE=4'b1000;
    defparam shift_srl_59_6_LC_19_11_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_59_6_LC_19_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71149),
            .lcout(shift_srl_59Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93230),
            .ce(N__73089),
            .sr(_gnd_net_));
    defparam shift_srl_59_7_LC_19_11_7.C_ON=1'b0;
    defparam shift_srl_59_7_LC_19_11_7.SEQ_MODE=4'b1000;
    defparam shift_srl_59_7_LC_19_11_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_59_7_LC_19_11_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71275),
            .lcout(shift_srl_59Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93230),
            .ce(N__73089),
            .sr(_gnd_net_));
    defparam shift_srl_44_10_LC_19_12_0.C_ON=1'b0;
    defparam shift_srl_44_10_LC_19_12_0.SEQ_MODE=4'b1000;
    defparam shift_srl_44_10_LC_19_12_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_44_10_LC_19_12_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71230),
            .lcout(shift_srl_44Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93211),
            .ce(N__71212),
            .sr(_gnd_net_));
    defparam shift_srl_44_11_LC_19_12_1.C_ON=1'b0;
    defparam shift_srl_44_11_LC_19_12_1.SEQ_MODE=4'b1000;
    defparam shift_srl_44_11_LC_19_12_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_44_11_LC_19_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71260),
            .lcout(shift_srl_44Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93211),
            .ce(N__71212),
            .sr(_gnd_net_));
    defparam shift_srl_44_12_LC_19_12_2.C_ON=1'b0;
    defparam shift_srl_44_12_LC_19_12_2.SEQ_MODE=4'b1000;
    defparam shift_srl_44_12_LC_19_12_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_44_12_LC_19_12_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71254),
            .lcout(shift_srl_44Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93211),
            .ce(N__71212),
            .sr(_gnd_net_));
    defparam shift_srl_44_13_LC_19_12_3.C_ON=1'b0;
    defparam shift_srl_44_13_LC_19_12_3.SEQ_MODE=4'b1000;
    defparam shift_srl_44_13_LC_19_12_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_44_13_LC_19_12_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71248),
            .lcout(shift_srl_44Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93211),
            .ce(N__71212),
            .sr(_gnd_net_));
    defparam shift_srl_44_14_LC_19_12_4.C_ON=1'b0;
    defparam shift_srl_44_14_LC_19_12_4.SEQ_MODE=4'b1000;
    defparam shift_srl_44_14_LC_19_12_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_44_14_LC_19_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71242),
            .lcout(shift_srl_44Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93211),
            .ce(N__71212),
            .sr(_gnd_net_));
    defparam shift_srl_44_15_LC_19_12_5.C_ON=1'b0;
    defparam shift_srl_44_15_LC_19_12_5.SEQ_MODE=4'b1000;
    defparam shift_srl_44_15_LC_19_12_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_44_15_LC_19_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71236),
            .lcout(shift_srl_44Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93211),
            .ce(N__71212),
            .sr(_gnd_net_));
    defparam shift_srl_44_9_LC_19_12_6.C_ON=1'b0;
    defparam shift_srl_44_9_LC_19_12_6.SEQ_MODE=4'b1000;
    defparam shift_srl_44_9_LC_19_12_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_44_9_LC_19_12_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71218),
            .lcout(shift_srl_44Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93211),
            .ce(N__71212),
            .sr(_gnd_net_));
    defparam shift_srl_44_8_LC_19_12_7.C_ON=1'b0;
    defparam shift_srl_44_8_LC_19_12_7.SEQ_MODE=4'b1000;
    defparam shift_srl_44_8_LC_19_12_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_44_8_LC_19_12_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71224),
            .lcout(shift_srl_44Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93211),
            .ce(N__71212),
            .sr(_gnd_net_));
    defparam shift_srl_48_11_LC_19_13_1.C_ON=1'b0;
    defparam shift_srl_48_11_LC_19_13_1.SEQ_MODE=4'b1000;
    defparam shift_srl_48_11_LC_19_13_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_48_11_LC_19_13_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71335),
            .lcout(shift_srl_48Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93191),
            .ce(N__73381),
            .sr(_gnd_net_));
    defparam shift_srl_48_9_LC_19_13_2.C_ON=1'b0;
    defparam shift_srl_48_9_LC_19_13_2.SEQ_MODE=4'b1000;
    defparam shift_srl_48_9_LC_19_13_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_48_9_LC_19_13_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71323),
            .lcout(shift_srl_48Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93191),
            .ce(N__73381),
            .sr(_gnd_net_));
    defparam shift_srl_48_8_LC_19_13_3.C_ON=1'b0;
    defparam shift_srl_48_8_LC_19_13_3.SEQ_MODE=4'b1000;
    defparam shift_srl_48_8_LC_19_13_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_48_8_LC_19_13_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71311),
            .lcout(shift_srl_48Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93191),
            .ce(N__73381),
            .sr(_gnd_net_));
    defparam shift_srl_48_7_LC_19_13_5.C_ON=1'b0;
    defparam shift_srl_48_7_LC_19_13_5.SEQ_MODE=4'b1000;
    defparam shift_srl_48_7_LC_19_13_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_48_7_LC_19_13_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71317),
            .lcout(shift_srl_48Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93191),
            .ce(N__73381),
            .sr(_gnd_net_));
    defparam shift_srl_39_RNIG4I71_15_LC_19_14_0.C_ON=1'b0;
    defparam shift_srl_39_RNIG4I71_15_LC_19_14_0.SEQ_MODE=4'b0000;
    defparam shift_srl_39_RNIG4I71_15_LC_19_14_0.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_39_RNIG4I71_15_LC_19_14_0 (
            .in0(N__79754),
            .in1(N__71499),
            .in2(N__81797),
            .in3(N__83791),
            .lcout(shift_srl_39_RNIG4I71Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_39_15_LC_19_14_1.C_ON=1'b0;
    defparam shift_srl_39_15_LC_19_14_1.SEQ_MODE=4'b1000;
    defparam shift_srl_39_15_LC_19_14_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_39_15_LC_19_14_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71299),
            .lcout(shift_srl_39Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93170),
            .ce(N__82030),
            .sr(_gnd_net_));
    defparam shift_srl_39_14_LC_19_14_2.C_ON=1'b0;
    defparam shift_srl_39_14_LC_19_14_2.SEQ_MODE=4'b1000;
    defparam shift_srl_39_14_LC_19_14_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_39_14_LC_19_14_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71293),
            .lcout(shift_srl_39Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93170),
            .ce(N__82030),
            .sr(_gnd_net_));
    defparam shift_srl_39_13_LC_19_14_3.C_ON=1'b0;
    defparam shift_srl_39_13_LC_19_14_3.SEQ_MODE=4'b1000;
    defparam shift_srl_39_13_LC_19_14_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_39_13_LC_19_14_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71287),
            .lcout(shift_srl_39Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93170),
            .ce(N__82030),
            .sr(_gnd_net_));
    defparam shift_srl_39_12_LC_19_14_4.C_ON=1'b0;
    defparam shift_srl_39_12_LC_19_14_4.SEQ_MODE=4'b1000;
    defparam shift_srl_39_12_LC_19_14_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_39_12_LC_19_14_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71281),
            .lcout(shift_srl_39Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93170),
            .ce(N__82030),
            .sr(_gnd_net_));
    defparam shift_srl_39_11_LC_19_14_5.C_ON=1'b0;
    defparam shift_srl_39_11_LC_19_14_5.SEQ_MODE=4'b1000;
    defparam shift_srl_39_11_LC_19_14_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_39_11_LC_19_14_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71377),
            .lcout(shift_srl_39Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93170),
            .ce(N__82030),
            .sr(_gnd_net_));
    defparam shift_srl_39_10_LC_19_14_6.C_ON=1'b0;
    defparam shift_srl_39_10_LC_19_14_6.SEQ_MODE=4'b1000;
    defparam shift_srl_39_10_LC_19_14_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_39_10_LC_19_14_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71371),
            .lcout(shift_srl_39Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93170),
            .ce(N__82030),
            .sr(_gnd_net_));
    defparam shift_srl_39_9_LC_19_14_7.C_ON=1'b0;
    defparam shift_srl_39_9_LC_19_14_7.SEQ_MODE=4'b1000;
    defparam shift_srl_39_9_LC_19_14_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_39_9_LC_19_14_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82045),
            .lcout(shift_srl_39Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93170),
            .ce(N__82030),
            .sr(_gnd_net_));
    defparam shift_srl_61_6_LC_19_15_0.C_ON=1'b0;
    defparam shift_srl_61_6_LC_19_15_0.SEQ_MODE=4'b1000;
    defparam shift_srl_61_6_LC_19_15_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_61_6_LC_19_15_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71341),
            .lcout(shift_srl_61Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93152),
            .ce(N__73417),
            .sr(_gnd_net_));
    defparam shift_srl_61_1_LC_19_15_1.C_ON=1'b0;
    defparam shift_srl_61_1_LC_19_15_1.SEQ_MODE=4'b1000;
    defparam shift_srl_61_1_LC_19_15_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_61_1_LC_19_15_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73321),
            .lcout(shift_srl_61Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93152),
            .ce(N__73417),
            .sr(_gnd_net_));
    defparam shift_srl_61_2_LC_19_15_2.C_ON=1'b0;
    defparam shift_srl_61_2_LC_19_15_2.SEQ_MODE=4'b1000;
    defparam shift_srl_61_2_LC_19_15_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_61_2_LC_19_15_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71365),
            .lcout(shift_srl_61Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93152),
            .ce(N__73417),
            .sr(_gnd_net_));
    defparam shift_srl_61_3_LC_19_15_3.C_ON=1'b0;
    defparam shift_srl_61_3_LC_19_15_3.SEQ_MODE=4'b1000;
    defparam shift_srl_61_3_LC_19_15_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_61_3_LC_19_15_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71359),
            .lcout(shift_srl_61Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93152),
            .ce(N__73417),
            .sr(_gnd_net_));
    defparam shift_srl_61_4_LC_19_15_4.C_ON=1'b0;
    defparam shift_srl_61_4_LC_19_15_4.SEQ_MODE=4'b1000;
    defparam shift_srl_61_4_LC_19_15_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_61_4_LC_19_15_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71353),
            .lcout(shift_srl_61Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93152),
            .ce(N__73417),
            .sr(_gnd_net_));
    defparam shift_srl_61_5_LC_19_15_5.C_ON=1'b0;
    defparam shift_srl_61_5_LC_19_15_5.SEQ_MODE=4'b1000;
    defparam shift_srl_61_5_LC_19_15_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_61_5_LC_19_15_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71347),
            .lcout(shift_srl_61Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93152),
            .ce(N__73417),
            .sr(_gnd_net_));
    defparam shift_srl_61_8_LC_19_15_6.C_ON=1'b0;
    defparam shift_srl_61_8_LC_19_15_6.SEQ_MODE=4'b1000;
    defparam shift_srl_61_8_LC_19_15_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_61_8_LC_19_15_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71575),
            .lcout(shift_srl_61Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93152),
            .ce(N__73417),
            .sr(_gnd_net_));
    defparam shift_srl_61_7_LC_19_15_7.C_ON=1'b0;
    defparam shift_srl_61_7_LC_19_15_7.SEQ_MODE=4'b1000;
    defparam shift_srl_61_7_LC_19_15_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_61_7_LC_19_15_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71581),
            .lcout(shift_srl_61Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93152),
            .ce(N__73417),
            .sr(_gnd_net_));
    defparam shift_srl_35_RNI6USP_15_LC_19_16_0.C_ON=1'b0;
    defparam shift_srl_35_RNI6USP_15_LC_19_16_0.SEQ_MODE=4'b0000;
    defparam shift_srl_35_RNI6USP_15_LC_19_16_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_35_RNI6USP_15_LC_19_16_0 (
            .in0(N__83348),
            .in1(N__85574),
            .in2(N__81910),
            .in3(N__87325),
            .lcout(rco_int_0_a2_0_a2_s_0_0_35),
            .ltout(rco_int_0_a2_0_a2_s_0_0_35_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_37_RNI1K6G3_15_LC_19_16_1.C_ON=1'b0;
    defparam shift_srl_37_RNI1K6G3_15_LC_19_16_1.SEQ_MODE=4'b0000;
    defparam shift_srl_37_RNI1K6G3_15_LC_19_16_1.LUT_INIT=16'b0000000000010000;
    LogicCell40 shift_srl_37_RNI1K6G3_15_LC_19_16_1 (
            .in0(N__71560),
            .in1(N__71566),
            .in2(N__71569),
            .in3(N__71395),
            .lcout(rco_int_0_a2_0_a2_0_0_37),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_31_RNI84161_0_15_LC_19_16_2.C_ON=1'b0;
    defparam shift_srl_31_RNI84161_0_15_LC_19_16_2.SEQ_MODE=4'b0000;
    defparam shift_srl_31_RNI84161_0_15_LC_19_16_2.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_31_RNI84161_0_15_LC_19_16_2 (
            .in0(N__83719),
            .in1(N__83884),
            .in2(N__83662),
            .in3(N__83840),
            .lcout(shift_srl_31_RNI84161_0Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_37_RNI973E_15_LC_19_16_3.C_ON=1'b0;
    defparam shift_srl_37_RNI973E_15_LC_19_16_3.SEQ_MODE=4'b0000;
    defparam shift_srl_37_RNI973E_15_LC_19_16_3.LUT_INIT=16'b0101010111111111;
    LogicCell40 shift_srl_37_RNI973E_15_LC_19_16_3 (
            .in0(N__83445),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83468),
            .lcout(shift_srl_37_RNI973EZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_36_15_LC_19_16_4.C_ON=1'b0;
    defparam shift_srl_36_15_LC_19_16_4.SEQ_MODE=4'b1000;
    defparam shift_srl_36_15_LC_19_16_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_36_15_LC_19_16_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__90964),
            .lcout(shift_srl_36Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93133),
            .ce(N__90942),
            .sr(_gnd_net_));
    defparam shift_srl_37_RNIG4IN_15_LC_19_16_5.C_ON=1'b0;
    defparam shift_srl_37_RNIG4IN_15_LC_19_16_5.SEQ_MODE=4'b0000;
    defparam shift_srl_37_RNIG4IN_15_LC_19_16_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_37_RNIG4IN_15_LC_19_16_5 (
            .in0(N__83469),
            .in1(N__71422),
            .in2(N__83446),
            .in3(N__71544),
            .lcout(rco_int_0_a2_0_a2_99_m6_0_a2_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_27_RNIAA521_0_15_LC_19_16_6.C_ON=1'b0;
    defparam shift_srl_27_RNIAA521_0_15_LC_19_16_6.SEQ_MODE=4'b0000;
    defparam shift_srl_27_RNIAA521_0_15_LC_19_16_6.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_27_RNIAA521_0_15_LC_19_16_6 (
            .in0(N__71545),
            .in1(N__71503),
            .in2(N__71430),
            .in3(N__83792),
            .lcout(shift_srl_27_RNIAA521_0Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_31_RNI84161_15_LC_19_16_7.C_ON=1'b0;
    defparam shift_srl_31_RNI84161_15_LC_19_16_7.SEQ_MODE=4'b0000;
    defparam shift_srl_31_RNI84161_15_LC_19_16_7.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_31_RNI84161_15_LC_19_16_7 (
            .in0(N__83841),
            .in1(N__83661),
            .in2(N__83892),
            .in3(N__83720),
            .lcout(rco_int_0_a2_0_a2_99_m6_0_a2_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_62_0_LC_19_17_0.C_ON=1'b0;
    defparam shift_srl_62_0_LC_19_17_0.SEQ_MODE=4'b1000;
    defparam shift_srl_62_0_LC_19_17_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_62_0_LC_19_17_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73516),
            .lcout(shift_srl_62Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93099),
            .ce(N__73486),
            .sr(_gnd_net_));
    defparam shift_srl_62_1_LC_19_17_1.C_ON=1'b0;
    defparam shift_srl_62_1_LC_19_17_1.SEQ_MODE=4'b1000;
    defparam shift_srl_62_1_LC_19_17_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_62_1_LC_19_17_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71623),
            .lcout(shift_srl_62Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93099),
            .ce(N__73486),
            .sr(_gnd_net_));
    defparam shift_srl_62_2_LC_19_17_2.C_ON=1'b0;
    defparam shift_srl_62_2_LC_19_17_2.SEQ_MODE=4'b1000;
    defparam shift_srl_62_2_LC_19_17_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_62_2_LC_19_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71617),
            .lcout(shift_srl_62Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93099),
            .ce(N__73486),
            .sr(_gnd_net_));
    defparam shift_srl_62_3_LC_19_17_3.C_ON=1'b0;
    defparam shift_srl_62_3_LC_19_17_3.SEQ_MODE=4'b1000;
    defparam shift_srl_62_3_LC_19_17_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_62_3_LC_19_17_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71611),
            .lcout(shift_srl_62Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93099),
            .ce(N__73486),
            .sr(_gnd_net_));
    defparam shift_srl_62_4_LC_19_17_4.C_ON=1'b0;
    defparam shift_srl_62_4_LC_19_17_4.SEQ_MODE=4'b1000;
    defparam shift_srl_62_4_LC_19_17_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_62_4_LC_19_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71605),
            .lcout(shift_srl_62Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93099),
            .ce(N__73486),
            .sr(_gnd_net_));
    defparam shift_srl_62_5_LC_19_17_5.C_ON=1'b0;
    defparam shift_srl_62_5_LC_19_17_5.SEQ_MODE=4'b1000;
    defparam shift_srl_62_5_LC_19_17_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_62_5_LC_19_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71599),
            .lcout(shift_srl_62Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93099),
            .ce(N__73486),
            .sr(_gnd_net_));
    defparam shift_srl_62_6_LC_19_17_6.C_ON=1'b0;
    defparam shift_srl_62_6_LC_19_17_6.SEQ_MODE=4'b1000;
    defparam shift_srl_62_6_LC_19_17_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_62_6_LC_19_17_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71593),
            .lcout(shift_srl_62Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93099),
            .ce(N__73486),
            .sr(_gnd_net_));
    defparam shift_srl_62_7_LC_19_17_7.C_ON=1'b0;
    defparam shift_srl_62_7_LC_19_17_7.SEQ_MODE=4'b1000;
    defparam shift_srl_62_7_LC_19_17_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_62_7_LC_19_17_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71587),
            .lcout(shift_srl_62Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93099),
            .ce(N__73486),
            .sr(_gnd_net_));
    defparam shift_srl_174_0_LC_19_18_0.C_ON=1'b0;
    defparam shift_srl_174_0_LC_19_18_0.SEQ_MODE=4'b1000;
    defparam shift_srl_174_0_LC_19_18_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_174_0_LC_19_18_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75990),
            .lcout(shift_srl_174Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93134),
            .ce(N__73563),
            .sr(_gnd_net_));
    defparam shift_srl_174_1_LC_19_18_1.C_ON=1'b0;
    defparam shift_srl_174_1_LC_19_18_1.SEQ_MODE=4'b1000;
    defparam shift_srl_174_1_LC_19_18_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_174_1_LC_19_18_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71725),
            .lcout(shift_srl_174Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93134),
            .ce(N__73563),
            .sr(_gnd_net_));
    defparam shift_srl_174_2_LC_19_18_2.C_ON=1'b0;
    defparam shift_srl_174_2_LC_19_18_2.SEQ_MODE=4'b1000;
    defparam shift_srl_174_2_LC_19_18_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_174_2_LC_19_18_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71719),
            .lcout(shift_srl_174Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93134),
            .ce(N__73563),
            .sr(_gnd_net_));
    defparam shift_srl_174_3_LC_19_18_3.C_ON=1'b0;
    defparam shift_srl_174_3_LC_19_18_3.SEQ_MODE=4'b1000;
    defparam shift_srl_174_3_LC_19_18_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_174_3_LC_19_18_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71713),
            .lcout(shift_srl_174Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93134),
            .ce(N__73563),
            .sr(_gnd_net_));
    defparam shift_srl_174_4_LC_19_18_4.C_ON=1'b0;
    defparam shift_srl_174_4_LC_19_18_4.SEQ_MODE=4'b1000;
    defparam shift_srl_174_4_LC_19_18_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_174_4_LC_19_18_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71707),
            .lcout(shift_srl_174Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93134),
            .ce(N__73563),
            .sr(_gnd_net_));
    defparam shift_srl_174_5_LC_19_18_5.C_ON=1'b0;
    defparam shift_srl_174_5_LC_19_18_5.SEQ_MODE=4'b1000;
    defparam shift_srl_174_5_LC_19_18_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_174_5_LC_19_18_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71701),
            .lcout(shift_srl_174Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93134),
            .ce(N__73563),
            .sr(_gnd_net_));
    defparam shift_srl_174_6_LC_19_18_6.C_ON=1'b0;
    defparam shift_srl_174_6_LC_19_18_6.SEQ_MODE=4'b1000;
    defparam shift_srl_174_6_LC_19_18_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_174_6_LC_19_18_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71695),
            .lcout(shift_srl_174Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93134),
            .ce(N__73563),
            .sr(_gnd_net_));
    defparam shift_srl_174_7_LC_19_18_7.C_ON=1'b0;
    defparam shift_srl_174_7_LC_19_18_7.SEQ_MODE=4'b1000;
    defparam shift_srl_174_7_LC_19_18_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_174_7_LC_19_18_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71689),
            .lcout(shift_srl_174Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93134),
            .ce(N__73563),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_166_LC_19_19_0.C_ON=1'b0;
    defparam rco_obuf_RNO_166_LC_19_19_0.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_166_LC_19_19_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 rco_obuf_RNO_166_LC_19_19_0 (
            .in0(N__83970),
            .in1(N__82415),
            .in2(N__87662),
            .in3(N__84011),
            .lcout(rco_c_166),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_159_RNIDDRE1_15_LC_19_19_1.C_ON=1'b0;
    defparam shift_srl_159_RNIDDRE1_15_LC_19_19_1.SEQ_MODE=4'b0000;
    defparam shift_srl_159_RNIDDRE1_15_LC_19_19_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_159_RNIDDRE1_15_LC_19_19_1 (
            .in0(N__77533),
            .in1(N__77280),
            .in2(N__77308),
            .in3(N__77898),
            .lcout(shift_srl_159_RNIDDRE1Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_165_RNI7STG91_15_LC_19_19_3.C_ON=1'b0;
    defparam shift_srl_165_RNI7STG91_15_LC_19_19_3.SEQ_MODE=4'b0000;
    defparam shift_srl_165_RNI7STG91_15_LC_19_19_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_165_RNI7STG91_15_LC_19_19_3 (
            .in0(N__90571),
            .in1(N__83969),
            .in2(N__82426),
            .in3(N__87635),
            .lcout(clk_en_166),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_173_RNIV9QIB1_15_LC_19_19_4.C_ON=1'b0;
    defparam shift_srl_173_RNIV9QIB1_15_LC_19_19_4.SEQ_MODE=4'b0000;
    defparam shift_srl_173_RNIV9QIB1_15_LC_19_19_4.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_173_RNIV9QIB1_15_LC_19_19_4 (
            .in0(N__87634),
            .in1(N__90569),
            .in2(N__84240),
            .in3(N__75969),
            .lcout(clk_en_174),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIE81AE1_15_LC_19_19_5.C_ON=1'b0;
    defparam shift_srl_0_RNIE81AE1_15_LC_19_19_5.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIE81AE1_15_LC_19_19_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNIE81AE1_15_LC_19_19_5 (
            .in0(N__86034),
            .in1(N__84230),
            .in2(N__90580),
            .in3(N__87633),
            .lcout(clk_en_184),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_162_RNIQ85P81_15_LC_19_19_6.C_ON=1'b0;
    defparam shift_srl_162_RNIQ85P81_15_LC_19_19_6.SEQ_MODE=4'b0000;
    defparam shift_srl_162_RNIQ85P81_15_LC_19_19_6.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_162_RNIQ85P81_15_LC_19_19_6 (
            .in0(N__82327),
            .in1(N__77764),
            .in2(N__88004),
            .in3(N__79390),
            .lcout(rco_c_162),
            .ltout(rco_c_162_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNI7LJSD1_15_LC_19_19_7.C_ON=1'b0;
    defparam shift_srl_0_RNI7LJSD1_15_LC_19_19_7.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNI7LJSD1_15_LC_19_19_7.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNI7LJSD1_15_LC_19_19_7 (
            .in0(N__90570),
            .in1(N__75837),
            .in2(N__71752),
            .in3(N__84234),
            .lcout(clk_en_183),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_184_0_LC_19_20_0.C_ON=1'b0;
    defparam shift_srl_184_0_LC_19_20_0.SEQ_MODE=4'b1000;
    defparam shift_srl_184_0_LC_19_20_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_184_0_LC_19_20_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__91689),
            .lcout(shift_srl_184Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93171),
            .ce(N__73935),
            .sr(_gnd_net_));
    defparam shift_srl_184_1_LC_19_20_1.C_ON=1'b0;
    defparam shift_srl_184_1_LC_19_20_1.SEQ_MODE=4'b1000;
    defparam shift_srl_184_1_LC_19_20_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_184_1_LC_19_20_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71749),
            .lcout(shift_srl_184Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93171),
            .ce(N__73935),
            .sr(_gnd_net_));
    defparam shift_srl_184_2_LC_19_20_2.C_ON=1'b0;
    defparam shift_srl_184_2_LC_19_20_2.SEQ_MODE=4'b1000;
    defparam shift_srl_184_2_LC_19_20_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_184_2_LC_19_20_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71743),
            .lcout(shift_srl_184Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93171),
            .ce(N__73935),
            .sr(_gnd_net_));
    defparam shift_srl_184_3_LC_19_20_3.C_ON=1'b0;
    defparam shift_srl_184_3_LC_19_20_3.SEQ_MODE=4'b1000;
    defparam shift_srl_184_3_LC_19_20_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_184_3_LC_19_20_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71737),
            .lcout(shift_srl_184Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93171),
            .ce(N__73935),
            .sr(_gnd_net_));
    defparam shift_srl_184_4_LC_19_20_4.C_ON=1'b0;
    defparam shift_srl_184_4_LC_19_20_4.SEQ_MODE=4'b1000;
    defparam shift_srl_184_4_LC_19_20_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_184_4_LC_19_20_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71731),
            .lcout(shift_srl_184Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93171),
            .ce(N__73935),
            .sr(_gnd_net_));
    defparam shift_srl_184_5_LC_19_20_5.C_ON=1'b0;
    defparam shift_srl_184_5_LC_19_20_5.SEQ_MODE=4'b1000;
    defparam shift_srl_184_5_LC_19_20_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_184_5_LC_19_20_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71806),
            .lcout(shift_srl_184Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93171),
            .ce(N__73935),
            .sr(_gnd_net_));
    defparam shift_srl_184_6_LC_19_20_6.C_ON=1'b0;
    defparam shift_srl_184_6_LC_19_20_6.SEQ_MODE=4'b1000;
    defparam shift_srl_184_6_LC_19_20_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_184_6_LC_19_20_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71800),
            .lcout(shift_srl_184Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93171),
            .ce(N__73935),
            .sr(_gnd_net_));
    defparam shift_srl_184_7_LC_19_20_7.C_ON=1'b0;
    defparam shift_srl_184_7_LC_19_20_7.SEQ_MODE=4'b1000;
    defparam shift_srl_184_7_LC_19_20_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_184_7_LC_19_20_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71794),
            .lcout(shift_srl_184Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93171),
            .ce(N__73935),
            .sr(_gnd_net_));
    defparam shift_srl_183_10_LC_19_21_0.C_ON=1'b0;
    defparam shift_srl_183_10_LC_19_21_0.SEQ_MODE=4'b1000;
    defparam shift_srl_183_10_LC_19_21_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_183_10_LC_19_21_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71758),
            .lcout(shift_srl_183Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93192),
            .ce(N__71864),
            .sr(_gnd_net_));
    defparam shift_srl_183_11_LC_19_21_1.C_ON=1'b0;
    defparam shift_srl_183_11_LC_19_21_1.SEQ_MODE=4'b1000;
    defparam shift_srl_183_11_LC_19_21_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_183_11_LC_19_21_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71788),
            .lcout(shift_srl_183Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93192),
            .ce(N__71864),
            .sr(_gnd_net_));
    defparam shift_srl_183_12_LC_19_21_2.C_ON=1'b0;
    defparam shift_srl_183_12_LC_19_21_2.SEQ_MODE=4'b1000;
    defparam shift_srl_183_12_LC_19_21_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_183_12_LC_19_21_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71782),
            .lcout(shift_srl_183Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93192),
            .ce(N__71864),
            .sr(_gnd_net_));
    defparam shift_srl_183_13_LC_19_21_3.C_ON=1'b0;
    defparam shift_srl_183_13_LC_19_21_3.SEQ_MODE=4'b1000;
    defparam shift_srl_183_13_LC_19_21_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_183_13_LC_19_21_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71776),
            .lcout(shift_srl_183Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93192),
            .ce(N__71864),
            .sr(_gnd_net_));
    defparam shift_srl_183_14_LC_19_21_4.C_ON=1'b0;
    defparam shift_srl_183_14_LC_19_21_4.SEQ_MODE=4'b1000;
    defparam shift_srl_183_14_LC_19_21_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_183_14_LC_19_21_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71770),
            .lcout(shift_srl_183Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93192),
            .ce(N__71864),
            .sr(_gnd_net_));
    defparam shift_srl_183_9_LC_19_21_5.C_ON=1'b0;
    defparam shift_srl_183_9_LC_19_21_5.SEQ_MODE=4'b1000;
    defparam shift_srl_183_9_LC_19_21_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_183_9_LC_19_21_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71917),
            .lcout(shift_srl_183Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93192),
            .ce(N__71864),
            .sr(_gnd_net_));
    defparam shift_srl_183_8_LC_19_21_6.C_ON=1'b0;
    defparam shift_srl_183_8_LC_19_21_6.SEQ_MODE=4'b1000;
    defparam shift_srl_183_8_LC_19_21_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_183_8_LC_19_21_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71911),
            .lcout(shift_srl_183Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93192),
            .ce(N__71864),
            .sr(_gnd_net_));
    defparam shift_srl_183_7_LC_19_21_7.C_ON=1'b0;
    defparam shift_srl_183_7_LC_19_21_7.SEQ_MODE=4'b1000;
    defparam shift_srl_183_7_LC_19_21_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_183_7_LC_19_21_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71875),
            .lcout(shift_srl_183Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93192),
            .ce(N__71864),
            .sr(_gnd_net_));
    defparam shift_srl_183_2_LC_19_22_0.C_ON=1'b0;
    defparam shift_srl_183_2_LC_19_22_0.SEQ_MODE=4'b1000;
    defparam shift_srl_183_2_LC_19_22_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_183_2_LC_19_22_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71905),
            .lcout(shift_srl_183Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93212),
            .ce(N__71865),
            .sr(_gnd_net_));
    defparam shift_srl_183_3_LC_19_22_1.C_ON=1'b0;
    defparam shift_srl_183_3_LC_19_22_1.SEQ_MODE=4'b1000;
    defparam shift_srl_183_3_LC_19_22_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_183_3_LC_19_22_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71899),
            .lcout(shift_srl_183Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93212),
            .ce(N__71865),
            .sr(_gnd_net_));
    defparam shift_srl_183_4_LC_19_22_2.C_ON=1'b0;
    defparam shift_srl_183_4_LC_19_22_2.SEQ_MODE=4'b1000;
    defparam shift_srl_183_4_LC_19_22_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_183_4_LC_19_22_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71893),
            .lcout(shift_srl_183Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93212),
            .ce(N__71865),
            .sr(_gnd_net_));
    defparam shift_srl_183_5_LC_19_22_3.C_ON=1'b0;
    defparam shift_srl_183_5_LC_19_22_3.SEQ_MODE=4'b1000;
    defparam shift_srl_183_5_LC_19_22_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_183_5_LC_19_22_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71887),
            .lcout(shift_srl_183Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93212),
            .ce(N__71865),
            .sr(_gnd_net_));
    defparam shift_srl_183_6_LC_19_22_4.C_ON=1'b0;
    defparam shift_srl_183_6_LC_19_22_4.SEQ_MODE=4'b1000;
    defparam shift_srl_183_6_LC_19_22_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_183_6_LC_19_22_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71881),
            .lcout(shift_srl_183Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93212),
            .ce(N__71865),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_181_LC_19_23_0.C_ON=1'b0;
    defparam rco_obuf_RNO_181_LC_19_23_0.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_181_LC_19_23_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 rco_obuf_RNO_181_LC_19_23_0 (
            .in0(N__75885),
            .in1(N__78162),
            .in2(N__85970),
            .in3(N__82753),
            .lcout(rco_c_181),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_180_LC_19_23_1.C_ON=1'b0;
    defparam rco_obuf_RNO_180_LC_19_23_1.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_180_LC_19_23_1.LUT_INIT=16'b1000100000000000;
    LogicCell40 rco_obuf_RNO_180_LC_19_23_1 (
            .in0(N__82752),
            .in1(N__78161),
            .in2(_gnd_net_),
            .in3(N__85948),
            .lcout(rco_c_180),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_181_RNITD9Q6_15_LC_19_23_2.C_ON=1'b0;
    defparam shift_srl_181_RNITD9Q6_15_LC_19_23_2.SEQ_MODE=4'b0000;
    defparam shift_srl_181_RNITD9Q6_15_LC_19_23_2.LUT_INIT=16'b1111111101111111;
    LogicCell40 shift_srl_181_RNITD9Q6_15_LC_19_23_2 (
            .in0(N__78160),
            .in1(N__82751),
            .in2(N__75886),
            .in3(N__84155),
            .lcout(),
            .ltout(clk_en_0_a3_0_a2_sx_182_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_181_RNI16CJD1_15_LC_19_23_3.C_ON=1'b0;
    defparam shift_srl_181_RNI16CJD1_15_LC_19_23_3.SEQ_MODE=4'b0000;
    defparam shift_srl_181_RNI16CJD1_15_LC_19_23_3.LUT_INIT=16'b0000010000000000;
    LogicCell40 shift_srl_181_RNI16CJD1_15_LC_19_23_3 (
            .in0(N__75177),
            .in1(N__77822),
            .in2(N__72115),
            .in3(N__75091),
            .lcout(clk_en_182),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_91_RNIQEMFF_15_LC_19_23_4.C_ON=1'b0;
    defparam shift_srl_91_RNIQEMFF_15_LC_19_23_4.SEQ_MODE=4'b0000;
    defparam shift_srl_91_RNIQEMFF_15_LC_19_23_4.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_91_RNIQEMFF_15_LC_19_23_4 (
            .in0(N__72112),
            .in1(N__85129),
            .in2(N__82341),
            .in3(N__72034),
            .lcout(rco_int_0_a2_0_a2_sx_153),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_145_RNIEG3VP_15_LC_19_23_5.C_ON=1'b0;
    defparam shift_srl_145_RNIEG3VP_15_LC_19_23_5.SEQ_MODE=4'b0000;
    defparam shift_srl_145_RNIEG3VP_15_LC_19_23_5.LUT_INIT=16'b1101111111111111;
    LogicCell40 shift_srl_145_RNIEG3VP_15_LC_19_23_5 (
            .in0(N__71976),
            .in1(N__71955),
            .in2(N__84235),
            .in3(N__75089),
            .lcout(),
            .ltout(rco_int_0_a3_0_a2_sx_183_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_183_RNIJS69E1_15_LC_19_23_6.C_ON=1'b0;
    defparam shift_srl_183_RNIJS69E1_15_LC_19_23_6.SEQ_MODE=4'b0000;
    defparam shift_srl_183_RNIJS69E1_15_LC_19_23_6.LUT_INIT=16'b0000000000001000;
    LogicCell40 shift_srl_183_RNIJS69E1_15_LC_19_23_6 (
            .in0(N__87992),
            .in1(N__86009),
            .in2(N__71932),
            .in3(N__75175),
            .lcout(rco_c_183),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIPRMFB1_15_LC_19_23_7.C_ON=1'b0;
    defparam shift_srl_0_RNIPRMFB1_15_LC_19_23_7.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIPRMFB1_15_LC_19_23_7.LUT_INIT=16'b0000010000000000;
    LogicCell40 shift_srl_0_RNIPRMFB1_15_LC_19_23_7 (
            .in0(N__75176),
            .in1(N__77821),
            .in2(N__84160),
            .in3(N__75090),
            .lcout(clk_en_173),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_195_10_LC_19_24_0.C_ON=1'b0;
    defparam shift_srl_195_10_LC_19_24_0.SEQ_MODE=4'b1000;
    defparam shift_srl_195_10_LC_19_24_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_195_10_LC_19_24_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72151),
            .lcout(shift_srl_195Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93252),
            .ce(N__73978),
            .sr(_gnd_net_));
    defparam shift_srl_195_11_LC_19_24_1.C_ON=1'b0;
    defparam shift_srl_195_11_LC_19_24_1.SEQ_MODE=4'b1000;
    defparam shift_srl_195_11_LC_19_24_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_195_11_LC_19_24_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71929),
            .lcout(shift_srl_195Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93252),
            .ce(N__73978),
            .sr(_gnd_net_));
    defparam shift_srl_195_12_LC_19_24_2.C_ON=1'b0;
    defparam shift_srl_195_12_LC_19_24_2.SEQ_MODE=4'b1000;
    defparam shift_srl_195_12_LC_19_24_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_195_12_LC_19_24_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71923),
            .lcout(shift_srl_195Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93252),
            .ce(N__73978),
            .sr(_gnd_net_));
    defparam shift_srl_195_13_LC_19_24_3.C_ON=1'b0;
    defparam shift_srl_195_13_LC_19_24_3.SEQ_MODE=4'b1000;
    defparam shift_srl_195_13_LC_19_24_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_195_13_LC_19_24_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72169),
            .lcout(shift_srl_195Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93252),
            .ce(N__73978),
            .sr(_gnd_net_));
    defparam shift_srl_195_14_LC_19_24_4.C_ON=1'b0;
    defparam shift_srl_195_14_LC_19_24_4.SEQ_MODE=4'b1000;
    defparam shift_srl_195_14_LC_19_24_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_195_14_LC_19_24_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72163),
            .lcout(shift_srl_195Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93252),
            .ce(N__73978),
            .sr(_gnd_net_));
    defparam shift_srl_195_15_LC_19_24_5.C_ON=1'b0;
    defparam shift_srl_195_15_LC_19_24_5.SEQ_MODE=4'b1000;
    defparam shift_srl_195_15_LC_19_24_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_195_15_LC_19_24_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72157),
            .lcout(shift_srl_195Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93252),
            .ce(N__73978),
            .sr(_gnd_net_));
    defparam shift_srl_195_9_LC_19_24_6.C_ON=1'b0;
    defparam shift_srl_195_9_LC_19_24_6.SEQ_MODE=4'b1000;
    defparam shift_srl_195_9_LC_19_24_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_195_9_LC_19_24_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72145),
            .lcout(shift_srl_195Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93252),
            .ce(N__73978),
            .sr(_gnd_net_));
    defparam shift_srl_195_8_LC_19_24_7.C_ON=1'b0;
    defparam shift_srl_195_8_LC_19_24_7.SEQ_MODE=4'b1000;
    defparam shift_srl_195_8_LC_19_24_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_195_8_LC_19_24_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73984),
            .lcout(shift_srl_195Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93252),
            .ce(N__73978),
            .sr(_gnd_net_));
    defparam shift_srl_185_0_LC_19_25_0.C_ON=1'b0;
    defparam shift_srl_185_0_LC_19_25_0.SEQ_MODE=4'b1000;
    defparam shift_srl_185_0_LC_19_25_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_185_0_LC_19_25_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__91736),
            .lcout(shift_srl_185Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93270),
            .ce(N__74055),
            .sr(_gnd_net_));
    defparam shift_srl_185_1_LC_19_25_1.C_ON=1'b0;
    defparam shift_srl_185_1_LC_19_25_1.SEQ_MODE=4'b1000;
    defparam shift_srl_185_1_LC_19_25_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_185_1_LC_19_25_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72139),
            .lcout(shift_srl_185Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93270),
            .ce(N__74055),
            .sr(_gnd_net_));
    defparam shift_srl_185_2_LC_19_25_2.C_ON=1'b0;
    defparam shift_srl_185_2_LC_19_25_2.SEQ_MODE=4'b1000;
    defparam shift_srl_185_2_LC_19_25_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_185_2_LC_19_25_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72133),
            .lcout(shift_srl_185Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93270),
            .ce(N__74055),
            .sr(_gnd_net_));
    defparam shift_srl_185_3_LC_19_25_3.C_ON=1'b0;
    defparam shift_srl_185_3_LC_19_25_3.SEQ_MODE=4'b1000;
    defparam shift_srl_185_3_LC_19_25_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_185_3_LC_19_25_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72127),
            .lcout(shift_srl_185Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93270),
            .ce(N__74055),
            .sr(_gnd_net_));
    defparam shift_srl_185_4_LC_19_25_4.C_ON=1'b0;
    defparam shift_srl_185_4_LC_19_25_4.SEQ_MODE=4'b1000;
    defparam shift_srl_185_4_LC_19_25_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_185_4_LC_19_25_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72121),
            .lcout(shift_srl_185Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93270),
            .ce(N__74055),
            .sr(_gnd_net_));
    defparam shift_srl_185_5_LC_19_25_5.C_ON=1'b0;
    defparam shift_srl_185_5_LC_19_25_5.SEQ_MODE=4'b1000;
    defparam shift_srl_185_5_LC_19_25_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_185_5_LC_19_25_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72283),
            .lcout(shift_srl_185Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93270),
            .ce(N__74055),
            .sr(_gnd_net_));
    defparam shift_srl_185_6_LC_19_25_6.C_ON=1'b0;
    defparam shift_srl_185_6_LC_19_25_6.SEQ_MODE=4'b1000;
    defparam shift_srl_185_6_LC_19_25_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_185_6_LC_19_25_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72277),
            .lcout(shift_srl_185Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93270),
            .ce(N__74055),
            .sr(_gnd_net_));
    defparam shift_srl_185_7_LC_19_25_7.C_ON=1'b0;
    defparam shift_srl_185_7_LC_19_25_7.SEQ_MODE=4'b1000;
    defparam shift_srl_185_7_LC_19_25_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_185_7_LC_19_25_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72271),
            .lcout(shift_srl_185Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93270),
            .ce(N__74055),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNI7PDOG1_15_LC_19_26_0.C_ON=1'b0;
    defparam shift_srl_0_RNI7PDOG1_15_LC_19_26_0.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNI7PDOG1_15_LC_19_26_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNI7PDOG1_15_LC_19_26_0 (
            .in0(N__90556),
            .in1(N__86036),
            .in2(N__85930),
            .in3(N__73857),
            .lcout(clk_en_194),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIH2AHH1_15_LC_19_26_1.C_ON=1'b0;
    defparam shift_srl_0_RNIH2AHH1_15_LC_19_26_1.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIH2AHH1_15_LC_19_26_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNIH2AHH1_15_LC_19_26_1 (
            .in0(N__86037),
            .in1(N__72234),
            .in2(N__90554),
            .in3(N__85899),
            .lcout(clk_en_198),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_184_RNIMVKBE1_15_LC_19_26_2.C_ON=1'b0;
    defparam shift_srl_184_RNIMVKBE1_15_LC_19_26_2.SEQ_MODE=4'b0000;
    defparam shift_srl_184_RNIMVKBE1_15_LC_19_26_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_184_RNIMVKBE1_15_LC_19_26_2 (
            .in0(N__90559),
            .in1(N__86035),
            .in2(N__85932),
            .in3(N__91690),
            .lcout(clk_en_185),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_172_RNIUFSEB1_15_LC_19_26_3.C_ON=1'b0;
    defparam shift_srl_172_RNIUFSEB1_15_LC_19_26_3.SEQ_MODE=4'b0000;
    defparam shift_srl_172_RNIUFSEB1_15_LC_19_26_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_172_RNIUFSEB1_15_LC_19_26_3 (
            .in0(N__84220),
            .in1(N__82342),
            .in2(N__88012),
            .in3(N__82202),
            .lcout(rco_c_172),
            .ltout(rco_c_172_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIKTK9F1_15_LC_19_26_4.C_ON=1'b0;
    defparam shift_srl_0_RNIKTK9F1_15_LC_19_26_4.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIKTK9F1_15_LC_19_26_4.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNIKTK9F1_15_LC_19_26_4 (
            .in0(N__80345),
            .in1(N__86038),
            .in2(N__72172),
            .in3(N__90494),
            .lcout(clk_en_188),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIOC4DG1_15_LC_19_26_5.C_ON=1'b0;
    defparam shift_srl_0_RNIOC4DG1_15_LC_19_26_5.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIOC4DG1_15_LC_19_26_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNIOC4DG1_15_LC_19_26_5 (
            .in0(N__86039),
            .in1(N__90557),
            .in2(N__74259),
            .in3(N__85895),
            .lcout(clk_en_192),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIQLF4H1_15_LC_19_26_6.C_ON=1'b0;
    defparam shift_srl_0_RNIQLF4H1_15_LC_19_26_6.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIQLF4H1_15_LC_19_26_6.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNIQLF4H1_15_LC_19_26_6 (
            .in0(N__90558),
            .in1(N__86040),
            .in2(N__85931),
            .in3(N__73822),
            .lcout(clk_en_196),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_174_RNI6S3QB1_15_LC_19_26_7.C_ON=1'b0;
    defparam shift_srl_174_RNI6S3QB1_15_LC_19_26_7.SEQ_MODE=4'b0000;
    defparam shift_srl_174_RNI6S3QB1_15_LC_19_26_7.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_174_RNI6S3QB1_15_LC_19_26_7 (
            .in0(N__76023),
            .in1(N__75952),
            .in2(N__90555),
            .in3(N__85900),
            .lcout(clk_en_175),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_196_0_LC_19_27_0.C_ON=1'b0;
    defparam shift_srl_196_0_LC_19_27_0.SEQ_MODE=4'b1000;
    defparam shift_srl_196_0_LC_19_27_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_196_0_LC_19_27_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72384),
            .lcout(shift_srl_196Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93303),
            .ce(N__72497),
            .sr(_gnd_net_));
    defparam shift_srl_196_1_LC_19_27_1.C_ON=1'b0;
    defparam shift_srl_196_1_LC_19_27_1.SEQ_MODE=4'b1000;
    defparam shift_srl_196_1_LC_19_27_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_196_1_LC_19_27_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72319),
            .lcout(shift_srl_196Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93303),
            .ce(N__72497),
            .sr(_gnd_net_));
    defparam shift_srl_196_2_LC_19_27_2.C_ON=1'b0;
    defparam shift_srl_196_2_LC_19_27_2.SEQ_MODE=4'b1000;
    defparam shift_srl_196_2_LC_19_27_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_196_2_LC_19_27_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72313),
            .lcout(shift_srl_196Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93303),
            .ce(N__72497),
            .sr(_gnd_net_));
    defparam shift_srl_196_3_LC_19_27_3.C_ON=1'b0;
    defparam shift_srl_196_3_LC_19_27_3.SEQ_MODE=4'b1000;
    defparam shift_srl_196_3_LC_19_27_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_196_3_LC_19_27_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72307),
            .lcout(shift_srl_196Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93303),
            .ce(N__72497),
            .sr(_gnd_net_));
    defparam shift_srl_196_4_LC_19_27_4.C_ON=1'b0;
    defparam shift_srl_196_4_LC_19_27_4.SEQ_MODE=4'b1000;
    defparam shift_srl_196_4_LC_19_27_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_196_4_LC_19_27_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72301),
            .lcout(shift_srl_196Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93303),
            .ce(N__72497),
            .sr(_gnd_net_));
    defparam shift_srl_196_5_LC_19_27_5.C_ON=1'b0;
    defparam shift_srl_196_5_LC_19_27_5.SEQ_MODE=4'b1000;
    defparam shift_srl_196_5_LC_19_27_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_196_5_LC_19_27_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72295),
            .lcout(shift_srl_196Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93303),
            .ce(N__72497),
            .sr(_gnd_net_));
    defparam shift_srl_196_6_LC_19_27_6.C_ON=1'b0;
    defparam shift_srl_196_6_LC_19_27_6.SEQ_MODE=4'b1000;
    defparam shift_srl_196_6_LC_19_27_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_196_6_LC_19_27_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72289),
            .lcout(shift_srl_196Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93303),
            .ce(N__72497),
            .sr(_gnd_net_));
    defparam shift_srl_196_7_LC_19_27_7.C_ON=1'b0;
    defparam shift_srl_196_7_LC_19_27_7.SEQ_MODE=4'b1000;
    defparam shift_srl_196_7_LC_19_27_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_196_7_LC_19_27_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72433),
            .lcout(shift_srl_196Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93303),
            .ce(N__72497),
            .sr(_gnd_net_));
    defparam shift_srl_196_8_LC_19_28_0.C_ON=1'b0;
    defparam shift_srl_196_8_LC_19_28_0.SEQ_MODE=4'b1000;
    defparam shift_srl_196_8_LC_19_28_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_196_8_LC_19_28_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72427),
            .lcout(shift_srl_196Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93324),
            .ce(N__72504),
            .sr(_gnd_net_));
    defparam shift_srl_196_9_LC_19_28_1.C_ON=1'b0;
    defparam shift_srl_196_9_LC_19_28_1.SEQ_MODE=4'b1000;
    defparam shift_srl_196_9_LC_19_28_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_196_9_LC_19_28_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72421),
            .lcout(shift_srl_196Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93324),
            .ce(N__72504),
            .sr(_gnd_net_));
    defparam shift_srl_196_10_LC_19_28_5.C_ON=1'b0;
    defparam shift_srl_196_10_LC_19_28_5.SEQ_MODE=4'b1000;
    defparam shift_srl_196_10_LC_19_28_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_196_10_LC_19_28_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72415),
            .lcout(shift_srl_196Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93324),
            .ce(N__72504),
            .sr(_gnd_net_));
    defparam shift_srl_196_RNI5QP8H1_15_LC_19_29_0.C_ON=1'b0;
    defparam shift_srl_196_RNI5QP8H1_15_LC_19_29_0.SEQ_MODE=4'b0000;
    defparam shift_srl_196_RNI5QP8H1_15_LC_19_29_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_196_RNI5QP8H1_15_LC_19_29_0 (
            .in0(N__90561),
            .in1(N__73832),
            .in2(N__72383),
            .in3(N__91478),
            .lcout(clk_en_197),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_196_15_LC_19_29_1.C_ON=1'b0;
    defparam shift_srl_196_15_LC_19_29_1.SEQ_MODE=4'b1000;
    defparam shift_srl_196_15_LC_19_29_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_196_15_LC_19_29_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72337),
            .lcout(shift_srl_196Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93346),
            .ce(N__72505),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_196_LC_19_29_2.C_ON=1'b0;
    defparam rco_obuf_RNO_196_LC_19_29_2.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_196_LC_19_29_2.LUT_INIT=16'b1000100000000000;
    LogicCell40 rco_obuf_RNO_196_LC_19_29_2 (
            .in0(N__72376),
            .in1(N__73833),
            .in2(_gnd_net_),
            .in3(N__91479),
            .lcout(rco_c_196),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_196_14_LC_19_29_3.C_ON=1'b0;
    defparam shift_srl_196_14_LC_19_29_3.SEQ_MODE=4'b1000;
    defparam shift_srl_196_14_LC_19_29_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_196_14_LC_19_29_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72331),
            .lcout(shift_srl_196Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93346),
            .ce(N__72505),
            .sr(_gnd_net_));
    defparam shift_srl_196_13_LC_19_29_4.C_ON=1'b0;
    defparam shift_srl_196_13_LC_19_29_4.SEQ_MODE=4'b1000;
    defparam shift_srl_196_13_LC_19_29_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_196_13_LC_19_29_4 (
            .in0(N__72325),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_196Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93346),
            .ce(N__72505),
            .sr(_gnd_net_));
    defparam shift_srl_196_12_LC_19_29_5.C_ON=1'b0;
    defparam shift_srl_196_12_LC_19_29_5.SEQ_MODE=4'b1000;
    defparam shift_srl_196_12_LC_19_29_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_196_12_LC_19_29_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72511),
            .lcout(shift_srl_196Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93346),
            .ce(N__72505),
            .sr(_gnd_net_));
    defparam shift_srl_196_11_LC_19_29_6.C_ON=1'b0;
    defparam shift_srl_196_11_LC_19_29_6.SEQ_MODE=4'b1000;
    defparam shift_srl_196_11_LC_19_29_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_196_11_LC_19_29_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72517),
            .lcout(shift_srl_196Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93346),
            .ce(N__72505),
            .sr(_gnd_net_));
    defparam shift_srl_182_10_LC_19_30_0.C_ON=1'b0;
    defparam shift_srl_182_10_LC_19_30_0.SEQ_MODE=4'b1000;
    defparam shift_srl_182_10_LC_19_30_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_182_10_LC_19_30_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72445),
            .lcout(shift_srl_182Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93364),
            .ce(N__72549),
            .sr(_gnd_net_));
    defparam shift_srl_182_11_LC_19_30_1.C_ON=1'b0;
    defparam shift_srl_182_11_LC_19_30_1.SEQ_MODE=4'b1000;
    defparam shift_srl_182_11_LC_19_30_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_182_11_LC_19_30_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72475),
            .lcout(shift_srl_182Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93364),
            .ce(N__72549),
            .sr(_gnd_net_));
    defparam shift_srl_182_12_LC_19_30_2.C_ON=1'b0;
    defparam shift_srl_182_12_LC_19_30_2.SEQ_MODE=4'b1000;
    defparam shift_srl_182_12_LC_19_30_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_182_12_LC_19_30_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72469),
            .lcout(shift_srl_182Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93364),
            .ce(N__72549),
            .sr(_gnd_net_));
    defparam shift_srl_182_13_LC_19_30_3.C_ON=1'b0;
    defparam shift_srl_182_13_LC_19_30_3.SEQ_MODE=4'b1000;
    defparam shift_srl_182_13_LC_19_30_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_182_13_LC_19_30_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72463),
            .lcout(shift_srl_182Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93364),
            .ce(N__72549),
            .sr(_gnd_net_));
    defparam shift_srl_182_14_LC_19_30_4.C_ON=1'b0;
    defparam shift_srl_182_14_LC_19_30_4.SEQ_MODE=4'b1000;
    defparam shift_srl_182_14_LC_19_30_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_182_14_LC_19_30_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72457),
            .lcout(shift_srl_182Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93364),
            .ce(N__72549),
            .sr(_gnd_net_));
    defparam shift_srl_182_15_LC_19_30_5.C_ON=1'b0;
    defparam shift_srl_182_15_LC_19_30_5.SEQ_MODE=4'b1000;
    defparam shift_srl_182_15_LC_19_30_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_182_15_LC_19_30_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72451),
            .lcout(shift_srl_182Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93364),
            .ce(N__72549),
            .sr(_gnd_net_));
    defparam shift_srl_182_9_LC_19_30_6.C_ON=1'b0;
    defparam shift_srl_182_9_LC_19_30_6.SEQ_MODE=4'b1000;
    defparam shift_srl_182_9_LC_19_30_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_182_9_LC_19_30_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72439),
            .lcout(shift_srl_182Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93364),
            .ce(N__72549),
            .sr(_gnd_net_));
    defparam shift_srl_182_8_LC_19_30_7.C_ON=1'b0;
    defparam shift_srl_182_8_LC_19_30_7.SEQ_MODE=4'b1000;
    defparam shift_srl_182_8_LC_19_30_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_182_8_LC_19_30_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72559),
            .lcout(shift_srl_182Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93364),
            .ce(N__72549),
            .sr(_gnd_net_));
    defparam shift_srl_182_0_LC_19_31_0.C_ON=1'b0;
    defparam shift_srl_182_0_LC_19_31_0.SEQ_MODE=4'b1000;
    defparam shift_srl_182_0_LC_19_31_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_182_0_LC_19_31_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75900),
            .lcout(shift_srl_182Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93381),
            .ce(N__72553),
            .sr(_gnd_net_));
    defparam shift_srl_182_1_LC_19_31_1.C_ON=1'b0;
    defparam shift_srl_182_1_LC_19_31_1.SEQ_MODE=4'b1000;
    defparam shift_srl_182_1_LC_19_31_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_182_1_LC_19_31_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72601),
            .lcout(shift_srl_182Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93381),
            .ce(N__72553),
            .sr(_gnd_net_));
    defparam shift_srl_182_2_LC_19_31_2.C_ON=1'b0;
    defparam shift_srl_182_2_LC_19_31_2.SEQ_MODE=4'b1000;
    defparam shift_srl_182_2_LC_19_31_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_182_2_LC_19_31_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72595),
            .lcout(shift_srl_182Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93381),
            .ce(N__72553),
            .sr(_gnd_net_));
    defparam shift_srl_182_3_LC_19_31_3.C_ON=1'b0;
    defparam shift_srl_182_3_LC_19_31_3.SEQ_MODE=4'b1000;
    defparam shift_srl_182_3_LC_19_31_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_182_3_LC_19_31_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72589),
            .lcout(shift_srl_182Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93381),
            .ce(N__72553),
            .sr(_gnd_net_));
    defparam shift_srl_182_4_LC_19_31_4.C_ON=1'b0;
    defparam shift_srl_182_4_LC_19_31_4.SEQ_MODE=4'b1000;
    defparam shift_srl_182_4_LC_19_31_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_182_4_LC_19_31_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72583),
            .lcout(shift_srl_182Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93381),
            .ce(N__72553),
            .sr(_gnd_net_));
    defparam shift_srl_182_5_LC_19_31_5.C_ON=1'b0;
    defparam shift_srl_182_5_LC_19_31_5.SEQ_MODE=4'b1000;
    defparam shift_srl_182_5_LC_19_31_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_182_5_LC_19_31_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72577),
            .lcout(shift_srl_182Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93381),
            .ce(N__72553),
            .sr(_gnd_net_));
    defparam shift_srl_182_6_LC_19_31_6.C_ON=1'b0;
    defparam shift_srl_182_6_LC_19_31_6.SEQ_MODE=4'b1000;
    defparam shift_srl_182_6_LC_19_31_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_182_6_LC_19_31_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72571),
            .lcout(shift_srl_182Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93381),
            .ce(N__72553),
            .sr(_gnd_net_));
    defparam shift_srl_182_7_LC_19_31_7.C_ON=1'b0;
    defparam shift_srl_182_7_LC_19_31_7.SEQ_MODE=4'b1000;
    defparam shift_srl_182_7_LC_19_31_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_182_7_LC_19_31_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72565),
            .lcout(shift_srl_182Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93381),
            .ce(N__72553),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_94_LC_20_4_0.C_ON=1'b0;
    defparam rco_obuf_RNO_94_LC_20_4_0.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_94_LC_20_4_0.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_94_LC_20_4_0 (
            .in0(N__72724),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72787),
            .lcout(rco_c_94),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_95_LC_20_4_1.C_ON=1'b0;
    defparam rco_obuf_RNO_95_LC_20_4_1.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_95_LC_20_4_1.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_95_LC_20_4_1 (
            .in0(N__72788),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72882),
            .lcout(rco_c_95),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_98_LC_20_4_2.C_ON=1'b0;
    defparam rco_obuf_RNO_98_LC_20_4_2.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_98_LC_20_4_2.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_98_LC_20_4_2 (
            .in0(N__72823),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72789),
            .lcout(rco_c_98),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_94_0_LC_20_4_3.C_ON=1'b0;
    defparam shift_srl_94_0_LC_20_4_3.SEQ_MODE=4'b1000;
    defparam shift_srl_94_0_LC_20_4_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_94_0_LC_20_4_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72723),
            .lcout(shift_srl_94Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93383),
            .ce(N__72655),
            .sr(_gnd_net_));
    defparam shift_srl_94_1_LC_20_4_4.C_ON=1'b0;
    defparam shift_srl_94_1_LC_20_4_4.SEQ_MODE=4'b1000;
    defparam shift_srl_94_1_LC_20_4_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_94_1_LC_20_4_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72688),
            .lcout(shift_srl_94Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93383),
            .ce(N__72655),
            .sr(_gnd_net_));
    defparam shift_srl_94_2_LC_20_4_5.C_ON=1'b0;
    defparam shift_srl_94_2_LC_20_4_5.SEQ_MODE=4'b1000;
    defparam shift_srl_94_2_LC_20_4_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_94_2_LC_20_4_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72682),
            .lcout(shift_srl_94Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93383),
            .ce(N__72655),
            .sr(_gnd_net_));
    defparam shift_srl_94_3_LC_20_4_6.C_ON=1'b0;
    defparam shift_srl_94_3_LC_20_4_6.SEQ_MODE=4'b1000;
    defparam shift_srl_94_3_LC_20_4_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_94_3_LC_20_4_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72676),
            .lcout(shift_srl_94Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93383),
            .ce(N__72655),
            .sr(_gnd_net_));
    defparam shift_srl_94_4_LC_20_4_7.C_ON=1'b0;
    defparam shift_srl_94_4_LC_20_4_7.SEQ_MODE=4'b1000;
    defparam shift_srl_94_4_LC_20_4_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_94_4_LC_20_4_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72670),
            .lcout(shift_srl_94Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93383),
            .ce(N__72655),
            .sr(_gnd_net_));
    defparam shift_srl_49_10_LC_20_5_0.C_ON=1'b0;
    defparam shift_srl_49_10_LC_20_5_0.SEQ_MODE=4'b1000;
    defparam shift_srl_49_10_LC_20_5_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_49_10_LC_20_5_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72607),
            .lcout(shift_srl_49Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93365),
            .ce(N__74431),
            .sr(_gnd_net_));
    defparam shift_srl_49_9_LC_20_5_1.C_ON=1'b0;
    defparam shift_srl_49_9_LC_20_5_1.SEQ_MODE=4'b1000;
    defparam shift_srl_49_9_LC_20_5_1.LUT_INIT=16'b1100110011001100;
    LogicCell40 shift_srl_49_9_LC_20_5_1 (
            .in0(_gnd_net_),
            .in1(N__72937),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_49Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93365),
            .ce(N__74431),
            .sr(_gnd_net_));
    defparam shift_srl_49_8_LC_20_6_0.C_ON=1'b0;
    defparam shift_srl_49_8_LC_20_6_0.SEQ_MODE=4'b1000;
    defparam shift_srl_49_8_LC_20_6_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_49_8_LC_20_6_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72931),
            .lcout(shift_srl_49Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93349),
            .ce(N__74426),
            .sr(_gnd_net_));
    defparam shift_srl_49_7_LC_20_6_1.C_ON=1'b0;
    defparam shift_srl_49_7_LC_20_6_1.SEQ_MODE=4'b1000;
    defparam shift_srl_49_7_LC_20_6_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_49_7_LC_20_6_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74509),
            .lcout(shift_srl_49Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93349),
            .ce(N__74426),
            .sr(_gnd_net_));
    defparam shift_srl_51_0_LC_20_7_0.C_ON=1'b0;
    defparam shift_srl_51_0_LC_20_7_0.SEQ_MODE=4'b1000;
    defparam shift_srl_51_0_LC_20_7_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_51_0_LC_20_7_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74627),
            .lcout(shift_srl_51Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93327),
            .ce(N__72981),
            .sr(_gnd_net_));
    defparam shift_srl_51_1_LC_20_7_1.C_ON=1'b0;
    defparam shift_srl_51_1_LC_20_7_1.SEQ_MODE=4'b1000;
    defparam shift_srl_51_1_LC_20_7_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_51_1_LC_20_7_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72925),
            .lcout(shift_srl_51Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93327),
            .ce(N__72981),
            .sr(_gnd_net_));
    defparam shift_srl_51_2_LC_20_7_2.C_ON=1'b0;
    defparam shift_srl_51_2_LC_20_7_2.SEQ_MODE=4'b1000;
    defparam shift_srl_51_2_LC_20_7_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_51_2_LC_20_7_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72919),
            .lcout(shift_srl_51Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93327),
            .ce(N__72981),
            .sr(_gnd_net_));
    defparam shift_srl_51_3_LC_20_7_3.C_ON=1'b0;
    defparam shift_srl_51_3_LC_20_7_3.SEQ_MODE=4'b1000;
    defparam shift_srl_51_3_LC_20_7_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_51_3_LC_20_7_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72913),
            .lcout(shift_srl_51Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93327),
            .ce(N__72981),
            .sr(_gnd_net_));
    defparam shift_srl_51_4_LC_20_7_4.C_ON=1'b0;
    defparam shift_srl_51_4_LC_20_7_4.SEQ_MODE=4'b1000;
    defparam shift_srl_51_4_LC_20_7_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_51_4_LC_20_7_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72907),
            .lcout(shift_srl_51Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93327),
            .ce(N__72981),
            .sr(_gnd_net_));
    defparam shift_srl_51_5_LC_20_7_5.C_ON=1'b0;
    defparam shift_srl_51_5_LC_20_7_5.SEQ_MODE=4'b1000;
    defparam shift_srl_51_5_LC_20_7_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_51_5_LC_20_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72901),
            .lcout(shift_srl_51Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93327),
            .ce(N__72981),
            .sr(_gnd_net_));
    defparam shift_srl_51_8_LC_20_7_6.C_ON=1'b0;
    defparam shift_srl_51_8_LC_20_7_6.SEQ_MODE=4'b1000;
    defparam shift_srl_51_8_LC_20_7_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_51_8_LC_20_7_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72889),
            .lcout(shift_srl_51Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93327),
            .ce(N__72981),
            .sr(_gnd_net_));
    defparam shift_srl_51_9_LC_20_7_7.C_ON=1'b0;
    defparam shift_srl_51_9_LC_20_7_7.SEQ_MODE=4'b1000;
    defparam shift_srl_51_9_LC_20_7_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_51_9_LC_20_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73021),
            .lcout(shift_srl_51Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93327),
            .ce(N__72981),
            .sr(_gnd_net_));
    defparam shift_srl_52_RNICF6KD_15_LC_20_8_0.C_ON=1'b0;
    defparam shift_srl_52_RNICF6KD_15_LC_20_8_0.SEQ_MODE=4'b0000;
    defparam shift_srl_52_RNICF6KD_15_LC_20_8_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_52_RNICF6KD_15_LC_20_8_0 (
            .in0(N__76441),
            .in1(N__74399),
            .in2(N__88320),
            .in3(N__74626),
            .lcout(clk_en_53),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_49_15_LC_20_8_1.C_ON=1'b0;
    defparam shift_srl_49_15_LC_20_8_1.SEQ_MODE=4'b1000;
    defparam shift_srl_49_15_LC_20_8_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_49_15_LC_20_8_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72970),
            .lcout(shift_srl_49Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93306),
            .ce(N__74427),
            .sr(_gnd_net_));
    defparam shift_srl_50_RNI869C_15_LC_20_8_2.C_ON=1'b0;
    defparam shift_srl_50_RNI869C_15_LC_20_8_2.SEQ_MODE=4'b0000;
    defparam shift_srl_50_RNI869C_15_LC_20_8_2.LUT_INIT=16'b1100110000000000;
    LogicCell40 shift_srl_50_RNI869C_15_LC_20_8_2 (
            .in0(_gnd_net_),
            .in1(N__93478),
            .in2(_gnd_net_),
            .in3(N__76346),
            .lcout(shift_srl_50_RNI869CZ0Z_15),
            .ltout(shift_srl_50_RNI869CZ0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNI9SN6D_15_LC_20_8_3.C_ON=1'b0;
    defparam shift_srl_0_RNI9SN6D_15_LC_20_8_3.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNI9SN6D_15_LC_20_8_3.LUT_INIT=16'b1010000000000000;
    LogicCell40 shift_srl_0_RNI9SN6D_15_LC_20_8_3 (
            .in0(N__89972),
            .in1(_gnd_net_),
            .in2(N__72985),
            .in3(N__93587),
            .lcout(clk_en_51),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_49_14_LC_20_8_4.C_ON=1'b0;
    defparam shift_srl_49_14_LC_20_8_4.SEQ_MODE=4'b1000;
    defparam shift_srl_49_14_LC_20_8_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_49_14_LC_20_8_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72964),
            .lcout(shift_srl_49Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93306),
            .ce(N__74427),
            .sr(_gnd_net_));
    defparam shift_srl_49_13_LC_20_8_5.C_ON=1'b0;
    defparam shift_srl_49_13_LC_20_8_5.SEQ_MODE=4'b1000;
    defparam shift_srl_49_13_LC_20_8_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_49_13_LC_20_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72958),
            .lcout(shift_srl_49Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93306),
            .ce(N__74427),
            .sr(_gnd_net_));
    defparam shift_srl_49_12_LC_20_8_6.C_ON=1'b0;
    defparam shift_srl_49_12_LC_20_8_6.SEQ_MODE=4'b1000;
    defparam shift_srl_49_12_LC_20_8_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_49_12_LC_20_8_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72943),
            .lcout(shift_srl_49Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93306),
            .ce(N__74427),
            .sr(_gnd_net_));
    defparam shift_srl_49_11_LC_20_8_7.C_ON=1'b0;
    defparam shift_srl_49_11_LC_20_8_7.SEQ_MODE=4'b1000;
    defparam shift_srl_49_11_LC_20_8_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_49_11_LC_20_8_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72952),
            .lcout(shift_srl_49Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93306),
            .ce(N__74427),
            .sr(_gnd_net_));
    defparam shift_srl_40_RNI5HIIA_15_LC_20_9_0.C_ON=1'b0;
    defparam shift_srl_40_RNI5HIIA_15_LC_20_9_0.SEQ_MODE=4'b0000;
    defparam shift_srl_40_RNI5HIIA_15_LC_20_9_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_40_RNI5HIIA_15_LC_20_9_0 (
            .in0(N__74710),
            .in1(N__74740),
            .in2(N__90243),
            .in3(N__81332),
            .lcout(clk_en_41),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_39_RNIDNRE_15_LC_20_9_1.C_ON=1'b0;
    defparam shift_srl_39_RNIDNRE_15_LC_20_9_1.SEQ_MODE=4'b0000;
    defparam shift_srl_39_RNIDNRE_15_LC_20_9_1.LUT_INIT=16'b1100110000000000;
    LogicCell40 shift_srl_39_RNIDNRE_15_LC_20_9_1 (
            .in0(_gnd_net_),
            .in1(N__81804),
            .in2(_gnd_net_),
            .in3(N__79761),
            .lcout(rco_int_0_a2_0_a2_0_39),
            .ltout(rco_int_0_a2_0_a2_0_39_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_41_RNIBS3L1_15_LC_20_9_2.C_ON=1'b0;
    defparam shift_srl_41_RNIBS3L1_15_LC_20_9_2.SEQ_MODE=4'b0000;
    defparam shift_srl_41_RNIBS3L1_15_LC_20_9_2.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_41_RNIBS3L1_15_LC_20_9_2 (
            .in0(N__74709),
            .in1(N__78779),
            .in2(N__73078),
            .in3(N__76841),
            .lcout(rco_int_0_a2_1_a2_1_48),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_41_RNIK8RU1_15_LC_20_9_3.C_ON=1'b0;
    defparam shift_srl_41_RNIK8RU1_15_LC_20_9_3.SEQ_MODE=4'b0000;
    defparam shift_srl_41_RNIK8RU1_15_LC_20_9_3.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_41_RNIK8RU1_15_LC_20_9_3 (
            .in0(N__78778),
            .in1(N__76608),
            .in2(N__74715),
            .in3(N__81526),
            .lcout(),
            .ltout(rco_int_0_a2_0_a2_83_m6_0_a2_3_sx_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_41_RNIM3K34_15_LC_20_9_4.C_ON=1'b0;
    defparam shift_srl_41_RNIM3K34_15_LC_20_9_4.SEQ_MODE=4'b0000;
    defparam shift_srl_41_RNIM3K34_15_LC_20_9_4.LUT_INIT=16'b0000100000000000;
    LogicCell40 shift_srl_41_RNIM3K34_15_LC_20_9_4 (
            .in0(N__75135),
            .in1(N__74739),
            .in2(N__73075),
            .in3(N__76842),
            .lcout(rco_int_0_a2_0_a2_83_m6_0_a2_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_53_RNI66TQ_15_LC_20_9_5.C_ON=1'b0;
    defparam shift_srl_53_RNI66TQ_15_LC_20_9_5.SEQ_MODE=4'b0000;
    defparam shift_srl_53_RNI66TQ_15_LC_20_9_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_53_RNI66TQ_15_LC_20_9_5 (
            .in0(N__76351),
            .in1(N__74628),
            .in2(N__76450),
            .in3(N__73041),
            .lcout(),
            .ltout(shift_srl_53_RNI66TQZ0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_49_RNIU8OU_15_LC_20_9_6.C_ON=1'b0;
    defparam shift_srl_49_RNIU8OU_15_LC_20_9_6.SEQ_MODE=4'b0000;
    defparam shift_srl_49_RNIU8OU_15_LC_20_9_6.LUT_INIT=16'b1110001011100010;
    LogicCell40 shift_srl_49_RNIU8OU_15_LC_20_9_6 (
            .in0(_gnd_net_),
            .in1(N__93477),
            .in2(N__73030),
            .in3(_gnd_net_),
            .lcout(rco_int_0_a2_1_a2_0_53),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_56_10_LC_20_10_0.C_ON=1'b0;
    defparam shift_srl_56_10_LC_20_10_0.SEQ_MODE=4'b1000;
    defparam shift_srl_56_10_LC_20_10_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_56_10_LC_20_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73120),
            .lcout(shift_srl_56Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93272),
            .ce(N__78828),
            .sr(_gnd_net_));
    defparam shift_srl_56_11_LC_20_10_1.C_ON=1'b0;
    defparam shift_srl_56_11_LC_20_10_1.SEQ_MODE=4'b1000;
    defparam shift_srl_56_11_LC_20_10_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_56_11_LC_20_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73027),
            .lcout(shift_srl_56Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93272),
            .ce(N__78828),
            .sr(_gnd_net_));
    defparam shift_srl_56_12_LC_20_10_2.C_ON=1'b0;
    defparam shift_srl_56_12_LC_20_10_2.SEQ_MODE=4'b1000;
    defparam shift_srl_56_12_LC_20_10_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_56_12_LC_20_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73144),
            .lcout(shift_srl_56Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93272),
            .ce(N__78828),
            .sr(_gnd_net_));
    defparam shift_srl_56_13_LC_20_10_3.C_ON=1'b0;
    defparam shift_srl_56_13_LC_20_10_3.SEQ_MODE=4'b1000;
    defparam shift_srl_56_13_LC_20_10_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_56_13_LC_20_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73138),
            .lcout(shift_srl_56Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93272),
            .ce(N__78828),
            .sr(_gnd_net_));
    defparam shift_srl_56_14_LC_20_10_4.C_ON=1'b0;
    defparam shift_srl_56_14_LC_20_10_4.SEQ_MODE=4'b1000;
    defparam shift_srl_56_14_LC_20_10_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_56_14_LC_20_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73132),
            .lcout(shift_srl_56Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93272),
            .ce(N__78828),
            .sr(_gnd_net_));
    defparam shift_srl_56_15_LC_20_10_5.C_ON=1'b0;
    defparam shift_srl_56_15_LC_20_10_5.SEQ_MODE=4'b1000;
    defparam shift_srl_56_15_LC_20_10_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_56_15_LC_20_10_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73126),
            .lcout(shift_srl_56Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93272),
            .ce(N__78828),
            .sr(_gnd_net_));
    defparam shift_srl_56_9_LC_20_10_6.C_ON=1'b0;
    defparam shift_srl_56_9_LC_20_10_6.SEQ_MODE=4'b1000;
    defparam shift_srl_56_9_LC_20_10_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_56_9_LC_20_10_6 (
            .in0(N__78838),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_56Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93272),
            .ce(N__78828),
            .sr(_gnd_net_));
    defparam shift_srl_56_0_LC_20_10_7.C_ON=1'b0;
    defparam shift_srl_56_0_LC_20_10_7.SEQ_MODE=4'b1000;
    defparam shift_srl_56_0_LC_20_10_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_56_0_LC_20_10_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76532),
            .lcout(shift_srl_56Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93272),
            .ce(N__78828),
            .sr(_gnd_net_));
    defparam shift_srl_58_RNIQMNU_15_LC_20_11_0.C_ON=1'b0;
    defparam shift_srl_58_RNIQMNU_15_LC_20_11_0.SEQ_MODE=4'b0000;
    defparam shift_srl_58_RNIQMNU_15_LC_20_11_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_58_RNIQMNU_15_LC_20_11_0 (
            .in0(N__76798),
            .in1(N__79006),
            .in2(N__74875),
            .in3(N__76526),
            .lcout(),
            .ltout(shift_srl_58_RNIQMNUZ0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_54_RNIEAU71_15_LC_20_11_1.C_ON=1'b0;
    defparam shift_srl_54_RNIEAU71_15_LC_20_11_1.SEQ_MODE=4'b0000;
    defparam shift_srl_54_RNIEAU71_15_LC_20_11_1.LUT_INIT=16'b1111000010101010;
    LogicCell40 shift_srl_54_RNIEAU71_15_LC_20_11_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__73114),
            .in3(N__77004),
            .lcout(shift_srl_54_RNIEAU71Z0Z_15),
            .ltout(shift_srl_54_RNIEAU71Z0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNID951F_15_LC_20_11_2.C_ON=1'b0;
    defparam shift_srl_0_RNID951F_15_LC_20_11_2.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNID951F_15_LC_20_11_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNID951F_15_LC_20_11_2 (
            .in0(N__81540),
            .in1(N__90013),
            .in2(N__73111),
            .in3(N__93565),
            .lcout(clk_en_59),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_55_15_LC_20_11_3.C_ON=1'b0;
    defparam shift_srl_55_15_LC_20_11_3.SEQ_MODE=4'b1000;
    defparam shift_srl_55_15_LC_20_11_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_55_15_LC_20_11_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73192),
            .lcout(shift_srl_55Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93253),
            .ce(N__74894),
            .sr(_gnd_net_));
    defparam shift_srl_55_14_LC_20_11_4.C_ON=1'b0;
    defparam shift_srl_55_14_LC_20_11_4.SEQ_MODE=4'b1000;
    defparam shift_srl_55_14_LC_20_11_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_55_14_LC_20_11_4 (
            .in0(N__73186),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_55Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93253),
            .ce(N__74894),
            .sr(_gnd_net_));
    defparam shift_srl_55_13_LC_20_11_5.C_ON=1'b0;
    defparam shift_srl_55_13_LC_20_11_5.SEQ_MODE=4'b1000;
    defparam shift_srl_55_13_LC_20_11_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_55_13_LC_20_11_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73180),
            .lcout(shift_srl_55Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93253),
            .ce(N__74894),
            .sr(_gnd_net_));
    defparam shift_srl_55_12_LC_20_11_6.C_ON=1'b0;
    defparam shift_srl_55_12_LC_20_11_6.SEQ_MODE=4'b1000;
    defparam shift_srl_55_12_LC_20_11_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_55_12_LC_20_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73174),
            .lcout(shift_srl_55Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93253),
            .ce(N__74894),
            .sr(_gnd_net_));
    defparam shift_srl_55_11_LC_20_11_7.C_ON=1'b0;
    defparam shift_srl_55_11_LC_20_11_7.SEQ_MODE=4'b1000;
    defparam shift_srl_55_11_LC_20_11_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_55_11_LC_20_11_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73351),
            .lcout(shift_srl_55Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93253),
            .ce(N__74894),
            .sr(_gnd_net_));
    defparam shift_srl_55_0_LC_20_12_0.C_ON=1'b0;
    defparam shift_srl_55_0_LC_20_12_0.SEQ_MODE=4'b1000;
    defparam shift_srl_55_0_LC_20_12_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_55_0_LC_20_12_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74874),
            .lcout(shift_srl_55Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93231),
            .ce(N__74901),
            .sr(_gnd_net_));
    defparam shift_srl_55_1_LC_20_12_1.C_ON=1'b0;
    defparam shift_srl_55_1_LC_20_12_1.SEQ_MODE=4'b1000;
    defparam shift_srl_55_1_LC_20_12_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_55_1_LC_20_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73168),
            .lcout(shift_srl_55Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93231),
            .ce(N__74901),
            .sr(_gnd_net_));
    defparam shift_srl_55_2_LC_20_12_2.C_ON=1'b0;
    defparam shift_srl_55_2_LC_20_12_2.SEQ_MODE=4'b1000;
    defparam shift_srl_55_2_LC_20_12_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_55_2_LC_20_12_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73162),
            .lcout(shift_srl_55Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93231),
            .ce(N__74901),
            .sr(_gnd_net_));
    defparam shift_srl_55_3_LC_20_12_3.C_ON=1'b0;
    defparam shift_srl_55_3_LC_20_12_3.SEQ_MODE=4'b1000;
    defparam shift_srl_55_3_LC_20_12_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_55_3_LC_20_12_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73156),
            .lcout(shift_srl_55Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93231),
            .ce(N__74901),
            .sr(_gnd_net_));
    defparam shift_srl_55_4_LC_20_12_4.C_ON=1'b0;
    defparam shift_srl_55_4_LC_20_12_4.SEQ_MODE=4'b1000;
    defparam shift_srl_55_4_LC_20_12_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_55_4_LC_20_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73150),
            .lcout(shift_srl_55Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93231),
            .ce(N__74901),
            .sr(_gnd_net_));
    defparam shift_srl_55_5_LC_20_12_5.C_ON=1'b0;
    defparam shift_srl_55_5_LC_20_12_5.SEQ_MODE=4'b1000;
    defparam shift_srl_55_5_LC_20_12_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_55_5_LC_20_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73309),
            .lcout(shift_srl_55Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93231),
            .ce(N__74901),
            .sr(_gnd_net_));
    defparam shift_srl_55_6_LC_20_12_6.C_ON=1'b0;
    defparam shift_srl_55_6_LC_20_12_6.SEQ_MODE=4'b1000;
    defparam shift_srl_55_6_LC_20_12_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_55_6_LC_20_12_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73303),
            .lcout(shift_srl_55Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93231),
            .ce(N__74901),
            .sr(_gnd_net_));
    defparam shift_srl_55_7_LC_20_12_7.C_ON=1'b0;
    defparam shift_srl_55_7_LC_20_12_7.SEQ_MODE=4'b1000;
    defparam shift_srl_55_7_LC_20_12_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_55_7_LC_20_12_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73297),
            .lcout(shift_srl_55Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93231),
            .ce(N__74901),
            .sr(_gnd_net_));
    defparam shift_srl_48_RNILVDK5_15_LC_20_13_0.C_ON=1'b0;
    defparam shift_srl_48_RNILVDK5_15_LC_20_13_0.SEQ_MODE=4'b0000;
    defparam shift_srl_48_RNILVDK5_15_LC_20_13_0.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_48_RNILVDK5_15_LC_20_13_0 (
            .in0(N__76594),
            .in1(N__76856),
            .in2(N__74480),
            .in3(N__81550),
            .lcout(rco_int_0_a2_1_a2_sx_53),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_48_RNISHHA7_15_LC_20_13_1.C_ON=1'b0;
    defparam shift_srl_48_RNISHHA7_15_LC_20_13_1.SEQ_MODE=4'b0000;
    defparam shift_srl_48_RNISHHA7_15_LC_20_13_1.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_48_RNISHHA7_15_LC_20_13_1 (
            .in0(N__76855),
            .in1(N__76593),
            .in2(N__81442),
            .in3(N__74469),
            .lcout(rco_int_0_a2_1_a2_sx_59),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_44_RNIMV201_15_LC_20_13_2.C_ON=1'b0;
    defparam shift_srl_44_RNIMV201_15_LC_20_13_2.SEQ_MODE=4'b0000;
    defparam shift_srl_44_RNIMV201_15_LC_20_13_2.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_44_RNIMV201_15_LC_20_13_2 (
            .in0(N__73290),
            .in1(N__73278),
            .in2(_gnd_net_),
            .in3(N__73238),
            .lcout(rco_int_0_a2_1_a2_0_44),
            .ltout(rco_int_0_a2_1_a2_0_44_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_48_RNIDUNF1_15_LC_20_13_3.C_ON=1'b0;
    defparam shift_srl_48_RNIDUNF1_15_LC_20_13_3.SEQ_MODE=4'b0000;
    defparam shift_srl_48_RNIDUNF1_15_LC_20_13_3.LUT_INIT=16'b0000111111111111;
    LogicCell40 shift_srl_48_RNIDUNF1_15_LC_20_13_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__73201),
            .in3(N__76592),
            .lcout(rco_int_0_a3_0_a2cf1_1_66),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_48_15_LC_20_13_4.C_ON=1'b0;
    defparam shift_srl_48_15_LC_20_13_4.SEQ_MODE=4'b1000;
    defparam shift_srl_48_15_LC_20_13_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_48_15_LC_20_13_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73198),
            .lcout(shift_srl_48Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93213),
            .ce(N__73380),
            .sr(_gnd_net_));
    defparam shift_srl_48_14_LC_20_13_5.C_ON=1'b0;
    defparam shift_srl_48_14_LC_20_13_5.SEQ_MODE=4'b1000;
    defparam shift_srl_48_14_LC_20_13_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_48_14_LC_20_13_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73399),
            .lcout(shift_srl_48Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93213),
            .ce(N__73380),
            .sr(_gnd_net_));
    defparam shift_srl_48_13_LC_20_13_6.C_ON=1'b0;
    defparam shift_srl_48_13_LC_20_13_6.SEQ_MODE=4'b1000;
    defparam shift_srl_48_13_LC_20_13_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_48_13_LC_20_13_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73387),
            .lcout(shift_srl_48Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93213),
            .ce(N__73380),
            .sr(_gnd_net_));
    defparam shift_srl_48_12_LC_20_13_7.C_ON=1'b0;
    defparam shift_srl_48_12_LC_20_13_7.SEQ_MODE=4'b1000;
    defparam shift_srl_48_12_LC_20_13_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_48_12_LC_20_13_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73393),
            .lcout(shift_srl_48Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93213),
            .ce(N__73380),
            .sr(_gnd_net_));
    defparam shift_srl_55_10_LC_20_14_0.C_ON=1'b0;
    defparam shift_srl_55_10_LC_20_14_0.SEQ_MODE=4'b1000;
    defparam shift_srl_55_10_LC_20_14_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_55_10_LC_20_14_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73342),
            .lcout(shift_srl_55Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93193),
            .ce(N__74902),
            .sr(_gnd_net_));
    defparam shift_srl_55_9_LC_20_14_1.C_ON=1'b0;
    defparam shift_srl_55_9_LC_20_14_1.SEQ_MODE=4'b1000;
    defparam shift_srl_55_9_LC_20_14_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_55_9_LC_20_14_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73327),
            .lcout(shift_srl_55Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93193),
            .ce(N__74902),
            .sr(_gnd_net_));
    defparam shift_srl_55_8_LC_20_14_2.C_ON=1'b0;
    defparam shift_srl_55_8_LC_20_14_2.SEQ_MODE=4'b1000;
    defparam shift_srl_55_8_LC_20_14_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_55_8_LC_20_14_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73336),
            .lcout(shift_srl_55Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93193),
            .ce(N__74902),
            .sr(_gnd_net_));
    defparam shift_srl_61_10_LC_20_15_0.C_ON=1'b0;
    defparam shift_srl_61_10_LC_20_15_0.SEQ_MODE=4'b1000;
    defparam shift_srl_61_10_LC_20_15_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_61_10_LC_20_15_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73444),
            .lcout(shift_srl_61Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93172),
            .ce(N__73416),
            .sr(_gnd_net_));
    defparam shift_srl_61_0_LC_20_15_1.C_ON=1'b0;
    defparam shift_srl_61_0_LC_20_15_1.SEQ_MODE=4'b1000;
    defparam shift_srl_61_0_LC_20_15_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_61_0_LC_20_15_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73435),
            .lcout(shift_srl_61Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93172),
            .ce(N__73416),
            .sr(_gnd_net_));
    defparam shift_srl_61_12_LC_20_15_2.C_ON=1'b0;
    defparam shift_srl_61_12_LC_20_15_2.SEQ_MODE=4'b1000;
    defparam shift_srl_61_12_LC_20_15_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_61_12_LC_20_15_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73456),
            .lcout(shift_srl_61Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93172),
            .ce(N__73416),
            .sr(_gnd_net_));
    defparam shift_srl_61_13_LC_20_15_3.C_ON=1'b0;
    defparam shift_srl_61_13_LC_20_15_3.SEQ_MODE=4'b1000;
    defparam shift_srl_61_13_LC_20_15_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_61_13_LC_20_15_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73315),
            .lcout(shift_srl_61Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93172),
            .ce(N__73416),
            .sr(_gnd_net_));
    defparam shift_srl_61_14_LC_20_15_4.C_ON=1'b0;
    defparam shift_srl_61_14_LC_20_15_4.SEQ_MODE=4'b1000;
    defparam shift_srl_61_14_LC_20_15_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_61_14_LC_20_15_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73474),
            .lcout(shift_srl_61Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93172),
            .ce(N__73416),
            .sr(_gnd_net_));
    defparam shift_srl_61_15_LC_20_15_5.C_ON=1'b0;
    defparam shift_srl_61_15_LC_20_15_5.SEQ_MODE=4'b1000;
    defparam shift_srl_61_15_LC_20_15_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_61_15_LC_20_15_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73468),
            .lcout(shift_srl_61Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93172),
            .ce(N__73416),
            .sr(_gnd_net_));
    defparam shift_srl_61_11_LC_20_15_6.C_ON=1'b0;
    defparam shift_srl_61_11_LC_20_15_6.SEQ_MODE=4'b1000;
    defparam shift_srl_61_11_LC_20_15_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_61_11_LC_20_15_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73462),
            .lcout(shift_srl_61Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93172),
            .ce(N__73416),
            .sr(_gnd_net_));
    defparam shift_srl_61_9_LC_20_15_7.C_ON=1'b0;
    defparam shift_srl_61_9_LC_20_15_7.SEQ_MODE=4'b1000;
    defparam shift_srl_61_9_LC_20_15_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_61_9_LC_20_15_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73450),
            .lcout(shift_srl_61Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93172),
            .ce(N__73416),
            .sr(_gnd_net_));
    defparam shift_srl_61_RNI3LM9_15_LC_20_16_1.C_ON=1'b0;
    defparam shift_srl_61_RNI3LM9_15_LC_20_16_1.SEQ_MODE=4'b0000;
    defparam shift_srl_61_RNI3LM9_15_LC_20_16_1.LUT_INIT=16'b1100110000000000;
    LogicCell40 shift_srl_61_RNI3LM9_15_LC_20_16_1 (
            .in0(_gnd_net_),
            .in1(N__73434),
            .in2(_gnd_net_),
            .in3(N__75331),
            .lcout(shift_srl_61_RNI3LM9Z0Z_15),
            .ltout(shift_srl_61_RNI3LM9Z0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNI961PF_15_LC_20_16_2.C_ON=1'b0;
    defparam shift_srl_0_RNI961PF_15_LC_20_16_2.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNI961PF_15_LC_20_16_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNI961PF_15_LC_20_16_2 (
            .in0(N__90585),
            .in1(N__81444),
            .in2(N__73438),
            .in3(N__93595),
            .lcout(clk_en_62),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_62_RNIM5RK_15_LC_20_16_3.C_ON=1'b0;
    defparam shift_srl_62_RNIM5RK_15_LC_20_16_3.SEQ_MODE=4'b0000;
    defparam shift_srl_62_RNIM5RK_15_LC_20_16_3.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_62_RNIM5RK_15_LC_20_16_3 (
            .in0(N__73515),
            .in1(N__73433),
            .in2(_gnd_net_),
            .in3(N__75330),
            .lcout(shift_srl_62_RNIM5RKZ0Z_15),
            .ltout(shift_srl_62_RNIM5RKZ0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_64_RNICGAR1_15_LC_20_16_4.C_ON=1'b0;
    defparam shift_srl_64_RNICGAR1_15_LC_20_16_4.SEQ_MODE=4'b0000;
    defparam shift_srl_64_RNICGAR1_15_LC_20_16_4.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_64_RNICGAR1_15_LC_20_16_4 (
            .in0(N__81092),
            .in1(N__81137),
            .in2(N__73420),
            .in3(N__75001),
            .lcout(rco_int_0_a3_0_a2_0_66),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_60_RNINP2IF_15_LC_20_16_6.C_ON=1'b0;
    defparam shift_srl_60_RNINP2IF_15_LC_20_16_6.SEQ_MODE=4'b0000;
    defparam shift_srl_60_RNINP2IF_15_LC_20_16_6.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_60_RNINP2IF_15_LC_20_16_6 (
            .in0(N__75332),
            .in1(N__81443),
            .in2(N__90586),
            .in3(N__93593),
            .lcout(clk_en_61),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNISM54G_15_LC_20_16_7.C_ON=1'b0;
    defparam shift_srl_0_RNISM54G_15_LC_20_16_7.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNISM54G_15_LC_20_16_7.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNISM54G_15_LC_20_16_7 (
            .in0(N__93594),
            .in1(N__90584),
            .in2(N__81032),
            .in3(N__81445),
            .lcout(clk_en_63),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_62_10_LC_20_17_0.C_ON=1'b0;
    defparam shift_srl_62_10_LC_20_17_0.SEQ_MODE=4'b1000;
    defparam shift_srl_62_10_LC_20_17_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_62_10_LC_20_17_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73504),
            .lcout(shift_srl_62Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93117),
            .ce(N__73485),
            .sr(_gnd_net_));
    defparam shift_srl_62_11_LC_20_17_1.C_ON=1'b0;
    defparam shift_srl_62_11_LC_20_17_1.SEQ_MODE=4'b1000;
    defparam shift_srl_62_11_LC_20_17_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_62_11_LC_20_17_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73546),
            .lcout(shift_srl_62Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93117),
            .ce(N__73485),
            .sr(_gnd_net_));
    defparam shift_srl_62_12_LC_20_17_2.C_ON=1'b0;
    defparam shift_srl_62_12_LC_20_17_2.SEQ_MODE=4'b1000;
    defparam shift_srl_62_12_LC_20_17_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_62_12_LC_20_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73540),
            .lcout(shift_srl_62Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93117),
            .ce(N__73485),
            .sr(_gnd_net_));
    defparam shift_srl_62_13_LC_20_17_3.C_ON=1'b0;
    defparam shift_srl_62_13_LC_20_17_3.SEQ_MODE=4'b1000;
    defparam shift_srl_62_13_LC_20_17_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_62_13_LC_20_17_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73534),
            .lcout(shift_srl_62Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93117),
            .ce(N__73485),
            .sr(_gnd_net_));
    defparam shift_srl_62_14_LC_20_17_4.C_ON=1'b0;
    defparam shift_srl_62_14_LC_20_17_4.SEQ_MODE=4'b1000;
    defparam shift_srl_62_14_LC_20_17_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_62_14_LC_20_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73528),
            .lcout(shift_srl_62Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93117),
            .ce(N__73485),
            .sr(_gnd_net_));
    defparam shift_srl_62_15_LC_20_17_5.C_ON=1'b0;
    defparam shift_srl_62_15_LC_20_17_5.SEQ_MODE=4'b1000;
    defparam shift_srl_62_15_LC_20_17_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_62_15_LC_20_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73522),
            .lcout(shift_srl_62Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93117),
            .ce(N__73485),
            .sr(_gnd_net_));
    defparam shift_srl_62_9_LC_20_17_6.C_ON=1'b0;
    defparam shift_srl_62_9_LC_20_17_6.SEQ_MODE=4'b1000;
    defparam shift_srl_62_9_LC_20_17_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_62_9_LC_20_17_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73492),
            .lcout(shift_srl_62Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93117),
            .ce(N__73485),
            .sr(_gnd_net_));
    defparam shift_srl_62_8_LC_20_17_7.C_ON=1'b0;
    defparam shift_srl_62_8_LC_20_17_7.SEQ_MODE=4'b1000;
    defparam shift_srl_62_8_LC_20_17_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_62_8_LC_20_17_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73498),
            .lcout(shift_srl_62Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93117),
            .ce(N__73485),
            .sr(_gnd_net_));
    defparam shift_srl_174_10_LC_20_18_0.C_ON=1'b0;
    defparam shift_srl_174_10_LC_20_18_0.SEQ_MODE=4'b1000;
    defparam shift_srl_174_10_LC_20_18_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_174_10_LC_20_18_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73585),
            .lcout(shift_srl_174Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93153),
            .ce(N__73567),
            .sr(_gnd_net_));
    defparam shift_srl_174_11_LC_20_18_1.C_ON=1'b0;
    defparam shift_srl_174_11_LC_20_18_1.SEQ_MODE=4'b1000;
    defparam shift_srl_174_11_LC_20_18_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_174_11_LC_20_18_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73615),
            .lcout(shift_srl_174Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93153),
            .ce(N__73567),
            .sr(_gnd_net_));
    defparam shift_srl_174_12_LC_20_18_2.C_ON=1'b0;
    defparam shift_srl_174_12_LC_20_18_2.SEQ_MODE=4'b1000;
    defparam shift_srl_174_12_LC_20_18_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_174_12_LC_20_18_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73609),
            .lcout(shift_srl_174Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93153),
            .ce(N__73567),
            .sr(_gnd_net_));
    defparam shift_srl_174_13_LC_20_18_3.C_ON=1'b0;
    defparam shift_srl_174_13_LC_20_18_3.SEQ_MODE=4'b1000;
    defparam shift_srl_174_13_LC_20_18_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_174_13_LC_20_18_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73603),
            .lcout(shift_srl_174Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93153),
            .ce(N__73567),
            .sr(_gnd_net_));
    defparam shift_srl_174_14_LC_20_18_4.C_ON=1'b0;
    defparam shift_srl_174_14_LC_20_18_4.SEQ_MODE=4'b1000;
    defparam shift_srl_174_14_LC_20_18_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_174_14_LC_20_18_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73597),
            .lcout(shift_srl_174Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93153),
            .ce(N__73567),
            .sr(_gnd_net_));
    defparam shift_srl_174_15_LC_20_18_5.C_ON=1'b0;
    defparam shift_srl_174_15_LC_20_18_5.SEQ_MODE=4'b1000;
    defparam shift_srl_174_15_LC_20_18_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_174_15_LC_20_18_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73591),
            .lcout(shift_srl_174Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93153),
            .ce(N__73567),
            .sr(_gnd_net_));
    defparam shift_srl_174_9_LC_20_18_6.C_ON=1'b0;
    defparam shift_srl_174_9_LC_20_18_6.SEQ_MODE=4'b1000;
    defparam shift_srl_174_9_LC_20_18_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_174_9_LC_20_18_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73573),
            .lcout(shift_srl_174Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93153),
            .ce(N__73567),
            .sr(_gnd_net_));
    defparam shift_srl_174_8_LC_20_18_7.C_ON=1'b0;
    defparam shift_srl_174_8_LC_20_18_7.SEQ_MODE=4'b1000;
    defparam shift_srl_174_8_LC_20_18_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_174_8_LC_20_18_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73579),
            .lcout(shift_srl_174Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93153),
            .ce(N__73567),
            .sr(_gnd_net_));
    defparam shift_srl_166_8_LC_20_19_0.C_ON=1'b0;
    defparam shift_srl_166_8_LC_20_19_0.SEQ_MODE=4'b1000;
    defparam shift_srl_166_8_LC_20_19_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_166_8_LC_20_19_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73633),
            .lcout(shift_srl_166Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93173),
            .ce(N__73698),
            .sr(_gnd_net_));
    defparam shift_srl_166_1_LC_20_19_1.C_ON=1'b0;
    defparam shift_srl_166_1_LC_20_19_1.SEQ_MODE=4'b1000;
    defparam shift_srl_166_1_LC_20_19_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_166_1_LC_20_19_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73705),
            .lcout(shift_srl_166Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93173),
            .ce(N__73698),
            .sr(_gnd_net_));
    defparam shift_srl_166_2_LC_20_19_2.C_ON=1'b0;
    defparam shift_srl_166_2_LC_20_19_2.SEQ_MODE=4'b1000;
    defparam shift_srl_166_2_LC_20_19_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_166_2_LC_20_19_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73669),
            .lcout(shift_srl_166Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93173),
            .ce(N__73698),
            .sr(_gnd_net_));
    defparam shift_srl_166_3_LC_20_19_3.C_ON=1'b0;
    defparam shift_srl_166_3_LC_20_19_3.SEQ_MODE=4'b1000;
    defparam shift_srl_166_3_LC_20_19_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_166_3_LC_20_19_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73663),
            .lcout(shift_srl_166Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93173),
            .ce(N__73698),
            .sr(_gnd_net_));
    defparam shift_srl_166_4_LC_20_19_4.C_ON=1'b0;
    defparam shift_srl_166_4_LC_20_19_4.SEQ_MODE=4'b1000;
    defparam shift_srl_166_4_LC_20_19_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_166_4_LC_20_19_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73657),
            .lcout(shift_srl_166Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93173),
            .ce(N__73698),
            .sr(_gnd_net_));
    defparam shift_srl_166_5_LC_20_19_5.C_ON=1'b0;
    defparam shift_srl_166_5_LC_20_19_5.SEQ_MODE=4'b1000;
    defparam shift_srl_166_5_LC_20_19_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_166_5_LC_20_19_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73651),
            .lcout(shift_srl_166Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93173),
            .ce(N__73698),
            .sr(_gnd_net_));
    defparam shift_srl_166_6_LC_20_19_6.C_ON=1'b0;
    defparam shift_srl_166_6_LC_20_19_6.SEQ_MODE=4'b1000;
    defparam shift_srl_166_6_LC_20_19_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_166_6_LC_20_19_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73645),
            .lcout(shift_srl_166Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93173),
            .ce(N__73698),
            .sr(_gnd_net_));
    defparam shift_srl_166_7_LC_20_19_7.C_ON=1'b0;
    defparam shift_srl_166_7_LC_20_19_7.SEQ_MODE=4'b1000;
    defparam shift_srl_166_7_LC_20_19_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_166_7_LC_20_19_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73639),
            .lcout(shift_srl_166Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93173),
            .ce(N__73698),
            .sr(_gnd_net_));
    defparam shift_srl_166_10_LC_20_20_0.C_ON=1'b0;
    defparam shift_srl_166_10_LC_20_20_0.SEQ_MODE=4'b1000;
    defparam shift_srl_166_10_LC_20_20_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_166_10_LC_20_20_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73711),
            .lcout(shift_srl_166Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93194),
            .ce(N__73699),
            .sr(_gnd_net_));
    defparam shift_srl_166_11_LC_20_20_1.C_ON=1'b0;
    defparam shift_srl_166_11_LC_20_20_1.SEQ_MODE=4'b1000;
    defparam shift_srl_166_11_LC_20_20_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_166_11_LC_20_20_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73627),
            .lcout(shift_srl_166Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93194),
            .ce(N__73699),
            .sr(_gnd_net_));
    defparam shift_srl_166_12_LC_20_20_2.C_ON=1'b0;
    defparam shift_srl_166_12_LC_20_20_2.SEQ_MODE=4'b1000;
    defparam shift_srl_166_12_LC_20_20_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_166_12_LC_20_20_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73621),
            .lcout(shift_srl_166Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93194),
            .ce(N__73699),
            .sr(_gnd_net_));
    defparam shift_srl_166_13_LC_20_20_3.C_ON=1'b0;
    defparam shift_srl_166_13_LC_20_20_3.SEQ_MODE=4'b1000;
    defparam shift_srl_166_13_LC_20_20_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_166_13_LC_20_20_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73735),
            .lcout(shift_srl_166Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93194),
            .ce(N__73699),
            .sr(_gnd_net_));
    defparam shift_srl_166_14_LC_20_20_4.C_ON=1'b0;
    defparam shift_srl_166_14_LC_20_20_4.SEQ_MODE=4'b1000;
    defparam shift_srl_166_14_LC_20_20_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_166_14_LC_20_20_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73729),
            .lcout(shift_srl_166Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93194),
            .ce(N__73699),
            .sr(_gnd_net_));
    defparam shift_srl_166_15_LC_20_20_5.C_ON=1'b0;
    defparam shift_srl_166_15_LC_20_20_5.SEQ_MODE=4'b1000;
    defparam shift_srl_166_15_LC_20_20_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_166_15_LC_20_20_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73723),
            .lcout(shift_srl_166Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93194),
            .ce(N__73699),
            .sr(_gnd_net_));
    defparam shift_srl_166_9_LC_20_20_6.C_ON=1'b0;
    defparam shift_srl_166_9_LC_20_20_6.SEQ_MODE=4'b1000;
    defparam shift_srl_166_9_LC_20_20_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_166_9_LC_20_20_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73717),
            .lcout(shift_srl_166Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93194),
            .ce(N__73699),
            .sr(_gnd_net_));
    defparam shift_srl_166_0_LC_20_20_7.C_ON=1'b0;
    defparam shift_srl_166_0_LC_20_20_7.SEQ_MODE=4'b1000;
    defparam shift_srl_166_0_LC_20_20_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_166_0_LC_20_20_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84010),
            .lcout(shift_srl_166Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93194),
            .ce(N__73699),
            .sr(_gnd_net_));
    defparam shift_srl_184_10_LC_20_21_0.C_ON=1'b0;
    defparam shift_srl_184_10_LC_20_21_0.SEQ_MODE=4'b1000;
    defparam shift_srl_184_10_LC_20_21_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_184_10_LC_20_21_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73783),
            .lcout(shift_srl_184Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93214),
            .ce(N__73934),
            .sr(_gnd_net_));
    defparam shift_srl_184_11_LC_20_21_1.C_ON=1'b0;
    defparam shift_srl_184_11_LC_20_21_1.SEQ_MODE=4'b1000;
    defparam shift_srl_184_11_LC_20_21_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_184_11_LC_20_21_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73687),
            .lcout(shift_srl_184Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93214),
            .ce(N__73934),
            .sr(_gnd_net_));
    defparam shift_srl_184_12_LC_20_21_2.C_ON=1'b0;
    defparam shift_srl_184_12_LC_20_21_2.SEQ_MODE=4'b1000;
    defparam shift_srl_184_12_LC_20_21_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_184_12_LC_20_21_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73681),
            .lcout(shift_srl_184Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93214),
            .ce(N__73934),
            .sr(_gnd_net_));
    defparam shift_srl_184_13_LC_20_21_3.C_ON=1'b0;
    defparam shift_srl_184_13_LC_20_21_3.SEQ_MODE=4'b1000;
    defparam shift_srl_184_13_LC_20_21_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_184_13_LC_20_21_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73675),
            .lcout(shift_srl_184Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93214),
            .ce(N__73934),
            .sr(_gnd_net_));
    defparam shift_srl_184_14_LC_20_21_4.C_ON=1'b0;
    defparam shift_srl_184_14_LC_20_21_4.SEQ_MODE=4'b1000;
    defparam shift_srl_184_14_LC_20_21_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_184_14_LC_20_21_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73789),
            .lcout(shift_srl_184Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93214),
            .ce(N__73934),
            .sr(_gnd_net_));
    defparam shift_srl_184_9_LC_20_21_5.C_ON=1'b0;
    defparam shift_srl_184_9_LC_20_21_5.SEQ_MODE=4'b1000;
    defparam shift_srl_184_9_LC_20_21_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_184_9_LC_20_21_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73771),
            .lcout(shift_srl_184Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93214),
            .ce(N__73934),
            .sr(_gnd_net_));
    defparam shift_srl_184_8_LC_20_21_6.C_ON=1'b0;
    defparam shift_srl_184_8_LC_20_21_6.SEQ_MODE=4'b1000;
    defparam shift_srl_184_8_LC_20_21_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_184_8_LC_20_21_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73777),
            .lcout(shift_srl_184Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93214),
            .ce(N__73934),
            .sr(_gnd_net_));
    defparam shift_srl_186_0_LC_20_22_0.C_ON=1'b0;
    defparam shift_srl_186_0_LC_20_22_0.SEQ_MODE=4'b1000;
    defparam shift_srl_186_0_LC_20_22_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_186_0_LC_20_22_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__91807),
            .lcout(shift_srl_186Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93232),
            .ce(N__75567),
            .sr(_gnd_net_));
    defparam shift_srl_186_1_LC_20_22_1.C_ON=1'b0;
    defparam shift_srl_186_1_LC_20_22_1.SEQ_MODE=4'b1000;
    defparam shift_srl_186_1_LC_20_22_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_186_1_LC_20_22_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73765),
            .lcout(shift_srl_186Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93232),
            .ce(N__75567),
            .sr(_gnd_net_));
    defparam shift_srl_186_2_LC_20_22_2.C_ON=1'b0;
    defparam shift_srl_186_2_LC_20_22_2.SEQ_MODE=4'b1000;
    defparam shift_srl_186_2_LC_20_22_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_186_2_LC_20_22_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73759),
            .lcout(shift_srl_186Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93232),
            .ce(N__75567),
            .sr(_gnd_net_));
    defparam shift_srl_186_3_LC_20_22_3.C_ON=1'b0;
    defparam shift_srl_186_3_LC_20_22_3.SEQ_MODE=4'b1000;
    defparam shift_srl_186_3_LC_20_22_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_186_3_LC_20_22_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73753),
            .lcout(shift_srl_186Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93232),
            .ce(N__75567),
            .sr(_gnd_net_));
    defparam shift_srl_186_4_LC_20_22_4.C_ON=1'b0;
    defparam shift_srl_186_4_LC_20_22_4.SEQ_MODE=4'b1000;
    defparam shift_srl_186_4_LC_20_22_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_186_4_LC_20_22_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73747),
            .lcout(shift_srl_186Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93232),
            .ce(N__75567),
            .sr(_gnd_net_));
    defparam shift_srl_186_5_LC_20_22_5.C_ON=1'b0;
    defparam shift_srl_186_5_LC_20_22_5.SEQ_MODE=4'b1000;
    defparam shift_srl_186_5_LC_20_22_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_186_5_LC_20_22_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73741),
            .lcout(shift_srl_186Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93232),
            .ce(N__75567),
            .sr(_gnd_net_));
    defparam shift_srl_186_6_LC_20_22_6.C_ON=1'b0;
    defparam shift_srl_186_6_LC_20_22_6.SEQ_MODE=4'b1000;
    defparam shift_srl_186_6_LC_20_22_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_186_6_LC_20_22_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73960),
            .lcout(shift_srl_186Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93232),
            .ce(N__75567),
            .sr(_gnd_net_));
    defparam shift_srl_186_7_LC_20_22_7.C_ON=1'b0;
    defparam shift_srl_186_7_LC_20_22_7.SEQ_MODE=4'b1000;
    defparam shift_srl_186_7_LC_20_22_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_186_7_LC_20_22_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73954),
            .lcout(shift_srl_186Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93232),
            .ce(N__75567),
            .sr(_gnd_net_));
    defparam shift_srl_185_RNIVQEHE1_15_LC_20_23_0.C_ON=1'b0;
    defparam shift_srl_185_RNIVQEHE1_15_LC_20_23_0.SEQ_MODE=4'b0000;
    defparam shift_srl_185_RNIVQEHE1_15_LC_20_23_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_185_RNIVQEHE1_15_LC_20_23_0 (
            .in0(N__91761),
            .in1(N__91647),
            .in2(N__90560),
            .in3(N__91457),
            .lcout(clk_en_186),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_184_15_LC_20_23_1.C_ON=1'b0;
    defparam shift_srl_184_15_LC_20_23_1.SEQ_MODE=4'b1000;
    defparam shift_srl_184_15_LC_20_23_1.LUT_INIT=16'b1100110011001100;
    LogicCell40 shift_srl_184_15_LC_20_23_1 (
            .in0(_gnd_net_),
            .in1(N__73948),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_184Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93254),
            .ce(N__73939),
            .sr(_gnd_net_));
    defparam shift_srl_187_RNI6LJV_15_LC_20_23_2.C_ON=1'b0;
    defparam shift_srl_187_RNI6LJV_15_LC_20_23_2.SEQ_MODE=4'b0000;
    defparam shift_srl_187_RNI6LJV_15_LC_20_23_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_187_RNI6LJV_15_LC_20_23_2 (
            .in0(N__91798),
            .in1(N__91742),
            .in2(N__86169),
            .in3(N__91646),
            .lcout(N_4173),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_191_RNI4FF31_15_LC_20_23_3.C_ON=1'b0;
    defparam shift_srl_191_RNI4FF31_15_LC_20_23_3.SEQ_MODE=4'b0000;
    defparam shift_srl_191_RNI4FF31_15_LC_20_23_3.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_191_RNI4FF31_15_LC_20_23_3 (
            .in0(N__91608),
            .in1(N__86136),
            .in2(N__85783),
            .in3(N__86103),
            .lcout(clk_en_0_a2_0_a2_0_sx_192),
            .ltout(clk_en_0_a2_0_a2_0_sx_192_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_193_RNIPGCE2_15_LC_20_23_4.C_ON=1'b0;
    defparam shift_srl_193_RNIPGCE2_15_LC_20_23_4.SEQ_MODE=4'b0000;
    defparam shift_srl_193_RNIPGCE2_15_LC_20_23_4.LUT_INIT=16'b0000100000000000;
    LogicCell40 shift_srl_193_RNIPGCE2_15_LC_20_23_4 (
            .in0(N__76105),
            .in1(N__74218),
            .in2(N__73909),
            .in3(N__80334),
            .lcout(N_4179),
            .ltout(N_4179_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_194_RNIGLB4H1_15_LC_20_23_5.C_ON=1'b0;
    defparam shift_srl_194_RNIGLB4H1_15_LC_20_23_5.SEQ_MODE=4'b0000;
    defparam shift_srl_194_RNIGLB4H1_15_LC_20_23_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_194_RNIGLB4H1_15_LC_20_23_5 (
            .in0(N__91458),
            .in1(N__73901),
            .in2(N__73906),
            .in3(N__90513),
            .lcout(clk_en_195),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_195_RNICDEQ2_15_LC_20_23_6.C_ON=1'b0;
    defparam shift_srl_195_RNICDEQ2_15_LC_20_23_6.SEQ_MODE=4'b0000;
    defparam shift_srl_195_RNICDEQ2_15_LC_20_23_6.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_195_RNICDEQ2_15_LC_20_23_6 (
            .in0(N__74037),
            .in1(N__73900),
            .in2(_gnd_net_),
            .in3(N__73845),
            .lcout(N_4181),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_191_RNIA4332_15_LC_20_23_7.C_ON=1'b0;
    defparam shift_srl_191_RNIA4332_15_LC_20_23_7.SEQ_MODE=4'b0000;
    defparam shift_srl_191_RNIA4332_15_LC_20_23_7.LUT_INIT=16'b0000000010101010;
    LogicCell40 shift_srl_191_RNIA4332_15_LC_20_23_7 (
            .in0(N__80335),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74044),
            .lcout(N_4177),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_195_0_LC_20_24_0.C_ON=1'b0;
    defparam shift_srl_195_0_LC_20_24_0.SEQ_MODE=4'b1000;
    defparam shift_srl_195_0_LC_20_24_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_195_0_LC_20_24_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74038),
            .lcout(shift_srl_195Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93273),
            .ce(N__73977),
            .sr(_gnd_net_));
    defparam shift_srl_195_1_LC_20_24_1.C_ON=1'b0;
    defparam shift_srl_195_1_LC_20_24_1.SEQ_MODE=4'b1000;
    defparam shift_srl_195_1_LC_20_24_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_195_1_LC_20_24_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74026),
            .lcout(shift_srl_195Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93273),
            .ce(N__73977),
            .sr(_gnd_net_));
    defparam shift_srl_195_2_LC_20_24_2.C_ON=1'b0;
    defparam shift_srl_195_2_LC_20_24_2.SEQ_MODE=4'b1000;
    defparam shift_srl_195_2_LC_20_24_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_195_2_LC_20_24_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74020),
            .lcout(shift_srl_195Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93273),
            .ce(N__73977),
            .sr(_gnd_net_));
    defparam shift_srl_195_3_LC_20_24_3.C_ON=1'b0;
    defparam shift_srl_195_3_LC_20_24_3.SEQ_MODE=4'b1000;
    defparam shift_srl_195_3_LC_20_24_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_195_3_LC_20_24_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74014),
            .lcout(shift_srl_195Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93273),
            .ce(N__73977),
            .sr(_gnd_net_));
    defparam shift_srl_195_4_LC_20_24_4.C_ON=1'b0;
    defparam shift_srl_195_4_LC_20_24_4.SEQ_MODE=4'b1000;
    defparam shift_srl_195_4_LC_20_24_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_195_4_LC_20_24_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74008),
            .lcout(shift_srl_195Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93273),
            .ce(N__73977),
            .sr(_gnd_net_));
    defparam shift_srl_195_5_LC_20_24_5.C_ON=1'b0;
    defparam shift_srl_195_5_LC_20_24_5.SEQ_MODE=4'b1000;
    defparam shift_srl_195_5_LC_20_24_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_195_5_LC_20_24_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74002),
            .lcout(shift_srl_195Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93273),
            .ce(N__73977),
            .sr(_gnd_net_));
    defparam shift_srl_195_6_LC_20_24_6.C_ON=1'b0;
    defparam shift_srl_195_6_LC_20_24_6.SEQ_MODE=4'b1000;
    defparam shift_srl_195_6_LC_20_24_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_195_6_LC_20_24_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73996),
            .lcout(shift_srl_195Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93273),
            .ce(N__73977),
            .sr(_gnd_net_));
    defparam shift_srl_195_7_LC_20_24_7.C_ON=1'b0;
    defparam shift_srl_195_7_LC_20_24_7.SEQ_MODE=4'b1000;
    defparam shift_srl_195_7_LC_20_24_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_195_7_LC_20_24_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73990),
            .lcout(shift_srl_195Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93273),
            .ce(N__73977),
            .sr(_gnd_net_));
    defparam shift_srl_185_10_LC_20_25_0.C_ON=1'b0;
    defparam shift_srl_185_10_LC_20_25_0.SEQ_MODE=4'b1000;
    defparam shift_srl_185_10_LC_20_25_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_185_10_LC_20_25_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74074),
            .lcout(shift_srl_185Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93289),
            .ce(N__74056),
            .sr(_gnd_net_));
    defparam shift_srl_185_11_LC_20_25_1.C_ON=1'b0;
    defparam shift_srl_185_11_LC_20_25_1.SEQ_MODE=4'b1000;
    defparam shift_srl_185_11_LC_20_25_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_185_11_LC_20_25_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74104),
            .lcout(shift_srl_185Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93289),
            .ce(N__74056),
            .sr(_gnd_net_));
    defparam shift_srl_185_12_LC_20_25_2.C_ON=1'b0;
    defparam shift_srl_185_12_LC_20_25_2.SEQ_MODE=4'b1000;
    defparam shift_srl_185_12_LC_20_25_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_185_12_LC_20_25_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74098),
            .lcout(shift_srl_185Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93289),
            .ce(N__74056),
            .sr(_gnd_net_));
    defparam shift_srl_185_13_LC_20_25_3.C_ON=1'b0;
    defparam shift_srl_185_13_LC_20_25_3.SEQ_MODE=4'b1000;
    defparam shift_srl_185_13_LC_20_25_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_185_13_LC_20_25_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74092),
            .lcout(shift_srl_185Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93289),
            .ce(N__74056),
            .sr(_gnd_net_));
    defparam shift_srl_185_14_LC_20_25_4.C_ON=1'b0;
    defparam shift_srl_185_14_LC_20_25_4.SEQ_MODE=4'b1000;
    defparam shift_srl_185_14_LC_20_25_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_185_14_LC_20_25_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74086),
            .lcout(shift_srl_185Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93289),
            .ce(N__74056),
            .sr(_gnd_net_));
    defparam shift_srl_185_15_LC_20_25_5.C_ON=1'b0;
    defparam shift_srl_185_15_LC_20_25_5.SEQ_MODE=4'b1000;
    defparam shift_srl_185_15_LC_20_25_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_185_15_LC_20_25_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74080),
            .lcout(shift_srl_185Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93289),
            .ce(N__74056),
            .sr(_gnd_net_));
    defparam shift_srl_185_9_LC_20_25_6.C_ON=1'b0;
    defparam shift_srl_185_9_LC_20_25_6.SEQ_MODE=4'b1000;
    defparam shift_srl_185_9_LC_20_25_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_185_9_LC_20_25_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74062),
            .lcout(shift_srl_185Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93289),
            .ce(N__74056),
            .sr(_gnd_net_));
    defparam shift_srl_185_8_LC_20_25_7.C_ON=1'b0;
    defparam shift_srl_185_8_LC_20_25_7.SEQ_MODE=4'b1000;
    defparam shift_srl_185_8_LC_20_25_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_185_8_LC_20_25_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74068),
            .lcout(shift_srl_185Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93289),
            .ce(N__74056),
            .sr(_gnd_net_));
    defparam shift_srl_175_10_LC_20_26_0.C_ON=1'b0;
    defparam shift_srl_175_10_LC_20_26_0.SEQ_MODE=4'b1000;
    defparam shift_srl_175_10_LC_20_26_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_175_10_LC_20_26_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74146),
            .lcout(shift_srl_175Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93305),
            .ce(N__74125),
            .sr(_gnd_net_));
    defparam shift_srl_175_11_LC_20_26_1.C_ON=1'b0;
    defparam shift_srl_175_11_LC_20_26_1.SEQ_MODE=4'b1000;
    defparam shift_srl_175_11_LC_20_26_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_175_11_LC_20_26_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74176),
            .lcout(shift_srl_175Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93305),
            .ce(N__74125),
            .sr(_gnd_net_));
    defparam shift_srl_175_12_LC_20_26_2.C_ON=1'b0;
    defparam shift_srl_175_12_LC_20_26_2.SEQ_MODE=4'b1000;
    defparam shift_srl_175_12_LC_20_26_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_175_12_LC_20_26_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74170),
            .lcout(shift_srl_175Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93305),
            .ce(N__74125),
            .sr(_gnd_net_));
    defparam shift_srl_175_13_LC_20_26_3.C_ON=1'b0;
    defparam shift_srl_175_13_LC_20_26_3.SEQ_MODE=4'b1000;
    defparam shift_srl_175_13_LC_20_26_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_175_13_LC_20_26_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74164),
            .lcout(shift_srl_175Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93305),
            .ce(N__74125),
            .sr(_gnd_net_));
    defparam shift_srl_175_14_LC_20_26_4.C_ON=1'b0;
    defparam shift_srl_175_14_LC_20_26_4.SEQ_MODE=4'b1000;
    defparam shift_srl_175_14_LC_20_26_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_175_14_LC_20_26_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74158),
            .lcout(shift_srl_175Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93305),
            .ce(N__74125),
            .sr(_gnd_net_));
    defparam shift_srl_175_15_LC_20_26_5.C_ON=1'b0;
    defparam shift_srl_175_15_LC_20_26_5.SEQ_MODE=4'b1000;
    defparam shift_srl_175_15_LC_20_26_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_175_15_LC_20_26_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74152),
            .lcout(shift_srl_175Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93305),
            .ce(N__74125),
            .sr(_gnd_net_));
    defparam shift_srl_175_9_LC_20_26_6.C_ON=1'b0;
    defparam shift_srl_175_9_LC_20_26_6.SEQ_MODE=4'b1000;
    defparam shift_srl_175_9_LC_20_26_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_175_9_LC_20_26_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74131),
            .lcout(shift_srl_175Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93305),
            .ce(N__74125),
            .sr(_gnd_net_));
    defparam shift_srl_175_8_LC_20_26_7.C_ON=1'b0;
    defparam shift_srl_175_8_LC_20_26_7.SEQ_MODE=4'b1000;
    defparam shift_srl_175_8_LC_20_26_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_175_8_LC_20_26_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74140),
            .lcout(shift_srl_175Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93305),
            .ce(N__74125),
            .sr(_gnd_net_));
    defparam shift_srl_192_0_LC_20_27_0.C_ON=1'b0;
    defparam shift_srl_192_0_LC_20_27_0.SEQ_MODE=4'b1000;
    defparam shift_srl_192_0_LC_20_27_0.LUT_INIT=16'b1100110011001100;
    LogicCell40 shift_srl_192_0_LC_20_27_0 (
            .in0(_gnd_net_),
            .in1(N__74217),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_192Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93326),
            .ce(N__80673),
            .sr(_gnd_net_));
    defparam shift_srl_192_1_LC_20_27_1.C_ON=1'b0;
    defparam shift_srl_192_1_LC_20_27_1.SEQ_MODE=4'b1000;
    defparam shift_srl_192_1_LC_20_27_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_192_1_LC_20_27_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74110),
            .lcout(shift_srl_192Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93326),
            .ce(N__80673),
            .sr(_gnd_net_));
    defparam shift_srl_192_2_LC_20_27_2.C_ON=1'b0;
    defparam shift_srl_192_2_LC_20_27_2.SEQ_MODE=4'b1000;
    defparam shift_srl_192_2_LC_20_27_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_192_2_LC_20_27_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74296),
            .lcout(shift_srl_192Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93326),
            .ce(N__80673),
            .sr(_gnd_net_));
    defparam shift_srl_192_3_LC_20_27_3.C_ON=1'b0;
    defparam shift_srl_192_3_LC_20_27_3.SEQ_MODE=4'b1000;
    defparam shift_srl_192_3_LC_20_27_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_192_3_LC_20_27_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74290),
            .lcout(shift_srl_192Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93326),
            .ce(N__80673),
            .sr(_gnd_net_));
    defparam shift_srl_192_4_LC_20_27_4.C_ON=1'b0;
    defparam shift_srl_192_4_LC_20_27_4.SEQ_MODE=4'b1000;
    defparam shift_srl_192_4_LC_20_27_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_192_4_LC_20_27_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74284),
            .lcout(shift_srl_192Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93326),
            .ce(N__80673),
            .sr(_gnd_net_));
    defparam shift_srl_192_5_LC_20_27_5.C_ON=1'b0;
    defparam shift_srl_192_5_LC_20_27_5.SEQ_MODE=4'b1000;
    defparam shift_srl_192_5_LC_20_27_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_192_5_LC_20_27_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74278),
            .lcout(shift_srl_192Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93326),
            .ce(N__80673),
            .sr(_gnd_net_));
    defparam shift_srl_192_6_LC_20_27_6.C_ON=1'b0;
    defparam shift_srl_192_6_LC_20_27_6.SEQ_MODE=4'b1000;
    defparam shift_srl_192_6_LC_20_27_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_192_6_LC_20_27_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74272),
            .lcout(shift_srl_192Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93326),
            .ce(N__80673),
            .sr(_gnd_net_));
    defparam shift_srl_192_7_LC_20_27_7.C_ON=1'b0;
    defparam shift_srl_192_7_LC_20_27_7.SEQ_MODE=4'b1000;
    defparam shift_srl_192_7_LC_20_27_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_192_7_LC_20_27_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74266),
            .lcout(shift_srl_192Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93326),
            .ce(N__80673),
            .sr(_gnd_net_));
    defparam shift_srl_192_RNIV0MGG1_15_LC_20_28_0.C_ON=1'b0;
    defparam shift_srl_192_RNIV0MGG1_15_LC_20_28_0.SEQ_MODE=4'b0000;
    defparam shift_srl_192_RNIV0MGG1_15_LC_20_28_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_192_RNIV0MGG1_15_LC_20_28_0 (
            .in0(N__90473),
            .in1(N__74215),
            .in2(N__74258),
            .in3(N__91511),
            .lcout(clk_en_193),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_192_15_LC_20_28_1.C_ON=1'b0;
    defparam shift_srl_192_15_LC_20_28_1.SEQ_MODE=4'b1000;
    defparam shift_srl_192_15_LC_20_28_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_192_15_LC_20_28_1 (
            .in0(N__74182),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_192Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93348),
            .ce(N__80672),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_192_LC_20_28_2.C_ON=1'b0;
    defparam rco_obuf_RNO_192_LC_20_28_2.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_192_LC_20_28_2.LUT_INIT=16'b1000100000000000;
    LogicCell40 rco_obuf_RNO_192_LC_20_28_2 (
            .in0(N__74251),
            .in1(N__74216),
            .in2(_gnd_net_),
            .in3(N__91512),
            .lcout(rco_c_192),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_192_14_LC_20_28_3.C_ON=1'b0;
    defparam shift_srl_192_14_LC_20_28_3.SEQ_MODE=4'b1000;
    defparam shift_srl_192_14_LC_20_28_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_192_14_LC_20_28_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74350),
            .lcout(shift_srl_192Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93348),
            .ce(N__80672),
            .sr(_gnd_net_));
    defparam shift_srl_192_13_LC_20_28_4.C_ON=1'b0;
    defparam shift_srl_192_13_LC_20_28_4.SEQ_MODE=4'b1000;
    defparam shift_srl_192_13_LC_20_28_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_192_13_LC_20_28_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74344),
            .lcout(shift_srl_192Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93348),
            .ce(N__80672),
            .sr(_gnd_net_));
    defparam shift_srl_192_12_LC_20_28_5.C_ON=1'b0;
    defparam shift_srl_192_12_LC_20_28_5.SEQ_MODE=4'b1000;
    defparam shift_srl_192_12_LC_20_28_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_192_12_LC_20_28_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74338),
            .lcout(shift_srl_192Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93348),
            .ce(N__80672),
            .sr(_gnd_net_));
    defparam shift_srl_192_11_LC_20_28_6.C_ON=1'b0;
    defparam shift_srl_192_11_LC_20_28_6.SEQ_MODE=4'b1000;
    defparam shift_srl_192_11_LC_20_28_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_192_11_LC_20_28_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74332),
            .lcout(shift_srl_192Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93348),
            .ce(N__80672),
            .sr(_gnd_net_));
    defparam shift_srl_192_10_LC_20_28_7.C_ON=1'b0;
    defparam shift_srl_192_10_LC_20_28_7.SEQ_MODE=4'b1000;
    defparam shift_srl_192_10_LC_20_28_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_192_10_LC_20_28_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80689),
            .lcout(shift_srl_192Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93348),
            .ce(N__80672),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_46_LC_21_4_5.C_ON=1'b0;
    defparam rco_obuf_RNO_46_LC_21_4_5.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_46_LC_21_4_5.LUT_INIT=16'b1000100000000000;
    LogicCell40 rco_obuf_RNO_46_LC_21_4_5 (
            .in0(N__74383),
            .in1(N__76906),
            .in2(_gnd_net_),
            .in3(N__76209),
            .lcout(rco_c_46),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_50_14_LC_21_5_7.C_ON=1'b0;
    defparam shift_srl_50_14_LC_21_5_7.SEQ_MODE=4'b1000;
    defparam shift_srl_50_14_LC_21_5_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_50_14_LC_21_5_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74560),
            .lcout(shift_srl_50Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93384),
            .ce(N__76486),
            .sr(_gnd_net_));
    defparam shift_srl_49_0_LC_21_6_0.C_ON=1'b0;
    defparam shift_srl_49_0_LC_21_6_0.SEQ_MODE=4'b1000;
    defparam shift_srl_49_0_LC_21_6_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_49_0_LC_21_6_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__93491),
            .lcout(shift_srl_49Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93367),
            .ce(N__74408),
            .sr(_gnd_net_));
    defparam shift_srl_49_1_LC_21_6_1.C_ON=1'b0;
    defparam shift_srl_49_1_LC_21_6_1.SEQ_MODE=4'b1000;
    defparam shift_srl_49_1_LC_21_6_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_49_1_LC_21_6_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74308),
            .lcout(shift_srl_49Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93367),
            .ce(N__74408),
            .sr(_gnd_net_));
    defparam shift_srl_49_2_LC_21_6_2.C_ON=1'b0;
    defparam shift_srl_49_2_LC_21_6_2.SEQ_MODE=4'b1000;
    defparam shift_srl_49_2_LC_21_6_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_49_2_LC_21_6_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74302),
            .lcout(shift_srl_49Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93367),
            .ce(N__74408),
            .sr(_gnd_net_));
    defparam shift_srl_49_3_LC_21_6_3.C_ON=1'b0;
    defparam shift_srl_49_3_LC_21_6_3.SEQ_MODE=4'b1000;
    defparam shift_srl_49_3_LC_21_6_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_49_3_LC_21_6_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74533),
            .lcout(shift_srl_49Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93367),
            .ce(N__74408),
            .sr(_gnd_net_));
    defparam shift_srl_49_4_LC_21_6_4.C_ON=1'b0;
    defparam shift_srl_49_4_LC_21_6_4.SEQ_MODE=4'b1000;
    defparam shift_srl_49_4_LC_21_6_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_49_4_LC_21_6_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74527),
            .lcout(shift_srl_49Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93367),
            .ce(N__74408),
            .sr(_gnd_net_));
    defparam shift_srl_49_5_LC_21_6_5.C_ON=1'b0;
    defparam shift_srl_49_5_LC_21_6_5.SEQ_MODE=4'b1000;
    defparam shift_srl_49_5_LC_21_6_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_49_5_LC_21_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74521),
            .lcout(shift_srl_49Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93367),
            .ce(N__74408),
            .sr(_gnd_net_));
    defparam shift_srl_49_6_LC_21_6_6.C_ON=1'b0;
    defparam shift_srl_49_6_LC_21_6_6.SEQ_MODE=4'b1000;
    defparam shift_srl_49_6_LC_21_6_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_49_6_LC_21_6_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74515),
            .lcout(shift_srl_49Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93367),
            .ce(N__74408),
            .sr(_gnd_net_));
    defparam shift_srl_41_RNIG75KB_15_LC_21_7_1.C_ON=1'b0;
    defparam shift_srl_41_RNIG75KB_15_LC_21_7_1.SEQ_MODE=4'b0000;
    defparam shift_srl_41_RNIG75KB_15_LC_21_7_1.LUT_INIT=16'b0000110000000000;
    LogicCell40 shift_srl_41_RNIG75KB_15_LC_21_7_1 (
            .in0(_gnd_net_),
            .in1(N__85195),
            .in2(N__85267),
            .in3(N__74500),
            .lcout(rco_c_44),
            .ltout(rco_c_44_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_46_RNIKSAVB_15_LC_21_7_2.C_ON=1'b0;
    defparam shift_srl_46_RNIKSAVB_15_LC_21_7_2.SEQ_MODE=4'b0000;
    defparam shift_srl_46_RNIKSAVB_15_LC_21_7_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_46_RNIKSAVB_15_LC_21_7_2 (
            .in0(N__76202),
            .in1(N__90224),
            .in2(N__74503),
            .in3(N__74382),
            .lcout(clk_en_47),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_48_RNII2GM4_15_LC_21_7_3.C_ON=1'b0;
    defparam shift_srl_48_RNII2GM4_15_LC_21_7_3.SEQ_MODE=4'b0000;
    defparam shift_srl_48_RNII2GM4_15_LC_21_7_3.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_48_RNII2GM4_15_LC_21_7_3 (
            .in0(N__76618),
            .in1(N__74499),
            .in2(N__90432),
            .in3(N__76832),
            .lcout(),
            .ltout(clk_en_0_a3_0_a2_sx_49_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_48_RNI1MEQC_15_LC_21_7_4.C_ON=1'b0;
    defparam shift_srl_48_RNI1MEQC_15_LC_21_7_4.SEQ_MODE=4'b0000;
    defparam shift_srl_48_RNI1MEQC_15_LC_21_7_4.LUT_INIT=16'b0000001000000010;
    LogicCell40 shift_srl_48_RNI1MEQC_15_LC_21_7_4 (
            .in0(N__85196),
            .in1(N__85261),
            .in2(N__74434),
            .in3(_gnd_net_),
            .lcout(clk_en_49),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_47_RNIV3QL_15_LC_21_7_6.C_ON=1'b0;
    defparam shift_srl_47_RNIV3QL_15_LC_21_7_6.SEQ_MODE=4'b0000;
    defparam shift_srl_47_RNIV3QL_15_LC_21_7_6.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_47_RNIV3QL_15_LC_21_7_6 (
            .in0(N__76201),
            .in1(N__76320),
            .in2(_gnd_net_),
            .in3(N__74381),
            .lcout(shift_srl_47_RNIV3QLZ0Z_15),
            .ltout(shift_srl_47_RNIV3QLZ0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_47_LC_21_7_7.C_ON=1'b0;
    defparam rco_obuf_RNO_47_LC_21_7_7.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_47_LC_21_7_7.LUT_INIT=16'b1010000010100000;
    LogicCell40 rco_obuf_RNO_47_LC_21_7_7 (
            .in0(N__76893),
            .in1(_gnd_net_),
            .in2(N__74602),
            .in3(_gnd_net_),
            .lcout(rco_c_47),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_50_11_LC_21_8_0.C_ON=1'b0;
    defparam shift_srl_50_11_LC_21_8_0.SEQ_MODE=4'b1000;
    defparam shift_srl_50_11_LC_21_8_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_50_11_LC_21_8_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76387),
            .lcout(shift_srl_50Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93329),
            .ce(N__76482),
            .sr(_gnd_net_));
    defparam shift_srl_50_15_LC_21_8_1.C_ON=1'b0;
    defparam shift_srl_50_15_LC_21_8_1.SEQ_MODE=4'b1000;
    defparam shift_srl_50_15_LC_21_8_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_50_15_LC_21_8_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74581),
            .lcout(shift_srl_50Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93329),
            .ce(N__76482),
            .sr(_gnd_net_));
    defparam shift_srl_50_12_LC_21_8_3.C_ON=1'b0;
    defparam shift_srl_50_12_LC_21_8_3.SEQ_MODE=4'b1000;
    defparam shift_srl_50_12_LC_21_8_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_50_12_LC_21_8_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74572),
            .lcout(shift_srl_50Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93329),
            .ce(N__76482),
            .sr(_gnd_net_));
    defparam shift_srl_50_13_LC_21_8_5.C_ON=1'b0;
    defparam shift_srl_50_13_LC_21_8_5.SEQ_MODE=4'b1000;
    defparam shift_srl_50_13_LC_21_8_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_50_13_LC_21_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74566),
            .lcout(shift_srl_50Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93329),
            .ce(N__76482),
            .sr(_gnd_net_));
    defparam shift_srl_52_10_LC_21_9_0.C_ON=1'b0;
    defparam shift_srl_52_10_LC_21_9_0.SEQ_MODE=4'b1000;
    defparam shift_srl_52_10_LC_21_9_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_52_10_LC_21_9_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74818),
            .lcout(shift_srl_52Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93308),
            .ce(N__76689),
            .sr(_gnd_net_));
    defparam shift_srl_52_11_LC_21_9_1.C_ON=1'b0;
    defparam shift_srl_52_11_LC_21_9_1.SEQ_MODE=4'b1000;
    defparam shift_srl_52_11_LC_21_9_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_52_11_LC_21_9_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74551),
            .lcout(shift_srl_52Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93308),
            .ce(N__76689),
            .sr(_gnd_net_));
    defparam shift_srl_52_12_LC_21_9_2.C_ON=1'b0;
    defparam shift_srl_52_12_LC_21_9_2.SEQ_MODE=4'b1000;
    defparam shift_srl_52_12_LC_21_9_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_52_12_LC_21_9_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74545),
            .lcout(shift_srl_52Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93308),
            .ce(N__76689),
            .sr(_gnd_net_));
    defparam shift_srl_52_13_LC_21_9_3.C_ON=1'b0;
    defparam shift_srl_52_13_LC_21_9_3.SEQ_MODE=4'b1000;
    defparam shift_srl_52_13_LC_21_9_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_52_13_LC_21_9_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74539),
            .lcout(shift_srl_52Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93308),
            .ce(N__76689),
            .sr(_gnd_net_));
    defparam shift_srl_52_14_LC_21_9_4.C_ON=1'b0;
    defparam shift_srl_52_14_LC_21_9_4.SEQ_MODE=4'b1000;
    defparam shift_srl_52_14_LC_21_9_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_52_14_LC_21_9_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74830),
            .lcout(shift_srl_52Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93308),
            .ce(N__76689),
            .sr(_gnd_net_));
    defparam shift_srl_52_15_LC_21_9_5.C_ON=1'b0;
    defparam shift_srl_52_15_LC_21_9_5.SEQ_MODE=4'b1000;
    defparam shift_srl_52_15_LC_21_9_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_52_15_LC_21_9_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74824),
            .lcout(shift_srl_52Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93308),
            .ce(N__76689),
            .sr(_gnd_net_));
    defparam shift_srl_52_9_LC_21_9_6.C_ON=1'b0;
    defparam shift_srl_52_9_LC_21_9_6.SEQ_MODE=4'b1000;
    defparam shift_srl_52_9_LC_21_9_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_52_9_LC_21_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74812),
            .lcout(shift_srl_52Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93308),
            .ce(N__76689),
            .sr(_gnd_net_));
    defparam shift_srl_52_8_LC_21_9_7.C_ON=1'b0;
    defparam shift_srl_52_8_LC_21_9_7.SEQ_MODE=4'b1000;
    defparam shift_srl_52_8_LC_21_9_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_52_8_LC_21_9_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76696),
            .lcout(shift_srl_52Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93308),
            .ce(N__76689),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_52_LC_21_10_0.C_ON=1'b0;
    defparam rco_obuf_RNO_52_LC_21_10_0.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_52_LC_21_10_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 rco_obuf_RNO_52_LC_21_10_0 (
            .in0(N__74638),
            .in1(N__88325),
            .in2(N__93576),
            .in3(N__76449),
            .lcout(rco_c_52),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_51_LC_21_10_1.C_ON=1'b0;
    defparam rco_obuf_RNO_51_LC_21_10_1.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_51_LC_21_10_1.LUT_INIT=16'b1000100000000000;
    LogicCell40 rco_obuf_RNO_51_LC_21_10_1 (
            .in0(N__88324),
            .in1(N__93557),
            .in2(_gnd_net_),
            .in3(N__74637),
            .lcout(rco_c_51),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_41_RNI2OCV1_15_LC_21_10_2.C_ON=1'b0;
    defparam shift_srl_41_RNI2OCV1_15_LC_21_10_2.SEQ_MODE=4'b0000;
    defparam shift_srl_41_RNI2OCV1_15_LC_21_10_2.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_41_RNI2OCV1_15_LC_21_10_2 (
            .in0(N__74741),
            .in1(N__75137),
            .in2(N__74716),
            .in3(N__78793),
            .lcout(rco_int_0_a2_1_a2_sx_44),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_51_RNIQ3CJD_15_LC_21_10_3.C_ON=1'b0;
    defparam shift_srl_51_RNIQ3CJD_15_LC_21_10_3.SEQ_MODE=4'b0000;
    defparam shift_srl_51_RNIQ3CJD_15_LC_21_10_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_51_RNIQ3CJD_15_LC_21_10_3 (
            .in0(N__90226),
            .in1(N__93556),
            .in2(N__88329),
            .in3(N__74636),
            .lcout(clk_en_52),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNI8AQFE_15_LC_21_10_4.C_ON=1'b0;
    defparam shift_srl_0_RNI8AQFE_15_LC_21_10_4.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNI8AQFE_15_LC_21_10_4.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNI8AQFE_15_LC_21_10_4 (
            .in0(N__93555),
            .in1(N__76928),
            .in2(N__90433),
            .in3(N__81532),
            .lcout(clk_en_56),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNI6HAFF_15_LC_21_10_5.C_ON=1'b0;
    defparam shift_srl_0_RNI6HAFF_15_LC_21_10_5.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNI6HAFF_15_LC_21_10_5.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_0_RNI6HAFF_15_LC_21_10_5 (
            .in0(N__90225),
            .in1(N__81440),
            .in2(_gnd_net_),
            .in3(N__93554),
            .lcout(clk_en_60),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_48_RNI6AKPC_15_LC_21_10_6.C_ON=1'b0;
    defparam shift_srl_48_RNI6AKPC_15_LC_21_10_6.SEQ_MODE=4'b0000;
    defparam shift_srl_48_RNI6AKPC_15_LC_21_10_6.LUT_INIT=16'b0000100000000000;
    LogicCell40 shift_srl_48_RNI6AKPC_15_LC_21_10_6 (
            .in0(N__76613),
            .in1(N__75136),
            .in2(N__81363),
            .in3(N__81323),
            .lcout(rco_c_48),
            .ltout(rco_c_48_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_59_RNI6SV1J_15_LC_21_10_7.C_ON=1'b0;
    defparam shift_srl_59_RNI6SV1J_15_LC_21_10_7.SEQ_MODE=4'b0000;
    defparam shift_srl_59_RNI6SV1J_15_LC_21_10_7.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_59_RNI6SV1J_15_LC_21_10_7 (
            .in0(N__86815),
            .in1(N__81441),
            .in2(N__74905),
            .in3(N__84999),
            .lcout(rco_c_74),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_54_RNIJID2E_15_LC_21_11_0.C_ON=1'b0;
    defparam shift_srl_54_RNIJID2E_15_LC_21_11_0.SEQ_MODE=4'b0000;
    defparam shift_srl_54_RNIJID2E_15_LC_21_11_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_54_RNIJID2E_15_LC_21_11_0 (
            .in0(N__93566),
            .in1(N__77006),
            .in2(N__90285),
            .in3(N__81539),
            .lcout(clk_en_55),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_54_15_LC_21_11_1.C_ON=1'b0;
    defparam shift_srl_54_15_LC_21_11_1.SEQ_MODE=4'b1000;
    defparam shift_srl_54_15_LC_21_11_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_54_15_LC_21_11_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74854),
            .lcout(shift_srl_54Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93274),
            .ce(N__87170),
            .sr(_gnd_net_));
    defparam shift_srl_55_RNI9BJM_15_LC_21_11_2.C_ON=1'b0;
    defparam shift_srl_55_RNI9BJM_15_LC_21_11_2.SEQ_MODE=4'b0000;
    defparam shift_srl_55_RNI9BJM_15_LC_21_11_2.LUT_INIT=16'b1100110000000000;
    LogicCell40 shift_srl_55_RNI9BJM_15_LC_21_11_2 (
            .in0(_gnd_net_),
            .in1(N__77005),
            .in2(_gnd_net_),
            .in3(N__74873),
            .lcout(shift_srl_55_RNI9BJMZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_54_14_LC_21_11_3.C_ON=1'b0;
    defparam shift_srl_54_14_LC_21_11_3.SEQ_MODE=4'b1000;
    defparam shift_srl_54_14_LC_21_11_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_54_14_LC_21_11_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74848),
            .lcout(shift_srl_54Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93274),
            .ce(N__87170),
            .sr(_gnd_net_));
    defparam shift_srl_54_13_LC_21_11_4.C_ON=1'b0;
    defparam shift_srl_54_13_LC_21_11_4.SEQ_MODE=4'b1000;
    defparam shift_srl_54_13_LC_21_11_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_54_13_LC_21_11_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74842),
            .lcout(shift_srl_54Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93274),
            .ce(N__87170),
            .sr(_gnd_net_));
    defparam shift_srl_54_12_LC_21_11_5.C_ON=1'b0;
    defparam shift_srl_54_12_LC_21_11_5.SEQ_MODE=4'b1000;
    defparam shift_srl_54_12_LC_21_11_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_54_12_LC_21_11_5 (
            .in0(N__74836),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_54Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93274),
            .ce(N__87170),
            .sr(_gnd_net_));
    defparam shift_srl_54_11_LC_21_11_6.C_ON=1'b0;
    defparam shift_srl_54_11_LC_21_11_6.SEQ_MODE=4'b1000;
    defparam shift_srl_54_11_LC_21_11_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_54_11_LC_21_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74953),
            .lcout(shift_srl_54Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93274),
            .ce(N__87170),
            .sr(_gnd_net_));
    defparam shift_srl_54_10_LC_21_11_7.C_ON=1'b0;
    defparam shift_srl_54_10_LC_21_11_7.SEQ_MODE=4'b1000;
    defparam shift_srl_54_10_LC_21_11_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_54_10_LC_21_11_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87202),
            .lcout(shift_srl_54Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93274),
            .ce(N__87170),
            .sr(_gnd_net_));
    defparam shift_srl_57_10_LC_21_12_0.C_ON=1'b0;
    defparam shift_srl_57_10_LC_21_12_0.SEQ_MODE=4'b1000;
    defparam shift_srl_57_10_LC_21_12_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_57_10_LC_21_12_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74917),
            .lcout(shift_srl_57Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93255),
            .ce(N__76726),
            .sr(_gnd_net_));
    defparam shift_srl_57_11_LC_21_12_1.C_ON=1'b0;
    defparam shift_srl_57_11_LC_21_12_1.SEQ_MODE=4'b1000;
    defparam shift_srl_57_11_LC_21_12_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_57_11_LC_21_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74947),
            .lcout(shift_srl_57Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93255),
            .ce(N__76726),
            .sr(_gnd_net_));
    defparam shift_srl_57_12_LC_21_12_2.C_ON=1'b0;
    defparam shift_srl_57_12_LC_21_12_2.SEQ_MODE=4'b1000;
    defparam shift_srl_57_12_LC_21_12_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_57_12_LC_21_12_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74941),
            .lcout(shift_srl_57Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93255),
            .ce(N__76726),
            .sr(_gnd_net_));
    defparam shift_srl_57_13_LC_21_12_3.C_ON=1'b0;
    defparam shift_srl_57_13_LC_21_12_3.SEQ_MODE=4'b1000;
    defparam shift_srl_57_13_LC_21_12_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_57_13_LC_21_12_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74935),
            .lcout(shift_srl_57Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93255),
            .ce(N__76726),
            .sr(_gnd_net_));
    defparam shift_srl_57_14_LC_21_12_4.C_ON=1'b0;
    defparam shift_srl_57_14_LC_21_12_4.SEQ_MODE=4'b1000;
    defparam shift_srl_57_14_LC_21_12_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_57_14_LC_21_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74929),
            .lcout(shift_srl_57Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93255),
            .ce(N__76726),
            .sr(_gnd_net_));
    defparam shift_srl_57_15_LC_21_12_5.C_ON=1'b0;
    defparam shift_srl_57_15_LC_21_12_5.SEQ_MODE=4'b1000;
    defparam shift_srl_57_15_LC_21_12_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_57_15_LC_21_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74923),
            .lcout(shift_srl_57Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93255),
            .ce(N__76726),
            .sr(_gnd_net_));
    defparam shift_srl_57_9_LC_21_12_6.C_ON=1'b0;
    defparam shift_srl_57_9_LC_21_12_6.SEQ_MODE=4'b1000;
    defparam shift_srl_57_9_LC_21_12_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_57_9_LC_21_12_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74911),
            .lcout(shift_srl_57Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93255),
            .ce(N__76726),
            .sr(_gnd_net_));
    defparam shift_srl_57_8_LC_21_12_7.C_ON=1'b0;
    defparam shift_srl_57_8_LC_21_12_7.SEQ_MODE=4'b1000;
    defparam shift_srl_57_8_LC_21_12_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_57_8_LC_21_12_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76732),
            .lcout(shift_srl_57Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93255),
            .ce(N__76726),
            .sr(_gnd_net_));
    defparam shift_srl_60_10_LC_21_13_0.C_ON=1'b0;
    defparam shift_srl_60_10_LC_21_13_0.SEQ_MODE=4'b1000;
    defparam shift_srl_60_10_LC_21_13_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_60_10_LC_21_13_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74971),
            .lcout(shift_srl_60Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93233),
            .ce(N__79080),
            .sr(_gnd_net_));
    defparam shift_srl_60_11_LC_21_13_1.C_ON=1'b0;
    defparam shift_srl_60_11_LC_21_13_1.SEQ_MODE=4'b1000;
    defparam shift_srl_60_11_LC_21_13_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_60_11_LC_21_13_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74995),
            .lcout(shift_srl_60Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93233),
            .ce(N__79080),
            .sr(_gnd_net_));
    defparam shift_srl_60_12_LC_21_13_2.C_ON=1'b0;
    defparam shift_srl_60_12_LC_21_13_2.SEQ_MODE=4'b1000;
    defparam shift_srl_60_12_LC_21_13_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_60_12_LC_21_13_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74989),
            .lcout(shift_srl_60Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93233),
            .ce(N__79080),
            .sr(_gnd_net_));
    defparam shift_srl_60_13_LC_21_13_3.C_ON=1'b0;
    defparam shift_srl_60_13_LC_21_13_3.SEQ_MODE=4'b1000;
    defparam shift_srl_60_13_LC_21_13_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_60_13_LC_21_13_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74983),
            .lcout(shift_srl_60Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93233),
            .ce(N__79080),
            .sr(_gnd_net_));
    defparam shift_srl_60_14_LC_21_13_4.C_ON=1'b0;
    defparam shift_srl_60_14_LC_21_13_4.SEQ_MODE=4'b1000;
    defparam shift_srl_60_14_LC_21_13_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_60_14_LC_21_13_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74977),
            .lcout(shift_srl_60Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93233),
            .ce(N__79080),
            .sr(_gnd_net_));
    defparam shift_srl_60_9_LC_21_13_5.C_ON=1'b0;
    defparam shift_srl_60_9_LC_21_13_5.SEQ_MODE=4'b1000;
    defparam shift_srl_60_9_LC_21_13_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_60_9_LC_21_13_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74965),
            .lcout(shift_srl_60Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93233),
            .ce(N__79080),
            .sr(_gnd_net_));
    defparam shift_srl_60_8_LC_21_13_6.C_ON=1'b0;
    defparam shift_srl_60_8_LC_21_13_6.SEQ_MODE=4'b1000;
    defparam shift_srl_60_8_LC_21_13_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_60_8_LC_21_13_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75193),
            .lcout(shift_srl_60Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93233),
            .ce(N__79080),
            .sr(_gnd_net_));
    defparam shift_srl_60_15_LC_21_13_7.C_ON=1'b0;
    defparam shift_srl_60_15_LC_21_13_7.SEQ_MODE=4'b1000;
    defparam shift_srl_60_15_LC_21_13_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_60_15_LC_21_13_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74959),
            .lcout(shift_srl_60Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93233),
            .ce(N__79080),
            .sr(_gnd_net_));
    defparam shift_srl_60_4_LC_21_14_0.C_ON=1'b0;
    defparam shift_srl_60_4_LC_21_14_0.SEQ_MODE=4'b1000;
    defparam shift_srl_60_4_LC_21_14_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_60_4_LC_21_14_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75286),
            .lcout(shift_srl_60Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93215),
            .ce(N__79075),
            .sr(_gnd_net_));
    defparam shift_srl_60_5_LC_21_14_1.C_ON=1'b0;
    defparam shift_srl_60_5_LC_21_14_1.SEQ_MODE=4'b1000;
    defparam shift_srl_60_5_LC_21_14_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_60_5_LC_21_14_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75211),
            .lcout(shift_srl_60Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93215),
            .ce(N__79075),
            .sr(_gnd_net_));
    defparam shift_srl_60_6_LC_21_14_2.C_ON=1'b0;
    defparam shift_srl_60_6_LC_21_14_2.SEQ_MODE=4'b1000;
    defparam shift_srl_60_6_LC_21_14_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_60_6_LC_21_14_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75205),
            .lcout(shift_srl_60Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93215),
            .ce(N__79075),
            .sr(_gnd_net_));
    defparam shift_srl_60_7_LC_21_14_5.C_ON=1'b0;
    defparam shift_srl_60_7_LC_21_14_5.SEQ_MODE=4'b1000;
    defparam shift_srl_60_7_LC_21_14_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_60_7_LC_21_14_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75199),
            .lcout(shift_srl_60Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93215),
            .ce(N__79075),
            .sr(_gnd_net_));
    defparam shift_srl_178_RNI8L486_15_LC_21_15_2.C_ON=1'b0;
    defparam shift_srl_178_RNI8L486_15_LC_21_15_2.SEQ_MODE=4'b0000;
    defparam shift_srl_178_RNI8L486_15_LC_21_15_2.LUT_INIT=16'b1111111101111111;
    LogicCell40 shift_srl_178_RNI8L486_15_LC_21_15_2 (
            .in0(N__80415),
            .in1(N__80476),
            .in2(N__80539),
            .in3(N__84154),
            .lcout(),
            .ltout(clk_en_0_a3_0_a2_sx_179_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_178_RNICD71D1_15_LC_21_15_3.C_ON=1'b0;
    defparam shift_srl_178_RNICD71D1_15_LC_21_15_3.SEQ_MODE=4'b0000;
    defparam shift_srl_178_RNICD71D1_15_LC_21_15_3.LUT_INIT=16'b0000010000000000;
    LogicCell40 shift_srl_178_RNICD71D1_15_LC_21_15_3 (
            .in0(N__75187),
            .in1(N__77830),
            .in2(N__75160),
            .in3(N__75035),
            .lcout(clk_en_179),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_59_RNISPG43_15_LC_21_15_4.C_ON=1'b0;
    defparam shift_srl_59_RNISPG43_15_LC_21_15_4.SEQ_MODE=4'b0000;
    defparam shift_srl_59_RNISPG43_15_LC_21_15_4.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_59_RNISPG43_15_LC_21_15_4 (
            .in0(N__81588),
            .in1(N__76601),
            .in2(N__81489),
            .in3(N__81549),
            .lcout(),
            .ltout(rco_int_0_a2_0_a2_93_m6_0_a2_4_7_4_sx_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_40_fast_RNIKUQC5_15_LC_21_15_5.C_ON=1'b0;
    defparam shift_srl_40_fast_RNIKUQC5_15_LC_21_15_5.SEQ_MODE=4'b0000;
    defparam shift_srl_40_fast_RNIKUQC5_15_LC_21_15_5.LUT_INIT=16'b0000100000000000;
    LogicCell40 shift_srl_40_fast_RNIKUQC5_15_LC_21_15_5 (
            .in0(N__75157),
            .in1(N__75145),
            .in2(N__75097),
            .in3(N__76854),
            .lcout(),
            .ltout(rco_int_0_a2_0_a2_93_m6_0_a2_4_7_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_83_RNIU84BB_15_LC_21_15_6.C_ON=1'b0;
    defparam shift_srl_83_RNIU84BB_15_LC_21_15_6.SEQ_MODE=4'b0000;
    defparam shift_srl_83_RNIU84BB_15_LC_21_15_6.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_83_RNIU84BB_15_LC_21_15_6 (
            .in0(N__86811),
            .in1(N__84951),
            .in2(N__75094),
            .in3(N__80775),
            .lcout(rco_int_0_a2_0_a2_93_m6_0_a2_4_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_66_RNIDTJJ_15_LC_21_15_7.C_ON=1'b0;
    defparam shift_srl_66_RNIDTJJ_15_LC_21_15_7.SEQ_MODE=4'b0000;
    defparam shift_srl_66_RNIDTJJ_15_LC_21_15_7.LUT_INIT=16'b1100110000000000;
    LogicCell40 shift_srl_66_RNIDTJJ_15_LC_21_15_7 (
            .in0(_gnd_net_),
            .in1(N__81721),
            .in2(_gnd_net_),
            .in3(N__80990),
            .lcout(rco_int_0_a3_0_a2_0_0_66),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_63_0_LC_21_16_0.C_ON=1'b0;
    defparam shift_srl_63_0_LC_21_16_0.SEQ_MODE=4'b1000;
    defparam shift_srl_63_0_LC_21_16_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_63_0_LC_21_16_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81138),
            .lcout(shift_srl_63Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93174),
            .ce(N__79184),
            .sr(_gnd_net_));
    defparam shift_srl_63_1_LC_21_16_1.C_ON=1'b0;
    defparam shift_srl_63_1_LC_21_16_1.SEQ_MODE=4'b1000;
    defparam shift_srl_63_1_LC_21_16_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_63_1_LC_21_16_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75277),
            .lcout(shift_srl_63Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93174),
            .ce(N__79184),
            .sr(_gnd_net_));
    defparam shift_srl_63_2_LC_21_16_2.C_ON=1'b0;
    defparam shift_srl_63_2_LC_21_16_2.SEQ_MODE=4'b1000;
    defparam shift_srl_63_2_LC_21_16_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_63_2_LC_21_16_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75271),
            .lcout(shift_srl_63Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93174),
            .ce(N__79184),
            .sr(_gnd_net_));
    defparam shift_srl_63_3_LC_21_16_3.C_ON=1'b0;
    defparam shift_srl_63_3_LC_21_16_3.SEQ_MODE=4'b1000;
    defparam shift_srl_63_3_LC_21_16_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_63_3_LC_21_16_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75265),
            .lcout(shift_srl_63Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93174),
            .ce(N__79184),
            .sr(_gnd_net_));
    defparam shift_srl_63_4_LC_21_16_4.C_ON=1'b0;
    defparam shift_srl_63_4_LC_21_16_4.SEQ_MODE=4'b1000;
    defparam shift_srl_63_4_LC_21_16_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_63_4_LC_21_16_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75259),
            .lcout(shift_srl_63Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93174),
            .ce(N__79184),
            .sr(_gnd_net_));
    defparam shift_srl_63_5_LC_21_16_5.C_ON=1'b0;
    defparam shift_srl_63_5_LC_21_16_5.SEQ_MODE=4'b1000;
    defparam shift_srl_63_5_LC_21_16_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_63_5_LC_21_16_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75253),
            .lcout(shift_srl_63Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93174),
            .ce(N__79184),
            .sr(_gnd_net_));
    defparam shift_srl_63_6_LC_21_16_6.C_ON=1'b0;
    defparam shift_srl_63_6_LC_21_16_6.SEQ_MODE=4'b1000;
    defparam shift_srl_63_6_LC_21_16_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_63_6_LC_21_16_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75247),
            .lcout(shift_srl_63Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93174),
            .ce(N__79184),
            .sr(_gnd_net_));
    defparam shift_srl_63_7_LC_21_16_7.C_ON=1'b0;
    defparam shift_srl_63_7_LC_21_16_7.SEQ_MODE=4'b1000;
    defparam shift_srl_63_7_LC_21_16_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_63_7_LC_21_16_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75241),
            .lcout(shift_srl_63Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93174),
            .ce(N__79184),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_60_LC_21_17_0.C_ON=1'b0;
    defparam rco_obuf_RNO_60_LC_21_17_0.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_60_LC_21_17_0.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_60_LC_21_17_0 (
            .in0(N__75334),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84922),
            .lcout(rco_c_60),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_61_LC_21_17_1.C_ON=1'b0;
    defparam rco_obuf_RNO_61_LC_21_17_1.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_61_LC_21_17_1.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_61_LC_21_17_1 (
            .in0(N__84923),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75217),
            .lcout(rco_c_61),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_62_LC_21_17_2.C_ON=1'b0;
    defparam rco_obuf_RNO_62_LC_21_17_2.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_62_LC_21_17_2.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_62_LC_21_17_2 (
            .in0(N__81028),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84924),
            .lcout(rco_c_62),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_65_LC_21_17_3.C_ON=1'b0;
    defparam rco_obuf_RNO_65_LC_21_17_3.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_65_LC_21_17_3.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_65_LC_21_17_3 (
            .in0(N__84925),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80974),
            .lcout(rco_c_65),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_60_0_LC_21_17_4.C_ON=1'b0;
    defparam shift_srl_60_0_LC_21_17_4.SEQ_MODE=4'b1000;
    defparam shift_srl_60_0_LC_21_17_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_60_0_LC_21_17_4 (
            .in0(N__75333),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_60Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93136),
            .ce(N__79081),
            .sr(_gnd_net_));
    defparam shift_srl_60_1_LC_21_17_5.C_ON=1'b0;
    defparam shift_srl_60_1_LC_21_17_5.SEQ_MODE=4'b1000;
    defparam shift_srl_60_1_LC_21_17_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_60_1_LC_21_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75304),
            .lcout(shift_srl_60Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93136),
            .ce(N__79081),
            .sr(_gnd_net_));
    defparam shift_srl_60_2_LC_21_17_6.C_ON=1'b0;
    defparam shift_srl_60_2_LC_21_17_6.SEQ_MODE=4'b1000;
    defparam shift_srl_60_2_LC_21_17_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_60_2_LC_21_17_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75298),
            .lcout(shift_srl_60Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93136),
            .ce(N__79081),
            .sr(_gnd_net_));
    defparam shift_srl_60_3_LC_21_17_7.C_ON=1'b0;
    defparam shift_srl_60_3_LC_21_17_7.SEQ_MODE=4'b1000;
    defparam shift_srl_60_3_LC_21_17_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_60_3_LC_21_17_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75292),
            .lcout(shift_srl_60Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93136),
            .ce(N__79081),
            .sr(_gnd_net_));
    defparam shift_srl_159_11_LC_21_18_0.C_ON=1'b0;
    defparam shift_srl_159_11_LC_21_18_0.SEQ_MODE=4'b1000;
    defparam shift_srl_159_11_LC_21_18_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_159_11_LC_21_18_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75442),
            .lcout(shift_srl_159Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93175),
            .ce(N__77707),
            .sr(_gnd_net_));
    defparam shift_srl_159_13_LC_21_18_1.C_ON=1'b0;
    defparam shift_srl_159_13_LC_21_18_1.SEQ_MODE=4'b1000;
    defparam shift_srl_159_13_LC_21_18_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_159_13_LC_21_18_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75424),
            .lcout(shift_srl_159Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93175),
            .ce(N__77707),
            .sr(_gnd_net_));
    defparam shift_srl_159_5_LC_21_18_2.C_ON=1'b0;
    defparam shift_srl_159_5_LC_21_18_2.SEQ_MODE=4'b1000;
    defparam shift_srl_159_5_LC_21_18_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_159_5_LC_21_18_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75496),
            .lcout(shift_srl_159Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93175),
            .ce(N__77707),
            .sr(_gnd_net_));
    defparam shift_srl_159_10_LC_21_18_3.C_ON=1'b0;
    defparam shift_srl_159_10_LC_21_18_3.SEQ_MODE=4'b1000;
    defparam shift_srl_159_10_LC_21_18_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_159_10_LC_21_18_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75436),
            .lcout(shift_srl_159Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93175),
            .ce(N__77707),
            .sr(_gnd_net_));
    defparam shift_srl_159_9_LC_21_18_4.C_ON=1'b0;
    defparam shift_srl_159_9_LC_21_18_4.SEQ_MODE=4'b1000;
    defparam shift_srl_159_9_LC_21_18_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_159_9_LC_21_18_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75484),
            .lcout(shift_srl_159Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93175),
            .ce(N__77707),
            .sr(_gnd_net_));
    defparam shift_srl_159_12_LC_21_18_5.C_ON=1'b0;
    defparam shift_srl_159_12_LC_21_18_5.SEQ_MODE=4'b1000;
    defparam shift_srl_159_12_LC_21_18_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_159_12_LC_21_18_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75430),
            .lcout(shift_srl_159Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93175),
            .ce(N__77707),
            .sr(_gnd_net_));
    defparam shift_srl_159_6_LC_21_18_6.C_ON=1'b0;
    defparam shift_srl_159_6_LC_21_18_6.SEQ_MODE=4'b1000;
    defparam shift_srl_159_6_LC_21_18_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_159_6_LC_21_18_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75418),
            .lcout(shift_srl_159Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93175),
            .ce(N__77707),
            .sr(_gnd_net_));
    defparam shift_srl_159_14_LC_21_18_7.C_ON=1'b0;
    defparam shift_srl_159_14_LC_21_18_7.SEQ_MODE=4'b1000;
    defparam shift_srl_159_14_LC_21_18_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_159_14_LC_21_18_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75412),
            .lcout(shift_srl_159Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93175),
            .ce(N__77707),
            .sr(_gnd_net_));
    defparam shift_srl_159_3_LC_21_19_0.C_ON=1'b0;
    defparam shift_srl_159_3_LC_21_19_0.SEQ_MODE=4'b1000;
    defparam shift_srl_159_3_LC_21_19_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_159_3_LC_21_19_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75472),
            .lcout(shift_srl_159Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93195),
            .ce(N__77702),
            .sr(_gnd_net_));
    defparam shift_srl_159_0_LC_21_19_2.C_ON=1'b0;
    defparam shift_srl_159_0_LC_21_19_2.SEQ_MODE=4'b1000;
    defparam shift_srl_159_0_LC_21_19_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_159_0_LC_21_19_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77304),
            .lcout(shift_srl_159Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93195),
            .ce(N__77702),
            .sr(_gnd_net_));
    defparam shift_srl_159_1_LC_21_19_3.C_ON=1'b0;
    defparam shift_srl_159_1_LC_21_19_3.SEQ_MODE=4'b1000;
    defparam shift_srl_159_1_LC_21_19_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_159_1_LC_21_19_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75406),
            .lcout(shift_srl_159Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93195),
            .ce(N__77702),
            .sr(_gnd_net_));
    defparam shift_srl_159_7_LC_21_19_4.C_ON=1'b0;
    defparam shift_srl_159_7_LC_21_19_4.SEQ_MODE=4'b1000;
    defparam shift_srl_159_7_LC_21_19_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_159_7_LC_21_19_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75400),
            .lcout(shift_srl_159Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93195),
            .ce(N__77702),
            .sr(_gnd_net_));
    defparam shift_srl_159_4_LC_21_19_5.C_ON=1'b0;
    defparam shift_srl_159_4_LC_21_19_5.SEQ_MODE=4'b1000;
    defparam shift_srl_159_4_LC_21_19_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_159_4_LC_21_19_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75502),
            .lcout(shift_srl_159Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93195),
            .ce(N__77702),
            .sr(_gnd_net_));
    defparam shift_srl_159_8_LC_21_19_6.C_ON=1'b0;
    defparam shift_srl_159_8_LC_21_19_6.SEQ_MODE=4'b1000;
    defparam shift_srl_159_8_LC_21_19_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_159_8_LC_21_19_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75490),
            .lcout(shift_srl_159Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93195),
            .ce(N__77702),
            .sr(_gnd_net_));
    defparam shift_srl_159_2_LC_21_19_7.C_ON=1'b0;
    defparam shift_srl_159_2_LC_21_19_7.SEQ_MODE=4'b1000;
    defparam shift_srl_159_2_LC_21_19_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_159_2_LC_21_19_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75478),
            .lcout(shift_srl_159Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93195),
            .ce(N__77702),
            .sr(_gnd_net_));
    defparam shift_srl_171_0_LC_21_20_0.C_ON=1'b0;
    defparam shift_srl_171_0_LC_21_20_0.SEQ_MODE=4'b1000;
    defparam shift_srl_171_0_LC_21_20_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_171_0_LC_21_20_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87494),
            .lcout(shift_srl_171Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93216),
            .ce(N__77956),
            .sr(_gnd_net_));
    defparam shift_srl_171_6_LC_21_20_1.C_ON=1'b0;
    defparam shift_srl_171_6_LC_21_20_1.SEQ_MODE=4'b1000;
    defparam shift_srl_171_6_LC_21_20_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_171_6_LC_21_20_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75448),
            .lcout(shift_srl_171Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93216),
            .ce(N__77956),
            .sr(_gnd_net_));
    defparam shift_srl_171_2_LC_21_20_2.C_ON=1'b0;
    defparam shift_srl_171_2_LC_21_20_2.SEQ_MODE=4'b1000;
    defparam shift_srl_171_2_LC_21_20_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_171_2_LC_21_20_2 (
            .in0(N__77962),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_171Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93216),
            .ce(N__77956),
            .sr(_gnd_net_));
    defparam shift_srl_171_3_LC_21_20_3.C_ON=1'b0;
    defparam shift_srl_171_3_LC_21_20_3.SEQ_MODE=4'b1000;
    defparam shift_srl_171_3_LC_21_20_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_171_3_LC_21_20_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75466),
            .lcout(shift_srl_171Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93216),
            .ce(N__77956),
            .sr(_gnd_net_));
    defparam shift_srl_171_4_LC_21_20_4.C_ON=1'b0;
    defparam shift_srl_171_4_LC_21_20_4.SEQ_MODE=4'b1000;
    defparam shift_srl_171_4_LC_21_20_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_171_4_LC_21_20_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75460),
            .lcout(shift_srl_171Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93216),
            .ce(N__77956),
            .sr(_gnd_net_));
    defparam shift_srl_171_5_LC_21_20_5.C_ON=1'b0;
    defparam shift_srl_171_5_LC_21_20_5.SEQ_MODE=4'b1000;
    defparam shift_srl_171_5_LC_21_20_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_171_5_LC_21_20_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75454),
            .lcout(shift_srl_171Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93216),
            .ce(N__77956),
            .sr(_gnd_net_));
    defparam shift_srl_171_8_LC_21_20_6.C_ON=1'b0;
    defparam shift_srl_171_8_LC_21_20_6.SEQ_MODE=4'b1000;
    defparam shift_srl_171_8_LC_21_20_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_171_8_LC_21_20_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75544),
            .lcout(shift_srl_171Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93216),
            .ce(N__77956),
            .sr(_gnd_net_));
    defparam shift_srl_171_7_LC_21_20_7.C_ON=1'b0;
    defparam shift_srl_171_7_LC_21_20_7.SEQ_MODE=4'b1000;
    defparam shift_srl_171_7_LC_21_20_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_171_7_LC_21_20_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75550),
            .lcout(shift_srl_171Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93216),
            .ce(N__77956),
            .sr(_gnd_net_));
    defparam shift_srl_179_0_LC_21_21_0.C_ON=1'b0;
    defparam shift_srl_179_0_LC_21_21_0.SEQ_MODE=4'b1000;
    defparam shift_srl_179_0_LC_21_21_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_179_0_LC_21_21_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78131),
            .lcout(shift_srl_179Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93234),
            .ce(N__78060),
            .sr(_gnd_net_));
    defparam shift_srl_179_1_LC_21_21_1.C_ON=1'b0;
    defparam shift_srl_179_1_LC_21_21_1.SEQ_MODE=4'b1000;
    defparam shift_srl_179_1_LC_21_21_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_179_1_LC_21_21_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75538),
            .lcout(shift_srl_179Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93234),
            .ce(N__78060),
            .sr(_gnd_net_));
    defparam shift_srl_179_2_LC_21_21_2.C_ON=1'b0;
    defparam shift_srl_179_2_LC_21_21_2.SEQ_MODE=4'b1000;
    defparam shift_srl_179_2_LC_21_21_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_179_2_LC_21_21_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75532),
            .lcout(shift_srl_179Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93234),
            .ce(N__78060),
            .sr(_gnd_net_));
    defparam shift_srl_179_3_LC_21_21_3.C_ON=1'b0;
    defparam shift_srl_179_3_LC_21_21_3.SEQ_MODE=4'b1000;
    defparam shift_srl_179_3_LC_21_21_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_179_3_LC_21_21_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75526),
            .lcout(shift_srl_179Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93234),
            .ce(N__78060),
            .sr(_gnd_net_));
    defparam shift_srl_179_4_LC_21_21_4.C_ON=1'b0;
    defparam shift_srl_179_4_LC_21_21_4.SEQ_MODE=4'b1000;
    defparam shift_srl_179_4_LC_21_21_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_179_4_LC_21_21_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75520),
            .lcout(shift_srl_179Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93234),
            .ce(N__78060),
            .sr(_gnd_net_));
    defparam shift_srl_179_5_LC_21_21_5.C_ON=1'b0;
    defparam shift_srl_179_5_LC_21_21_5.SEQ_MODE=4'b1000;
    defparam shift_srl_179_5_LC_21_21_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_179_5_LC_21_21_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75514),
            .lcout(shift_srl_179Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93234),
            .ce(N__78060),
            .sr(_gnd_net_));
    defparam shift_srl_179_6_LC_21_21_6.C_ON=1'b0;
    defparam shift_srl_179_6_LC_21_21_6.SEQ_MODE=4'b1000;
    defparam shift_srl_179_6_LC_21_21_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_179_6_LC_21_21_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75508),
            .lcout(shift_srl_179Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93234),
            .ce(N__78060),
            .sr(_gnd_net_));
    defparam shift_srl_179_7_LC_21_21_7.C_ON=1'b0;
    defparam shift_srl_179_7_LC_21_21_7.SEQ_MODE=4'b1000;
    defparam shift_srl_179_7_LC_21_21_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_179_7_LC_21_21_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75628),
            .lcout(shift_srl_179Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93234),
            .ce(N__78060),
            .sr(_gnd_net_));
    defparam shift_srl_186_10_LC_21_22_0.C_ON=1'b0;
    defparam shift_srl_186_10_LC_21_22_0.SEQ_MODE=4'b1000;
    defparam shift_srl_186_10_LC_21_22_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_186_10_LC_21_22_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75592),
            .lcout(shift_srl_186Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93256),
            .ce(N__75574),
            .sr(_gnd_net_));
    defparam shift_srl_186_11_LC_21_22_1.C_ON=1'b0;
    defparam shift_srl_186_11_LC_21_22_1.SEQ_MODE=4'b1000;
    defparam shift_srl_186_11_LC_21_22_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_186_11_LC_21_22_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75622),
            .lcout(shift_srl_186Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93256),
            .ce(N__75574),
            .sr(_gnd_net_));
    defparam shift_srl_186_12_LC_21_22_2.C_ON=1'b0;
    defparam shift_srl_186_12_LC_21_22_2.SEQ_MODE=4'b1000;
    defparam shift_srl_186_12_LC_21_22_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_186_12_LC_21_22_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75616),
            .lcout(shift_srl_186Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93256),
            .ce(N__75574),
            .sr(_gnd_net_));
    defparam shift_srl_186_13_LC_21_22_3.C_ON=1'b0;
    defparam shift_srl_186_13_LC_21_22_3.SEQ_MODE=4'b1000;
    defparam shift_srl_186_13_LC_21_22_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_186_13_LC_21_22_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75610),
            .lcout(shift_srl_186Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93256),
            .ce(N__75574),
            .sr(_gnd_net_));
    defparam shift_srl_186_14_LC_21_22_4.C_ON=1'b0;
    defparam shift_srl_186_14_LC_21_22_4.SEQ_MODE=4'b1000;
    defparam shift_srl_186_14_LC_21_22_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_186_14_LC_21_22_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75604),
            .lcout(shift_srl_186Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93256),
            .ce(N__75574),
            .sr(_gnd_net_));
    defparam shift_srl_186_15_LC_21_22_5.C_ON=1'b0;
    defparam shift_srl_186_15_LC_21_22_5.SEQ_MODE=4'b1000;
    defparam shift_srl_186_15_LC_21_22_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_186_15_LC_21_22_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75598),
            .lcout(shift_srl_186Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93256),
            .ce(N__75574),
            .sr(_gnd_net_));
    defparam shift_srl_186_9_LC_21_22_6.C_ON=1'b0;
    defparam shift_srl_186_9_LC_21_22_6.SEQ_MODE=4'b1000;
    defparam shift_srl_186_9_LC_21_22_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_186_9_LC_21_22_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75580),
            .lcout(shift_srl_186Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93256),
            .ce(N__75574),
            .sr(_gnd_net_));
    defparam shift_srl_186_8_LC_21_22_7.C_ON=1'b0;
    defparam shift_srl_186_8_LC_21_22_7.SEQ_MODE=4'b1000;
    defparam shift_srl_186_8_LC_21_22_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_186_8_LC_21_22_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75586),
            .lcout(shift_srl_186Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93256),
            .ce(N__75574),
            .sr(_gnd_net_));
    defparam shift_srl_178_0_LC_21_23_0.C_ON=1'b0;
    defparam shift_srl_178_0_LC_21_23_0.SEQ_MODE=4'b1000;
    defparam shift_srl_178_0_LC_21_23_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_178_0_LC_21_23_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80405),
            .lcout(shift_srl_178Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93275),
            .ce(N__78102),
            .sr(_gnd_net_));
    defparam shift_srl_178_1_LC_21_23_1.C_ON=1'b0;
    defparam shift_srl_178_1_LC_21_23_1.SEQ_MODE=4'b1000;
    defparam shift_srl_178_1_LC_21_23_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_178_1_LC_21_23_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75664),
            .lcout(shift_srl_178Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93275),
            .ce(N__78102),
            .sr(_gnd_net_));
    defparam shift_srl_178_2_LC_21_23_2.C_ON=1'b0;
    defparam shift_srl_178_2_LC_21_23_2.SEQ_MODE=4'b1000;
    defparam shift_srl_178_2_LC_21_23_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_178_2_LC_21_23_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75658),
            .lcout(shift_srl_178Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93275),
            .ce(N__78102),
            .sr(_gnd_net_));
    defparam shift_srl_178_3_LC_21_23_3.C_ON=1'b0;
    defparam shift_srl_178_3_LC_21_23_3.SEQ_MODE=4'b1000;
    defparam shift_srl_178_3_LC_21_23_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_178_3_LC_21_23_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75652),
            .lcout(shift_srl_178Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93275),
            .ce(N__78102),
            .sr(_gnd_net_));
    defparam shift_srl_178_4_LC_21_23_4.C_ON=1'b0;
    defparam shift_srl_178_4_LC_21_23_4.SEQ_MODE=4'b1000;
    defparam shift_srl_178_4_LC_21_23_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_178_4_LC_21_23_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75646),
            .lcout(shift_srl_178Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93275),
            .ce(N__78102),
            .sr(_gnd_net_));
    defparam shift_srl_178_5_LC_21_23_5.C_ON=1'b0;
    defparam shift_srl_178_5_LC_21_23_5.SEQ_MODE=4'b1000;
    defparam shift_srl_178_5_LC_21_23_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_178_5_LC_21_23_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75640),
            .lcout(shift_srl_178Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93275),
            .ce(N__78102),
            .sr(_gnd_net_));
    defparam shift_srl_178_10_LC_21_23_6.C_ON=1'b0;
    defparam shift_srl_178_10_LC_21_23_6.SEQ_MODE=4'b1000;
    defparam shift_srl_178_10_LC_21_23_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_178_10_LC_21_23_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75634),
            .lcout(shift_srl_178Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93275),
            .ce(N__78102),
            .sr(_gnd_net_));
    defparam shift_srl_178_9_LC_21_23_7.C_ON=1'b0;
    defparam shift_srl_178_9_LC_21_23_7.SEQ_MODE=4'b1000;
    defparam shift_srl_178_9_LC_21_23_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_178_9_LC_21_23_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77986),
            .lcout(shift_srl_178Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93275),
            .ce(N__78102),
            .sr(_gnd_net_));
    defparam shift_srl_181_15_LC_21_24_0.C_ON=1'b0;
    defparam shift_srl_181_15_LC_21_24_0.SEQ_MODE=4'b1000;
    defparam shift_srl_181_15_LC_21_24_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_181_15_LC_21_24_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78235),
            .lcout(shift_srl_181Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93290),
            .ce(N__78211),
            .sr(_gnd_net_));
    defparam shift_srl_181_1_LC_21_24_1.C_ON=1'b0;
    defparam shift_srl_181_1_LC_21_24_1.SEQ_MODE=4'b1000;
    defparam shift_srl_181_1_LC_21_24_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_181_1_LC_21_24_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75682),
            .lcout(shift_srl_181Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93290),
            .ce(N__78211),
            .sr(_gnd_net_));
    defparam shift_srl_181_2_LC_21_24_2.C_ON=1'b0;
    defparam shift_srl_181_2_LC_21_24_2.SEQ_MODE=4'b1000;
    defparam shift_srl_181_2_LC_21_24_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_181_2_LC_21_24_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75712),
            .lcout(shift_srl_181Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93290),
            .ce(N__78211),
            .sr(_gnd_net_));
    defparam shift_srl_181_3_LC_21_24_3.C_ON=1'b0;
    defparam shift_srl_181_3_LC_21_24_3.SEQ_MODE=4'b1000;
    defparam shift_srl_181_3_LC_21_24_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_181_3_LC_21_24_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75706),
            .lcout(shift_srl_181Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93290),
            .ce(N__78211),
            .sr(_gnd_net_));
    defparam shift_srl_181_4_LC_21_24_4.C_ON=1'b0;
    defparam shift_srl_181_4_LC_21_24_4.SEQ_MODE=4'b1000;
    defparam shift_srl_181_4_LC_21_24_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_181_4_LC_21_24_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75700),
            .lcout(shift_srl_181Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93290),
            .ce(N__78211),
            .sr(_gnd_net_));
    defparam shift_srl_181_5_LC_21_24_5.C_ON=1'b0;
    defparam shift_srl_181_5_LC_21_24_5.SEQ_MODE=4'b1000;
    defparam shift_srl_181_5_LC_21_24_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_181_5_LC_21_24_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75694),
            .lcout(shift_srl_181Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93290),
            .ce(N__78211),
            .sr(_gnd_net_));
    defparam shift_srl_181_6_LC_21_24_6.C_ON=1'b0;
    defparam shift_srl_181_6_LC_21_24_6.SEQ_MODE=4'b1000;
    defparam shift_srl_181_6_LC_21_24_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_181_6_LC_21_24_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75688),
            .lcout(shift_srl_181Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93290),
            .ce(N__78211),
            .sr(_gnd_net_));
    defparam shift_srl_181_0_LC_21_24_7.C_ON=1'b0;
    defparam shift_srl_181_0_LC_21_24_7.SEQ_MODE=4'b1000;
    defparam shift_srl_181_0_LC_21_24_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_181_0_LC_21_24_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75875),
            .lcout(shift_srl_181Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93290),
            .ce(N__78211),
            .sr(_gnd_net_));
    defparam shift_srl_176_10_LC_21_25_0.C_ON=1'b0;
    defparam shift_srl_176_10_LC_21_25_0.SEQ_MODE=4'b1000;
    defparam shift_srl_176_10_LC_21_25_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_176_10_LC_21_25_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75760),
            .lcout(shift_srl_176Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93307),
            .ce(N__78531),
            .sr(_gnd_net_));
    defparam shift_srl_176_11_LC_21_25_1.C_ON=1'b0;
    defparam shift_srl_176_11_LC_21_25_1.SEQ_MODE=4'b1000;
    defparam shift_srl_176_11_LC_21_25_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_176_11_LC_21_25_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75676),
            .lcout(shift_srl_176Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93307),
            .ce(N__78531),
            .sr(_gnd_net_));
    defparam shift_srl_176_12_LC_21_25_2.C_ON=1'b0;
    defparam shift_srl_176_12_LC_21_25_2.SEQ_MODE=4'b1000;
    defparam shift_srl_176_12_LC_21_25_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_176_12_LC_21_25_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75670),
            .lcout(shift_srl_176Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93307),
            .ce(N__78531),
            .sr(_gnd_net_));
    defparam shift_srl_176_13_LC_21_25_3.C_ON=1'b0;
    defparam shift_srl_176_13_LC_21_25_3.SEQ_MODE=4'b1000;
    defparam shift_srl_176_13_LC_21_25_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_176_13_LC_21_25_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75778),
            .lcout(shift_srl_176Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93307),
            .ce(N__78531),
            .sr(_gnd_net_));
    defparam shift_srl_176_14_LC_21_25_4.C_ON=1'b0;
    defparam shift_srl_176_14_LC_21_25_4.SEQ_MODE=4'b1000;
    defparam shift_srl_176_14_LC_21_25_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_176_14_LC_21_25_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75772),
            .lcout(shift_srl_176Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93307),
            .ce(N__78531),
            .sr(_gnd_net_));
    defparam shift_srl_176_15_LC_21_25_5.C_ON=1'b0;
    defparam shift_srl_176_15_LC_21_25_5.SEQ_MODE=4'b1000;
    defparam shift_srl_176_15_LC_21_25_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_176_15_LC_21_25_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75766),
            .lcout(shift_srl_176Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93307),
            .ce(N__78531),
            .sr(_gnd_net_));
    defparam shift_srl_176_9_LC_21_25_6.C_ON=1'b0;
    defparam shift_srl_176_9_LC_21_25_6.SEQ_MODE=4'b1000;
    defparam shift_srl_176_9_LC_21_25_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_176_9_LC_21_25_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75754),
            .lcout(shift_srl_176Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93307),
            .ce(N__78531),
            .sr(_gnd_net_));
    defparam shift_srl_176_8_LC_21_25_7.C_ON=1'b0;
    defparam shift_srl_176_8_LC_21_25_7.SEQ_MODE=4'b1000;
    defparam shift_srl_176_8_LC_21_25_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_176_8_LC_21_25_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78541),
            .lcout(shift_srl_176Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93307),
            .ce(N__78531),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_175_LC_21_26_0.C_ON=1'b0;
    defparam rco_obuf_RNO_175_LC_21_26_0.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_175_LC_21_26_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 rco_obuf_RNO_175_LC_21_26_0 (
            .in0(N__76050),
            .in1(N__76015),
            .in2(N__85968),
            .in3(N__75939),
            .lcout(rco_c_175),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_174_LC_21_26_1.C_ON=1'b0;
    defparam rco_obuf_RNO_174_LC_21_26_1.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_174_LC_21_26_1.LUT_INIT=16'b1000100000000000;
    LogicCell40 rco_obuf_RNO_174_LC_21_26_1 (
            .in0(N__75938),
            .in1(N__76024),
            .in2(_gnd_net_),
            .in3(N__85941),
            .lcout(rco_c_174),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_175_RNILMSL_15_LC_21_26_2.C_ON=1'b0;
    defparam shift_srl_175_RNILMSL_15_LC_21_26_2.SEQ_MODE=4'b0000;
    defparam shift_srl_175_RNILMSL_15_LC_21_26_2.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_175_RNILMSL_15_LC_21_26_2 (
            .in0(N__76049),
            .in1(N__76014),
            .in2(_gnd_net_),
            .in3(N__75937),
            .lcout(),
            .ltout(clk_en_0_a3_0_a2cf1_176_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_175_RNIEIJ5C1_15_LC_21_26_3.C_ON=1'b0;
    defparam shift_srl_175_RNIEIJ5C1_15_LC_21_26_3.SEQ_MODE=4'b0000;
    defparam shift_srl_175_RNIEIJ5C1_15_LC_21_26_3.LUT_INIT=16'b0011000000000000;
    LogicCell40 shift_srl_175_RNIEIJ5C1_15_LC_21_26_3 (
            .in0(_gnd_net_),
            .in1(N__84159),
            .in2(N__75715),
            .in3(N__87900),
            .lcout(clk_en_176),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_173_15_LC_21_26_4.C_ON=1'b0;
    defparam shift_srl_173_15_LC_21_26_4.SEQ_MODE=4'b1000;
    defparam shift_srl_173_15_LC_21_26_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_173_15_LC_21_26_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80623),
            .lcout(shift_srl_173Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93328),
            .ce(N__80583),
            .sr(_gnd_net_));
    defparam shift_srl_176_RNIUGI51_0_15_LC_21_26_5.C_ON=1'b0;
    defparam shift_srl_176_RNIUGI51_0_15_LC_21_26_5.SEQ_MODE=4'b0000;
    defparam shift_srl_176_RNIUGI51_0_15_LC_21_26_5.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_176_RNIUGI51_0_15_LC_21_26_5 (
            .in0(N__75936),
            .in1(N__78350),
            .in2(N__76022),
            .in3(N__76048),
            .lcout(rco_int_0_a2_1_a2_0_sx_179),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_176_RNIUGI51_15_LC_21_26_6.C_ON=1'b0;
    defparam shift_srl_176_RNIUGI51_15_LC_21_26_6.SEQ_MODE=4'b0000;
    defparam shift_srl_176_RNIUGI51_15_LC_21_26_6.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_176_RNIUGI51_15_LC_21_26_6 (
            .in0(N__76047),
            .in1(N__76010),
            .in2(N__78352),
            .in3(N__75935),
            .lcout(shift_srl_176_RNIUGI51Z0Z_15),
            .ltout(shift_srl_176_RNIUGI51Z0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_182_RNIEPSC2_15_LC_21_26_7.C_ON=1'b0;
    defparam shift_srl_182_RNIEPSC2_15_LC_21_26_7.SEQ_MODE=4'b0000;
    defparam shift_srl_182_RNIEPSC2_15_LC_21_26_7.LUT_INIT=16'b0000000010000000;
    LogicCell40 shift_srl_182_RNIEPSC2_15_LC_21_26_7 (
            .in0(N__75904),
            .in1(N__75876),
            .in2(N__75853),
            .in3(N__78115),
            .lcout(shift_srl_182_RNIEPSC2Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_193_10_LC_21_27_0.C_ON=1'b0;
    defparam shift_srl_193_10_LC_21_27_0.SEQ_MODE=4'b1000;
    defparam shift_srl_193_10_LC_21_27_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_193_10_LC_21_27_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76117),
            .lcout(shift_srl_193Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93350),
            .ce(N__76231),
            .sr(_gnd_net_));
    defparam shift_srl_193_11_LC_21_27_1.C_ON=1'b0;
    defparam shift_srl_193_11_LC_21_27_1.SEQ_MODE=4'b1000;
    defparam shift_srl_193_11_LC_21_27_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_193_11_LC_21_27_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75802),
            .lcout(shift_srl_193Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93350),
            .ce(N__76231),
            .sr(_gnd_net_));
    defparam shift_srl_193_12_LC_21_27_2.C_ON=1'b0;
    defparam shift_srl_193_12_LC_21_27_2.SEQ_MODE=4'b1000;
    defparam shift_srl_193_12_LC_21_27_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_193_12_LC_21_27_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75796),
            .lcout(shift_srl_193Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93350),
            .ce(N__76231),
            .sr(_gnd_net_));
    defparam shift_srl_193_13_LC_21_27_3.C_ON=1'b0;
    defparam shift_srl_193_13_LC_21_27_3.SEQ_MODE=4'b1000;
    defparam shift_srl_193_13_LC_21_27_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_193_13_LC_21_27_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75790),
            .lcout(shift_srl_193Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93350),
            .ce(N__76231),
            .sr(_gnd_net_));
    defparam shift_srl_193_14_LC_21_27_4.C_ON=1'b0;
    defparam shift_srl_193_14_LC_21_27_4.SEQ_MODE=4'b1000;
    defparam shift_srl_193_14_LC_21_27_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_193_14_LC_21_27_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75784),
            .lcout(shift_srl_193Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93350),
            .ce(N__76231),
            .sr(_gnd_net_));
    defparam shift_srl_193_15_LC_21_27_5.C_ON=1'b0;
    defparam shift_srl_193_15_LC_21_27_5.SEQ_MODE=4'b1000;
    defparam shift_srl_193_15_LC_21_27_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_193_15_LC_21_27_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76123),
            .lcout(shift_srl_193Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93350),
            .ce(N__76231),
            .sr(_gnd_net_));
    defparam shift_srl_193_9_LC_21_27_6.C_ON=1'b0;
    defparam shift_srl_193_9_LC_21_27_6.SEQ_MODE=4'b1000;
    defparam shift_srl_193_9_LC_21_27_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_193_9_LC_21_27_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76111),
            .lcout(shift_srl_193Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93350),
            .ce(N__76231),
            .sr(_gnd_net_));
    defparam shift_srl_193_8_LC_21_27_7.C_ON=1'b0;
    defparam shift_srl_193_8_LC_21_27_7.SEQ_MODE=4'b1000;
    defparam shift_srl_193_8_LC_21_27_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_193_8_LC_21_27_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76237),
            .lcout(shift_srl_193Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93350),
            .ce(N__76231),
            .sr(_gnd_net_));
    defparam shift_srl_193_0_LC_21_28_0.C_ON=1'b0;
    defparam shift_srl_193_0_LC_21_28_0.SEQ_MODE=4'b1000;
    defparam shift_srl_193_0_LC_21_28_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_193_0_LC_21_28_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76101),
            .lcout(shift_srl_193Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93366),
            .ce(N__76224),
            .sr(_gnd_net_));
    defparam shift_srl_193_1_LC_21_28_1.C_ON=1'b0;
    defparam shift_srl_193_1_LC_21_28_1.SEQ_MODE=4'b1000;
    defparam shift_srl_193_1_LC_21_28_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_193_1_LC_21_28_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76087),
            .lcout(shift_srl_193Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93366),
            .ce(N__76224),
            .sr(_gnd_net_));
    defparam shift_srl_193_2_LC_21_28_2.C_ON=1'b0;
    defparam shift_srl_193_2_LC_21_28_2.SEQ_MODE=4'b1000;
    defparam shift_srl_193_2_LC_21_28_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_193_2_LC_21_28_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76081),
            .lcout(shift_srl_193Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93366),
            .ce(N__76224),
            .sr(_gnd_net_));
    defparam shift_srl_193_3_LC_21_28_3.C_ON=1'b0;
    defparam shift_srl_193_3_LC_21_28_3.SEQ_MODE=4'b1000;
    defparam shift_srl_193_3_LC_21_28_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_193_3_LC_21_28_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76075),
            .lcout(shift_srl_193Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93366),
            .ce(N__76224),
            .sr(_gnd_net_));
    defparam shift_srl_193_4_LC_21_28_4.C_ON=1'b0;
    defparam shift_srl_193_4_LC_21_28_4.SEQ_MODE=4'b1000;
    defparam shift_srl_193_4_LC_21_28_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_193_4_LC_21_28_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76069),
            .lcout(shift_srl_193Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93366),
            .ce(N__76224),
            .sr(_gnd_net_));
    defparam shift_srl_193_5_LC_21_28_5.C_ON=1'b0;
    defparam shift_srl_193_5_LC_21_28_5.SEQ_MODE=4'b1000;
    defparam shift_srl_193_5_LC_21_28_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_193_5_LC_21_28_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76063),
            .lcout(shift_srl_193Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93366),
            .ce(N__76224),
            .sr(_gnd_net_));
    defparam shift_srl_193_6_LC_21_28_6.C_ON=1'b0;
    defparam shift_srl_193_6_LC_21_28_6.SEQ_MODE=4'b1000;
    defparam shift_srl_193_6_LC_21_28_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_193_6_LC_21_28_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76057),
            .lcout(shift_srl_193Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93366),
            .ce(N__76224),
            .sr(_gnd_net_));
    defparam shift_srl_193_7_LC_21_28_7.C_ON=1'b0;
    defparam shift_srl_193_7_LC_21_28_7.SEQ_MODE=4'b1000;
    defparam shift_srl_193_7_LC_21_28_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_193_7_LC_21_28_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76243),
            .lcout(shift_srl_193Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93366),
            .ce(N__76224),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_45_LC_22_4_4.C_ON=1'b0;
    defparam rco_obuf_RNO_45_LC_22_4_4.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_45_LC_22_4_4.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_45_LC_22_4_4 (
            .in0(N__76907),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76210),
            .lcout(rco_c_45),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_47_0_LC_22_6_0.C_ON=1'b0;
    defparam shift_srl_47_0_LC_22_6_0.SEQ_MODE=4'b1000;
    defparam shift_srl_47_0_LC_22_6_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_47_0_LC_22_6_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76321),
            .lcout(shift_srl_47Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93385),
            .ce(N__76255),
            .sr(_gnd_net_));
    defparam shift_srl_47_1_LC_22_6_1.C_ON=1'b0;
    defparam shift_srl_47_1_LC_22_6_1.SEQ_MODE=4'b1000;
    defparam shift_srl_47_1_LC_22_6_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_47_1_LC_22_6_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76159),
            .lcout(shift_srl_47Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93385),
            .ce(N__76255),
            .sr(_gnd_net_));
    defparam shift_srl_47_2_LC_22_6_2.C_ON=1'b0;
    defparam shift_srl_47_2_LC_22_6_2.SEQ_MODE=4'b1000;
    defparam shift_srl_47_2_LC_22_6_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_47_2_LC_22_6_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76153),
            .lcout(shift_srl_47Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93385),
            .ce(N__76255),
            .sr(_gnd_net_));
    defparam shift_srl_47_3_LC_22_6_3.C_ON=1'b0;
    defparam shift_srl_47_3_LC_22_6_3.SEQ_MODE=4'b1000;
    defparam shift_srl_47_3_LC_22_6_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_47_3_LC_22_6_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76147),
            .lcout(shift_srl_47Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93385),
            .ce(N__76255),
            .sr(_gnd_net_));
    defparam shift_srl_47_4_LC_22_6_4.C_ON=1'b0;
    defparam shift_srl_47_4_LC_22_6_4.SEQ_MODE=4'b1000;
    defparam shift_srl_47_4_LC_22_6_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_47_4_LC_22_6_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76141),
            .lcout(shift_srl_47Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93385),
            .ce(N__76255),
            .sr(_gnd_net_));
    defparam shift_srl_47_5_LC_22_6_5.C_ON=1'b0;
    defparam shift_srl_47_5_LC_22_6_5.SEQ_MODE=4'b1000;
    defparam shift_srl_47_5_LC_22_6_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_47_5_LC_22_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76135),
            .lcout(shift_srl_47Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93385),
            .ce(N__76255),
            .sr(_gnd_net_));
    defparam shift_srl_47_6_LC_22_6_6.C_ON=1'b0;
    defparam shift_srl_47_6_LC_22_6_6.SEQ_MODE=4'b1000;
    defparam shift_srl_47_6_LC_22_6_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_47_6_LC_22_6_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76129),
            .lcout(shift_srl_47Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93385),
            .ce(N__76255),
            .sr(_gnd_net_));
    defparam shift_srl_47_15_LC_22_6_7.C_ON=1'b0;
    defparam shift_srl_47_15_LC_22_6_7.SEQ_MODE=4'b1000;
    defparam shift_srl_47_15_LC_22_6_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_47_15_LC_22_6_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76285),
            .lcout(shift_srl_47Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93385),
            .ce(N__76255),
            .sr(_gnd_net_));
    defparam shift_srl_47_10_LC_22_7_0.C_ON=1'b0;
    defparam shift_srl_47_10_LC_22_7_0.SEQ_MODE=4'b1000;
    defparam shift_srl_47_10_LC_22_7_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_47_10_LC_22_7_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76273),
            .lcout(shift_srl_47Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93369),
            .ce(N__76254),
            .sr(_gnd_net_));
    defparam shift_srl_47_11_LC_22_7_1.C_ON=1'b0;
    defparam shift_srl_47_11_LC_22_7_1.SEQ_MODE=4'b1000;
    defparam shift_srl_47_11_LC_22_7_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_47_11_LC_22_7_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76309),
            .lcout(shift_srl_47Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93369),
            .ce(N__76254),
            .sr(_gnd_net_));
    defparam shift_srl_47_12_LC_22_7_2.C_ON=1'b0;
    defparam shift_srl_47_12_LC_22_7_2.SEQ_MODE=4'b1000;
    defparam shift_srl_47_12_LC_22_7_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_47_12_LC_22_7_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76303),
            .lcout(shift_srl_47Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93369),
            .ce(N__76254),
            .sr(_gnd_net_));
    defparam shift_srl_47_13_LC_22_7_3.C_ON=1'b0;
    defparam shift_srl_47_13_LC_22_7_3.SEQ_MODE=4'b1000;
    defparam shift_srl_47_13_LC_22_7_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_47_13_LC_22_7_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76297),
            .lcout(shift_srl_47Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93369),
            .ce(N__76254),
            .sr(_gnd_net_));
    defparam shift_srl_47_14_LC_22_7_4.C_ON=1'b0;
    defparam shift_srl_47_14_LC_22_7_4.SEQ_MODE=4'b1000;
    defparam shift_srl_47_14_LC_22_7_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_47_14_LC_22_7_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76291),
            .lcout(shift_srl_47Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93369),
            .ce(N__76254),
            .sr(_gnd_net_));
    defparam shift_srl_47_7_LC_22_7_5.C_ON=1'b0;
    defparam shift_srl_47_7_LC_22_7_5.SEQ_MODE=4'b1000;
    defparam shift_srl_47_7_LC_22_7_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_47_7_LC_22_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76279),
            .lcout(shift_srl_47Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93369),
            .ce(N__76254),
            .sr(_gnd_net_));
    defparam shift_srl_47_9_LC_22_7_6.C_ON=1'b0;
    defparam shift_srl_47_9_LC_22_7_6.SEQ_MODE=4'b1000;
    defparam shift_srl_47_9_LC_22_7_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_47_9_LC_22_7_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76261),
            .lcout(shift_srl_47Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93369),
            .ce(N__76254),
            .sr(_gnd_net_));
    defparam shift_srl_47_8_LC_22_7_7.C_ON=1'b0;
    defparam shift_srl_47_8_LC_22_7_7.SEQ_MODE=4'b1000;
    defparam shift_srl_47_8_LC_22_7_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_47_8_LC_22_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76267),
            .lcout(shift_srl_47Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93369),
            .ce(N__76254),
            .sr(_gnd_net_));
    defparam shift_srl_50_10_LC_22_8_0.C_ON=1'b0;
    defparam shift_srl_50_10_LC_22_8_0.SEQ_MODE=4'b1000;
    defparam shift_srl_50_10_LC_22_8_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_50_10_LC_22_8_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76369),
            .lcout(shift_srl_50Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93352),
            .ce(N__76475),
            .sr(_gnd_net_));
    defparam shift_srl_50_5_LC_22_8_2.C_ON=1'b0;
    defparam shift_srl_50_5_LC_22_8_2.SEQ_MODE=4'b1000;
    defparam shift_srl_50_5_LC_22_8_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_50_5_LC_22_8_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76492),
            .lcout(shift_srl_50Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93352),
            .ce(N__76475),
            .sr(_gnd_net_));
    defparam shift_srl_50_6_LC_22_8_4.C_ON=1'b0;
    defparam shift_srl_50_6_LC_22_8_4.SEQ_MODE=4'b1000;
    defparam shift_srl_50_6_LC_22_8_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_50_6_LC_22_8_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76381),
            .lcout(shift_srl_50Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93352),
            .ce(N__76475),
            .sr(_gnd_net_));
    defparam shift_srl_50_7_LC_22_8_5.C_ON=1'b0;
    defparam shift_srl_50_7_LC_22_8_5.SEQ_MODE=4'b1000;
    defparam shift_srl_50_7_LC_22_8_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_50_7_LC_22_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76375),
            .lcout(shift_srl_50Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93352),
            .ce(N__76475),
            .sr(_gnd_net_));
    defparam shift_srl_50_9_LC_22_8_6.C_ON=1'b0;
    defparam shift_srl_50_9_LC_22_8_6.SEQ_MODE=4'b1000;
    defparam shift_srl_50_9_LC_22_8_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_50_9_LC_22_8_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76357),
            .lcout(shift_srl_50Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93352),
            .ce(N__76475),
            .sr(_gnd_net_));
    defparam shift_srl_50_8_LC_22_8_7.C_ON=1'b0;
    defparam shift_srl_50_8_LC_22_8_7.SEQ_MODE=4'b1000;
    defparam shift_srl_50_8_LC_22_8_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_50_8_LC_22_8_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76363),
            .lcout(shift_srl_50Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93352),
            .ce(N__76475),
            .sr(_gnd_net_));
    defparam shift_srl_49_RNIPO9UC_15_LC_22_9_0.C_ON=1'b0;
    defparam shift_srl_49_RNIPO9UC_15_LC_22_9_0.SEQ_MODE=4'b0000;
    defparam shift_srl_49_RNIPO9UC_15_LC_22_9_0.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_49_RNIPO9UC_15_LC_22_9_0 (
            .in0(N__90227),
            .in1(N__93564),
            .in2(_gnd_net_),
            .in3(N__93495),
            .lcout(clk_en_50),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_50_0_LC_22_9_2.C_ON=1'b0;
    defparam shift_srl_50_0_LC_22_9_2.SEQ_MODE=4'b1000;
    defparam shift_srl_50_0_LC_22_9_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_50_0_LC_22_9_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76347),
            .lcout(shift_srl_50Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93331),
            .ce(N__76474),
            .sr(_gnd_net_));
    defparam shift_srl_50_1_LC_22_9_3.C_ON=1'b0;
    defparam shift_srl_50_1_LC_22_9_3.SEQ_MODE=4'b1000;
    defparam shift_srl_50_1_LC_22_9_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_50_1_LC_22_9_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76327),
            .lcout(shift_srl_50Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93331),
            .ce(N__76474),
            .sr(_gnd_net_));
    defparam shift_srl_50_2_LC_22_9_4.C_ON=1'b0;
    defparam shift_srl_50_2_LC_22_9_4.SEQ_MODE=4'b1000;
    defparam shift_srl_50_2_LC_22_9_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_50_2_LC_22_9_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76510),
            .lcout(shift_srl_50Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93331),
            .ce(N__76474),
            .sr(_gnd_net_));
    defparam shift_srl_50_3_LC_22_9_5.C_ON=1'b0;
    defparam shift_srl_50_3_LC_22_9_5.SEQ_MODE=4'b1000;
    defparam shift_srl_50_3_LC_22_9_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_50_3_LC_22_9_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76504),
            .lcout(shift_srl_50Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93331),
            .ce(N__76474),
            .sr(_gnd_net_));
    defparam shift_srl_50_4_LC_22_9_6.C_ON=1'b0;
    defparam shift_srl_50_4_LC_22_9_6.SEQ_MODE=4'b1000;
    defparam shift_srl_50_4_LC_22_9_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_50_4_LC_22_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76498),
            .lcout(shift_srl_50Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93331),
            .ce(N__76474),
            .sr(_gnd_net_));
    defparam shift_srl_52_0_LC_22_10_0.C_ON=1'b0;
    defparam shift_srl_52_0_LC_22_10_0.SEQ_MODE=4'b1000;
    defparam shift_srl_52_0_LC_22_10_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_52_0_LC_22_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76442),
            .lcout(shift_srl_52Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93309),
            .ce(N__76690),
            .sr(_gnd_net_));
    defparam shift_srl_52_1_LC_22_10_1.C_ON=1'b0;
    defparam shift_srl_52_1_LC_22_10_1.SEQ_MODE=4'b1000;
    defparam shift_srl_52_1_LC_22_10_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_52_1_LC_22_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76417),
            .lcout(shift_srl_52Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93309),
            .ce(N__76690),
            .sr(_gnd_net_));
    defparam shift_srl_52_2_LC_22_10_2.C_ON=1'b0;
    defparam shift_srl_52_2_LC_22_10_2.SEQ_MODE=4'b1000;
    defparam shift_srl_52_2_LC_22_10_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_52_2_LC_22_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76411),
            .lcout(shift_srl_52Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93309),
            .ce(N__76690),
            .sr(_gnd_net_));
    defparam shift_srl_52_3_LC_22_10_3.C_ON=1'b0;
    defparam shift_srl_52_3_LC_22_10_3.SEQ_MODE=4'b1000;
    defparam shift_srl_52_3_LC_22_10_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_52_3_LC_22_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76405),
            .lcout(shift_srl_52Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93309),
            .ce(N__76690),
            .sr(_gnd_net_));
    defparam shift_srl_52_4_LC_22_10_4.C_ON=1'b0;
    defparam shift_srl_52_4_LC_22_10_4.SEQ_MODE=4'b1000;
    defparam shift_srl_52_4_LC_22_10_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_52_4_LC_22_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76399),
            .lcout(shift_srl_52Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93309),
            .ce(N__76690),
            .sr(_gnd_net_));
    defparam shift_srl_52_5_LC_22_10_5.C_ON=1'b0;
    defparam shift_srl_52_5_LC_22_10_5.SEQ_MODE=4'b1000;
    defparam shift_srl_52_5_LC_22_10_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_52_5_LC_22_10_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76393),
            .lcout(shift_srl_52Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93309),
            .ce(N__76690),
            .sr(_gnd_net_));
    defparam shift_srl_52_6_LC_22_10_6.C_ON=1'b0;
    defparam shift_srl_52_6_LC_22_10_6.SEQ_MODE=4'b1000;
    defparam shift_srl_52_6_LC_22_10_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_52_6_LC_22_10_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76708),
            .lcout(shift_srl_52Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93309),
            .ce(N__76690),
            .sr(_gnd_net_));
    defparam shift_srl_52_7_LC_22_10_7.C_ON=1'b0;
    defparam shift_srl_52_7_LC_22_10_7.SEQ_MODE=4'b1000;
    defparam shift_srl_52_7_LC_22_10_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_52_7_LC_22_10_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76702),
            .lcout(shift_srl_52Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93309),
            .ce(N__76690),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_57_LC_22_11_0.C_ON=1'b0;
    defparam rco_obuf_RNO_57_LC_22_11_0.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_57_LC_22_11_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 rco_obuf_RNO_57_LC_22_11_0 (
            .in0(N__76796),
            .in1(N__77048),
            .in2(N__76945),
            .in3(N__76548),
            .lcout(rco_c_57),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_56_LC_22_11_1.C_ON=1'b0;
    defparam rco_obuf_RNO_56_LC_22_11_1.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_56_LC_22_11_1.LUT_INIT=16'b1000100000000000;
    LogicCell40 rco_obuf_RNO_56_LC_22_11_1 (
            .in0(N__77047),
            .in1(N__76546),
            .in2(_gnd_net_),
            .in3(N__76941),
            .lcout(rco_c_56),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIVU6PD_15_LC_22_11_2.C_ON=1'b0;
    defparam shift_srl_0_RNIVU6PD_15_LC_22_11_2.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIVU6PD_15_LC_22_11_2.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_0_RNIVU6PD_15_LC_22_11_2 (
            .in0(N__93553),
            .in1(N__89658),
            .in2(_gnd_net_),
            .in3(N__81553),
            .lcout(clk_en_54),
            .ltout(clk_en_54_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_57_RNIL56NE_15_LC_22_11_3.C_ON=1'b0;
    defparam shift_srl_57_RNIL56NE_15_LC_22_11_3.SEQ_MODE=4'b0000;
    defparam shift_srl_57_RNIL56NE_15_LC_22_11_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_57_RNIL56NE_15_LC_22_11_3 (
            .in0(N__76547),
            .in1(N__76939),
            .in2(N__76642),
            .in3(N__76795),
            .lcout(clk_en_58),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_55_LC_22_11_4.C_ON=1'b0;
    defparam rco_obuf_RNO_55_LC_22_11_4.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_55_LC_22_11_4.LUT_INIT=16'b1000100010001000;
    LogicCell40 rco_obuf_RNO_55_LC_22_11_4 (
            .in0(N__76940),
            .in1(N__77046),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(rco_c_55),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNII1LAH_15_LC_22_11_5.C_ON=1'b0;
    defparam shift_srl_0_RNII1LAH_15_LC_22_11_5.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNII1LAH_15_LC_22_11_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNII1LAH_15_LC_22_11_5 (
            .in0(N__81423),
            .in1(N__93552),
            .in2(N__89946),
            .in3(N__85004),
            .lcout(clk_en_67),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_56_RNI6FQG1_15_LC_22_11_6.C_ON=1'b0;
    defparam shift_srl_56_RNI6FQG1_15_LC_22_11_6.SEQ_MODE=4'b0000;
    defparam shift_srl_56_RNI6FQG1_15_LC_22_11_6.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_56_RNI6FQG1_15_LC_22_11_6 (
            .in0(N__76617),
            .in1(N__81552),
            .in2(N__76549),
            .in3(N__89659),
            .lcout(),
            .ltout(clk_en_0_a3_0_a2_sx_57_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_56_RNIU5DHE_15_LC_22_11_7.C_ON=1'b0;
    defparam shift_srl_56_RNIU5DHE_15_LC_22_11_7.SEQ_MODE=4'b0000;
    defparam shift_srl_56_RNIU5DHE_15_LC_22_11_7.LUT_INIT=16'b0000100000000000;
    LogicCell40 shift_srl_56_RNIU5DHE_15_LC_22_11_7 (
            .in0(N__76929),
            .in1(N__76911),
            .in2(N__76864),
            .in3(N__76857),
            .lcout(clk_en_57),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_57_0_LC_22_12_0.C_ON=1'b0;
    defparam shift_srl_57_0_LC_22_12_0.SEQ_MODE=4'b1000;
    defparam shift_srl_57_0_LC_22_12_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_57_0_LC_22_12_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76797),
            .lcout(shift_srl_57Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93276),
            .ce(N__76725),
            .sr(_gnd_net_));
    defparam shift_srl_57_1_LC_22_12_1.C_ON=1'b0;
    defparam shift_srl_57_1_LC_22_12_1.SEQ_MODE=4'b1000;
    defparam shift_srl_57_1_LC_22_12_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_57_1_LC_22_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76774),
            .lcout(shift_srl_57Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93276),
            .ce(N__76725),
            .sr(_gnd_net_));
    defparam shift_srl_57_2_LC_22_12_2.C_ON=1'b0;
    defparam shift_srl_57_2_LC_22_12_2.SEQ_MODE=4'b1000;
    defparam shift_srl_57_2_LC_22_12_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_57_2_LC_22_12_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76768),
            .lcout(shift_srl_57Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93276),
            .ce(N__76725),
            .sr(_gnd_net_));
    defparam shift_srl_57_3_LC_22_12_3.C_ON=1'b0;
    defparam shift_srl_57_3_LC_22_12_3.SEQ_MODE=4'b1000;
    defparam shift_srl_57_3_LC_22_12_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_57_3_LC_22_12_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76762),
            .lcout(shift_srl_57Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93276),
            .ce(N__76725),
            .sr(_gnd_net_));
    defparam shift_srl_57_4_LC_22_12_4.C_ON=1'b0;
    defparam shift_srl_57_4_LC_22_12_4.SEQ_MODE=4'b1000;
    defparam shift_srl_57_4_LC_22_12_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_57_4_LC_22_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76756),
            .lcout(shift_srl_57Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93276),
            .ce(N__76725),
            .sr(_gnd_net_));
    defparam shift_srl_57_5_LC_22_12_5.C_ON=1'b0;
    defparam shift_srl_57_5_LC_22_12_5.SEQ_MODE=4'b1000;
    defparam shift_srl_57_5_LC_22_12_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_57_5_LC_22_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76750),
            .lcout(shift_srl_57Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93276),
            .ce(N__76725),
            .sr(_gnd_net_));
    defparam shift_srl_57_6_LC_22_12_6.C_ON=1'b0;
    defparam shift_srl_57_6_LC_22_12_6.SEQ_MODE=4'b1000;
    defparam shift_srl_57_6_LC_22_12_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_57_6_LC_22_12_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76744),
            .lcout(shift_srl_57Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93276),
            .ce(N__76725),
            .sr(_gnd_net_));
    defparam shift_srl_57_7_LC_22_12_7.C_ON=1'b0;
    defparam shift_srl_57_7_LC_22_12_7.SEQ_MODE=4'b1000;
    defparam shift_srl_57_7_LC_22_12_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_57_7_LC_22_12_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76738),
            .lcout(shift_srl_57Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93276),
            .ce(N__76725),
            .sr(_gnd_net_));
    defparam shift_srl_48_RNI4JCOD_15_LC_22_13_0.C_ON=1'b0;
    defparam shift_srl_48_RNI4JCOD_15_LC_22_13_0.SEQ_MODE=4'b0000;
    defparam shift_srl_48_RNI4JCOD_15_LC_22_13_0.LUT_INIT=16'b0000000000100010;
    LogicCell40 shift_srl_48_RNI4JCOD_15_LC_22_13_0 (
            .in0(N__85215),
            .in1(N__77098),
            .in2(_gnd_net_),
            .in3(N__85265),
            .lcout(rco_c_53),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_54_0_LC_22_13_3.C_ON=1'b0;
    defparam shift_srl_54_0_LC_22_13_3.SEQ_MODE=4'b1000;
    defparam shift_srl_54_0_LC_22_13_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_54_0_LC_22_13_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77013),
            .lcout(shift_srl_54Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93257),
            .ce(N__87187),
            .sr(_gnd_net_));
    defparam shift_srl_54_1_LC_22_13_4.C_ON=1'b0;
    defparam shift_srl_54_1_LC_22_13_4.SEQ_MODE=4'b1000;
    defparam shift_srl_54_1_LC_22_13_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_54_1_LC_22_13_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76981),
            .lcout(shift_srl_54Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93257),
            .ce(N__87187),
            .sr(_gnd_net_));
    defparam shift_srl_54_2_LC_22_13_5.C_ON=1'b0;
    defparam shift_srl_54_2_LC_22_13_5.SEQ_MODE=4'b1000;
    defparam shift_srl_54_2_LC_22_13_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_54_2_LC_22_13_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76975),
            .lcout(shift_srl_54Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93257),
            .ce(N__87187),
            .sr(_gnd_net_));
    defparam shift_srl_54_3_LC_22_13_6.C_ON=1'b0;
    defparam shift_srl_54_3_LC_22_13_6.SEQ_MODE=4'b1000;
    defparam shift_srl_54_3_LC_22_13_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_54_3_LC_22_13_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76969),
            .lcout(shift_srl_54Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93257),
            .ce(N__87187),
            .sr(_gnd_net_));
    defparam shift_srl_54_4_LC_22_13_7.C_ON=1'b0;
    defparam shift_srl_54_4_LC_22_13_7.SEQ_MODE=4'b1000;
    defparam shift_srl_54_4_LC_22_13_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_54_4_LC_22_13_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76963),
            .lcout(shift_srl_54Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93257),
            .ce(N__87187),
            .sr(_gnd_net_));
    defparam shift_srl_64_10_LC_22_14_0.C_ON=1'b0;
    defparam shift_srl_64_10_LC_22_14_0.SEQ_MODE=4'b1000;
    defparam shift_srl_64_10_LC_22_14_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_64_10_LC_22_14_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77128),
            .lcout(shift_srl_64Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93235),
            .ce(N__79102),
            .sr(_gnd_net_));
    defparam shift_srl_64_11_LC_22_14_1.C_ON=1'b0;
    defparam shift_srl_64_11_LC_22_14_1.SEQ_MODE=4'b1000;
    defparam shift_srl_64_11_LC_22_14_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_64_11_LC_22_14_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76957),
            .lcout(shift_srl_64Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93235),
            .ce(N__79102),
            .sr(_gnd_net_));
    defparam shift_srl_64_12_LC_22_14_2.C_ON=1'b0;
    defparam shift_srl_64_12_LC_22_14_2.SEQ_MODE=4'b1000;
    defparam shift_srl_64_12_LC_22_14_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_64_12_LC_22_14_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76951),
            .lcout(shift_srl_64Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93235),
            .ce(N__79102),
            .sr(_gnd_net_));
    defparam shift_srl_64_13_LC_22_14_3.C_ON=1'b0;
    defparam shift_srl_64_13_LC_22_14_3.SEQ_MODE=4'b1000;
    defparam shift_srl_64_13_LC_22_14_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_64_13_LC_22_14_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77146),
            .lcout(shift_srl_64Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93235),
            .ce(N__79102),
            .sr(_gnd_net_));
    defparam shift_srl_64_14_LC_22_14_4.C_ON=1'b0;
    defparam shift_srl_64_14_LC_22_14_4.SEQ_MODE=4'b1000;
    defparam shift_srl_64_14_LC_22_14_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_64_14_LC_22_14_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77140),
            .lcout(shift_srl_64Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93235),
            .ce(N__79102),
            .sr(_gnd_net_));
    defparam shift_srl_64_15_LC_22_14_5.C_ON=1'b0;
    defparam shift_srl_64_15_LC_22_14_5.SEQ_MODE=4'b1000;
    defparam shift_srl_64_15_LC_22_14_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_64_15_LC_22_14_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77134),
            .lcout(shift_srl_64Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93235),
            .ce(N__79102),
            .sr(_gnd_net_));
    defparam shift_srl_64_9_LC_22_14_6.C_ON=1'b0;
    defparam shift_srl_64_9_LC_22_14_6.SEQ_MODE=4'b1000;
    defparam shift_srl_64_9_LC_22_14_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_64_9_LC_22_14_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77122),
            .lcout(shift_srl_64Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93235),
            .ce(N__79102),
            .sr(_gnd_net_));
    defparam shift_srl_64_8_LC_22_14_7.C_ON=1'b0;
    defparam shift_srl_64_8_LC_22_14_7.SEQ_MODE=4'b1000;
    defparam shift_srl_64_8_LC_22_14_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_64_8_LC_22_14_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79108),
            .lcout(shift_srl_64Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93235),
            .ce(N__79102),
            .sr(_gnd_net_));
    defparam shift_srl_65_10_LC_22_15_0.C_ON=1'b0;
    defparam shift_srl_65_10_LC_22_15_0.SEQ_MODE=4'b1000;
    defparam shift_srl_65_10_LC_22_15_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_65_10_LC_22_15_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77182),
            .lcout(shift_srl_65Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93217),
            .ce(N__79786),
            .sr(_gnd_net_));
    defparam shift_srl_65_11_LC_22_15_1.C_ON=1'b0;
    defparam shift_srl_65_11_LC_22_15_1.SEQ_MODE=4'b1000;
    defparam shift_srl_65_11_LC_22_15_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_65_11_LC_22_15_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77116),
            .lcout(shift_srl_65Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93217),
            .ce(N__79786),
            .sr(_gnd_net_));
    defparam shift_srl_65_12_LC_22_15_2.C_ON=1'b0;
    defparam shift_srl_65_12_LC_22_15_2.SEQ_MODE=4'b1000;
    defparam shift_srl_65_12_LC_22_15_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_65_12_LC_22_15_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77110),
            .lcout(shift_srl_65Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93217),
            .ce(N__79786),
            .sr(_gnd_net_));
    defparam shift_srl_65_13_LC_22_15_3.C_ON=1'b0;
    defparam shift_srl_65_13_LC_22_15_3.SEQ_MODE=4'b1000;
    defparam shift_srl_65_13_LC_22_15_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_65_13_LC_22_15_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77104),
            .lcout(shift_srl_65Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93217),
            .ce(N__79786),
            .sr(_gnd_net_));
    defparam shift_srl_65_14_LC_22_15_4.C_ON=1'b0;
    defparam shift_srl_65_14_LC_22_15_4.SEQ_MODE=4'b1000;
    defparam shift_srl_65_14_LC_22_15_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_65_14_LC_22_15_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77194),
            .lcout(shift_srl_65Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93217),
            .ce(N__79786),
            .sr(_gnd_net_));
    defparam shift_srl_65_15_LC_22_15_5.C_ON=1'b0;
    defparam shift_srl_65_15_LC_22_15_5.SEQ_MODE=4'b1000;
    defparam shift_srl_65_15_LC_22_15_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_65_15_LC_22_15_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77188),
            .lcout(shift_srl_65Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93217),
            .ce(N__79786),
            .sr(_gnd_net_));
    defparam shift_srl_65_9_LC_22_15_6.C_ON=1'b0;
    defparam shift_srl_65_9_LC_22_15_6.SEQ_MODE=4'b1000;
    defparam shift_srl_65_9_LC_22_15_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_65_9_LC_22_15_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77176),
            .lcout(shift_srl_65Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93217),
            .ce(N__79786),
            .sr(_gnd_net_));
    defparam shift_srl_65_8_LC_22_15_7.C_ON=1'b0;
    defparam shift_srl_65_8_LC_22_15_7.SEQ_MODE=4'b1000;
    defparam shift_srl_65_8_LC_22_15_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_65_8_LC_22_15_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79792),
            .lcout(shift_srl_65Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93217),
            .ce(N__79786),
            .sr(_gnd_net_));
    defparam shift_srl_63_8_LC_22_16_0.C_ON=1'b0;
    defparam shift_srl_63_8_LC_22_16_0.SEQ_MODE=4'b1000;
    defparam shift_srl_63_8_LC_22_16_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_63_8_LC_22_16_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77170),
            .lcout(shift_srl_63Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93196),
            .ce(N__79191),
            .sr(_gnd_net_));
    defparam shift_srl_63_9_LC_22_16_1.C_ON=1'b0;
    defparam shift_srl_63_9_LC_22_16_1.SEQ_MODE=4'b1000;
    defparam shift_srl_63_9_LC_22_16_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_63_9_LC_22_16_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77164),
            .lcout(shift_srl_63Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93196),
            .ce(N__79191),
            .sr(_gnd_net_));
    defparam shift_srl_31_0_LC_22_17_0.C_ON=1'b0;
    defparam shift_srl_31_0_LC_22_17_0.SEQ_MODE=4'b1000;
    defparam shift_srl_31_0_LC_22_17_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_31_0_LC_22_17_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83651),
            .lcout(shift_srl_31Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93154),
            .ce(N__79893),
            .sr(_gnd_net_));
    defparam shift_srl_31_1_LC_22_17_1.C_ON=1'b0;
    defparam shift_srl_31_1_LC_22_17_1.SEQ_MODE=4'b1000;
    defparam shift_srl_31_1_LC_22_17_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_31_1_LC_22_17_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77158),
            .lcout(shift_srl_31Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93154),
            .ce(N__79893),
            .sr(_gnd_net_));
    defparam shift_srl_31_2_LC_22_17_2.C_ON=1'b0;
    defparam shift_srl_31_2_LC_22_17_2.SEQ_MODE=4'b1000;
    defparam shift_srl_31_2_LC_22_17_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_31_2_LC_22_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77152),
            .lcout(shift_srl_31Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93154),
            .ce(N__79893),
            .sr(_gnd_net_));
    defparam shift_srl_31_3_LC_22_17_3.C_ON=1'b0;
    defparam shift_srl_31_3_LC_22_17_3.SEQ_MODE=4'b1000;
    defparam shift_srl_31_3_LC_22_17_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_31_3_LC_22_17_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77248),
            .lcout(shift_srl_31Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93154),
            .ce(N__79893),
            .sr(_gnd_net_));
    defparam shift_srl_31_4_LC_22_17_4.C_ON=1'b0;
    defparam shift_srl_31_4_LC_22_17_4.SEQ_MODE=4'b1000;
    defparam shift_srl_31_4_LC_22_17_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_31_4_LC_22_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77242),
            .lcout(shift_srl_31Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93154),
            .ce(N__79893),
            .sr(_gnd_net_));
    defparam shift_srl_31_5_LC_22_17_5.C_ON=1'b0;
    defparam shift_srl_31_5_LC_22_17_5.SEQ_MODE=4'b1000;
    defparam shift_srl_31_5_LC_22_17_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_31_5_LC_22_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77236),
            .lcout(shift_srl_31Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93154),
            .ce(N__79893),
            .sr(_gnd_net_));
    defparam shift_srl_31_6_LC_22_17_6.C_ON=1'b0;
    defparam shift_srl_31_6_LC_22_17_6.SEQ_MODE=4'b1000;
    defparam shift_srl_31_6_LC_22_17_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_31_6_LC_22_17_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77230),
            .lcout(shift_srl_31Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93154),
            .ce(N__79893),
            .sr(_gnd_net_));
    defparam shift_srl_31_7_LC_22_17_7.C_ON=1'b0;
    defparam shift_srl_31_7_LC_22_17_7.SEQ_MODE=4'b1000;
    defparam shift_srl_31_7_LC_22_17_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_31_7_LC_22_17_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77224),
            .lcout(shift_srl_31Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93154),
            .ce(N__79893),
            .sr(_gnd_net_));
    defparam shift_srl_31_10_LC_22_18_0.C_ON=1'b0;
    defparam shift_srl_31_10_LC_22_18_0.SEQ_MODE=4'b1000;
    defparam shift_srl_31_10_LC_22_18_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_31_10_LC_22_18_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77455),
            .lcout(shift_srl_31Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93197),
            .ce(N__79897),
            .sr(_gnd_net_));
    defparam shift_srl_31_11_LC_22_18_1.C_ON=1'b0;
    defparam shift_srl_31_11_LC_22_18_1.SEQ_MODE=4'b1000;
    defparam shift_srl_31_11_LC_22_18_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_31_11_LC_22_18_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77218),
            .lcout(shift_srl_31Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93197),
            .ce(N__79897),
            .sr(_gnd_net_));
    defparam shift_srl_31_12_LC_22_18_2.C_ON=1'b0;
    defparam shift_srl_31_12_LC_22_18_2.SEQ_MODE=4'b1000;
    defparam shift_srl_31_12_LC_22_18_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_31_12_LC_22_18_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77212),
            .lcout(shift_srl_31Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93197),
            .ce(N__79897),
            .sr(_gnd_net_));
    defparam shift_srl_31_13_LC_22_18_3.C_ON=1'b0;
    defparam shift_srl_31_13_LC_22_18_3.SEQ_MODE=4'b1000;
    defparam shift_srl_31_13_LC_22_18_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_31_13_LC_22_18_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77206),
            .lcout(shift_srl_31Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93197),
            .ce(N__79897),
            .sr(_gnd_net_));
    defparam shift_srl_31_14_LC_22_18_4.C_ON=1'b0;
    defparam shift_srl_31_14_LC_22_18_4.SEQ_MODE=4'b1000;
    defparam shift_srl_31_14_LC_22_18_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_31_14_LC_22_18_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77200),
            .lcout(shift_srl_31Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93197),
            .ce(N__79897),
            .sr(_gnd_net_));
    defparam shift_srl_31_15_LC_22_18_5.C_ON=1'b0;
    defparam shift_srl_31_15_LC_22_18_5.SEQ_MODE=4'b1000;
    defparam shift_srl_31_15_LC_22_18_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_31_15_LC_22_18_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77461),
            .lcout(shift_srl_31Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93197),
            .ce(N__79897),
            .sr(_gnd_net_));
    defparam shift_srl_31_9_LC_22_18_6.C_ON=1'b0;
    defparam shift_srl_31_9_LC_22_18_6.SEQ_MODE=4'b1000;
    defparam shift_srl_31_9_LC_22_18_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_31_9_LC_22_18_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77443),
            .lcout(shift_srl_31Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93197),
            .ce(N__79897),
            .sr(_gnd_net_));
    defparam shift_srl_31_8_LC_22_18_7.C_ON=1'b0;
    defparam shift_srl_31_8_LC_22_18_7.SEQ_MODE=4'b1000;
    defparam shift_srl_31_8_LC_22_18_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_31_8_LC_22_18_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77449),
            .lcout(shift_srl_31Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93197),
            .ce(N__79897),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNI0BOF91_15_LC_22_19_0.C_ON=1'b0;
    defparam shift_srl_0_RNI0BOF91_15_LC_22_19_0.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNI0BOF91_15_LC_22_19_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNI0BOF91_15_LC_22_19_0 (
            .in0(N__90389),
            .in1(N__87960),
            .in2(N__82425),
            .in3(N__87879),
            .lcout(clk_en_165),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_159_RNIT5G61_15_LC_22_19_1.C_ON=1'b0;
    defparam shift_srl_159_RNIT5G61_15_LC_22_19_1.SEQ_MODE=4'b0000;
    defparam shift_srl_159_RNIT5G61_15_LC_22_19_1.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_159_RNIT5G61_15_LC_22_19_1 (
            .in0(N__77300),
            .in1(N__77279),
            .in2(N__77437),
            .in3(N__77872),
            .lcout(),
            .ltout(rco_int_0_a3_0_a2_0_sx_162_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_162_RNIMG202_15_LC_22_19_2.C_ON=1'b0;
    defparam shift_srl_162_RNIMG202_15_LC_22_19_2.SEQ_MODE=4'b0000;
    defparam shift_srl_162_RNIMG202_15_LC_22_19_2.LUT_INIT=16'b0000100000000000;
    LogicCell40 shift_srl_162_RNIMG202_15_LC_22_19_2 (
            .in0(N__77398),
            .in1(N__77376),
            .in2(N__77323),
            .in3(N__77519),
            .lcout(rco_int_0_a3_0_a2_0_162),
            .ltout(rco_int_0_a3_0_a2_0_162_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIGB2MA1_15_LC_22_19_3.C_ON=1'b0;
    defparam shift_srl_0_RNIGB2MA1_15_LC_22_19_3.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIGB2MA1_15_LC_22_19_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNIGB2MA1_15_LC_22_19_3 (
            .in0(N__87880),
            .in1(N__90391),
            .in2(N__77320),
            .in3(N__87466),
            .lcout(clk_en_171),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_159_15_LC_22_19_4.C_ON=1'b0;
    defparam shift_srl_159_15_LC_22_19_4.SEQ_MODE=4'b1000;
    defparam shift_srl_159_15_LC_22_19_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_159_15_LC_22_19_4 (
            .in0(N__77317),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_159Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93218),
            .ce(N__77706),
            .sr(_gnd_net_));
    defparam shift_srl_158_RNIKL9G2_15_LC_22_19_5.C_ON=1'b0;
    defparam shift_srl_158_RNIKL9G2_15_LC_22_19_5.SEQ_MODE=4'b0000;
    defparam shift_srl_158_RNIKL9G2_15_LC_22_19_5.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_158_RNIKL9G2_15_LC_22_19_5 (
            .in0(N__77284),
            .in1(N__90390),
            .in2(N__77908),
            .in3(N__82340),
            .lcout(),
            .ltout(clk_en_0_a3_0_a2_sx_159_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_158_RNI2L4181_15_LC_22_19_6.C_ON=1'b0;
    defparam shift_srl_158_RNI2L4181_15_LC_22_19_6.SEQ_MODE=4'b0000;
    defparam shift_srl_158_RNI2L4181_15_LC_22_19_6.LUT_INIT=16'b0000100000000000;
    LogicCell40 shift_srl_158_RNI2L4181_15_LC_22_19_6 (
            .in0(N__77529),
            .in1(N__77804),
            .in2(N__77710),
            .in3(N__79391),
            .lcout(clk_en_159),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_156_RNII4IK_15_LC_22_19_7.C_ON=1'b0;
    defparam shift_srl_156_RNII4IK_15_LC_22_19_7.SEQ_MODE=4'b0000;
    defparam shift_srl_156_RNII4IK_15_LC_22_19_7.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_156_RNII4IK_15_LC_22_19_7 (
            .in0(N__77674),
            .in1(N__77651),
            .in2(_gnd_net_),
            .in3(N__77607),
            .lcout(shift_srl_156_RNII4IKZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_171_10_LC_22_20_0.C_ON=1'b0;
    defparam shift_srl_171_10_LC_22_20_0.SEQ_MODE=4'b1000;
    defparam shift_srl_171_10_LC_22_20_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_171_10_LC_22_20_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77974),
            .lcout(shift_srl_171Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93236),
            .ce(N__77955),
            .sr(_gnd_net_));
    defparam shift_srl_171_11_LC_22_20_1.C_ON=1'b0;
    defparam shift_srl_171_11_LC_22_20_1.SEQ_MODE=4'b1000;
    defparam shift_srl_171_11_LC_22_20_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_171_11_LC_22_20_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77491),
            .lcout(shift_srl_171Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93236),
            .ce(N__77955),
            .sr(_gnd_net_));
    defparam shift_srl_171_12_LC_22_20_2.C_ON=1'b0;
    defparam shift_srl_171_12_LC_22_20_2.SEQ_MODE=4'b1000;
    defparam shift_srl_171_12_LC_22_20_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_171_12_LC_22_20_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77485),
            .lcout(shift_srl_171Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93236),
            .ce(N__77955),
            .sr(_gnd_net_));
    defparam shift_srl_171_13_LC_22_20_3.C_ON=1'b0;
    defparam shift_srl_171_13_LC_22_20_3.SEQ_MODE=4'b1000;
    defparam shift_srl_171_13_LC_22_20_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_171_13_LC_22_20_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77479),
            .lcout(shift_srl_171Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93236),
            .ce(N__77955),
            .sr(_gnd_net_));
    defparam shift_srl_171_14_LC_22_20_4.C_ON=1'b0;
    defparam shift_srl_171_14_LC_22_20_4.SEQ_MODE=4'b1000;
    defparam shift_srl_171_14_LC_22_20_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_171_14_LC_22_20_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77473),
            .lcout(shift_srl_171Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93236),
            .ce(N__77955),
            .sr(_gnd_net_));
    defparam shift_srl_171_15_LC_22_20_5.C_ON=1'b0;
    defparam shift_srl_171_15_LC_22_20_5.SEQ_MODE=4'b1000;
    defparam shift_srl_171_15_LC_22_20_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_171_15_LC_22_20_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77467),
            .lcout(shift_srl_171Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93236),
            .ce(N__77955),
            .sr(_gnd_net_));
    defparam shift_srl_171_9_LC_22_20_6.C_ON=1'b0;
    defparam shift_srl_171_9_LC_22_20_6.SEQ_MODE=4'b1000;
    defparam shift_srl_171_9_LC_22_20_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_171_9_LC_22_20_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77980),
            .lcout(shift_srl_171Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93236),
            .ce(N__77955),
            .sr(_gnd_net_));
    defparam shift_srl_171_1_LC_22_20_7.C_ON=1'b0;
    defparam shift_srl_171_1_LC_22_20_7.SEQ_MODE=4'b1000;
    defparam shift_srl_171_1_LC_22_20_7.LUT_INIT=16'b1100110011001100;
    LogicCell40 shift_srl_171_1_LC_22_20_7 (
            .in0(_gnd_net_),
            .in1(N__77968),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_171Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93236),
            .ce(N__77955),
            .sr(_gnd_net_));
    defparam shift_srl_179_10_LC_22_21_0.C_ON=1'b0;
    defparam shift_srl_179_10_LC_22_21_0.SEQ_MODE=4'b1000;
    defparam shift_srl_179_10_LC_22_21_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_179_10_LC_22_21_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77914),
            .lcout(shift_srl_179Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93258),
            .ce(N__78061),
            .sr(_gnd_net_));
    defparam shift_srl_179_11_LC_22_21_1.C_ON=1'b0;
    defparam shift_srl_179_11_LC_22_21_1.SEQ_MODE=4'b1000;
    defparam shift_srl_179_11_LC_22_21_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_179_11_LC_22_21_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77944),
            .lcout(shift_srl_179Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93258),
            .ce(N__78061),
            .sr(_gnd_net_));
    defparam shift_srl_179_12_LC_22_21_2.C_ON=1'b0;
    defparam shift_srl_179_12_LC_22_21_2.SEQ_MODE=4'b1000;
    defparam shift_srl_179_12_LC_22_21_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_179_12_LC_22_21_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77938),
            .lcout(shift_srl_179Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93258),
            .ce(N__78061),
            .sr(_gnd_net_));
    defparam shift_srl_179_13_LC_22_21_3.C_ON=1'b0;
    defparam shift_srl_179_13_LC_22_21_3.SEQ_MODE=4'b1000;
    defparam shift_srl_179_13_LC_22_21_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_179_13_LC_22_21_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77932),
            .lcout(shift_srl_179Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93258),
            .ce(N__78061),
            .sr(_gnd_net_));
    defparam shift_srl_179_14_LC_22_21_4.C_ON=1'b0;
    defparam shift_srl_179_14_LC_22_21_4.SEQ_MODE=4'b1000;
    defparam shift_srl_179_14_LC_22_21_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_179_14_LC_22_21_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77926),
            .lcout(shift_srl_179Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93258),
            .ce(N__78061),
            .sr(_gnd_net_));
    defparam shift_srl_179_15_LC_22_21_5.C_ON=1'b0;
    defparam shift_srl_179_15_LC_22_21_5.SEQ_MODE=4'b1000;
    defparam shift_srl_179_15_LC_22_21_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_179_15_LC_22_21_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77920),
            .lcout(shift_srl_179Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93258),
            .ce(N__78061),
            .sr(_gnd_net_));
    defparam shift_srl_179_9_LC_22_21_6.C_ON=1'b0;
    defparam shift_srl_179_9_LC_22_21_6.SEQ_MODE=4'b1000;
    defparam shift_srl_179_9_LC_22_21_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_179_9_LC_22_21_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78067),
            .lcout(shift_srl_179Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93258),
            .ce(N__78061),
            .sr(_gnd_net_));
    defparam shift_srl_179_8_LC_22_21_7.C_ON=1'b0;
    defparam shift_srl_179_8_LC_22_21_7.SEQ_MODE=4'b1000;
    defparam shift_srl_179_8_LC_22_21_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_179_8_LC_22_21_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78073),
            .lcout(shift_srl_179Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93258),
            .ce(N__78061),
            .sr(_gnd_net_));
    defparam shift_srl_178_6_LC_22_22_0.C_ON=1'b0;
    defparam shift_srl_178_6_LC_22_22_0.SEQ_MODE=4'b1000;
    defparam shift_srl_178_6_LC_22_22_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_178_6_LC_22_22_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78034),
            .lcout(shift_srl_178Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93277),
            .ce(N__78106),
            .sr(_gnd_net_));
    defparam shift_srl_178_11_LC_22_22_1.C_ON=1'b0;
    defparam shift_srl_178_11_LC_22_22_1.SEQ_MODE=4'b1000;
    defparam shift_srl_178_11_LC_22_22_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_178_11_LC_22_22_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78028),
            .lcout(shift_srl_178Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93277),
            .ce(N__78106),
            .sr(_gnd_net_));
    defparam shift_srl_178_12_LC_22_22_2.C_ON=1'b0;
    defparam shift_srl_178_12_LC_22_22_2.SEQ_MODE=4'b1000;
    defparam shift_srl_178_12_LC_22_22_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_178_12_LC_22_22_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78022),
            .lcout(shift_srl_178Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93277),
            .ce(N__78106),
            .sr(_gnd_net_));
    defparam shift_srl_178_13_LC_22_22_3.C_ON=1'b0;
    defparam shift_srl_178_13_LC_22_22_3.SEQ_MODE=4'b1000;
    defparam shift_srl_178_13_LC_22_22_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_178_13_LC_22_22_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78016),
            .lcout(shift_srl_178Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93277),
            .ce(N__78106),
            .sr(_gnd_net_));
    defparam shift_srl_178_7_LC_22_22_4.C_ON=1'b0;
    defparam shift_srl_178_7_LC_22_22_4.SEQ_MODE=4'b1000;
    defparam shift_srl_178_7_LC_22_22_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_178_7_LC_22_22_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78010),
            .lcout(shift_srl_178Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93277),
            .ce(N__78106),
            .sr(_gnd_net_));
    defparam shift_srl_178_15_LC_22_22_5.C_ON=1'b0;
    defparam shift_srl_178_15_LC_22_22_5.SEQ_MODE=4'b1000;
    defparam shift_srl_178_15_LC_22_22_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_178_15_LC_22_22_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77998),
            .lcout(shift_srl_178Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93277),
            .ce(N__78106),
            .sr(_gnd_net_));
    defparam shift_srl_178_14_LC_22_22_6.C_ON=1'b0;
    defparam shift_srl_178_14_LC_22_22_6.SEQ_MODE=4'b1000;
    defparam shift_srl_178_14_LC_22_22_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_178_14_LC_22_22_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78004),
            .lcout(shift_srl_178Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93277),
            .ce(N__78106),
            .sr(_gnd_net_));
    defparam shift_srl_178_8_LC_22_22_7.C_ON=1'b0;
    defparam shift_srl_178_8_LC_22_22_7.SEQ_MODE=4'b1000;
    defparam shift_srl_178_8_LC_22_22_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_178_8_LC_22_22_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77992),
            .lcout(shift_srl_178Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93277),
            .ce(N__78106),
            .sr(_gnd_net_));
    defparam shift_srl_179_RNIVNOT1_15_LC_22_23_0.C_ON=1'b0;
    defparam shift_srl_179_RNIVNOT1_15_LC_22_23_0.SEQ_MODE=4'b0000;
    defparam shift_srl_179_RNIVNOT1_15_LC_22_23_0.LUT_INIT=16'b0000100000000000;
    LogicCell40 shift_srl_179_RNIVNOT1_15_LC_22_23_0 (
            .in0(N__78133),
            .in1(N__80401),
            .in2(N__78187),
            .in3(N__80450),
            .lcout(shift_srl_179_RNIVNOT1Z0Z_15),
            .ltout(shift_srl_179_RNIVNOT1Z0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIOJFDD1_15_LC_22_23_1.C_ON=1'b0;
    defparam shift_srl_0_RNIOJFDD1_15_LC_22_23_1.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIOJFDD1_15_LC_22_23_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNIOJFDD1_15_LC_22_23_1 (
            .in0(N__84212),
            .in1(N__90452),
            .in2(N__78175),
            .in3(N__87670),
            .lcout(clk_en_180),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNINC9LC1_15_LC_22_23_2.C_ON=1'b0;
    defparam shift_srl_0_RNINC9LC1_15_LC_22_23_2.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNINC9LC1_15_LC_22_23_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNINC9LC1_15_LC_22_23_2 (
            .in0(N__90450),
            .in1(N__84211),
            .in2(N__80543),
            .in3(N__87669),
            .lcout(clk_en_177),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_180_RNISQAED1_15_LC_22_23_3.C_ON=1'b0;
    defparam shift_srl_180_RNISQAED1_15_LC_22_23_3.SEQ_MODE=4'b0000;
    defparam shift_srl_180_RNISQAED1_15_LC_22_23_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_180_RNISQAED1_15_LC_22_23_3 (
            .in0(N__90141),
            .in1(N__78159),
            .in2(N__85985),
            .in3(N__82742),
            .lcout(clk_en_181),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_179_RNI5E1P_15_LC_22_23_4.C_ON=1'b0;
    defparam shift_srl_179_RNI5E1P_15_LC_22_23_4.SEQ_MODE=4'b0000;
    defparam shift_srl_179_RNI5E1P_15_LC_22_23_4.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_179_RNI5E1P_15_LC_22_23_4 (
            .in0(N__78132),
            .in1(N__80400),
            .in2(N__82750),
            .in3(N__80449),
            .lcout(rco_int_0_a2_1_a2_0_sx_182),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_177_15_LC_22_23_5.C_ON=1'b0;
    defparam shift_srl_177_15_LC_22_23_5.SEQ_MODE=4'b1000;
    defparam shift_srl_177_15_LC_22_23_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_177_15_LC_22_23_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78085),
            .lcout(shift_srl_177Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93291),
            .ce(N__82598),
            .sr(_gnd_net_));
    defparam shift_srl_177_RNI1B5PC1_15_LC_22_23_6.C_ON=1'b0;
    defparam shift_srl_177_RNI1B5PC1_15_LC_22_23_6.SEQ_MODE=4'b0000;
    defparam shift_srl_177_RNI1B5PC1_15_LC_22_23_6.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_177_RNI1B5PC1_15_LC_22_23_6 (
            .in0(N__90451),
            .in1(N__80451),
            .in2(N__80544),
            .in3(N__85964),
            .lcout(clk_en_178),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_177_14_LC_22_23_7.C_ON=1'b0;
    defparam shift_srl_177_14_LC_22_23_7.SEQ_MODE=4'b1000;
    defparam shift_srl_177_14_LC_22_23_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_177_14_LC_22_23_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80257),
            .lcout(shift_srl_177Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93291),
            .ce(N__82598),
            .sr(_gnd_net_));
    defparam shift_srl_181_10_LC_22_24_0.C_ON=1'b0;
    defparam shift_srl_181_10_LC_22_24_0.SEQ_MODE=4'b1000;
    defparam shift_srl_181_10_LC_22_24_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_181_10_LC_22_24_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78229),
            .lcout(shift_srl_181Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93310),
            .ce(N__78210),
            .sr(_gnd_net_));
    defparam shift_srl_181_11_LC_22_24_1.C_ON=1'b0;
    defparam shift_srl_181_11_LC_22_24_1.SEQ_MODE=4'b1000;
    defparam shift_srl_181_11_LC_22_24_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_181_11_LC_22_24_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78079),
            .lcout(shift_srl_181Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93310),
            .ce(N__78210),
            .sr(_gnd_net_));
    defparam shift_srl_181_12_LC_22_24_2.C_ON=1'b0;
    defparam shift_srl_181_12_LC_22_24_2.SEQ_MODE=4'b1000;
    defparam shift_srl_181_12_LC_22_24_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_181_12_LC_22_24_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78259),
            .lcout(shift_srl_181Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93310),
            .ce(N__78210),
            .sr(_gnd_net_));
    defparam shift_srl_181_13_LC_22_24_3.C_ON=1'b0;
    defparam shift_srl_181_13_LC_22_24_3.SEQ_MODE=4'b1000;
    defparam shift_srl_181_13_LC_22_24_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_181_13_LC_22_24_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78253),
            .lcout(shift_srl_181Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93310),
            .ce(N__78210),
            .sr(_gnd_net_));
    defparam shift_srl_181_7_LC_22_24_4.C_ON=1'b0;
    defparam shift_srl_181_7_LC_22_24_4.SEQ_MODE=4'b1000;
    defparam shift_srl_181_7_LC_22_24_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_181_7_LC_22_24_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78247),
            .lcout(shift_srl_181Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93310),
            .ce(N__78210),
            .sr(_gnd_net_));
    defparam shift_srl_181_14_LC_22_24_5.C_ON=1'b0;
    defparam shift_srl_181_14_LC_22_24_5.SEQ_MODE=4'b1000;
    defparam shift_srl_181_14_LC_22_24_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_181_14_LC_22_24_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78241),
            .lcout(shift_srl_181Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93310),
            .ce(N__78210),
            .sr(_gnd_net_));
    defparam shift_srl_181_9_LC_22_24_6.C_ON=1'b0;
    defparam shift_srl_181_9_LC_22_24_6.SEQ_MODE=4'b1000;
    defparam shift_srl_181_9_LC_22_24_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_181_9_LC_22_24_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78217),
            .lcout(shift_srl_181Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93310),
            .ce(N__78210),
            .sr(_gnd_net_));
    defparam shift_srl_181_8_LC_22_24_7.C_ON=1'b0;
    defparam shift_srl_181_8_LC_22_24_7.SEQ_MODE=4'b1000;
    defparam shift_srl_181_8_LC_22_24_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_181_8_LC_22_24_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78223),
            .lcout(shift_srl_181Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93310),
            .ce(N__78210),
            .sr(_gnd_net_));
    defparam shift_srl_189_10_LC_22_25_0.C_ON=1'b0;
    defparam shift_srl_189_10_LC_22_25_0.SEQ_MODE=4'b1000;
    defparam shift_srl_189_10_LC_22_25_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_189_10_LC_22_25_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78289),
            .lcout(shift_srl_189Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93330),
            .ce(N__82846),
            .sr(_gnd_net_));
    defparam shift_srl_189_11_LC_22_25_1.C_ON=1'b0;
    defparam shift_srl_189_11_LC_22_25_1.SEQ_MODE=4'b1000;
    defparam shift_srl_189_11_LC_22_25_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_189_11_LC_22_25_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78199),
            .lcout(shift_srl_189Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93330),
            .ce(N__82846),
            .sr(_gnd_net_));
    defparam shift_srl_189_12_LC_22_25_2.C_ON=1'b0;
    defparam shift_srl_189_12_LC_22_25_2.SEQ_MODE=4'b1000;
    defparam shift_srl_189_12_LC_22_25_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_189_12_LC_22_25_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78193),
            .lcout(shift_srl_189Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93330),
            .ce(N__82846),
            .sr(_gnd_net_));
    defparam shift_srl_189_13_LC_22_25_3.C_ON=1'b0;
    defparam shift_srl_189_13_LC_22_25_3.SEQ_MODE=4'b1000;
    defparam shift_srl_189_13_LC_22_25_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_189_13_LC_22_25_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78307),
            .lcout(shift_srl_189Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93330),
            .ce(N__82846),
            .sr(_gnd_net_));
    defparam shift_srl_189_14_LC_22_25_4.C_ON=1'b0;
    defparam shift_srl_189_14_LC_22_25_4.SEQ_MODE=4'b1000;
    defparam shift_srl_189_14_LC_22_25_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_189_14_LC_22_25_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78301),
            .lcout(shift_srl_189Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93330),
            .ce(N__82846),
            .sr(_gnd_net_));
    defparam shift_srl_189_15_LC_22_25_5.C_ON=1'b0;
    defparam shift_srl_189_15_LC_22_25_5.SEQ_MODE=4'b1000;
    defparam shift_srl_189_15_LC_22_25_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_189_15_LC_22_25_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78295),
            .lcout(shift_srl_189Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93330),
            .ce(N__82846),
            .sr(_gnd_net_));
    defparam shift_srl_189_9_LC_22_25_6.C_ON=1'b0;
    defparam shift_srl_189_9_LC_22_25_6.SEQ_MODE=4'b1000;
    defparam shift_srl_189_9_LC_22_25_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_189_9_LC_22_25_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78283),
            .lcout(shift_srl_189Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93330),
            .ce(N__82846),
            .sr(_gnd_net_));
    defparam shift_srl_189_8_LC_22_25_7.C_ON=1'b0;
    defparam shift_srl_189_8_LC_22_25_7.SEQ_MODE=4'b1000;
    defparam shift_srl_189_8_LC_22_25_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_189_8_LC_22_25_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82855),
            .lcout(shift_srl_189Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93330),
            .ce(N__82846),
            .sr(_gnd_net_));
    defparam shift_srl_188_0_LC_22_26_0.C_ON=1'b0;
    defparam shift_srl_188_0_LC_22_26_0.SEQ_MODE=4'b1000;
    defparam shift_srl_188_0_LC_22_26_0.LUT_INIT=16'b1100110011001100;
    LogicCell40 shift_srl_188_0_LC_22_26_0 (
            .in0(_gnd_net_),
            .in1(N__86096),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_188Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93351),
            .ce(N__82797),
            .sr(_gnd_net_));
    defparam shift_srl_188_1_LC_22_26_1.C_ON=1'b0;
    defparam shift_srl_188_1_LC_22_26_1.SEQ_MODE=4'b1000;
    defparam shift_srl_188_1_LC_22_26_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_188_1_LC_22_26_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78277),
            .lcout(shift_srl_188Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93351),
            .ce(N__82797),
            .sr(_gnd_net_));
    defparam shift_srl_188_2_LC_22_26_2.C_ON=1'b0;
    defparam shift_srl_188_2_LC_22_26_2.SEQ_MODE=4'b1000;
    defparam shift_srl_188_2_LC_22_26_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_188_2_LC_22_26_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78271),
            .lcout(shift_srl_188Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93351),
            .ce(N__82797),
            .sr(_gnd_net_));
    defparam shift_srl_188_3_LC_22_26_3.C_ON=1'b0;
    defparam shift_srl_188_3_LC_22_26_3.SEQ_MODE=4'b1000;
    defparam shift_srl_188_3_LC_22_26_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_188_3_LC_22_26_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78265),
            .lcout(shift_srl_188Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93351),
            .ce(N__82797),
            .sr(_gnd_net_));
    defparam shift_srl_188_4_LC_22_26_4.C_ON=1'b0;
    defparam shift_srl_188_4_LC_22_26_4.SEQ_MODE=4'b1000;
    defparam shift_srl_188_4_LC_22_26_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_188_4_LC_22_26_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78376),
            .lcout(shift_srl_188Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93351),
            .ce(N__82797),
            .sr(_gnd_net_));
    defparam shift_srl_188_5_LC_22_26_5.C_ON=1'b0;
    defparam shift_srl_188_5_LC_22_26_5.SEQ_MODE=4'b1000;
    defparam shift_srl_188_5_LC_22_26_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_188_5_LC_22_26_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78370),
            .lcout(shift_srl_188Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93351),
            .ce(N__82797),
            .sr(_gnd_net_));
    defparam shift_srl_188_6_LC_22_26_6.C_ON=1'b0;
    defparam shift_srl_188_6_LC_22_26_6.SEQ_MODE=4'b1000;
    defparam shift_srl_188_6_LC_22_26_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_188_6_LC_22_26_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78364),
            .lcout(shift_srl_188Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93351),
            .ce(N__82797),
            .sr(_gnd_net_));
    defparam shift_srl_188_7_LC_22_26_7.C_ON=1'b0;
    defparam shift_srl_188_7_LC_22_26_7.SEQ_MODE=4'b1000;
    defparam shift_srl_188_7_LC_22_26_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_188_7_LC_22_26_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78358),
            .lcout(shift_srl_188Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93351),
            .ce(N__82797),
            .sr(_gnd_net_));
    defparam shift_srl_176_0_LC_22_27_0.C_ON=1'b0;
    defparam shift_srl_176_0_LC_22_27_0.SEQ_MODE=4'b1000;
    defparam shift_srl_176_0_LC_22_27_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_176_0_LC_22_27_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78351),
            .lcout(shift_srl_176Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93368),
            .ce(N__78532),
            .sr(_gnd_net_));
    defparam shift_srl_176_1_LC_22_27_1.C_ON=1'b0;
    defparam shift_srl_176_1_LC_22_27_1.SEQ_MODE=4'b1000;
    defparam shift_srl_176_1_LC_22_27_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_176_1_LC_22_27_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78331),
            .lcout(shift_srl_176Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93368),
            .ce(N__78532),
            .sr(_gnd_net_));
    defparam shift_srl_176_2_LC_22_27_2.C_ON=1'b0;
    defparam shift_srl_176_2_LC_22_27_2.SEQ_MODE=4'b1000;
    defparam shift_srl_176_2_LC_22_27_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_176_2_LC_22_27_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78325),
            .lcout(shift_srl_176Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93368),
            .ce(N__78532),
            .sr(_gnd_net_));
    defparam shift_srl_176_3_LC_22_27_3.C_ON=1'b0;
    defparam shift_srl_176_3_LC_22_27_3.SEQ_MODE=4'b1000;
    defparam shift_srl_176_3_LC_22_27_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_176_3_LC_22_27_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78319),
            .lcout(shift_srl_176Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93368),
            .ce(N__78532),
            .sr(_gnd_net_));
    defparam shift_srl_176_4_LC_22_27_4.C_ON=1'b0;
    defparam shift_srl_176_4_LC_22_27_4.SEQ_MODE=4'b1000;
    defparam shift_srl_176_4_LC_22_27_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_176_4_LC_22_27_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78313),
            .lcout(shift_srl_176Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93368),
            .ce(N__78532),
            .sr(_gnd_net_));
    defparam shift_srl_176_5_LC_22_27_5.C_ON=1'b0;
    defparam shift_srl_176_5_LC_22_27_5.SEQ_MODE=4'b1000;
    defparam shift_srl_176_5_LC_22_27_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_176_5_LC_22_27_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78559),
            .lcout(shift_srl_176Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93368),
            .ce(N__78532),
            .sr(_gnd_net_));
    defparam shift_srl_176_6_LC_22_27_6.C_ON=1'b0;
    defparam shift_srl_176_6_LC_22_27_6.SEQ_MODE=4'b1000;
    defparam shift_srl_176_6_LC_22_27_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_176_6_LC_22_27_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78553),
            .lcout(shift_srl_176Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93368),
            .ce(N__78532),
            .sr(_gnd_net_));
    defparam shift_srl_176_7_LC_22_27_7.C_ON=1'b0;
    defparam shift_srl_176_7_LC_22_27_7.SEQ_MODE=4'b1000;
    defparam shift_srl_176_7_LC_22_27_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_176_7_LC_22_27_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78547),
            .lcout(shift_srl_176Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93368),
            .ce(N__78532),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_121_LC_22_28_4.C_ON=1'b0;
    defparam rco_obuf_RNO_121_LC_22_28_4.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_121_LC_22_28_4.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_121_LC_22_28_4 (
            .in0(N__78520),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78478),
            .lcout(rco_c_121),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_177_LC_22_29_4.C_ON=1'b0;
    defparam rco_obuf_RNO_177_LC_22_29_4.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_177_LC_22_29_4.LUT_INIT=16'b1000100000000000;
    LogicCell40 rco_obuf_RNO_177_LC_22_29_4 (
            .in0(N__85969),
            .in1(N__80522),
            .in2(_gnd_net_),
            .in3(N__80474),
            .lcout(rco_c_177),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_83_4_LC_23_5_1.C_ON=1'b0;
    defparam shift_srl_83_4_LC_23_5_1.SEQ_MODE=4'b1000;
    defparam shift_srl_83_4_LC_23_5_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_83_4_LC_23_5_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78577),
            .lcout(shift_srl_83Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93403),
            .ce(N__80872),
            .sr(_gnd_net_));
    defparam shift_srl_83_12_LC_23_5_2.C_ON=1'b0;
    defparam shift_srl_83_12_LC_23_5_2.SEQ_MODE=4'b1000;
    defparam shift_srl_83_12_LC_23_5_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_83_12_LC_23_5_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78601),
            .lcout(shift_srl_83Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93403),
            .ce(N__80872),
            .sr(_gnd_net_));
    defparam shift_srl_83_13_LC_23_5_3.C_ON=1'b0;
    defparam shift_srl_83_13_LC_23_5_3.SEQ_MODE=4'b1000;
    defparam shift_srl_83_13_LC_23_5_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_83_13_LC_23_5_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78388),
            .lcout(shift_srl_83Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93403),
            .ce(N__80872),
            .sr(_gnd_net_));
    defparam shift_srl_83_14_LC_23_5_4.C_ON=1'b0;
    defparam shift_srl_83_14_LC_23_5_4.SEQ_MODE=4'b1000;
    defparam shift_srl_83_14_LC_23_5_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_83_14_LC_23_5_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78382),
            .lcout(shift_srl_83Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93403),
            .ce(N__80872),
            .sr(_gnd_net_));
    defparam shift_srl_83_15_LC_23_5_5.C_ON=1'b0;
    defparam shift_srl_83_15_LC_23_5_5.SEQ_MODE=4'b1000;
    defparam shift_srl_83_15_LC_23_5_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_83_15_LC_23_5_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78607),
            .lcout(shift_srl_83Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93403),
            .ce(N__80872),
            .sr(_gnd_net_));
    defparam shift_srl_83_11_LC_23_5_6.C_ON=1'b0;
    defparam shift_srl_83_11_LC_23_5_6.SEQ_MODE=4'b1000;
    defparam shift_srl_83_11_LC_23_5_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_83_11_LC_23_5_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80749),
            .lcout(shift_srl_83Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93403),
            .ce(N__80872),
            .sr(_gnd_net_));
    defparam shift_srl_83_8_LC_23_5_7.C_ON=1'b0;
    defparam shift_srl_83_8_LC_23_5_7.SEQ_MODE=4'b1000;
    defparam shift_srl_83_8_LC_23_5_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_83_8_LC_23_5_7 (
            .in0(N__78571),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_83Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93403),
            .ce(N__80872),
            .sr(_gnd_net_));
    defparam shift_srl_83_0_LC_23_6_0.C_ON=1'b0;
    defparam shift_srl_83_0_LC_23_6_0.SEQ_MODE=4'b1000;
    defparam shift_srl_83_0_LC_23_6_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_83_0_LC_23_6_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80799),
            .lcout(shift_srl_83Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93396),
            .ce(N__80864),
            .sr(_gnd_net_));
    defparam shift_srl_83_1_LC_23_6_1.C_ON=1'b0;
    defparam shift_srl_83_1_LC_23_6_1.SEQ_MODE=4'b1000;
    defparam shift_srl_83_1_LC_23_6_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_83_1_LC_23_6_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78595),
            .lcout(shift_srl_83Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93396),
            .ce(N__80864),
            .sr(_gnd_net_));
    defparam shift_srl_83_2_LC_23_6_2.C_ON=1'b0;
    defparam shift_srl_83_2_LC_23_6_2.SEQ_MODE=4'b1000;
    defparam shift_srl_83_2_LC_23_6_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_83_2_LC_23_6_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78589),
            .lcout(shift_srl_83Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93396),
            .ce(N__80864),
            .sr(_gnd_net_));
    defparam shift_srl_83_3_LC_23_6_3.C_ON=1'b0;
    defparam shift_srl_83_3_LC_23_6_3.SEQ_MODE=4'b1000;
    defparam shift_srl_83_3_LC_23_6_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_83_3_LC_23_6_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78583),
            .lcout(shift_srl_83Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93396),
            .ce(N__80864),
            .sr(_gnd_net_));
    defparam shift_srl_83_7_LC_23_6_4.C_ON=1'b0;
    defparam shift_srl_83_7_LC_23_6_4.SEQ_MODE=4'b1000;
    defparam shift_srl_83_7_LC_23_6_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_83_7_LC_23_6_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78655),
            .lcout(shift_srl_83Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93396),
            .ce(N__80864),
            .sr(_gnd_net_));
    defparam shift_srl_83_5_LC_23_6_5.C_ON=1'b0;
    defparam shift_srl_83_5_LC_23_6_5.SEQ_MODE=4'b1000;
    defparam shift_srl_83_5_LC_23_6_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_83_5_LC_23_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78565),
            .lcout(shift_srl_83Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93396),
            .ce(N__80864),
            .sr(_gnd_net_));
    defparam shift_srl_83_6_LC_23_6_6.C_ON=1'b0;
    defparam shift_srl_83_6_LC_23_6_6.SEQ_MODE=4'b1000;
    defparam shift_srl_83_6_LC_23_6_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_83_6_LC_23_6_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78661),
            .lcout(shift_srl_83Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93396),
            .ce(N__80864),
            .sr(_gnd_net_));
    defparam shift_srl_82_0_LC_23_7_0.C_ON=1'b0;
    defparam shift_srl_82_0_LC_23_7_0.SEQ_MODE=4'b1000;
    defparam shift_srl_82_0_LC_23_7_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_82_0_LC_23_7_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80821),
            .lcout(shift_srl_82Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93387),
            .ce(N__80841),
            .sr(_gnd_net_));
    defparam shift_srl_82_1_LC_23_7_1.C_ON=1'b0;
    defparam shift_srl_82_1_LC_23_7_1.SEQ_MODE=4'b1000;
    defparam shift_srl_82_1_LC_23_7_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_82_1_LC_23_7_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78649),
            .lcout(shift_srl_82Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93387),
            .ce(N__80841),
            .sr(_gnd_net_));
    defparam shift_srl_82_2_LC_23_7_2.C_ON=1'b0;
    defparam shift_srl_82_2_LC_23_7_2.SEQ_MODE=4'b1000;
    defparam shift_srl_82_2_LC_23_7_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_82_2_LC_23_7_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78643),
            .lcout(shift_srl_82Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93387),
            .ce(N__80841),
            .sr(_gnd_net_));
    defparam shift_srl_82_3_LC_23_7_3.C_ON=1'b0;
    defparam shift_srl_82_3_LC_23_7_3.SEQ_MODE=4'b1000;
    defparam shift_srl_82_3_LC_23_7_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_82_3_LC_23_7_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78637),
            .lcout(shift_srl_82Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93387),
            .ce(N__80841),
            .sr(_gnd_net_));
    defparam shift_srl_82_4_LC_23_7_4.C_ON=1'b0;
    defparam shift_srl_82_4_LC_23_7_4.SEQ_MODE=4'b1000;
    defparam shift_srl_82_4_LC_23_7_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_82_4_LC_23_7_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78631),
            .lcout(shift_srl_82Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93387),
            .ce(N__80841),
            .sr(_gnd_net_));
    defparam shift_srl_82_5_LC_23_7_5.C_ON=1'b0;
    defparam shift_srl_82_5_LC_23_7_5.SEQ_MODE=4'b1000;
    defparam shift_srl_82_5_LC_23_7_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_82_5_LC_23_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78625),
            .lcout(shift_srl_82Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93387),
            .ce(N__80841),
            .sr(_gnd_net_));
    defparam shift_srl_82_6_LC_23_7_6.C_ON=1'b0;
    defparam shift_srl_82_6_LC_23_7_6.SEQ_MODE=4'b1000;
    defparam shift_srl_82_6_LC_23_7_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_82_6_LC_23_7_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78619),
            .lcout(shift_srl_82Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93387),
            .ce(N__80841),
            .sr(_gnd_net_));
    defparam shift_srl_82_7_LC_23_7_7.C_ON=1'b0;
    defparam shift_srl_82_7_LC_23_7_7.SEQ_MODE=4'b1000;
    defparam shift_srl_82_7_LC_23_7_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_82_7_LC_23_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78613),
            .lcout(shift_srl_82Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93387),
            .ce(N__80841),
            .sr(_gnd_net_));
    defparam shift_srl_41_0_LC_23_9_0.C_ON=1'b0;
    defparam shift_srl_41_0_LC_23_9_0.SEQ_MODE=4'b1000;
    defparam shift_srl_41_0_LC_23_9_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_41_0_LC_23_9_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78799),
            .lcout(shift_srl_41Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93354),
            .ce(N__78691),
            .sr(_gnd_net_));
    defparam shift_srl_41_1_LC_23_9_1.C_ON=1'b0;
    defparam shift_srl_41_1_LC_23_9_1.SEQ_MODE=4'b1000;
    defparam shift_srl_41_1_LC_23_9_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_41_1_LC_23_9_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78745),
            .lcout(shift_srl_41Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93354),
            .ce(N__78691),
            .sr(_gnd_net_));
    defparam shift_srl_41_2_LC_23_9_2.C_ON=1'b0;
    defparam shift_srl_41_2_LC_23_9_2.SEQ_MODE=4'b1000;
    defparam shift_srl_41_2_LC_23_9_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_41_2_LC_23_9_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78739),
            .lcout(shift_srl_41Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93354),
            .ce(N__78691),
            .sr(_gnd_net_));
    defparam shift_srl_41_3_LC_23_9_3.C_ON=1'b0;
    defparam shift_srl_41_3_LC_23_9_3.SEQ_MODE=4'b1000;
    defparam shift_srl_41_3_LC_23_9_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_41_3_LC_23_9_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78733),
            .lcout(shift_srl_41Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93354),
            .ce(N__78691),
            .sr(_gnd_net_));
    defparam shift_srl_41_4_LC_23_9_4.C_ON=1'b0;
    defparam shift_srl_41_4_LC_23_9_4.SEQ_MODE=4'b1000;
    defparam shift_srl_41_4_LC_23_9_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_41_4_LC_23_9_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78727),
            .lcout(shift_srl_41Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93354),
            .ce(N__78691),
            .sr(_gnd_net_));
    defparam shift_srl_41_5_LC_23_9_5.C_ON=1'b0;
    defparam shift_srl_41_5_LC_23_9_5.SEQ_MODE=4'b1000;
    defparam shift_srl_41_5_LC_23_9_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_41_5_LC_23_9_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78721),
            .lcout(shift_srl_41Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93354),
            .ce(N__78691),
            .sr(_gnd_net_));
    defparam shift_srl_41_6_LC_23_9_6.C_ON=1'b0;
    defparam shift_srl_41_6_LC_23_9_6.SEQ_MODE=4'b1000;
    defparam shift_srl_41_6_LC_23_9_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_41_6_LC_23_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78715),
            .lcout(shift_srl_41Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93354),
            .ce(N__78691),
            .sr(_gnd_net_));
    defparam shift_srl_41_7_LC_23_9_7.C_ON=1'b0;
    defparam shift_srl_41_7_LC_23_9_7.SEQ_MODE=4'b1000;
    defparam shift_srl_41_7_LC_23_9_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_41_7_LC_23_9_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78709),
            .lcout(shift_srl_41Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93354),
            .ce(N__78691),
            .sr(_gnd_net_));
    defparam shift_srl_56_1_LC_23_10_0.C_ON=1'b0;
    defparam shift_srl_56_1_LC_23_10_0.SEQ_MODE=4'b1000;
    defparam shift_srl_56_1_LC_23_10_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_56_1_LC_23_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78670),
            .lcout(shift_srl_56Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93332),
            .ce(N__78829),
            .sr(_gnd_net_));
    defparam shift_srl_56_7_LC_23_10_1.C_ON=1'b0;
    defparam shift_srl_56_7_LC_23_10_1.SEQ_MODE=4'b1000;
    defparam shift_srl_56_7_LC_23_10_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_56_7_LC_23_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78874),
            .lcout(shift_srl_56Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93332),
            .ce(N__78829),
            .sr(_gnd_net_));
    defparam shift_srl_56_2_LC_23_10_2.C_ON=1'b0;
    defparam shift_srl_56_2_LC_23_10_2.SEQ_MODE=4'b1000;
    defparam shift_srl_56_2_LC_23_10_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_56_2_LC_23_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78880),
            .lcout(shift_srl_56Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93332),
            .ce(N__78829),
            .sr(_gnd_net_));
    defparam shift_srl_56_6_LC_23_10_3.C_ON=1'b0;
    defparam shift_srl_56_6_LC_23_10_3.SEQ_MODE=4'b1000;
    defparam shift_srl_56_6_LC_23_10_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_56_6_LC_23_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78862),
            .lcout(shift_srl_56Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93332),
            .ce(N__78829),
            .sr(_gnd_net_));
    defparam shift_srl_56_3_LC_23_10_4.C_ON=1'b0;
    defparam shift_srl_56_3_LC_23_10_4.SEQ_MODE=4'b1000;
    defparam shift_srl_56_3_LC_23_10_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_56_3_LC_23_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78868),
            .lcout(shift_srl_56Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93332),
            .ce(N__78829),
            .sr(_gnd_net_));
    defparam shift_srl_56_5_LC_23_10_5.C_ON=1'b0;
    defparam shift_srl_56_5_LC_23_10_5.SEQ_MODE=4'b1000;
    defparam shift_srl_56_5_LC_23_10_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_56_5_LC_23_10_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78850),
            .lcout(shift_srl_56Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93332),
            .ce(N__78829),
            .sr(_gnd_net_));
    defparam shift_srl_56_4_LC_23_10_6.C_ON=1'b0;
    defparam shift_srl_56_4_LC_23_10_6.SEQ_MODE=4'b1000;
    defparam shift_srl_56_4_LC_23_10_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_56_4_LC_23_10_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78856),
            .lcout(shift_srl_56Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93332),
            .ce(N__78829),
            .sr(_gnd_net_));
    defparam shift_srl_56_8_LC_23_10_7.C_ON=1'b0;
    defparam shift_srl_56_8_LC_23_10_7.SEQ_MODE=4'b1000;
    defparam shift_srl_56_8_LC_23_10_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_56_8_LC_23_10_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78844),
            .lcout(shift_srl_56Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93332),
            .ce(N__78829),
            .sr(_gnd_net_));
    defparam shift_srl_58_0_LC_23_11_0.C_ON=1'b0;
    defparam shift_srl_58_0_LC_23_11_0.SEQ_MODE=4'b1000;
    defparam shift_srl_58_0_LC_23_11_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_58_0_LC_23_11_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79002),
            .lcout(shift_srl_58Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93311),
            .ce(N__78969),
            .sr(_gnd_net_));
    defparam shift_srl_58_1_LC_23_11_1.C_ON=1'b0;
    defparam shift_srl_58_1_LC_23_11_1.SEQ_MODE=4'b1000;
    defparam shift_srl_58_1_LC_23_11_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_58_1_LC_23_11_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78805),
            .lcout(shift_srl_58Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93311),
            .ce(N__78969),
            .sr(_gnd_net_));
    defparam shift_srl_58_2_LC_23_11_2.C_ON=1'b0;
    defparam shift_srl_58_2_LC_23_11_2.SEQ_MODE=4'b1000;
    defparam shift_srl_58_2_LC_23_11_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_58_2_LC_23_11_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78934),
            .lcout(shift_srl_58Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93311),
            .ce(N__78969),
            .sr(_gnd_net_));
    defparam shift_srl_58_3_LC_23_11_3.C_ON=1'b0;
    defparam shift_srl_58_3_LC_23_11_3.SEQ_MODE=4'b1000;
    defparam shift_srl_58_3_LC_23_11_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_58_3_LC_23_11_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78928),
            .lcout(shift_srl_58Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93311),
            .ce(N__78969),
            .sr(_gnd_net_));
    defparam shift_srl_58_4_LC_23_11_4.C_ON=1'b0;
    defparam shift_srl_58_4_LC_23_11_4.SEQ_MODE=4'b1000;
    defparam shift_srl_58_4_LC_23_11_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_58_4_LC_23_11_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78922),
            .lcout(shift_srl_58Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93311),
            .ce(N__78969),
            .sr(_gnd_net_));
    defparam shift_srl_58_5_LC_23_11_5.C_ON=1'b0;
    defparam shift_srl_58_5_LC_23_11_5.SEQ_MODE=4'b1000;
    defparam shift_srl_58_5_LC_23_11_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_58_5_LC_23_11_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78916),
            .lcout(shift_srl_58Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93311),
            .ce(N__78969),
            .sr(_gnd_net_));
    defparam shift_srl_58_6_LC_23_11_6.C_ON=1'b0;
    defparam shift_srl_58_6_LC_23_11_6.SEQ_MODE=4'b1000;
    defparam shift_srl_58_6_LC_23_11_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_58_6_LC_23_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78910),
            .lcout(shift_srl_58Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93311),
            .ce(N__78969),
            .sr(_gnd_net_));
    defparam shift_srl_58_7_LC_23_11_7.C_ON=1'b0;
    defparam shift_srl_58_7_LC_23_11_7.SEQ_MODE=4'b1000;
    defparam shift_srl_58_7_LC_23_11_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_58_7_LC_23_11_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78904),
            .lcout(shift_srl_58Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93311),
            .ce(N__78969),
            .sr(_gnd_net_));
    defparam shift_srl_58_10_LC_23_12_0.C_ON=1'b0;
    defparam shift_srl_58_10_LC_23_12_0.SEQ_MODE=4'b1000;
    defparam shift_srl_58_10_LC_23_12_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_58_10_LC_23_12_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78988),
            .lcout(shift_srl_58Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93292),
            .ce(N__78970),
            .sr(_gnd_net_));
    defparam shift_srl_58_11_LC_23_12_1.C_ON=1'b0;
    defparam shift_srl_58_11_LC_23_12_1.SEQ_MODE=4'b1000;
    defparam shift_srl_58_11_LC_23_12_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_58_11_LC_23_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78898),
            .lcout(shift_srl_58Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93292),
            .ce(N__78970),
            .sr(_gnd_net_));
    defparam shift_srl_58_12_LC_23_12_2.C_ON=1'b0;
    defparam shift_srl_58_12_LC_23_12_2.SEQ_MODE=4'b1000;
    defparam shift_srl_58_12_LC_23_12_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_58_12_LC_23_12_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78892),
            .lcout(shift_srl_58Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93292),
            .ce(N__78970),
            .sr(_gnd_net_));
    defparam shift_srl_58_13_LC_23_12_3.C_ON=1'b0;
    defparam shift_srl_58_13_LC_23_12_3.SEQ_MODE=4'b1000;
    defparam shift_srl_58_13_LC_23_12_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_58_13_LC_23_12_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78886),
            .lcout(shift_srl_58Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93292),
            .ce(N__78970),
            .sr(_gnd_net_));
    defparam shift_srl_58_14_LC_23_12_4.C_ON=1'b0;
    defparam shift_srl_58_14_LC_23_12_4.SEQ_MODE=4'b1000;
    defparam shift_srl_58_14_LC_23_12_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_58_14_LC_23_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79018),
            .lcout(shift_srl_58Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93292),
            .ce(N__78970),
            .sr(_gnd_net_));
    defparam shift_srl_58_15_LC_23_12_5.C_ON=1'b0;
    defparam shift_srl_58_15_LC_23_12_5.SEQ_MODE=4'b1000;
    defparam shift_srl_58_15_LC_23_12_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_58_15_LC_23_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79012),
            .lcout(shift_srl_58Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93292),
            .ce(N__78970),
            .sr(_gnd_net_));
    defparam shift_srl_58_9_LC_23_12_6.C_ON=1'b0;
    defparam shift_srl_58_9_LC_23_12_6.SEQ_MODE=4'b1000;
    defparam shift_srl_58_9_LC_23_12_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_58_9_LC_23_12_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78976),
            .lcout(shift_srl_58Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93292),
            .ce(N__78970),
            .sr(_gnd_net_));
    defparam shift_srl_58_8_LC_23_12_7.C_ON=1'b0;
    defparam shift_srl_58_8_LC_23_12_7.SEQ_MODE=4'b1000;
    defparam shift_srl_58_8_LC_23_12_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_58_8_LC_23_12_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78982),
            .lcout(shift_srl_58Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93292),
            .ce(N__78970),
            .sr(_gnd_net_));
    defparam shift_srl_64_0_LC_23_13_0.C_ON=1'b0;
    defparam shift_srl_64_0_LC_23_13_0.SEQ_MODE=4'b1000;
    defparam shift_srl_64_0_LC_23_13_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_64_0_LC_23_13_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81083),
            .lcout(shift_srl_64Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93278),
            .ce(N__79101),
            .sr(_gnd_net_));
    defparam shift_srl_64_1_LC_23_13_1.C_ON=1'b0;
    defparam shift_srl_64_1_LC_23_13_1.SEQ_MODE=4'b1000;
    defparam shift_srl_64_1_LC_23_13_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_64_1_LC_23_13_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78958),
            .lcout(shift_srl_64Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93278),
            .ce(N__79101),
            .sr(_gnd_net_));
    defparam shift_srl_64_2_LC_23_13_2.C_ON=1'b0;
    defparam shift_srl_64_2_LC_23_13_2.SEQ_MODE=4'b1000;
    defparam shift_srl_64_2_LC_23_13_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_64_2_LC_23_13_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78952),
            .lcout(shift_srl_64Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93278),
            .ce(N__79101),
            .sr(_gnd_net_));
    defparam shift_srl_64_3_LC_23_13_3.C_ON=1'b0;
    defparam shift_srl_64_3_LC_23_13_3.SEQ_MODE=4'b1000;
    defparam shift_srl_64_3_LC_23_13_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_64_3_LC_23_13_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78946),
            .lcout(shift_srl_64Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93278),
            .ce(N__79101),
            .sr(_gnd_net_));
    defparam shift_srl_64_4_LC_23_13_4.C_ON=1'b0;
    defparam shift_srl_64_4_LC_23_13_4.SEQ_MODE=4'b1000;
    defparam shift_srl_64_4_LC_23_13_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_64_4_LC_23_13_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78940),
            .lcout(shift_srl_64Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93278),
            .ce(N__79101),
            .sr(_gnd_net_));
    defparam shift_srl_64_5_LC_23_13_5.C_ON=1'b0;
    defparam shift_srl_64_5_LC_23_13_5.SEQ_MODE=4'b1000;
    defparam shift_srl_64_5_LC_23_13_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_64_5_LC_23_13_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79126),
            .lcout(shift_srl_64Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93278),
            .ce(N__79101),
            .sr(_gnd_net_));
    defparam shift_srl_64_6_LC_23_13_6.C_ON=1'b0;
    defparam shift_srl_64_6_LC_23_13_6.SEQ_MODE=4'b1000;
    defparam shift_srl_64_6_LC_23_13_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_64_6_LC_23_13_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79120),
            .lcout(shift_srl_64Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93278),
            .ce(N__79101),
            .sr(_gnd_net_));
    defparam shift_srl_64_7_LC_23_13_7.C_ON=1'b0;
    defparam shift_srl_64_7_LC_23_13_7.SEQ_MODE=4'b1000;
    defparam shift_srl_64_7_LC_23_13_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_64_7_LC_23_13_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79114),
            .lcout(shift_srl_64Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93278),
            .ce(N__79101),
            .sr(_gnd_net_));
    defparam shift_srl_63_RNIGBGJG_15_LC_23_14_0.C_ON=1'b0;
    defparam shift_srl_63_RNIGBGJG_15_LC_23_14_0.SEQ_MODE=4'b0000;
    defparam shift_srl_63_RNIGBGJG_15_LC_23_14_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_63_RNIGBGJG_15_LC_23_14_0 (
            .in0(N__84903),
            .in1(N__90278),
            .in2(N__81056),
            .in3(N__81124),
            .lcout(clk_en_64),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_63_15_LC_23_14_1.C_ON=1'b0;
    defparam shift_srl_63_15_LC_23_14_1.SEQ_MODE=4'b1000;
    defparam shift_srl_63_15_LC_23_14_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_63_15_LC_23_14_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79036),
            .lcout(shift_srl_63Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93259),
            .ce(N__79192),
            .sr(_gnd_net_));
    defparam shift_srl_64_RNI541NG_15_LC_23_14_2.C_ON=1'b0;
    defparam shift_srl_64_RNI541NG_15_LC_23_14_2.SEQ_MODE=4'b0000;
    defparam shift_srl_64_RNI541NG_15_LC_23_14_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_64_RNI541NG_15_LC_23_14_2 (
            .in0(N__81082),
            .in1(N__81125),
            .in2(N__81057),
            .in3(N__79079),
            .lcout(clk_en_65),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_63_14_LC_23_14_3.C_ON=1'b0;
    defparam shift_srl_63_14_LC_23_14_3.SEQ_MODE=4'b1000;
    defparam shift_srl_63_14_LC_23_14_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_63_14_LC_23_14_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79030),
            .lcout(shift_srl_63Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93259),
            .ce(N__79192),
            .sr(_gnd_net_));
    defparam shift_srl_63_13_LC_23_14_4.C_ON=1'b0;
    defparam shift_srl_63_13_LC_23_14_4.SEQ_MODE=4'b1000;
    defparam shift_srl_63_13_LC_23_14_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_63_13_LC_23_14_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79024),
            .lcout(shift_srl_63Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93259),
            .ce(N__79192),
            .sr(_gnd_net_));
    defparam shift_srl_63_12_LC_23_14_5.C_ON=1'b0;
    defparam shift_srl_63_12_LC_23_14_5.SEQ_MODE=4'b1000;
    defparam shift_srl_63_12_LC_23_14_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_63_12_LC_23_14_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79213),
            .lcout(shift_srl_63Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93259),
            .ce(N__79192),
            .sr(_gnd_net_));
    defparam shift_srl_63_11_LC_23_14_6.C_ON=1'b0;
    defparam shift_srl_63_11_LC_23_14_6.SEQ_MODE=4'b1000;
    defparam shift_srl_63_11_LC_23_14_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_63_11_LC_23_14_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79198),
            .lcout(shift_srl_63Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93259),
            .ce(N__79192),
            .sr(_gnd_net_));
    defparam shift_srl_63_10_LC_23_14_7.C_ON=1'b0;
    defparam shift_srl_63_10_LC_23_14_7.SEQ_MODE=4'b1000;
    defparam shift_srl_63_10_LC_23_14_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_63_10_LC_23_14_7 (
            .in0(N__79207),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_63Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93259),
            .ce(N__79192),
            .sr(_gnd_net_));
    defparam shift_srl_65_0_LC_23_15_0.C_ON=1'b0;
    defparam shift_srl_65_0_LC_23_15_0.SEQ_MODE=4'b1000;
    defparam shift_srl_65_0_LC_23_15_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_65_0_LC_23_15_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80994),
            .lcout(shift_srl_65Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93237),
            .ce(N__79785),
            .sr(_gnd_net_));
    defparam shift_srl_65_1_LC_23_15_1.C_ON=1'b0;
    defparam shift_srl_65_1_LC_23_15_1.SEQ_MODE=4'b1000;
    defparam shift_srl_65_1_LC_23_15_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_65_1_LC_23_15_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79162),
            .lcout(shift_srl_65Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93237),
            .ce(N__79785),
            .sr(_gnd_net_));
    defparam shift_srl_65_2_LC_23_15_2.C_ON=1'b0;
    defparam shift_srl_65_2_LC_23_15_2.SEQ_MODE=4'b1000;
    defparam shift_srl_65_2_LC_23_15_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_65_2_LC_23_15_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79156),
            .lcout(shift_srl_65Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93237),
            .ce(N__79785),
            .sr(_gnd_net_));
    defparam shift_srl_65_3_LC_23_15_3.C_ON=1'b0;
    defparam shift_srl_65_3_LC_23_15_3.SEQ_MODE=4'b1000;
    defparam shift_srl_65_3_LC_23_15_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_65_3_LC_23_15_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79150),
            .lcout(shift_srl_65Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93237),
            .ce(N__79785),
            .sr(_gnd_net_));
    defparam shift_srl_65_4_LC_23_15_4.C_ON=1'b0;
    defparam shift_srl_65_4_LC_23_15_4.SEQ_MODE=4'b1000;
    defparam shift_srl_65_4_LC_23_15_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_65_4_LC_23_15_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79144),
            .lcout(shift_srl_65Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93237),
            .ce(N__79785),
            .sr(_gnd_net_));
    defparam shift_srl_65_5_LC_23_15_5.C_ON=1'b0;
    defparam shift_srl_65_5_LC_23_15_5.SEQ_MODE=4'b1000;
    defparam shift_srl_65_5_LC_23_15_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_65_5_LC_23_15_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79138),
            .lcout(shift_srl_65Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93237),
            .ce(N__79785),
            .sr(_gnd_net_));
    defparam shift_srl_65_6_LC_23_15_6.C_ON=1'b0;
    defparam shift_srl_65_6_LC_23_15_6.SEQ_MODE=4'b1000;
    defparam shift_srl_65_6_LC_23_15_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_65_6_LC_23_15_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79132),
            .lcout(shift_srl_65Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93237),
            .ce(N__79785),
            .sr(_gnd_net_));
    defparam shift_srl_65_7_LC_23_15_7.C_ON=1'b0;
    defparam shift_srl_65_7_LC_23_15_7.SEQ_MODE=4'b1000;
    defparam shift_srl_65_7_LC_23_15_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_65_7_LC_23_15_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79798),
            .lcout(shift_srl_65Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93237),
            .ce(N__79785),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNITUO18_15_LC_23_16_0.C_ON=1'b0;
    defparam shift_srl_0_RNITUO18_15_LC_23_16_0.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNITUO18_15_LC_23_16_0.LUT_INIT=16'b1010101000000000;
    LogicCell40 shift_srl_0_RNITUO18_15_LC_23_16_0 (
            .in0(N__90265),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79916),
            .lcout(clk_en_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_30_7_LC_23_16_1.C_ON=1'b0;
    defparam shift_srl_30_7_LC_23_16_1.SEQ_MODE=4'b1000;
    defparam shift_srl_30_7_LC_23_16_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_30_7_LC_23_16_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79774),
            .lcout(shift_srl_30Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93219),
            .ce(N__79823),
            .sr(_gnd_net_));
    defparam shift_srl_38_RNI493Q9_15_LC_23_16_2.C_ON=1'b0;
    defparam shift_srl_38_RNI493Q9_15_LC_23_16_2.SEQ_MODE=4'b0000;
    defparam shift_srl_38_RNI493Q9_15_LC_23_16_2.LUT_INIT=16'b1100110000000000;
    LogicCell40 shift_srl_38_RNI493Q9_15_LC_23_16_2 (
            .in0(_gnd_net_),
            .in1(N__79762),
            .in2(_gnd_net_),
            .in3(N__81333),
            .lcout(rco_c_38),
            .ltout(rco_c_38_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIVKTQ9_15_LC_23_16_3.C_ON=1'b0;
    defparam shift_srl_0_RNIVKTQ9_15_LC_23_16_3.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIVKTQ9_15_LC_23_16_3.LUT_INIT=16'b1111000000000000;
    LogicCell40 shift_srl_0_RNIVKTQ9_15_LC_23_16_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__79702),
            .in3(N__90264),
            .lcout(clk_en_39),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_30_8_LC_23_16_4.C_ON=1'b0;
    defparam shift_srl_30_8_LC_23_16_4.SEQ_MODE=4'b1000;
    defparam shift_srl_30_8_LC_23_16_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_30_8_LC_23_16_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79699),
            .lcout(shift_srl_30Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93219),
            .ce(N__79823),
            .sr(_gnd_net_));
    defparam shift_srl_100_RNICPACP_15_LC_23_16_5.C_ON=1'b0;
    defparam shift_srl_100_RNICPACP_15_LC_23_16_5.SEQ_MODE=4'b0000;
    defparam shift_srl_100_RNICPACP_15_LC_23_16_5.LUT_INIT=16'b1010101000000000;
    LogicCell40 shift_srl_100_RNICPACP_15_LC_23_16_5 (
            .in0(N__79525),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79693),
            .lcout(rco_c_100),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_102_RNI6TFFQ_15_LC_23_16_6.C_ON=1'b0;
    defparam shift_srl_102_RNI6TFFQ_15_LC_23_16_6.SEQ_MODE=4'b0000;
    defparam shift_srl_102_RNI6TFFQ_15_LC_23_16_6.LUT_INIT=16'b1010101000000000;
    LogicCell40 shift_srl_102_RNI6TFFQ_15_LC_23_16_6 (
            .in0(N__79606),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79526),
            .lcout(rco_c_104),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_164_RNIBMOL_15_LC_23_16_7.C_ON=1'b0;
    defparam shift_srl_164_RNIBMOL_15_LC_23_16_7.SEQ_MODE=4'b0000;
    defparam shift_srl_164_RNIBMOL_15_LC_23_16_7.LUT_INIT=16'b1100110000000000;
    LogicCell40 shift_srl_164_RNIBMOL_15_LC_23_16_7 (
            .in0(_gnd_net_),
            .in1(N__87763),
            .in2(_gnd_net_),
            .in3(N__87255),
            .lcout(shift_srl_164_RNIBMOLZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_30_RNIBOI58_15_LC_23_17_0.C_ON=1'b0;
    defparam shift_srl_30_RNIBOI58_15_LC_23_17_0.SEQ_MODE=4'b0000;
    defparam shift_srl_30_RNIBOI58_15_LC_23_17_0.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_30_RNIBOI58_15_LC_23_17_0 (
            .in0(N__90263),
            .in1(N__79929),
            .in2(_gnd_net_),
            .in3(N__83699),
            .lcout(clk_en_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_30_15_LC_23_17_1.C_ON=1'b0;
    defparam shift_srl_30_15_LC_23_17_1.SEQ_MODE=4'b1000;
    defparam shift_srl_30_15_LC_23_17_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_30_15_LC_23_17_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79876),
            .lcout(shift_srl_30Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93176),
            .ce(N__79830),
            .sr(_gnd_net_));
    defparam shift_srl_30_14_LC_23_17_2.C_ON=1'b0;
    defparam shift_srl_30_14_LC_23_17_2.SEQ_MODE=4'b1000;
    defparam shift_srl_30_14_LC_23_17_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_30_14_LC_23_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79870),
            .lcout(shift_srl_30Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93176),
            .ce(N__79830),
            .sr(_gnd_net_));
    defparam shift_srl_30_13_LC_23_17_3.C_ON=1'b0;
    defparam shift_srl_30_13_LC_23_17_3.SEQ_MODE=4'b1000;
    defparam shift_srl_30_13_LC_23_17_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_30_13_LC_23_17_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79864),
            .lcout(shift_srl_30Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93176),
            .ce(N__79830),
            .sr(_gnd_net_));
    defparam shift_srl_30_12_LC_23_17_4.C_ON=1'b0;
    defparam shift_srl_30_12_LC_23_17_4.SEQ_MODE=4'b1000;
    defparam shift_srl_30_12_LC_23_17_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_30_12_LC_23_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79858),
            .lcout(shift_srl_30Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93176),
            .ce(N__79830),
            .sr(_gnd_net_));
    defparam shift_srl_30_11_LC_23_17_5.C_ON=1'b0;
    defparam shift_srl_30_11_LC_23_17_5.SEQ_MODE=4'b1000;
    defparam shift_srl_30_11_LC_23_17_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_30_11_LC_23_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79852),
            .lcout(shift_srl_30Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93176),
            .ce(N__79830),
            .sr(_gnd_net_));
    defparam shift_srl_30_10_LC_23_17_6.C_ON=1'b0;
    defparam shift_srl_30_10_LC_23_17_6.SEQ_MODE=4'b1000;
    defparam shift_srl_30_10_LC_23_17_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_30_10_LC_23_17_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79840),
            .lcout(shift_srl_30Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93176),
            .ce(N__79830),
            .sr(_gnd_net_));
    defparam shift_srl_30_9_LC_23_17_7.C_ON=1'b0;
    defparam shift_srl_30_9_LC_23_17_7.SEQ_MODE=4'b1000;
    defparam shift_srl_30_9_LC_23_17_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_30_9_LC_23_17_7 (
            .in0(N__79846),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_30Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93176),
            .ce(N__79830),
            .sr(_gnd_net_));
    defparam shift_srl_165_10_LC_23_18_0.C_ON=1'b0;
    defparam shift_srl_165_10_LC_23_18_0.SEQ_MODE=4'b1000;
    defparam shift_srl_165_10_LC_23_18_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_165_10_LC_23_18_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79954),
            .lcout(shift_srl_165Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93220),
            .ce(N__80017),
            .sr(_gnd_net_));
    defparam shift_srl_165_11_LC_23_18_1.C_ON=1'b0;
    defparam shift_srl_165_11_LC_23_18_1.SEQ_MODE=4'b1000;
    defparam shift_srl_165_11_LC_23_18_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_165_11_LC_23_18_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79984),
            .lcout(shift_srl_165Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93220),
            .ce(N__80017),
            .sr(_gnd_net_));
    defparam shift_srl_165_12_LC_23_18_2.C_ON=1'b0;
    defparam shift_srl_165_12_LC_23_18_2.SEQ_MODE=4'b1000;
    defparam shift_srl_165_12_LC_23_18_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_165_12_LC_23_18_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79978),
            .lcout(shift_srl_165Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93220),
            .ce(N__80017),
            .sr(_gnd_net_));
    defparam shift_srl_165_13_LC_23_18_3.C_ON=1'b0;
    defparam shift_srl_165_13_LC_23_18_3.SEQ_MODE=4'b1000;
    defparam shift_srl_165_13_LC_23_18_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_165_13_LC_23_18_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79972),
            .lcout(shift_srl_165Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93220),
            .ce(N__80017),
            .sr(_gnd_net_));
    defparam shift_srl_165_14_LC_23_18_4.C_ON=1'b0;
    defparam shift_srl_165_14_LC_23_18_4.SEQ_MODE=4'b1000;
    defparam shift_srl_165_14_LC_23_18_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_165_14_LC_23_18_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79966),
            .lcout(shift_srl_165Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93220),
            .ce(N__80017),
            .sr(_gnd_net_));
    defparam shift_srl_165_15_LC_23_18_5.C_ON=1'b0;
    defparam shift_srl_165_15_LC_23_18_5.SEQ_MODE=4'b1000;
    defparam shift_srl_165_15_LC_23_18_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_165_15_LC_23_18_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79960),
            .lcout(shift_srl_165Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93220),
            .ce(N__80017),
            .sr(_gnd_net_));
    defparam shift_srl_165_9_LC_23_18_6.C_ON=1'b0;
    defparam shift_srl_165_9_LC_23_18_6.SEQ_MODE=4'b1000;
    defparam shift_srl_165_9_LC_23_18_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_165_9_LC_23_18_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79948),
            .lcout(shift_srl_165Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93220),
            .ce(N__80017),
            .sr(_gnd_net_));
    defparam shift_srl_165_8_LC_23_18_7.C_ON=1'b0;
    defparam shift_srl_165_8_LC_23_18_7.SEQ_MODE=4'b1000;
    defparam shift_srl_165_8_LC_23_18_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_165_8_LC_23_18_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80023),
            .lcout(shift_srl_165Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93220),
            .ce(N__80017),
            .sr(_gnd_net_));
    defparam shift_srl_165_0_LC_23_19_0.C_ON=1'b0;
    defparam shift_srl_165_0_LC_23_19_0.SEQ_MODE=4'b1000;
    defparam shift_srl_165_0_LC_23_19_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_165_0_LC_23_19_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83949),
            .lcout(shift_srl_165Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93238),
            .ce(N__80010),
            .sr(_gnd_net_));
    defparam shift_srl_165_1_LC_23_19_1.C_ON=1'b0;
    defparam shift_srl_165_1_LC_23_19_1.SEQ_MODE=4'b1000;
    defparam shift_srl_165_1_LC_23_19_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_165_1_LC_23_19_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79942),
            .lcout(shift_srl_165Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93238),
            .ce(N__80010),
            .sr(_gnd_net_));
    defparam shift_srl_165_2_LC_23_19_2.C_ON=1'b0;
    defparam shift_srl_165_2_LC_23_19_2.SEQ_MODE=4'b1000;
    defparam shift_srl_165_2_LC_23_19_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_165_2_LC_23_19_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80059),
            .lcout(shift_srl_165Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93238),
            .ce(N__80010),
            .sr(_gnd_net_));
    defparam shift_srl_165_3_LC_23_19_3.C_ON=1'b0;
    defparam shift_srl_165_3_LC_23_19_3.SEQ_MODE=4'b1000;
    defparam shift_srl_165_3_LC_23_19_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_165_3_LC_23_19_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80053),
            .lcout(shift_srl_165Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93238),
            .ce(N__80010),
            .sr(_gnd_net_));
    defparam shift_srl_165_4_LC_23_19_4.C_ON=1'b0;
    defparam shift_srl_165_4_LC_23_19_4.SEQ_MODE=4'b1000;
    defparam shift_srl_165_4_LC_23_19_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_165_4_LC_23_19_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80047),
            .lcout(shift_srl_165Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93238),
            .ce(N__80010),
            .sr(_gnd_net_));
    defparam shift_srl_165_5_LC_23_19_5.C_ON=1'b0;
    defparam shift_srl_165_5_LC_23_19_5.SEQ_MODE=4'b1000;
    defparam shift_srl_165_5_LC_23_19_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_165_5_LC_23_19_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80041),
            .lcout(shift_srl_165Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93238),
            .ce(N__80010),
            .sr(_gnd_net_));
    defparam shift_srl_165_6_LC_23_19_6.C_ON=1'b0;
    defparam shift_srl_165_6_LC_23_19_6.SEQ_MODE=4'b1000;
    defparam shift_srl_165_6_LC_23_19_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_165_6_LC_23_19_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80035),
            .lcout(shift_srl_165Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93238),
            .ce(N__80010),
            .sr(_gnd_net_));
    defparam shift_srl_165_7_LC_23_19_7.C_ON=1'b0;
    defparam shift_srl_165_7_LC_23_19_7.SEQ_MODE=4'b1000;
    defparam shift_srl_165_7_LC_23_19_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_165_7_LC_23_19_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80029),
            .lcout(shift_srl_165Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93238),
            .ce(N__80010),
            .sr(_gnd_net_));
    defparam shift_srl_167_10_LC_23_20_0.C_ON=1'b0;
    defparam shift_srl_167_10_LC_23_20_0.SEQ_MODE=4'b1000;
    defparam shift_srl_167_10_LC_23_20_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_167_10_LC_23_20_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80089),
            .lcout(shift_srl_167Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93260),
            .ce(N__82366),
            .sr(_gnd_net_));
    defparam shift_srl_167_11_LC_23_20_1.C_ON=1'b0;
    defparam shift_srl_167_11_LC_23_20_1.SEQ_MODE=4'b1000;
    defparam shift_srl_167_11_LC_23_20_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_167_11_LC_23_20_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79996),
            .lcout(shift_srl_167Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93260),
            .ce(N__82366),
            .sr(_gnd_net_));
    defparam shift_srl_167_12_LC_23_20_2.C_ON=1'b0;
    defparam shift_srl_167_12_LC_23_20_2.SEQ_MODE=4'b1000;
    defparam shift_srl_167_12_LC_23_20_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_167_12_LC_23_20_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79990),
            .lcout(shift_srl_167Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93260),
            .ce(N__82366),
            .sr(_gnd_net_));
    defparam shift_srl_167_13_LC_23_20_3.C_ON=1'b0;
    defparam shift_srl_167_13_LC_23_20_3.SEQ_MODE=4'b1000;
    defparam shift_srl_167_13_LC_23_20_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_167_13_LC_23_20_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80107),
            .lcout(shift_srl_167Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93260),
            .ce(N__82366),
            .sr(_gnd_net_));
    defparam shift_srl_167_14_LC_23_20_4.C_ON=1'b0;
    defparam shift_srl_167_14_LC_23_20_4.SEQ_MODE=4'b1000;
    defparam shift_srl_167_14_LC_23_20_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_167_14_LC_23_20_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80101),
            .lcout(shift_srl_167Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93260),
            .ce(N__82366),
            .sr(_gnd_net_));
    defparam shift_srl_167_15_LC_23_20_5.C_ON=1'b0;
    defparam shift_srl_167_15_LC_23_20_5.SEQ_MODE=4'b1000;
    defparam shift_srl_167_15_LC_23_20_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_167_15_LC_23_20_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80095),
            .lcout(shift_srl_167Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93260),
            .ce(N__82366),
            .sr(_gnd_net_));
    defparam shift_srl_167_9_LC_23_20_6.C_ON=1'b0;
    defparam shift_srl_167_9_LC_23_20_6.SEQ_MODE=4'b1000;
    defparam shift_srl_167_9_LC_23_20_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_167_9_LC_23_20_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80083),
            .lcout(shift_srl_167Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93260),
            .ce(N__82366),
            .sr(_gnd_net_));
    defparam shift_srl_167_8_LC_23_20_7.C_ON=1'b0;
    defparam shift_srl_167_8_LC_23_20_7.SEQ_MODE=4'b1000;
    defparam shift_srl_167_8_LC_23_20_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_167_8_LC_23_20_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80143),
            .lcout(shift_srl_167Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93260),
            .ce(N__82366),
            .sr(_gnd_net_));
    defparam shift_srl_167_0_LC_23_21_0.C_ON=1'b0;
    defparam shift_srl_167_0_LC_23_21_0.SEQ_MODE=4'b1000;
    defparam shift_srl_167_0_LC_23_21_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_167_0_LC_23_21_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83910),
            .lcout(shift_srl_167Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93279),
            .ce(N__82362),
            .sr(_gnd_net_));
    defparam shift_srl_167_1_LC_23_21_1.C_ON=1'b0;
    defparam shift_srl_167_1_LC_23_21_1.SEQ_MODE=4'b1000;
    defparam shift_srl_167_1_LC_23_21_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_167_1_LC_23_21_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80077),
            .lcout(shift_srl_167Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93279),
            .ce(N__82362),
            .sr(_gnd_net_));
    defparam shift_srl_167_2_LC_23_21_2.C_ON=1'b0;
    defparam shift_srl_167_2_LC_23_21_2.SEQ_MODE=4'b1000;
    defparam shift_srl_167_2_LC_23_21_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_167_2_LC_23_21_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80071),
            .lcout(shift_srl_167Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93279),
            .ce(N__82362),
            .sr(_gnd_net_));
    defparam shift_srl_167_3_LC_23_21_3.C_ON=1'b0;
    defparam shift_srl_167_3_LC_23_21_3.SEQ_MODE=4'b1000;
    defparam shift_srl_167_3_LC_23_21_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_167_3_LC_23_21_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80065),
            .lcout(shift_srl_167Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93279),
            .ce(N__82362),
            .sr(_gnd_net_));
    defparam shift_srl_167_4_LC_23_21_4.C_ON=1'b0;
    defparam shift_srl_167_4_LC_23_21_4.SEQ_MODE=4'b1000;
    defparam shift_srl_167_4_LC_23_21_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_167_4_LC_23_21_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80167),
            .lcout(shift_srl_167Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93279),
            .ce(N__82362),
            .sr(_gnd_net_));
    defparam shift_srl_167_5_LC_23_21_5.C_ON=1'b0;
    defparam shift_srl_167_5_LC_23_21_5.SEQ_MODE=4'b1000;
    defparam shift_srl_167_5_LC_23_21_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_167_5_LC_23_21_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80161),
            .lcout(shift_srl_167Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93279),
            .ce(N__82362),
            .sr(_gnd_net_));
    defparam shift_srl_167_6_LC_23_21_6.C_ON=1'b0;
    defparam shift_srl_167_6_LC_23_21_6.SEQ_MODE=4'b1000;
    defparam shift_srl_167_6_LC_23_21_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_167_6_LC_23_21_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80155),
            .lcout(shift_srl_167Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93279),
            .ce(N__82362),
            .sr(_gnd_net_));
    defparam shift_srl_167_7_LC_23_21_7.C_ON=1'b0;
    defparam shift_srl_167_7_LC_23_21_7.SEQ_MODE=4'b1000;
    defparam shift_srl_167_7_LC_23_21_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_167_7_LC_23_21_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80149),
            .lcout(shift_srl_167Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93279),
            .ce(N__82362),
            .sr(_gnd_net_));
    defparam shift_srl_170_0_LC_23_22_0.C_ON=1'b0;
    defparam shift_srl_170_0_LC_23_22_0.SEQ_MODE=4'b1000;
    defparam shift_srl_170_0_LC_23_22_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_170_0_LC_23_22_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84288),
            .lcout(shift_srl_170Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93293),
            .ce(N__82480),
            .sr(_gnd_net_));
    defparam shift_srl_170_1_LC_23_22_1.C_ON=1'b0;
    defparam shift_srl_170_1_LC_23_22_1.SEQ_MODE=4'b1000;
    defparam shift_srl_170_1_LC_23_22_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_170_1_LC_23_22_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80137),
            .lcout(shift_srl_170Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93293),
            .ce(N__82480),
            .sr(_gnd_net_));
    defparam shift_srl_170_2_LC_23_22_2.C_ON=1'b0;
    defparam shift_srl_170_2_LC_23_22_2.SEQ_MODE=4'b1000;
    defparam shift_srl_170_2_LC_23_22_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_170_2_LC_23_22_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80131),
            .lcout(shift_srl_170Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93293),
            .ce(N__82480),
            .sr(_gnd_net_));
    defparam shift_srl_170_3_LC_23_22_3.C_ON=1'b0;
    defparam shift_srl_170_3_LC_23_22_3.SEQ_MODE=4'b1000;
    defparam shift_srl_170_3_LC_23_22_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_170_3_LC_23_22_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80125),
            .lcout(shift_srl_170Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93293),
            .ce(N__82480),
            .sr(_gnd_net_));
    defparam shift_srl_170_4_LC_23_22_4.C_ON=1'b0;
    defparam shift_srl_170_4_LC_23_22_4.SEQ_MODE=4'b1000;
    defparam shift_srl_170_4_LC_23_22_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_170_4_LC_23_22_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80119),
            .lcout(shift_srl_170Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93293),
            .ce(N__82480),
            .sr(_gnd_net_));
    defparam shift_srl_170_5_LC_23_22_5.C_ON=1'b0;
    defparam shift_srl_170_5_LC_23_22_5.SEQ_MODE=4'b1000;
    defparam shift_srl_170_5_LC_23_22_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_170_5_LC_23_22_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80113),
            .lcout(shift_srl_170Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93293),
            .ce(N__82480),
            .sr(_gnd_net_));
    defparam shift_srl_170_6_LC_23_22_6.C_ON=1'b0;
    defparam shift_srl_170_6_LC_23_22_6.SEQ_MODE=4'b1000;
    defparam shift_srl_170_6_LC_23_22_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_170_6_LC_23_22_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80215),
            .lcout(shift_srl_170Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93293),
            .ce(N__82480),
            .sr(_gnd_net_));
    defparam shift_srl_170_7_LC_23_22_7.C_ON=1'b0;
    defparam shift_srl_170_7_LC_23_22_7.SEQ_MODE=4'b1000;
    defparam shift_srl_170_7_LC_23_22_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_170_7_LC_23_22_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80209),
            .lcout(shift_srl_170Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93293),
            .ce(N__82480),
            .sr(_gnd_net_));
    defparam shift_srl_177_0_LC_23_23_0.C_ON=1'b0;
    defparam shift_srl_177_0_LC_23_23_0.SEQ_MODE=4'b1000;
    defparam shift_srl_177_0_LC_23_23_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_177_0_LC_23_23_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80455),
            .lcout(shift_srl_177Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93312),
            .ce(N__82599),
            .sr(_gnd_net_));
    defparam shift_srl_177_1_LC_23_23_1.C_ON=1'b0;
    defparam shift_srl_177_1_LC_23_23_1.SEQ_MODE=4'b1000;
    defparam shift_srl_177_1_LC_23_23_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_177_1_LC_23_23_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80203),
            .lcout(shift_srl_177Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93312),
            .ce(N__82599),
            .sr(_gnd_net_));
    defparam shift_srl_177_2_LC_23_23_2.C_ON=1'b0;
    defparam shift_srl_177_2_LC_23_23_2.SEQ_MODE=4'b1000;
    defparam shift_srl_177_2_LC_23_23_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_177_2_LC_23_23_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80197),
            .lcout(shift_srl_177Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93312),
            .ce(N__82599),
            .sr(_gnd_net_));
    defparam shift_srl_177_3_LC_23_23_3.C_ON=1'b0;
    defparam shift_srl_177_3_LC_23_23_3.SEQ_MODE=4'b1000;
    defparam shift_srl_177_3_LC_23_23_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_177_3_LC_23_23_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80191),
            .lcout(shift_srl_177Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93312),
            .ce(N__82599),
            .sr(_gnd_net_));
    defparam shift_srl_177_4_LC_23_23_4.C_ON=1'b0;
    defparam shift_srl_177_4_LC_23_23_4.SEQ_MODE=4'b1000;
    defparam shift_srl_177_4_LC_23_23_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_177_4_LC_23_23_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80185),
            .lcout(shift_srl_177Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93312),
            .ce(N__82599),
            .sr(_gnd_net_));
    defparam shift_srl_177_5_LC_23_23_5.C_ON=1'b0;
    defparam shift_srl_177_5_LC_23_23_5.SEQ_MODE=4'b1000;
    defparam shift_srl_177_5_LC_23_23_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_177_5_LC_23_23_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80179),
            .lcout(shift_srl_177Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93312),
            .ce(N__82599),
            .sr(_gnd_net_));
    defparam shift_srl_177_6_LC_23_23_6.C_ON=1'b0;
    defparam shift_srl_177_6_LC_23_23_6.SEQ_MODE=4'b1000;
    defparam shift_srl_177_6_LC_23_23_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_177_6_LC_23_23_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80173),
            .lcout(shift_srl_177Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93312),
            .ce(N__82599),
            .sr(_gnd_net_));
    defparam shift_srl_177_13_LC_23_23_7.C_ON=1'b0;
    defparam shift_srl_177_13_LC_23_23_7.SEQ_MODE=4'b1000;
    defparam shift_srl_177_13_LC_23_23_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_177_13_LC_23_23_7 (
            .in0(N__82636),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_177Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93312),
            .ce(N__82599),
            .sr(_gnd_net_));
    defparam shift_srl_180_0_LC_23_24_0.C_ON=1'b0;
    defparam shift_srl_180_0_LC_23_24_0.SEQ_MODE=4'b1000;
    defparam shift_srl_180_0_LC_23_24_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_180_0_LC_23_24_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82730),
            .lcout(shift_srl_180Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93333),
            .ce(N__82689),
            .sr(_gnd_net_));
    defparam shift_srl_180_1_LC_23_24_1.C_ON=1'b0;
    defparam shift_srl_180_1_LC_23_24_1.SEQ_MODE=4'b1000;
    defparam shift_srl_180_1_LC_23_24_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_180_1_LC_23_24_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80251),
            .lcout(shift_srl_180Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93333),
            .ce(N__82689),
            .sr(_gnd_net_));
    defparam shift_srl_180_2_LC_23_24_2.C_ON=1'b0;
    defparam shift_srl_180_2_LC_23_24_2.SEQ_MODE=4'b1000;
    defparam shift_srl_180_2_LC_23_24_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_180_2_LC_23_24_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80245),
            .lcout(shift_srl_180Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93333),
            .ce(N__82689),
            .sr(_gnd_net_));
    defparam shift_srl_180_3_LC_23_24_3.C_ON=1'b0;
    defparam shift_srl_180_3_LC_23_24_3.SEQ_MODE=4'b1000;
    defparam shift_srl_180_3_LC_23_24_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_180_3_LC_23_24_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80239),
            .lcout(shift_srl_180Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93333),
            .ce(N__82689),
            .sr(_gnd_net_));
    defparam shift_srl_180_4_LC_23_24_4.C_ON=1'b0;
    defparam shift_srl_180_4_LC_23_24_4.SEQ_MODE=4'b1000;
    defparam shift_srl_180_4_LC_23_24_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_180_4_LC_23_24_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80233),
            .lcout(shift_srl_180Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93333),
            .ce(N__82689),
            .sr(_gnd_net_));
    defparam shift_srl_180_7_LC_23_24_5.C_ON=1'b0;
    defparam shift_srl_180_7_LC_23_24_5.SEQ_MODE=4'b1000;
    defparam shift_srl_180_7_LC_23_24_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_180_7_LC_23_24_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80221),
            .lcout(shift_srl_180Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93333),
            .ce(N__82689),
            .sr(_gnd_net_));
    defparam shift_srl_180_8_LC_23_24_6.C_ON=1'b0;
    defparam shift_srl_180_8_LC_23_24_6.SEQ_MODE=4'b1000;
    defparam shift_srl_180_8_LC_23_24_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_180_8_LC_23_24_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80227),
            .lcout(shift_srl_180Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93333),
            .ce(N__82689),
            .sr(_gnd_net_));
    defparam shift_srl_180_6_LC_23_24_7.C_ON=1'b0;
    defparam shift_srl_180_6_LC_23_24_7.SEQ_MODE=4'b1000;
    defparam shift_srl_180_6_LC_23_24_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_180_6_LC_23_24_7 (
            .in0(N__82570),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_180Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93333),
            .ce(N__82689),
            .sr(_gnd_net_));
    defparam shift_srl_188_RNI051CF1_15_LC_23_25_0.C_ON=1'b0;
    defparam shift_srl_188_RNI051CF1_15_LC_23_25_0.SEQ_MODE=4'b0000;
    defparam shift_srl_188_RNI051CF1_15_LC_23_25_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_188_RNI051CF1_15_LC_23_25_0 (
            .in0(N__86094),
            .in1(N__80354),
            .in2(N__90546),
            .in3(N__91525),
            .lcout(clk_en_189),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_188_15_LC_23_25_1.C_ON=1'b0;
    defparam shift_srl_188_15_LC_23_25_1.SEQ_MODE=4'b1000;
    defparam shift_srl_188_15_LC_23_25_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_188_15_LC_23_25_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80299),
            .lcout(shift_srl_188Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93353),
            .ce(N__82804),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_188_LC_23_25_2.C_ON=1'b0;
    defparam rco_obuf_RNO_188_LC_23_25_2.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_188_LC_23_25_2.LUT_INIT=16'b1000100000000000;
    LogicCell40 rco_obuf_RNO_188_LC_23_25_2 (
            .in0(N__86095),
            .in1(N__80355),
            .in2(_gnd_net_),
            .in3(N__91526),
            .lcout(rco_c_188),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_188_14_LC_23_25_3.C_ON=1'b0;
    defparam shift_srl_188_14_LC_23_25_3.SEQ_MODE=4'b1000;
    defparam shift_srl_188_14_LC_23_25_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_188_14_LC_23_25_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80293),
            .lcout(shift_srl_188Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93353),
            .ce(N__82804),
            .sr(_gnd_net_));
    defparam shift_srl_188_13_LC_23_25_4.C_ON=1'b0;
    defparam shift_srl_188_13_LC_23_25_4.SEQ_MODE=4'b1000;
    defparam shift_srl_188_13_LC_23_25_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_188_13_LC_23_25_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80287),
            .lcout(shift_srl_188Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93353),
            .ce(N__82804),
            .sr(_gnd_net_));
    defparam shift_srl_188_12_LC_23_25_5.C_ON=1'b0;
    defparam shift_srl_188_12_LC_23_25_5.SEQ_MODE=4'b1000;
    defparam shift_srl_188_12_LC_23_25_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_188_12_LC_23_25_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80281),
            .lcout(shift_srl_188Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93353),
            .ce(N__82804),
            .sr(_gnd_net_));
    defparam shift_srl_188_11_LC_23_25_6.C_ON=1'b0;
    defparam shift_srl_188_11_LC_23_25_6.SEQ_MODE=4'b1000;
    defparam shift_srl_188_11_LC_23_25_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_188_11_LC_23_25_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80275),
            .lcout(shift_srl_188Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93353),
            .ce(N__82804),
            .sr(_gnd_net_));
    defparam shift_srl_188_10_LC_23_25_7.C_ON=1'b0;
    defparam shift_srl_188_10_LC_23_25_7.SEQ_MODE=4'b1000;
    defparam shift_srl_188_10_LC_23_25_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_188_10_LC_23_25_7 (
            .in0(N__82810),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_188Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93353),
            .ce(N__82804),
            .sr(_gnd_net_));
    defparam shift_srl_192_8_LC_23_26_0.C_ON=1'b0;
    defparam shift_srl_192_8_LC_23_26_0.SEQ_MODE=4'b1000;
    defparam shift_srl_192_8_LC_23_26_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_192_8_LC_23_26_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80269),
            .lcout(shift_srl_192Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93370),
            .ce(N__80677),
            .sr(_gnd_net_));
    defparam shift_srl_192_9_LC_23_26_1.C_ON=1'b0;
    defparam shift_srl_192_9_LC_23_26_1.SEQ_MODE=4'b1000;
    defparam shift_srl_192_9_LC_23_26_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_192_9_LC_23_26_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80695),
            .lcout(shift_srl_192Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93370),
            .ce(N__80677),
            .sr(_gnd_net_));
    defparam shift_srl_173_10_LC_23_27_0.C_ON=1'b0;
    defparam shift_srl_173_10_LC_23_27_0.SEQ_MODE=4'b1000;
    defparam shift_srl_173_10_LC_23_27_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_173_10_LC_23_27_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80611),
            .lcout(shift_srl_173Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93386),
            .ce(N__80584),
            .sr(_gnd_net_));
    defparam shift_srl_173_11_LC_23_27_1.C_ON=1'b0;
    defparam shift_srl_173_11_LC_23_27_1.SEQ_MODE=4'b1000;
    defparam shift_srl_173_11_LC_23_27_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_173_11_LC_23_27_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80647),
            .lcout(shift_srl_173Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93386),
            .ce(N__80584),
            .sr(_gnd_net_));
    defparam shift_srl_173_12_LC_23_27_2.C_ON=1'b0;
    defparam shift_srl_173_12_LC_23_27_2.SEQ_MODE=4'b1000;
    defparam shift_srl_173_12_LC_23_27_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_173_12_LC_23_27_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80641),
            .lcout(shift_srl_173Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93386),
            .ce(N__80584),
            .sr(_gnd_net_));
    defparam shift_srl_173_13_LC_23_27_3.C_ON=1'b0;
    defparam shift_srl_173_13_LC_23_27_3.SEQ_MODE=4'b1000;
    defparam shift_srl_173_13_LC_23_27_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_173_13_LC_23_27_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80635),
            .lcout(shift_srl_173Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93386),
            .ce(N__80584),
            .sr(_gnd_net_));
    defparam shift_srl_173_14_LC_23_27_4.C_ON=1'b0;
    defparam shift_srl_173_14_LC_23_27_4.SEQ_MODE=4'b1000;
    defparam shift_srl_173_14_LC_23_27_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_173_14_LC_23_27_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80629),
            .lcout(shift_srl_173Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93386),
            .ce(N__80584),
            .sr(_gnd_net_));
    defparam shift_srl_173_9_LC_23_27_5.C_ON=1'b0;
    defparam shift_srl_173_9_LC_23_27_5.SEQ_MODE=4'b1000;
    defparam shift_srl_173_9_LC_23_27_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_173_9_LC_23_27_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80590),
            .lcout(shift_srl_173Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93386),
            .ce(N__80584),
            .sr(_gnd_net_));
    defparam shift_srl_173_8_LC_23_27_6.C_ON=1'b0;
    defparam shift_srl_173_8_LC_23_27_6.SEQ_MODE=4'b1000;
    defparam shift_srl_173_8_LC_23_27_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_173_8_LC_23_27_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80605),
            .lcout(shift_srl_173Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93386),
            .ce(N__80584),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_178_LC_23_28_3.C_ON=1'b0;
    defparam rco_obuf_RNO_178_LC_23_28_3.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_178_LC_23_28_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 rco_obuf_RNO_178_LC_23_28_3 (
            .in0(N__80538),
            .in1(N__80475),
            .in2(N__80419),
            .in3(N__85971),
            .lcout(rco_c_178),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_83_10_LC_24_5_1.C_ON=1'b0;
    defparam shift_srl_83_10_LC_24_5_1.SEQ_MODE=4'b1000;
    defparam shift_srl_83_10_LC_24_5_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_83_10_LC_24_5_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80737),
            .lcout(shift_srl_83Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93411),
            .ce(N__80868),
            .sr(_gnd_net_));
    defparam shift_srl_83_9_LC_24_5_4.C_ON=1'b0;
    defparam shift_srl_83_9_LC_24_5_4.SEQ_MODE=4'b1000;
    defparam shift_srl_83_9_LC_24_5_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_83_9_LC_24_5_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80743),
            .lcout(shift_srl_83Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93411),
            .ce(N__80868),
            .sr(_gnd_net_));
    defparam shift_srl_82_10_LC_24_6_0.C_ON=1'b0;
    defparam shift_srl_82_10_LC_24_6_0.SEQ_MODE=4'b1000;
    defparam shift_srl_82_10_LC_24_6_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_82_10_LC_24_6_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80701),
            .lcout(shift_srl_82Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93404),
            .ce(N__80845),
            .sr(_gnd_net_));
    defparam shift_srl_82_11_LC_24_6_1.C_ON=1'b0;
    defparam shift_srl_82_11_LC_24_6_1.SEQ_MODE=4'b1000;
    defparam shift_srl_82_11_LC_24_6_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_82_11_LC_24_6_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80731),
            .lcout(shift_srl_82Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93404),
            .ce(N__80845),
            .sr(_gnd_net_));
    defparam shift_srl_82_12_LC_24_6_2.C_ON=1'b0;
    defparam shift_srl_82_12_LC_24_6_2.SEQ_MODE=4'b1000;
    defparam shift_srl_82_12_LC_24_6_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_82_12_LC_24_6_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80725),
            .lcout(shift_srl_82Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93404),
            .ce(N__80845),
            .sr(_gnd_net_));
    defparam shift_srl_82_13_LC_24_6_3.C_ON=1'b0;
    defparam shift_srl_82_13_LC_24_6_3.SEQ_MODE=4'b1000;
    defparam shift_srl_82_13_LC_24_6_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_82_13_LC_24_6_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80719),
            .lcout(shift_srl_82Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93404),
            .ce(N__80845),
            .sr(_gnd_net_));
    defparam shift_srl_82_14_LC_24_6_4.C_ON=1'b0;
    defparam shift_srl_82_14_LC_24_6_4.SEQ_MODE=4'b1000;
    defparam shift_srl_82_14_LC_24_6_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_82_14_LC_24_6_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80713),
            .lcout(shift_srl_82Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93404),
            .ce(N__80845),
            .sr(_gnd_net_));
    defparam shift_srl_82_15_LC_24_6_5.C_ON=1'b0;
    defparam shift_srl_82_15_LC_24_6_5.SEQ_MODE=4'b1000;
    defparam shift_srl_82_15_LC_24_6_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_82_15_LC_24_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80707),
            .lcout(shift_srl_82Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93404),
            .ce(N__80845),
            .sr(_gnd_net_));
    defparam shift_srl_82_9_LC_24_6_6.C_ON=1'b0;
    defparam shift_srl_82_9_LC_24_6_6.SEQ_MODE=4'b1000;
    defparam shift_srl_82_9_LC_24_6_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_82_9_LC_24_6_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80899),
            .lcout(shift_srl_82Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93404),
            .ce(N__80845),
            .sr(_gnd_net_));
    defparam shift_srl_82_8_LC_24_6_7.C_ON=1'b0;
    defparam shift_srl_82_8_LC_24_6_7.SEQ_MODE=4'b1000;
    defparam shift_srl_82_8_LC_24_6_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_82_8_LC_24_6_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80905),
            .lcout(shift_srl_82Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93404),
            .ce(N__80845),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_82_LC_24_7_0.C_ON=1'b0;
    defparam rco_obuf_RNO_82_LC_24_7_0.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_82_LC_24_7_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 rco_obuf_RNO_82_LC_24_7_0 (
            .in0(N__88509),
            .in1(N__88438),
            .in2(N__86353),
            .in3(N__80824),
            .lcout(N_3998_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_80_RNIG3FB1_15_LC_24_7_1.C_ON=1'b0;
    defparam shift_srl_80_RNIG3FB1_15_LC_24_7_1.SEQ_MODE=4'b0000;
    defparam shift_srl_80_RNIG3FB1_15_LC_24_7_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_80_RNIG3FB1_15_LC_24_7_1 (
            .in0(N__86476),
            .in1(N__84508),
            .in2(N__84682),
            .in3(N__88585),
            .lcout(shift_srl_80_RNIG3FB1Z0Z_15),
            .ltout(shift_srl_80_RNIG3FB1Z0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_82_RNIK0L72_15_LC_24_7_2.C_ON=1'b0;
    defparam shift_srl_82_RNIK0L72_15_LC_24_7_2.SEQ_MODE=4'b0000;
    defparam shift_srl_82_RNIK0L72_15_LC_24_7_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_82_RNIK0L72_15_LC_24_7_2 (
            .in0(N__89950),
            .in1(N__80823),
            .in2(N__80878),
            .in3(N__86348),
            .lcout(),
            .ltout(clk_en_0_a3_0_a2_0_83_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_82_RNIQSK9L_15_LC_24_7_3.C_ON=1'b0;
    defparam shift_srl_82_RNIQSK9L_15_LC_24_7_3.SEQ_MODE=4'b0000;
    defparam shift_srl_82_RNIQSK9L_15_LC_24_7_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_82_RNIQSK9L_15_LC_24_7_3 (
            .in0(N__84902),
            .in1(N__86817),
            .in2(N__80875),
            .in3(N__84998),
            .lcout(clk_en_83),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_81_RNI52SPK_15_LC_24_7_5.C_ON=1'b0;
    defparam shift_srl_81_RNI52SPK_15_LC_24_7_5.SEQ_MODE=4'b0000;
    defparam shift_srl_81_RNI52SPK_15_LC_24_7_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_81_RNI52SPK_15_LC_24_7_5 (
            .in0(N__86349),
            .in1(N__89951),
            .in2(N__88447),
            .in3(N__88508),
            .lcout(N_787),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_83_RNIFJPA2_15_LC_24_7_7.C_ON=1'b0;
    defparam shift_srl_83_RNIFJPA2_15_LC_24_7_7.SEQ_MODE=4'b0000;
    defparam shift_srl_83_RNIFJPA2_15_LC_24_7_7.LUT_INIT=16'b0010000000000000;
    LogicCell40 shift_srl_83_RNIFJPA2_15_LC_24_7_7 (
            .in0(N__80822),
            .in1(N__84475),
            .in2(N__80803),
            .in3(N__88584),
            .lcout(rco_int_0_a2_0_a2_0_83),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_77_RNI8HLI_15_LC_24_8_5.C_ON=1'b0;
    defparam shift_srl_77_RNI8HLI_15_LC_24_8_5.SEQ_MODE=4'b0000;
    defparam shift_srl_77_RNI8HLI_15_LC_24_8_5.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_77_RNI8HLI_15_LC_24_8_5 (
            .in0(N__88278),
            .in1(N__84572),
            .in2(_gnd_net_),
            .in3(N__88394),
            .lcout(shift_srl_77_RNI8HLIZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_76_10_LC_24_9_0.C_ON=1'b0;
    defparam shift_srl_76_10_LC_24_9_0.SEQ_MODE=4'b1000;
    defparam shift_srl_76_10_LC_24_9_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_76_10_LC_24_9_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80929),
            .lcout(shift_srl_76Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93372),
            .ce(N__81247),
            .sr(_gnd_net_));
    defparam shift_srl_76_11_LC_24_9_1.C_ON=1'b0;
    defparam shift_srl_76_11_LC_24_9_1.SEQ_MODE=4'b1000;
    defparam shift_srl_76_11_LC_24_9_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_76_11_LC_24_9_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80959),
            .lcout(shift_srl_76Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93372),
            .ce(N__81247),
            .sr(_gnd_net_));
    defparam shift_srl_76_12_LC_24_9_2.C_ON=1'b0;
    defparam shift_srl_76_12_LC_24_9_2.SEQ_MODE=4'b1000;
    defparam shift_srl_76_12_LC_24_9_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_76_12_LC_24_9_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80953),
            .lcout(shift_srl_76Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93372),
            .ce(N__81247),
            .sr(_gnd_net_));
    defparam shift_srl_76_13_LC_24_9_3.C_ON=1'b0;
    defparam shift_srl_76_13_LC_24_9_3.SEQ_MODE=4'b1000;
    defparam shift_srl_76_13_LC_24_9_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_76_13_LC_24_9_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80947),
            .lcout(shift_srl_76Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93372),
            .ce(N__81247),
            .sr(_gnd_net_));
    defparam shift_srl_76_14_LC_24_9_4.C_ON=1'b0;
    defparam shift_srl_76_14_LC_24_9_4.SEQ_MODE=4'b1000;
    defparam shift_srl_76_14_LC_24_9_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_76_14_LC_24_9_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80941),
            .lcout(shift_srl_76Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93372),
            .ce(N__81247),
            .sr(_gnd_net_));
    defparam shift_srl_76_15_LC_24_9_5.C_ON=1'b0;
    defparam shift_srl_76_15_LC_24_9_5.SEQ_MODE=4'b1000;
    defparam shift_srl_76_15_LC_24_9_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_76_15_LC_24_9_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80935),
            .lcout(shift_srl_76Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93372),
            .ce(N__81247),
            .sr(_gnd_net_));
    defparam shift_srl_76_9_LC_24_9_6.C_ON=1'b0;
    defparam shift_srl_76_9_LC_24_9_6.SEQ_MODE=4'b1000;
    defparam shift_srl_76_9_LC_24_9_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_76_9_LC_24_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80923),
            .lcout(shift_srl_76Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93372),
            .ce(N__81247),
            .sr(_gnd_net_));
    defparam shift_srl_76_8_LC_24_9_7.C_ON=1'b0;
    defparam shift_srl_76_8_LC_24_9_7.SEQ_MODE=4'b1000;
    defparam shift_srl_76_8_LC_24_9_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_76_8_LC_24_9_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81181),
            .lcout(shift_srl_76Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93372),
            .ce(N__81247),
            .sr(_gnd_net_));
    defparam shift_srl_76_0_LC_24_10_0.C_ON=1'b0;
    defparam shift_srl_76_0_LC_24_10_0.SEQ_MODE=4'b1000;
    defparam shift_srl_76_0_LC_24_10_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_76_0_LC_24_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84576),
            .lcout(shift_srl_76Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93355),
            .ce(N__81246),
            .sr(_gnd_net_));
    defparam shift_srl_76_1_LC_24_10_1.C_ON=1'b0;
    defparam shift_srl_76_1_LC_24_10_1.SEQ_MODE=4'b1000;
    defparam shift_srl_76_1_LC_24_10_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_76_1_LC_24_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80917),
            .lcout(shift_srl_76Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93355),
            .ce(N__81246),
            .sr(_gnd_net_));
    defparam shift_srl_76_2_LC_24_10_2.C_ON=1'b0;
    defparam shift_srl_76_2_LC_24_10_2.SEQ_MODE=4'b1000;
    defparam shift_srl_76_2_LC_24_10_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_76_2_LC_24_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80911),
            .lcout(shift_srl_76Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93355),
            .ce(N__81246),
            .sr(_gnd_net_));
    defparam shift_srl_76_3_LC_24_10_3.C_ON=1'b0;
    defparam shift_srl_76_3_LC_24_10_3.SEQ_MODE=4'b1000;
    defparam shift_srl_76_3_LC_24_10_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_76_3_LC_24_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81211),
            .lcout(shift_srl_76Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93355),
            .ce(N__81246),
            .sr(_gnd_net_));
    defparam shift_srl_76_4_LC_24_10_4.C_ON=1'b0;
    defparam shift_srl_76_4_LC_24_10_4.SEQ_MODE=4'b1000;
    defparam shift_srl_76_4_LC_24_10_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_76_4_LC_24_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81205),
            .lcout(shift_srl_76Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93355),
            .ce(N__81246),
            .sr(_gnd_net_));
    defparam shift_srl_76_5_LC_24_10_5.C_ON=1'b0;
    defparam shift_srl_76_5_LC_24_10_5.SEQ_MODE=4'b1000;
    defparam shift_srl_76_5_LC_24_10_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_76_5_LC_24_10_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81199),
            .lcout(shift_srl_76Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93355),
            .ce(N__81246),
            .sr(_gnd_net_));
    defparam shift_srl_76_6_LC_24_10_6.C_ON=1'b0;
    defparam shift_srl_76_6_LC_24_10_6.SEQ_MODE=4'b1000;
    defparam shift_srl_76_6_LC_24_10_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_76_6_LC_24_10_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81193),
            .lcout(shift_srl_76Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93355),
            .ce(N__81246),
            .sr(_gnd_net_));
    defparam shift_srl_76_7_LC_24_10_7.C_ON=1'b0;
    defparam shift_srl_76_7_LC_24_10_7.SEQ_MODE=4'b1000;
    defparam shift_srl_76_7_LC_24_10_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_76_7_LC_24_10_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81187),
            .lcout(shift_srl_76Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93355),
            .ce(N__81246),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_64_LC_24_11_0.C_ON=1'b0;
    defparam rco_obuf_RNO_64_LC_24_11_0.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_64_LC_24_11_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 rco_obuf_RNO_64_LC_24_11_0 (
            .in0(N__81055),
            .in1(N__84905),
            .in2(N__81139),
            .in3(N__81094),
            .lcout(rco_c_64),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_63_LC_24_11_1.C_ON=1'b0;
    defparam rco_obuf_RNO_63_LC_24_11_1.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_63_LC_24_11_1.LUT_INIT=16'b1000100000000000;
    LogicCell40 rco_obuf_RNO_63_LC_24_11_1 (
            .in0(N__84904),
            .in1(N__81054),
            .in2(_gnd_net_),
            .in3(N__81133),
            .lcout(rco_c_63),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_65_RNILFDF1_15_LC_24_11_2.C_ON=1'b0;
    defparam shift_srl_65_RNILFDF1_15_LC_24_11_2.SEQ_MODE=4'b0000;
    defparam shift_srl_65_RNILFDF1_15_LC_24_11_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_65_RNILFDF1_15_LC_24_11_2 (
            .in0(N__81132),
            .in1(N__81093),
            .in2(N__81058),
            .in3(N__80998),
            .lcout(shift_srl_65_RNILFDF1Z0Z_15),
            .ltout(shift_srl_65_RNILFDF1Z0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIR0OUG_15_LC_24_11_3.C_ON=1'b0;
    defparam shift_srl_0_RNIR0OUG_15_LC_24_11_3.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIR0OUG_15_LC_24_11_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNIR0OUG_15_LC_24_11_3 (
            .in0(N__81414),
            .in1(N__90460),
            .in2(N__81592),
            .in3(N__93596),
            .lcout(clk_en_66),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_59_RNI5RRK2_15_LC_24_11_4.C_ON=1'b0;
    defparam shift_srl_59_RNI5RRK2_15_LC_24_11_4.SEQ_MODE=4'b0000;
    defparam shift_srl_59_RNI5RRK2_15_LC_24_11_4.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_59_RNI5RRK2_15_LC_24_11_4 (
            .in0(N__81589),
            .in1(N__81551),
            .in2(_gnd_net_),
            .in3(N__81478),
            .lcout(rco_int_0_a2_1_a2_0_0_59),
            .ltout(rco_int_0_a2_1_a2_0_0_59_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_48_RNI962L7_15_LC_24_11_5.C_ON=1'b0;
    defparam shift_srl_48_RNI962L7_15_LC_24_11_5.SEQ_MODE=4'b0000;
    defparam shift_srl_48_RNI962L7_15_LC_24_11_5.LUT_INIT=16'b0001000000000000;
    LogicCell40 shift_srl_48_RNI962L7_15_LC_24_11_5 (
            .in0(N__81382),
            .in1(N__81367),
            .in2(N__81346),
            .in3(N__84997),
            .lcout(),
            .ltout(rco_int_0_a3_0_a2cf1_66_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_48_RNINLQ9H_15_LC_24_11_6.C_ON=1'b0;
    defparam shift_srl_48_RNINLQ9H_15_LC_24_11_6.SEQ_MODE=4'b0000;
    defparam shift_srl_48_RNINLQ9H_15_LC_24_11_6.LUT_INIT=16'b1111000000000000;
    LogicCell40 shift_srl_48_RNINLQ9H_15_LC_24_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__81343),
            .in3(N__81327),
            .lcout(rco_c_66),
            .ltout(rco_c_66_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_75_RNIO9R4J_15_LC_24_11_7.C_ON=1'b0;
    defparam shift_srl_75_RNIO9R4J_15_LC_24_11_7.SEQ_MODE=4'b0000;
    defparam shift_srl_75_RNIO9R4J_15_LC_24_11_7.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_75_RNIO9R4J_15_LC_24_11_7 (
            .in0(N__90459),
            .in1(N__86800),
            .in2(N__81250),
            .in3(N__88403),
            .lcout(clk_en_76),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_66_0_LC_24_12_0.C_ON=1'b0;
    defparam shift_srl_66_0_LC_24_12_0.SEQ_MODE=4'b1000;
    defparam shift_srl_66_0_LC_24_12_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_66_0_LC_24_12_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81717),
            .lcout(shift_srl_66Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93313),
            .ce(N__81681),
            .sr(_gnd_net_));
    defparam shift_srl_66_1_LC_24_12_1.C_ON=1'b0;
    defparam shift_srl_66_1_LC_24_12_1.SEQ_MODE=4'b1000;
    defparam shift_srl_66_1_LC_24_12_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_66_1_LC_24_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81229),
            .lcout(shift_srl_66Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93313),
            .ce(N__81681),
            .sr(_gnd_net_));
    defparam shift_srl_66_2_LC_24_12_2.C_ON=1'b0;
    defparam shift_srl_66_2_LC_24_12_2.SEQ_MODE=4'b1000;
    defparam shift_srl_66_2_LC_24_12_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_66_2_LC_24_12_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81223),
            .lcout(shift_srl_66Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93313),
            .ce(N__81681),
            .sr(_gnd_net_));
    defparam shift_srl_66_3_LC_24_12_3.C_ON=1'b0;
    defparam shift_srl_66_3_LC_24_12_3.SEQ_MODE=4'b1000;
    defparam shift_srl_66_3_LC_24_12_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_66_3_LC_24_12_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81217),
            .lcout(shift_srl_66Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93313),
            .ce(N__81681),
            .sr(_gnd_net_));
    defparam shift_srl_66_4_LC_24_12_4.C_ON=1'b0;
    defparam shift_srl_66_4_LC_24_12_4.SEQ_MODE=4'b1000;
    defparam shift_srl_66_4_LC_24_12_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_66_4_LC_24_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81640),
            .lcout(shift_srl_66Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93313),
            .ce(N__81681),
            .sr(_gnd_net_));
    defparam shift_srl_66_5_LC_24_12_5.C_ON=1'b0;
    defparam shift_srl_66_5_LC_24_12_5.SEQ_MODE=4'b1000;
    defparam shift_srl_66_5_LC_24_12_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_66_5_LC_24_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81634),
            .lcout(shift_srl_66Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93313),
            .ce(N__81681),
            .sr(_gnd_net_));
    defparam shift_srl_66_6_LC_24_12_6.C_ON=1'b0;
    defparam shift_srl_66_6_LC_24_12_6.SEQ_MODE=4'b1000;
    defparam shift_srl_66_6_LC_24_12_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_66_6_LC_24_12_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81628),
            .lcout(shift_srl_66Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93313),
            .ce(N__81681),
            .sr(_gnd_net_));
    defparam shift_srl_66_7_LC_24_12_7.C_ON=1'b0;
    defparam shift_srl_66_7_LC_24_12_7.SEQ_MODE=4'b1000;
    defparam shift_srl_66_7_LC_24_12_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_66_7_LC_24_12_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81622),
            .lcout(shift_srl_66Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93313),
            .ce(N__81681),
            .sr(_gnd_net_));
    defparam shift_srl_66_10_LC_24_13_0.C_ON=1'b0;
    defparam shift_srl_66_10_LC_24_13_0.SEQ_MODE=4'b1000;
    defparam shift_srl_66_10_LC_24_13_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_66_10_LC_24_13_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81703),
            .lcout(shift_srl_66Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93294),
            .ce(N__81685),
            .sr(_gnd_net_));
    defparam shift_srl_66_11_LC_24_13_1.C_ON=1'b0;
    defparam shift_srl_66_11_LC_24_13_1.SEQ_MODE=4'b1000;
    defparam shift_srl_66_11_LC_24_13_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_66_11_LC_24_13_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81616),
            .lcout(shift_srl_66Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93294),
            .ce(N__81685),
            .sr(_gnd_net_));
    defparam shift_srl_66_12_LC_24_13_2.C_ON=1'b0;
    defparam shift_srl_66_12_LC_24_13_2.SEQ_MODE=4'b1000;
    defparam shift_srl_66_12_LC_24_13_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_66_12_LC_24_13_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81610),
            .lcout(shift_srl_66Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93294),
            .ce(N__81685),
            .sr(_gnd_net_));
    defparam shift_srl_66_13_LC_24_13_3.C_ON=1'b0;
    defparam shift_srl_66_13_LC_24_13_3.SEQ_MODE=4'b1000;
    defparam shift_srl_66_13_LC_24_13_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_66_13_LC_24_13_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81604),
            .lcout(shift_srl_66Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93294),
            .ce(N__81685),
            .sr(_gnd_net_));
    defparam shift_srl_66_14_LC_24_13_4.C_ON=1'b0;
    defparam shift_srl_66_14_LC_24_13_4.SEQ_MODE=4'b1000;
    defparam shift_srl_66_14_LC_24_13_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_66_14_LC_24_13_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81598),
            .lcout(shift_srl_66Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93294),
            .ce(N__81685),
            .sr(_gnd_net_));
    defparam shift_srl_66_15_LC_24_13_5.C_ON=1'b0;
    defparam shift_srl_66_15_LC_24_13_5.SEQ_MODE=4'b1000;
    defparam shift_srl_66_15_LC_24_13_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_66_15_LC_24_13_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81727),
            .lcout(shift_srl_66Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93294),
            .ce(N__81685),
            .sr(_gnd_net_));
    defparam shift_srl_66_9_LC_24_13_6.C_ON=1'b0;
    defparam shift_srl_66_9_LC_24_13_6.SEQ_MODE=4'b1000;
    defparam shift_srl_66_9_LC_24_13_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_66_9_LC_24_13_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81691),
            .lcout(shift_srl_66Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93294),
            .ce(N__81685),
            .sr(_gnd_net_));
    defparam shift_srl_66_8_LC_24_13_7.C_ON=1'b0;
    defparam shift_srl_66_8_LC_24_13_7.SEQ_MODE=4'b1000;
    defparam shift_srl_66_8_LC_24_13_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_66_8_LC_24_13_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81697),
            .lcout(shift_srl_66Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93294),
            .ce(N__81685),
            .sr(_gnd_net_));
    defparam shift_srl_35_10_LC_24_14_0.C_ON=1'b0;
    defparam shift_srl_35_10_LC_24_14_0.SEQ_MODE=4'b1000;
    defparam shift_srl_35_10_LC_24_14_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_35_10_LC_24_14_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81775),
            .lcout(shift_srl_35Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93280),
            .ce(N__81822),
            .sr(_gnd_net_));
    defparam shift_srl_35_11_LC_24_14_1.C_ON=1'b0;
    defparam shift_srl_35_11_LC_24_14_1.SEQ_MODE=4'b1000;
    defparam shift_srl_35_11_LC_24_14_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_35_11_LC_24_14_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81670),
            .lcout(shift_srl_35Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93280),
            .ce(N__81822),
            .sr(_gnd_net_));
    defparam shift_srl_35_12_LC_24_14_2.C_ON=1'b0;
    defparam shift_srl_35_12_LC_24_14_2.SEQ_MODE=4'b1000;
    defparam shift_srl_35_12_LC_24_14_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_35_12_LC_24_14_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81664),
            .lcout(shift_srl_35Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93280),
            .ce(N__81822),
            .sr(_gnd_net_));
    defparam shift_srl_35_13_LC_24_14_3.C_ON=1'b0;
    defparam shift_srl_35_13_LC_24_14_3.SEQ_MODE=4'b1000;
    defparam shift_srl_35_13_LC_24_14_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_35_13_LC_24_14_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81658),
            .lcout(shift_srl_35Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93280),
            .ce(N__81822),
            .sr(_gnd_net_));
    defparam shift_srl_35_14_LC_24_14_4.C_ON=1'b0;
    defparam shift_srl_35_14_LC_24_14_4.SEQ_MODE=4'b1000;
    defparam shift_srl_35_14_LC_24_14_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_35_14_LC_24_14_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81652),
            .lcout(shift_srl_35Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93280),
            .ce(N__81822),
            .sr(_gnd_net_));
    defparam shift_srl_35_15_LC_24_14_5.C_ON=1'b0;
    defparam shift_srl_35_15_LC_24_14_5.SEQ_MODE=4'b1000;
    defparam shift_srl_35_15_LC_24_14_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_35_15_LC_24_14_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81646),
            .lcout(shift_srl_35Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93280),
            .ce(N__81822),
            .sr(_gnd_net_));
    defparam shift_srl_35_9_LC_24_14_6.C_ON=1'b0;
    defparam shift_srl_35_9_LC_24_14_6.SEQ_MODE=4'b1000;
    defparam shift_srl_35_9_LC_24_14_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_35_9_LC_24_14_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81769),
            .lcout(shift_srl_35Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93280),
            .ce(N__81822),
            .sr(_gnd_net_));
    defparam shift_srl_35_8_LC_24_14_7.C_ON=1'b0;
    defparam shift_srl_35_8_LC_24_14_7.SEQ_MODE=4'b1000;
    defparam shift_srl_35_8_LC_24_14_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_35_8_LC_24_14_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81835),
            .lcout(shift_srl_35Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93280),
            .ce(N__81822),
            .sr(_gnd_net_));
    defparam shift_srl_34_RNID6NU8_15_LC_24_15_0.C_ON=1'b0;
    defparam shift_srl_34_RNID6NU8_15_LC_24_15_0.SEQ_MODE=4'b0000;
    defparam shift_srl_34_RNID6NU8_15_LC_24_15_0.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_34_RNID6NU8_15_LC_24_15_0 (
            .in0(N__90458),
            .in1(N__83616),
            .in2(_gnd_net_),
            .in3(N__83338),
            .lcout(clk_en_35),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_34_15_LC_24_15_1.C_ON=1'b0;
    defparam shift_srl_34_15_LC_24_15_1.SEQ_MODE=4'b1000;
    defparam shift_srl_34_15_LC_24_15_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_34_15_LC_24_15_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81763),
            .lcout(shift_srl_34Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93261),
            .ce(N__87131),
            .sr(_gnd_net_));
    defparam shift_srl_34_14_LC_24_15_2.C_ON=1'b0;
    defparam shift_srl_34_14_LC_24_15_2.SEQ_MODE=4'b1000;
    defparam shift_srl_34_14_LC_24_15_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_34_14_LC_24_15_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81757),
            .lcout(shift_srl_34Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93261),
            .ce(N__87131),
            .sr(_gnd_net_));
    defparam shift_srl_34_13_LC_24_15_3.C_ON=1'b0;
    defparam shift_srl_34_13_LC_24_15_3.SEQ_MODE=4'b1000;
    defparam shift_srl_34_13_LC_24_15_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_34_13_LC_24_15_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81751),
            .lcout(shift_srl_34Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93261),
            .ce(N__87131),
            .sr(_gnd_net_));
    defparam shift_srl_34_12_LC_24_15_4.C_ON=1'b0;
    defparam shift_srl_34_12_LC_24_15_4.SEQ_MODE=4'b1000;
    defparam shift_srl_34_12_LC_24_15_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_34_12_LC_24_15_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81745),
            .lcout(shift_srl_34Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93261),
            .ce(N__87131),
            .sr(_gnd_net_));
    defparam shift_srl_34_11_LC_24_15_5.C_ON=1'b0;
    defparam shift_srl_34_11_LC_24_15_5.SEQ_MODE=4'b1000;
    defparam shift_srl_34_11_LC_24_15_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_34_11_LC_24_15_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81739),
            .lcout(shift_srl_34Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93261),
            .ce(N__87131),
            .sr(_gnd_net_));
    defparam shift_srl_34_10_LC_24_15_6.C_ON=1'b0;
    defparam shift_srl_34_10_LC_24_15_6.SEQ_MODE=4'b1000;
    defparam shift_srl_34_10_LC_24_15_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_34_10_LC_24_15_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81733),
            .lcout(shift_srl_34Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93261),
            .ce(N__87131),
            .sr(_gnd_net_));
    defparam shift_srl_34_9_LC_24_15_7.C_ON=1'b0;
    defparam shift_srl_34_9_LC_24_15_7.SEQ_MODE=4'b1000;
    defparam shift_srl_34_9_LC_24_15_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_34_9_LC_24_15_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87145),
            .lcout(shift_srl_34Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93261),
            .ce(N__87131),
            .sr(_gnd_net_));
    defparam shift_srl_35_0_LC_24_16_0.C_ON=1'b0;
    defparam shift_srl_35_0_LC_24_16_0.SEQ_MODE=4'b1000;
    defparam shift_srl_35_0_LC_24_16_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_35_0_LC_24_16_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81902),
            .lcout(shift_srl_35Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93239),
            .ce(N__81826),
            .sr(_gnd_net_));
    defparam shift_srl_35_1_LC_24_16_1.C_ON=1'b0;
    defparam shift_srl_35_1_LC_24_16_1.SEQ_MODE=4'b1000;
    defparam shift_srl_35_1_LC_24_16_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_35_1_LC_24_16_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81877),
            .lcout(shift_srl_35Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93239),
            .ce(N__81826),
            .sr(_gnd_net_));
    defparam shift_srl_35_2_LC_24_16_2.C_ON=1'b0;
    defparam shift_srl_35_2_LC_24_16_2.SEQ_MODE=4'b1000;
    defparam shift_srl_35_2_LC_24_16_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_35_2_LC_24_16_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81871),
            .lcout(shift_srl_35Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93239),
            .ce(N__81826),
            .sr(_gnd_net_));
    defparam shift_srl_35_3_LC_24_16_3.C_ON=1'b0;
    defparam shift_srl_35_3_LC_24_16_3.SEQ_MODE=4'b1000;
    defparam shift_srl_35_3_LC_24_16_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_35_3_LC_24_16_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81865),
            .lcout(shift_srl_35Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93239),
            .ce(N__81826),
            .sr(_gnd_net_));
    defparam shift_srl_35_4_LC_24_16_4.C_ON=1'b0;
    defparam shift_srl_35_4_LC_24_16_4.SEQ_MODE=4'b1000;
    defparam shift_srl_35_4_LC_24_16_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_35_4_LC_24_16_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81859),
            .lcout(shift_srl_35Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93239),
            .ce(N__81826),
            .sr(_gnd_net_));
    defparam shift_srl_35_5_LC_24_16_5.C_ON=1'b0;
    defparam shift_srl_35_5_LC_24_16_5.SEQ_MODE=4'b1000;
    defparam shift_srl_35_5_LC_24_16_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_35_5_LC_24_16_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81853),
            .lcout(shift_srl_35Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93239),
            .ce(N__81826),
            .sr(_gnd_net_));
    defparam shift_srl_35_6_LC_24_16_6.C_ON=1'b0;
    defparam shift_srl_35_6_LC_24_16_6.SEQ_MODE=4'b1000;
    defparam shift_srl_35_6_LC_24_16_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_35_6_LC_24_16_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81847),
            .lcout(shift_srl_35Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93239),
            .ce(N__81826),
            .sr(_gnd_net_));
    defparam shift_srl_35_7_LC_24_16_7.C_ON=1'b0;
    defparam shift_srl_35_7_LC_24_16_7.SEQ_MODE=4'b1000;
    defparam shift_srl_35_7_LC_24_16_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_35_7_LC_24_16_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81841),
            .lcout(shift_srl_35Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93239),
            .ce(N__81826),
            .sr(_gnd_net_));
    defparam shift_srl_39_0_LC_24_17_0.C_ON=1'b0;
    defparam shift_srl_39_0_LC_24_17_0.SEQ_MODE=4'b1000;
    defparam shift_srl_39_0_LC_24_17_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_39_0_LC_24_17_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81808),
            .lcout(shift_srl_39Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93198),
            .ce(N__82016),
            .sr(_gnd_net_));
    defparam shift_srl_39_1_LC_24_17_1.C_ON=1'b0;
    defparam shift_srl_39_1_LC_24_17_1.SEQ_MODE=4'b1000;
    defparam shift_srl_39_1_LC_24_17_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_39_1_LC_24_17_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81958),
            .lcout(shift_srl_39Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93198),
            .ce(N__82016),
            .sr(_gnd_net_));
    defparam shift_srl_39_2_LC_24_17_2.C_ON=1'b0;
    defparam shift_srl_39_2_LC_24_17_2.SEQ_MODE=4'b1000;
    defparam shift_srl_39_2_LC_24_17_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_39_2_LC_24_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81952),
            .lcout(shift_srl_39Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93198),
            .ce(N__82016),
            .sr(_gnd_net_));
    defparam shift_srl_39_3_LC_24_17_3.C_ON=1'b0;
    defparam shift_srl_39_3_LC_24_17_3.SEQ_MODE=4'b1000;
    defparam shift_srl_39_3_LC_24_17_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_39_3_LC_24_17_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81946),
            .lcout(shift_srl_39Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93198),
            .ce(N__82016),
            .sr(_gnd_net_));
    defparam shift_srl_39_4_LC_24_17_4.C_ON=1'b0;
    defparam shift_srl_39_4_LC_24_17_4.SEQ_MODE=4'b1000;
    defparam shift_srl_39_4_LC_24_17_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_39_4_LC_24_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81940),
            .lcout(shift_srl_39Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93198),
            .ce(N__82016),
            .sr(_gnd_net_));
    defparam shift_srl_39_5_LC_24_17_5.C_ON=1'b0;
    defparam shift_srl_39_5_LC_24_17_5.SEQ_MODE=4'b1000;
    defparam shift_srl_39_5_LC_24_17_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_39_5_LC_24_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81934),
            .lcout(shift_srl_39Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93198),
            .ce(N__82016),
            .sr(_gnd_net_));
    defparam shift_srl_39_6_LC_24_17_6.C_ON=1'b0;
    defparam shift_srl_39_6_LC_24_17_6.SEQ_MODE=4'b1000;
    defparam shift_srl_39_6_LC_24_17_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_39_6_LC_24_17_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81928),
            .lcout(shift_srl_39Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93198),
            .ce(N__82016),
            .sr(_gnd_net_));
    defparam shift_srl_39_7_LC_24_17_7.C_ON=1'b0;
    defparam shift_srl_39_7_LC_24_17_7.SEQ_MODE=4'b1000;
    defparam shift_srl_39_7_LC_24_17_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_39_7_LC_24_17_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81922),
            .lcout(shift_srl_39Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93198),
            .ce(N__82016),
            .sr(_gnd_net_));
    defparam shift_srl_169_4_LC_24_18_0.C_ON=1'b0;
    defparam shift_srl_169_4_LC_24_18_0.SEQ_MODE=4'b1000;
    defparam shift_srl_169_4_LC_24_18_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_169_4_LC_24_18_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81976),
            .lcout(shift_srl_169Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93240),
            .ce(N__82549),
            .sr(_gnd_net_));
    defparam shift_srl_169_5_LC_24_18_1.C_ON=1'b0;
    defparam shift_srl_169_5_LC_24_18_1.SEQ_MODE=4'b1000;
    defparam shift_srl_169_5_LC_24_18_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_169_5_LC_24_18_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81916),
            .lcout(shift_srl_169Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93240),
            .ce(N__82549),
            .sr(_gnd_net_));
    defparam shift_srl_169_6_LC_24_18_2.C_ON=1'b0;
    defparam shift_srl_169_6_LC_24_18_2.SEQ_MODE=4'b1000;
    defparam shift_srl_169_6_LC_24_18_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_169_6_LC_24_18_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82066),
            .lcout(shift_srl_169Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93240),
            .ce(N__82549),
            .sr(_gnd_net_));
    defparam shift_srl_169_7_LC_24_18_3.C_ON=1'b0;
    defparam shift_srl_169_7_LC_24_18_3.SEQ_MODE=4'b1000;
    defparam shift_srl_169_7_LC_24_18_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_169_7_LC_24_18_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82060),
            .lcout(shift_srl_169Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93240),
            .ce(N__82549),
            .sr(_gnd_net_));
    defparam shift_srl_169_12_LC_24_18_5.C_ON=1'b0;
    defparam shift_srl_169_12_LC_24_18_5.SEQ_MODE=4'b1000;
    defparam shift_srl_169_12_LC_24_18_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_169_12_LC_24_18_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81994),
            .lcout(shift_srl_169Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93240),
            .ce(N__82549),
            .sr(_gnd_net_));
    defparam shift_srl_169_2_LC_24_18_7.C_ON=1'b0;
    defparam shift_srl_169_2_LC_24_18_7.SEQ_MODE=4'b1000;
    defparam shift_srl_169_2_LC_24_18_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_169_2_LC_24_18_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82558),
            .lcout(shift_srl_169Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93240),
            .ce(N__82549),
            .sr(_gnd_net_));
    defparam shift_srl_39_8_LC_24_19_0.C_ON=1'b0;
    defparam shift_srl_39_8_LC_24_19_0.SEQ_MODE=4'b1000;
    defparam shift_srl_39_8_LC_24_19_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_39_8_LC_24_19_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82054),
            .lcout(shift_srl_39Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93262),
            .ce(N__82023),
            .sr(_gnd_net_));
    defparam shift_srl_169_10_LC_24_20_0.C_ON=1'b0;
    defparam shift_srl_169_10_LC_24_20_0.SEQ_MODE=4'b1000;
    defparam shift_srl_169_10_LC_24_20_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_169_10_LC_24_20_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82456),
            .lcout(shift_srl_169Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93281),
            .ce(N__82545),
            .sr(_gnd_net_));
    defparam shift_srl_169_11_LC_24_20_1.C_ON=1'b0;
    defparam shift_srl_169_11_LC_24_20_1.SEQ_MODE=4'b1000;
    defparam shift_srl_169_11_LC_24_20_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_169_11_LC_24_20_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82000),
            .lcout(shift_srl_169Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93281),
            .ce(N__82545),
            .sr(_gnd_net_));
    defparam shift_srl_169_3_LC_24_20_2.C_ON=1'b0;
    defparam shift_srl_169_3_LC_24_20_2.SEQ_MODE=4'b1000;
    defparam shift_srl_169_3_LC_24_20_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_169_3_LC_24_20_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81985),
            .lcout(shift_srl_169Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93281),
            .ce(N__82545),
            .sr(_gnd_net_));
    defparam shift_srl_169_13_LC_24_20_3.C_ON=1'b0;
    defparam shift_srl_169_13_LC_24_20_3.SEQ_MODE=4'b1000;
    defparam shift_srl_169_13_LC_24_20_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_169_13_LC_24_20_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81967),
            .lcout(shift_srl_169Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93281),
            .ce(N__82545),
            .sr(_gnd_net_));
    defparam shift_srl_169_14_LC_24_20_4.C_ON=1'b0;
    defparam shift_srl_169_14_LC_24_20_4.SEQ_MODE=4'b1000;
    defparam shift_srl_169_14_LC_24_20_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_169_14_LC_24_20_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82468),
            .lcout(shift_srl_169Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93281),
            .ce(N__82545),
            .sr(_gnd_net_));
    defparam shift_srl_169_15_LC_24_20_5.C_ON=1'b0;
    defparam shift_srl_169_15_LC_24_20_5.SEQ_MODE=4'b1000;
    defparam shift_srl_169_15_LC_24_20_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_169_15_LC_24_20_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82462),
            .lcout(shift_srl_169Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93281),
            .ce(N__82545),
            .sr(_gnd_net_));
    defparam shift_srl_169_9_LC_24_20_6.C_ON=1'b0;
    defparam shift_srl_169_9_LC_24_20_6.SEQ_MODE=4'b1000;
    defparam shift_srl_169_9_LC_24_20_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_169_9_LC_24_20_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82441),
            .lcout(shift_srl_169Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93281),
            .ce(N__82545),
            .sr(_gnd_net_));
    defparam shift_srl_169_8_LC_24_20_7.C_ON=1'b0;
    defparam shift_srl_169_8_LC_24_20_7.SEQ_MODE=4'b1000;
    defparam shift_srl_169_8_LC_24_20_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_169_8_LC_24_20_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82450),
            .lcout(shift_srl_169Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93281),
            .ce(N__82545),
            .sr(_gnd_net_));
    defparam shift_srl_166_RNIFH9M91_15_LC_24_21_0.C_ON=1'b0;
    defparam shift_srl_166_RNIFH9M91_15_LC_24_21_0.SEQ_MODE=4'b0000;
    defparam shift_srl_166_RNIFH9M91_15_LC_24_21_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_166_RNIFH9M91_15_LC_24_21_0 (
            .in0(N__84016),
            .in1(N__83965),
            .in2(N__82427),
            .in3(N__85796),
            .lcout(clk_en_167),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNILKVP81_15_LC_24_21_1.C_ON=1'b0;
    defparam shift_srl_0_RNILKVP81_15_LC_24_21_1.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNILKVP81_15_LC_24_21_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNILKVP81_15_LC_24_21_1 (
            .in0(N__87996),
            .in1(N__82339),
            .in2(N__90493),
            .in3(N__82160),
            .lcout(clk_en_163),
            .ltout(clk_en_163_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_169_RNID9HFA1_15_LC_24_21_2.C_ON=1'b0;
    defparam shift_srl_169_RNID9HFA1_15_LC_24_21_2.SEQ_MODE=4'b0000;
    defparam shift_srl_169_RNID9HFA1_15_LC_24_21_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_169_RNID9HFA1_15_LC_24_21_2 (
            .in0(N__84271),
            .in1(N__89178),
            .in2(N__82069),
            .in3(N__87429),
            .lcout(clk_en_170),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_168_RNI28JDA1_15_LC_24_21_3.C_ON=1'b0;
    defparam shift_srl_168_RNI28JDA1_15_LC_24_21_3.SEQ_MODE=4'b0000;
    defparam shift_srl_168_RNI28JDA1_15_LC_24_21_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_168_RNI28JDA1_15_LC_24_21_3 (
            .in0(N__89179),
            .in1(N__90370),
            .in2(N__87430),
            .in3(N__87698),
            .lcout(clk_en_169),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_169_0_LC_24_21_4.C_ON=1'b0;
    defparam shift_srl_169_0_LC_24_21_4.SEQ_MODE=4'b1000;
    defparam shift_srl_169_0_LC_24_21_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_169_0_LC_24_21_4 (
            .in0(N__84272),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_169Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93295),
            .ce(N__82544),
            .sr(_gnd_net_));
    defparam shift_srl_169_1_LC_24_21_5.C_ON=1'b0;
    defparam shift_srl_169_1_LC_24_21_5.SEQ_MODE=4'b1000;
    defparam shift_srl_169_1_LC_24_21_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_169_1_LC_24_21_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82564),
            .lcout(shift_srl_169Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93295),
            .ce(N__82544),
            .sr(_gnd_net_));
    defparam shift_srl_170_10_LC_24_22_0.C_ON=1'b0;
    defparam shift_srl_170_10_LC_24_22_0.SEQ_MODE=4'b1000;
    defparam shift_srl_170_10_LC_24_22_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_170_10_LC_24_22_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82498),
            .lcout(shift_srl_170Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93314),
            .ce(N__82479),
            .sr(_gnd_net_));
    defparam shift_srl_170_11_LC_24_22_1.C_ON=1'b0;
    defparam shift_srl_170_11_LC_24_22_1.SEQ_MODE=4'b1000;
    defparam shift_srl_170_11_LC_24_22_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_170_11_LC_24_22_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82528),
            .lcout(shift_srl_170Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93314),
            .ce(N__82479),
            .sr(_gnd_net_));
    defparam shift_srl_170_12_LC_24_22_2.C_ON=1'b0;
    defparam shift_srl_170_12_LC_24_22_2.SEQ_MODE=4'b1000;
    defparam shift_srl_170_12_LC_24_22_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_170_12_LC_24_22_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82522),
            .lcout(shift_srl_170Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93314),
            .ce(N__82479),
            .sr(_gnd_net_));
    defparam shift_srl_170_13_LC_24_22_3.C_ON=1'b0;
    defparam shift_srl_170_13_LC_24_22_3.SEQ_MODE=4'b1000;
    defparam shift_srl_170_13_LC_24_22_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_170_13_LC_24_22_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82516),
            .lcout(shift_srl_170Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93314),
            .ce(N__82479),
            .sr(_gnd_net_));
    defparam shift_srl_170_14_LC_24_22_4.C_ON=1'b0;
    defparam shift_srl_170_14_LC_24_22_4.SEQ_MODE=4'b1000;
    defparam shift_srl_170_14_LC_24_22_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_170_14_LC_24_22_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82510),
            .lcout(shift_srl_170Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93314),
            .ce(N__82479),
            .sr(_gnd_net_));
    defparam shift_srl_170_15_LC_24_22_5.C_ON=1'b0;
    defparam shift_srl_170_15_LC_24_22_5.SEQ_MODE=4'b1000;
    defparam shift_srl_170_15_LC_24_22_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_170_15_LC_24_22_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82504),
            .lcout(shift_srl_170Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93314),
            .ce(N__82479),
            .sr(_gnd_net_));
    defparam shift_srl_170_9_LC_24_22_6.C_ON=1'b0;
    defparam shift_srl_170_9_LC_24_22_6.SEQ_MODE=4'b1000;
    defparam shift_srl_170_9_LC_24_22_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_170_9_LC_24_22_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82486),
            .lcout(shift_srl_170Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93314),
            .ce(N__82479),
            .sr(_gnd_net_));
    defparam shift_srl_170_8_LC_24_22_7.C_ON=1'b0;
    defparam shift_srl_170_8_LC_24_22_7.SEQ_MODE=4'b1000;
    defparam shift_srl_170_8_LC_24_22_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_170_8_LC_24_22_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82492),
            .lcout(shift_srl_170Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93314),
            .ce(N__82479),
            .sr(_gnd_net_));
    defparam shift_srl_177_10_LC_24_23_0.C_ON=1'b0;
    defparam shift_srl_177_10_LC_24_23_0.SEQ_MODE=4'b1000;
    defparam shift_srl_177_10_LC_24_23_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_177_10_LC_24_23_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82624),
            .lcout(shift_srl_177Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93334),
            .ce(N__82606),
            .sr(_gnd_net_));
    defparam shift_srl_177_11_LC_24_23_1.C_ON=1'b0;
    defparam shift_srl_177_11_LC_24_23_1.SEQ_MODE=4'b1000;
    defparam shift_srl_177_11_LC_24_23_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_177_11_LC_24_23_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82648),
            .lcout(shift_srl_177Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93334),
            .ce(N__82606),
            .sr(_gnd_net_));
    defparam shift_srl_177_12_LC_24_23_2.C_ON=1'b0;
    defparam shift_srl_177_12_LC_24_23_2.SEQ_MODE=4'b1000;
    defparam shift_srl_177_12_LC_24_23_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_177_12_LC_24_23_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82642),
            .lcout(shift_srl_177Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93334),
            .ce(N__82606),
            .sr(_gnd_net_));
    defparam shift_srl_177_7_LC_24_23_3.C_ON=1'b0;
    defparam shift_srl_177_7_LC_24_23_3.SEQ_MODE=4'b1000;
    defparam shift_srl_177_7_LC_24_23_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_177_7_LC_24_23_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82630),
            .lcout(shift_srl_177Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93334),
            .ce(N__82606),
            .sr(_gnd_net_));
    defparam shift_srl_177_9_LC_24_23_4.C_ON=1'b0;
    defparam shift_srl_177_9_LC_24_23_4.SEQ_MODE=4'b1000;
    defparam shift_srl_177_9_LC_24_23_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_177_9_LC_24_23_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82612),
            .lcout(shift_srl_177Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93334),
            .ce(N__82606),
            .sr(_gnd_net_));
    defparam shift_srl_177_8_LC_24_23_5.C_ON=1'b0;
    defparam shift_srl_177_8_LC_24_23_5.SEQ_MODE=4'b1000;
    defparam shift_srl_177_8_LC_24_23_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_177_8_LC_24_23_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82618),
            .lcout(shift_srl_177Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93334),
            .ce(N__82606),
            .sr(_gnd_net_));
    defparam shift_srl_180_10_LC_24_24_0.C_ON=1'b0;
    defparam shift_srl_180_10_LC_24_24_0.SEQ_MODE=4'b1000;
    defparam shift_srl_180_10_LC_24_24_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_180_10_LC_24_24_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82696),
            .lcout(shift_srl_180Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93356),
            .ce(N__82690),
            .sr(_gnd_net_));
    defparam shift_srl_180_11_LC_24_24_1.C_ON=1'b0;
    defparam shift_srl_180_11_LC_24_24_1.SEQ_MODE=4'b1000;
    defparam shift_srl_180_11_LC_24_24_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_180_11_LC_24_24_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82582),
            .lcout(shift_srl_180Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93356),
            .ce(N__82690),
            .sr(_gnd_net_));
    defparam shift_srl_180_5_LC_24_24_2.C_ON=1'b0;
    defparam shift_srl_180_5_LC_24_24_2.SEQ_MODE=4'b1000;
    defparam shift_srl_180_5_LC_24_24_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_180_5_LC_24_24_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82576),
            .lcout(shift_srl_180Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93356),
            .ce(N__82690),
            .sr(_gnd_net_));
    defparam shift_srl_180_13_LC_24_24_3.C_ON=1'b0;
    defparam shift_srl_180_13_LC_24_24_3.SEQ_MODE=4'b1000;
    defparam shift_srl_180_13_LC_24_24_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_180_13_LC_24_24_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82708),
            .lcout(shift_srl_180Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93356),
            .ce(N__82690),
            .sr(_gnd_net_));
    defparam shift_srl_180_14_LC_24_24_4.C_ON=1'b0;
    defparam shift_srl_180_14_LC_24_24_4.SEQ_MODE=4'b1000;
    defparam shift_srl_180_14_LC_24_24_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_180_14_LC_24_24_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82765),
            .lcout(shift_srl_180Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93356),
            .ce(N__82690),
            .sr(_gnd_net_));
    defparam shift_srl_180_15_LC_24_24_5.C_ON=1'b0;
    defparam shift_srl_180_15_LC_24_24_5.SEQ_MODE=4'b1000;
    defparam shift_srl_180_15_LC_24_24_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_180_15_LC_24_24_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82759),
            .lcout(shift_srl_180Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93356),
            .ce(N__82690),
            .sr(_gnd_net_));
    defparam shift_srl_180_12_LC_24_24_6.C_ON=1'b0;
    defparam shift_srl_180_12_LC_24_24_6.SEQ_MODE=4'b1000;
    defparam shift_srl_180_12_LC_24_24_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_180_12_LC_24_24_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82714),
            .lcout(shift_srl_180Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93356),
            .ce(N__82690),
            .sr(_gnd_net_));
    defparam shift_srl_180_9_LC_24_24_7.C_ON=1'b0;
    defparam shift_srl_180_9_LC_24_24_7.SEQ_MODE=4'b1000;
    defparam shift_srl_180_9_LC_24_24_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_180_9_LC_24_24_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82702),
            .lcout(shift_srl_180Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93356),
            .ce(N__82690),
            .sr(_gnd_net_));
    defparam shift_srl_189_0_LC_24_25_0.C_ON=1'b0;
    defparam shift_srl_189_0_LC_24_25_0.SEQ_MODE=4'b1000;
    defparam shift_srl_189_0_LC_24_25_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_189_0_LC_24_25_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86135),
            .lcout(shift_srl_189Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93371),
            .ce(N__82845),
            .sr(_gnd_net_));
    defparam shift_srl_189_1_LC_24_25_1.C_ON=1'b0;
    defparam shift_srl_189_1_LC_24_25_1.SEQ_MODE=4'b1000;
    defparam shift_srl_189_1_LC_24_25_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_189_1_LC_24_25_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82666),
            .lcout(shift_srl_189Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93371),
            .ce(N__82845),
            .sr(_gnd_net_));
    defparam shift_srl_189_2_LC_24_25_2.C_ON=1'b0;
    defparam shift_srl_189_2_LC_24_25_2.SEQ_MODE=4'b1000;
    defparam shift_srl_189_2_LC_24_25_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_189_2_LC_24_25_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82660),
            .lcout(shift_srl_189Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93371),
            .ce(N__82845),
            .sr(_gnd_net_));
    defparam shift_srl_189_3_LC_24_25_3.C_ON=1'b0;
    defparam shift_srl_189_3_LC_24_25_3.SEQ_MODE=4'b1000;
    defparam shift_srl_189_3_LC_24_25_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_189_3_LC_24_25_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82654),
            .lcout(shift_srl_189Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93371),
            .ce(N__82845),
            .sr(_gnd_net_));
    defparam shift_srl_189_4_LC_24_25_4.C_ON=1'b0;
    defparam shift_srl_189_4_LC_24_25_4.SEQ_MODE=4'b1000;
    defparam shift_srl_189_4_LC_24_25_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_189_4_LC_24_25_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82879),
            .lcout(shift_srl_189Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93371),
            .ce(N__82845),
            .sr(_gnd_net_));
    defparam shift_srl_189_5_LC_24_25_5.C_ON=1'b0;
    defparam shift_srl_189_5_LC_24_25_5.SEQ_MODE=4'b1000;
    defparam shift_srl_189_5_LC_24_25_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_189_5_LC_24_25_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82873),
            .lcout(shift_srl_189Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93371),
            .ce(N__82845),
            .sr(_gnd_net_));
    defparam shift_srl_189_6_LC_24_25_6.C_ON=1'b0;
    defparam shift_srl_189_6_LC_24_25_6.SEQ_MODE=4'b1000;
    defparam shift_srl_189_6_LC_24_25_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_189_6_LC_24_25_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82867),
            .lcout(shift_srl_189Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93371),
            .ce(N__82845),
            .sr(_gnd_net_));
    defparam shift_srl_189_7_LC_24_25_7.C_ON=1'b0;
    defparam shift_srl_189_7_LC_24_25_7.SEQ_MODE=4'b1000;
    defparam shift_srl_189_7_LC_24_25_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_189_7_LC_24_25_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82861),
            .lcout(shift_srl_189Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93371),
            .ce(N__82845),
            .sr(_gnd_net_));
    defparam shift_srl_188_8_LC_24_26_0.C_ON=1'b0;
    defparam shift_srl_188_8_LC_24_26_0.SEQ_MODE=4'b1000;
    defparam shift_srl_188_8_LC_24_26_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_188_8_LC_24_26_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82825),
            .lcout(shift_srl_188Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93388),
            .ce(N__82796),
            .sr(_gnd_net_));
    defparam shift_srl_188_9_LC_24_26_1.C_ON=1'b0;
    defparam shift_srl_188_9_LC_24_26_1.SEQ_MODE=4'b1000;
    defparam shift_srl_188_9_LC_24_26_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_188_9_LC_24_26_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82816),
            .lcout(shift_srl_188Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93388),
            .ce(N__82796),
            .sr(_gnd_net_));
    defparam shift_srl_80_8_LC_26_5_0.C_ON=1'b0;
    defparam shift_srl_80_8_LC_26_5_0.SEQ_MODE=4'b1000;
    defparam shift_srl_80_8_LC_26_5_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_80_8_LC_26_5_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82897),
            .lcout(shift_srl_80Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93421),
            .ce(N__84613),
            .sr(_gnd_net_));
    defparam shift_srl_80_0_LC_26_6_0.C_ON=1'b0;
    defparam shift_srl_80_0_LC_26_6_0.SEQ_MODE=4'b1000;
    defparam shift_srl_80_0_LC_26_6_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_80_0_LC_26_6_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84678),
            .lcout(shift_srl_80Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93416),
            .ce(N__84605),
            .sr(_gnd_net_));
    defparam shift_srl_80_1_LC_26_6_1.C_ON=1'b0;
    defparam shift_srl_80_1_LC_26_6_1.SEQ_MODE=4'b1000;
    defparam shift_srl_80_1_LC_26_6_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_80_1_LC_26_6_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82771),
            .lcout(shift_srl_80Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93416),
            .ce(N__84605),
            .sr(_gnd_net_));
    defparam shift_srl_80_2_LC_26_6_2.C_ON=1'b0;
    defparam shift_srl_80_2_LC_26_6_2.SEQ_MODE=4'b1000;
    defparam shift_srl_80_2_LC_26_6_2.LUT_INIT=16'b1100110011001100;
    LogicCell40 shift_srl_80_2_LC_26_6_2 (
            .in0(_gnd_net_),
            .in1(N__82933),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_80Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93416),
            .ce(N__84605),
            .sr(_gnd_net_));
    defparam shift_srl_80_3_LC_26_6_3.C_ON=1'b0;
    defparam shift_srl_80_3_LC_26_6_3.SEQ_MODE=4'b1000;
    defparam shift_srl_80_3_LC_26_6_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_80_3_LC_26_6_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82927),
            .lcout(shift_srl_80Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93416),
            .ce(N__84605),
            .sr(_gnd_net_));
    defparam shift_srl_80_4_LC_26_6_4.C_ON=1'b0;
    defparam shift_srl_80_4_LC_26_6_4.SEQ_MODE=4'b1000;
    defparam shift_srl_80_4_LC_26_6_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_80_4_LC_26_6_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82921),
            .lcout(shift_srl_80Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93416),
            .ce(N__84605),
            .sr(_gnd_net_));
    defparam shift_srl_80_5_LC_26_6_5.C_ON=1'b0;
    defparam shift_srl_80_5_LC_26_6_5.SEQ_MODE=4'b1000;
    defparam shift_srl_80_5_LC_26_6_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_80_5_LC_26_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82915),
            .lcout(shift_srl_80Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93416),
            .ce(N__84605),
            .sr(_gnd_net_));
    defparam shift_srl_80_6_LC_26_6_6.C_ON=1'b0;
    defparam shift_srl_80_6_LC_26_6_6.SEQ_MODE=4'b1000;
    defparam shift_srl_80_6_LC_26_6_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_80_6_LC_26_6_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82909),
            .lcout(shift_srl_80Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93416),
            .ce(N__84605),
            .sr(_gnd_net_));
    defparam shift_srl_80_7_LC_26_6_7.C_ON=1'b0;
    defparam shift_srl_80_7_LC_26_6_7.SEQ_MODE=4'b1000;
    defparam shift_srl_80_7_LC_26_6_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_80_7_LC_26_6_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82903),
            .lcout(shift_srl_80Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93416),
            .ce(N__84605),
            .sr(_gnd_net_));
    defparam shift_srl_78_10_LC_26_7_0.C_ON=1'b0;
    defparam shift_srl_78_10_LC_26_7_0.SEQ_MODE=4'b1000;
    defparam shift_srl_78_10_LC_26_7_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_78_10_LC_26_7_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82963),
            .lcout(shift_srl_78Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93412),
            .ce(N__84730),
            .sr(_gnd_net_));
    defparam shift_srl_78_11_LC_26_7_1.C_ON=1'b0;
    defparam shift_srl_78_11_LC_26_7_1.SEQ_MODE=4'b1000;
    defparam shift_srl_78_11_LC_26_7_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_78_11_LC_26_7_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82891),
            .lcout(shift_srl_78Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93412),
            .ce(N__84730),
            .sr(_gnd_net_));
    defparam shift_srl_78_12_LC_26_7_2.C_ON=1'b0;
    defparam shift_srl_78_12_LC_26_7_2.SEQ_MODE=4'b1000;
    defparam shift_srl_78_12_LC_26_7_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_78_12_LC_26_7_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82885),
            .lcout(shift_srl_78Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93412),
            .ce(N__84730),
            .sr(_gnd_net_));
    defparam shift_srl_78_13_LC_26_7_3.C_ON=1'b0;
    defparam shift_srl_78_13_LC_26_7_3.SEQ_MODE=4'b1000;
    defparam shift_srl_78_13_LC_26_7_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_78_13_LC_26_7_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82981),
            .lcout(shift_srl_78Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93412),
            .ce(N__84730),
            .sr(_gnd_net_));
    defparam shift_srl_78_14_LC_26_7_4.C_ON=1'b0;
    defparam shift_srl_78_14_LC_26_7_4.SEQ_MODE=4'b1000;
    defparam shift_srl_78_14_LC_26_7_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_78_14_LC_26_7_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82975),
            .lcout(shift_srl_78Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93412),
            .ce(N__84730),
            .sr(_gnd_net_));
    defparam shift_srl_78_15_LC_26_7_5.C_ON=1'b0;
    defparam shift_srl_78_15_LC_26_7_5.SEQ_MODE=4'b1000;
    defparam shift_srl_78_15_LC_26_7_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_78_15_LC_26_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82969),
            .lcout(shift_srl_78Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93412),
            .ce(N__84730),
            .sr(_gnd_net_));
    defparam shift_srl_78_9_LC_26_7_6.C_ON=1'b0;
    defparam shift_srl_78_9_LC_26_7_6.SEQ_MODE=4'b1000;
    defparam shift_srl_78_9_LC_26_7_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_78_9_LC_26_7_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82957),
            .lcout(shift_srl_78Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93412),
            .ce(N__84730),
            .sr(_gnd_net_));
    defparam shift_srl_78_8_LC_26_7_7.C_ON=1'b0;
    defparam shift_srl_78_8_LC_26_7_7.SEQ_MODE=4'b1000;
    defparam shift_srl_78_8_LC_26_7_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_78_8_LC_26_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83011),
            .lcout(shift_srl_78Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93412),
            .ce(N__84730),
            .sr(_gnd_net_));
    defparam shift_srl_78_0_LC_26_8_0.C_ON=1'b0;
    defparam shift_srl_78_0_LC_26_8_0.SEQ_MODE=4'b1000;
    defparam shift_srl_78_0_LC_26_8_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_78_0_LC_26_8_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84507),
            .lcout(shift_srl_78Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93405),
            .ce(N__84729),
            .sr(_gnd_net_));
    defparam shift_srl_78_1_LC_26_8_1.C_ON=1'b0;
    defparam shift_srl_78_1_LC_26_8_1.SEQ_MODE=4'b1000;
    defparam shift_srl_78_1_LC_26_8_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_78_1_LC_26_8_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82951),
            .lcout(shift_srl_78Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93405),
            .ce(N__84729),
            .sr(_gnd_net_));
    defparam shift_srl_78_2_LC_26_8_2.C_ON=1'b0;
    defparam shift_srl_78_2_LC_26_8_2.SEQ_MODE=4'b1000;
    defparam shift_srl_78_2_LC_26_8_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_78_2_LC_26_8_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82945),
            .lcout(shift_srl_78Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93405),
            .ce(N__84729),
            .sr(_gnd_net_));
    defparam shift_srl_78_3_LC_26_8_3.C_ON=1'b0;
    defparam shift_srl_78_3_LC_26_8_3.SEQ_MODE=4'b1000;
    defparam shift_srl_78_3_LC_26_8_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_78_3_LC_26_8_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82939),
            .lcout(shift_srl_78Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93405),
            .ce(N__84729),
            .sr(_gnd_net_));
    defparam shift_srl_78_4_LC_26_8_4.C_ON=1'b0;
    defparam shift_srl_78_4_LC_26_8_4.SEQ_MODE=4'b1000;
    defparam shift_srl_78_4_LC_26_8_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_78_4_LC_26_8_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83035),
            .lcout(shift_srl_78Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93405),
            .ce(N__84729),
            .sr(_gnd_net_));
    defparam shift_srl_78_5_LC_26_8_5.C_ON=1'b0;
    defparam shift_srl_78_5_LC_26_8_5.SEQ_MODE=4'b1000;
    defparam shift_srl_78_5_LC_26_8_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_78_5_LC_26_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83029),
            .lcout(shift_srl_78Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93405),
            .ce(N__84729),
            .sr(_gnd_net_));
    defparam shift_srl_78_6_LC_26_8_6.C_ON=1'b0;
    defparam shift_srl_78_6_LC_26_8_6.SEQ_MODE=4'b1000;
    defparam shift_srl_78_6_LC_26_8_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_78_6_LC_26_8_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83023),
            .lcout(shift_srl_78Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93405),
            .ce(N__84729),
            .sr(_gnd_net_));
    defparam shift_srl_78_7_LC_26_8_7.C_ON=1'b0;
    defparam shift_srl_78_7_LC_26_8_7.SEQ_MODE=4'b1000;
    defparam shift_srl_78_7_LC_26_8_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_78_7_LC_26_8_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83017),
            .lcout(shift_srl_78Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93405),
            .ce(N__84729),
            .sr(_gnd_net_));
    defparam shift_srl_69_0_LC_26_9_0.C_ON=1'b0;
    defparam shift_srl_69_0_LC_26_9_0.SEQ_MODE=4'b1000;
    defparam shift_srl_69_0_LC_26_9_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_69_0_LC_26_9_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86665),
            .lcout(shift_srl_69Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93397),
            .ce(N__85421),
            .sr(_gnd_net_));
    defparam shift_srl_69_1_LC_26_9_1.C_ON=1'b0;
    defparam shift_srl_69_1_LC_26_9_1.SEQ_MODE=4'b1000;
    defparam shift_srl_69_1_LC_26_9_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_69_1_LC_26_9_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83005),
            .lcout(shift_srl_69Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93397),
            .ce(N__85421),
            .sr(_gnd_net_));
    defparam shift_srl_69_2_LC_26_9_2.C_ON=1'b0;
    defparam shift_srl_69_2_LC_26_9_2.SEQ_MODE=4'b1000;
    defparam shift_srl_69_2_LC_26_9_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_69_2_LC_26_9_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82999),
            .lcout(shift_srl_69Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93397),
            .ce(N__85421),
            .sr(_gnd_net_));
    defparam shift_srl_69_3_LC_26_9_3.C_ON=1'b0;
    defparam shift_srl_69_3_LC_26_9_3.SEQ_MODE=4'b1000;
    defparam shift_srl_69_3_LC_26_9_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_69_3_LC_26_9_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82993),
            .lcout(shift_srl_69Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93397),
            .ce(N__85421),
            .sr(_gnd_net_));
    defparam shift_srl_69_4_LC_26_9_4.C_ON=1'b0;
    defparam shift_srl_69_4_LC_26_9_4.SEQ_MODE=4'b1000;
    defparam shift_srl_69_4_LC_26_9_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_69_4_LC_26_9_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82987),
            .lcout(shift_srl_69Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93397),
            .ce(N__85421),
            .sr(_gnd_net_));
    defparam shift_srl_69_5_LC_26_9_5.C_ON=1'b0;
    defparam shift_srl_69_5_LC_26_9_5.SEQ_MODE=4'b1000;
    defparam shift_srl_69_5_LC_26_9_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_69_5_LC_26_9_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83125),
            .lcout(shift_srl_69Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93397),
            .ce(N__85421),
            .sr(_gnd_net_));
    defparam shift_srl_69_6_LC_26_9_6.C_ON=1'b0;
    defparam shift_srl_69_6_LC_26_9_6.SEQ_MODE=4'b1000;
    defparam shift_srl_69_6_LC_26_9_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_69_6_LC_26_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83119),
            .lcout(shift_srl_69Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93397),
            .ce(N__85421),
            .sr(_gnd_net_));
    defparam shift_srl_67_10_LC_26_10_0.C_ON=1'b0;
    defparam shift_srl_67_10_LC_26_10_0.SEQ_MODE=4'b1000;
    defparam shift_srl_67_10_LC_26_10_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_67_10_LC_26_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83113),
            .lcout(shift_srl_67Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93389),
            .ce(N__86934),
            .sr(_gnd_net_));
    defparam shift_srl_67_9_LC_26_10_1.C_ON=1'b0;
    defparam shift_srl_67_9_LC_26_10_1.SEQ_MODE=4'b1000;
    defparam shift_srl_67_9_LC_26_10_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_67_9_LC_26_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83107),
            .lcout(shift_srl_67Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93389),
            .ce(N__86934),
            .sr(_gnd_net_));
    defparam shift_srl_67_8_LC_26_10_2.C_ON=1'b0;
    defparam shift_srl_67_8_LC_26_10_2.SEQ_MODE=4'b1000;
    defparam shift_srl_67_8_LC_26_10_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_67_8_LC_26_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83101),
            .lcout(shift_srl_67Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93389),
            .ce(N__86934),
            .sr(_gnd_net_));
    defparam shift_srl_67_7_LC_26_10_3.C_ON=1'b0;
    defparam shift_srl_67_7_LC_26_10_3.SEQ_MODE=4'b1000;
    defparam shift_srl_67_7_LC_26_10_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_67_7_LC_26_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83095),
            .lcout(shift_srl_67Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93389),
            .ce(N__86934),
            .sr(_gnd_net_));
    defparam shift_srl_67_6_LC_26_10_4.C_ON=1'b0;
    defparam shift_srl_67_6_LC_26_10_4.SEQ_MODE=4'b1000;
    defparam shift_srl_67_6_LC_26_10_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_67_6_LC_26_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83089),
            .lcout(shift_srl_67Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93389),
            .ce(N__86934),
            .sr(_gnd_net_));
    defparam shift_srl_67_5_LC_26_10_5.C_ON=1'b0;
    defparam shift_srl_67_5_LC_26_10_5.SEQ_MODE=4'b1000;
    defparam shift_srl_67_5_LC_26_10_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_67_5_LC_26_10_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83137),
            .lcout(shift_srl_67Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93389),
            .ce(N__86934),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_67_LC_26_11_0.C_ON=1'b0;
    defparam rco_obuf_RNO_67_LC_26_11_0.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_67_LC_26_11_0.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_67_LC_26_11_0 (
            .in0(N__86861),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__90694),
            .lcout(rco_c_67),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_68_LC_26_11_1.C_ON=1'b0;
    defparam rco_obuf_RNO_68_LC_26_11_1.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_68_LC_26_11_1.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_68_LC_26_11_1 (
            .in0(N__90695),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84832),
            .lcout(rco_c_68),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_69_LC_26_11_2.C_ON=1'b0;
    defparam rco_obuf_RNO_69_LC_26_11_2.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_69_LC_26_11_2.LUT_INIT=16'b1100110000000000;
    LogicCell40 rco_obuf_RNO_69_LC_26_11_2 (
            .in0(_gnd_net_),
            .in1(N__83191),
            .in2(_gnd_net_),
            .in3(N__90696),
            .lcout(rco_c_69),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_67_0_LC_26_11_3.C_ON=1'b0;
    defparam shift_srl_67_0_LC_26_11_3.SEQ_MODE=4'b1000;
    defparam shift_srl_67_0_LC_26_11_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_67_0_LC_26_11_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86860),
            .lcout(shift_srl_67Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93373),
            .ce(N__86927),
            .sr(_gnd_net_));
    defparam shift_srl_67_1_LC_26_11_4.C_ON=1'b0;
    defparam shift_srl_67_1_LC_26_11_4.SEQ_MODE=4'b1000;
    defparam shift_srl_67_1_LC_26_11_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_67_1_LC_26_11_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83161),
            .lcout(shift_srl_67Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93373),
            .ce(N__86927),
            .sr(_gnd_net_));
    defparam shift_srl_67_2_LC_26_11_5.C_ON=1'b0;
    defparam shift_srl_67_2_LC_26_11_5.SEQ_MODE=4'b1000;
    defparam shift_srl_67_2_LC_26_11_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_67_2_LC_26_11_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83155),
            .lcout(shift_srl_67Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93373),
            .ce(N__86927),
            .sr(_gnd_net_));
    defparam shift_srl_67_3_LC_26_11_6.C_ON=1'b0;
    defparam shift_srl_67_3_LC_26_11_6.SEQ_MODE=4'b1000;
    defparam shift_srl_67_3_LC_26_11_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_67_3_LC_26_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83149),
            .lcout(shift_srl_67Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93373),
            .ce(N__86927),
            .sr(_gnd_net_));
    defparam shift_srl_67_4_LC_26_11_7.C_ON=1'b0;
    defparam shift_srl_67_4_LC_26_11_7.SEQ_MODE=4'b1000;
    defparam shift_srl_67_4_LC_26_11_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_67_4_LC_26_11_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83143),
            .lcout(shift_srl_67Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93373),
            .ce(N__86927),
            .sr(_gnd_net_));
    defparam shift_srl_71_4_LC_26_12_0.C_ON=1'b0;
    defparam shift_srl_71_4_LC_26_12_0.SEQ_MODE=4'b1000;
    defparam shift_srl_71_4_LC_26_12_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_71_4_LC_26_12_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83224),
            .lcout(shift_srl_71Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93357),
            .ce(N__85300),
            .sr(_gnd_net_));
    defparam shift_srl_71_10_LC_26_12_1.C_ON=1'b0;
    defparam shift_srl_71_10_LC_26_12_1.SEQ_MODE=4'b1000;
    defparam shift_srl_71_10_LC_26_12_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_71_10_LC_26_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83218),
            .lcout(shift_srl_71Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93357),
            .ce(N__85300),
            .sr(_gnd_net_));
    defparam shift_srl_71_11_LC_26_12_2.C_ON=1'b0;
    defparam shift_srl_71_11_LC_26_12_2.SEQ_MODE=4'b1000;
    defparam shift_srl_71_11_LC_26_12_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_71_11_LC_26_12_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83131),
            .lcout(shift_srl_71Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93357),
            .ce(N__85300),
            .sr(_gnd_net_));
    defparam shift_srl_71_3_LC_26_12_3.C_ON=1'b0;
    defparam shift_srl_71_3_LC_26_12_3.SEQ_MODE=4'b1000;
    defparam shift_srl_71_3_LC_26_12_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_71_3_LC_26_12_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83200),
            .lcout(shift_srl_71Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93357),
            .ce(N__85300),
            .sr(_gnd_net_));
    defparam shift_srl_71_9_LC_26_12_4.C_ON=1'b0;
    defparam shift_srl_71_9_LC_26_12_4.SEQ_MODE=4'b1000;
    defparam shift_srl_71_9_LC_26_12_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_71_9_LC_26_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85306),
            .lcout(shift_srl_71Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93357),
            .ce(N__85300),
            .sr(_gnd_net_));
    defparam shift_srl_71_1_LC_26_12_5.C_ON=1'b0;
    defparam shift_srl_71_1_LC_26_12_5.SEQ_MODE=4'b1000;
    defparam shift_srl_71_1_LC_26_12_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_71_1_LC_26_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83212),
            .lcout(shift_srl_71Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93357),
            .ce(N__85300),
            .sr(_gnd_net_));
    defparam shift_srl_71_0_LC_26_12_6.C_ON=1'b0;
    defparam shift_srl_71_0_LC_26_12_6.SEQ_MODE=4'b1000;
    defparam shift_srl_71_0_LC_26_12_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_71_0_LC_26_12_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86718),
            .lcout(shift_srl_71Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93357),
            .ce(N__85300),
            .sr(_gnd_net_));
    defparam shift_srl_71_2_LC_26_12_7.C_ON=1'b0;
    defparam shift_srl_71_2_LC_26_12_7.SEQ_MODE=4'b1000;
    defparam shift_srl_71_2_LC_26_12_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_71_2_LC_26_12_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83206),
            .lcout(shift_srl_71Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93357),
            .ce(N__85300),
            .sr(_gnd_net_));
    defparam shift_srl_68_RNIHDC4_15_LC_26_13_0.C_ON=1'b0;
    defparam shift_srl_68_RNIHDC4_15_LC_26_13_0.SEQ_MODE=4'b0000;
    defparam shift_srl_68_RNIHDC4_15_LC_26_13_0.LUT_INIT=16'b1100110000000000;
    LogicCell40 shift_srl_68_RNIHDC4_15_LC_26_13_0 (
            .in0(_gnd_net_),
            .in1(N__86896),
            .in2(_gnd_net_),
            .in3(N__86856),
            .lcout(shift_srl_68_RNIHDC4Z0Z_15),
            .ltout(shift_srl_68_RNIHDC4Z0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_69_RNIBQRC_15_LC_26_13_1.C_ON=1'b0;
    defparam shift_srl_69_RNIBQRC_15_LC_26_13_1.SEQ_MODE=4'b0000;
    defparam shift_srl_69_RNIBQRC_15_LC_26_13_1.LUT_INIT=16'b1111000000000000;
    LogicCell40 shift_srl_69_RNIBQRC_15_LC_26_13_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__83194),
            .in3(N__86664),
            .lcout(shift_srl_69_RNIBQRCZ0Z_15),
            .ltout(shift_srl_69_RNIBQRCZ0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNITRGNH_15_LC_26_13_2.C_ON=1'b0;
    defparam shift_srl_0_RNITRGNH_15_LC_26_13_2.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNITRGNH_15_LC_26_13_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNITRGNH_15_LC_26_13_2 (
            .in0(N__84895),
            .in1(N__90321),
            .in2(N__83182),
            .in3(N__85008),
            .lcout(clk_en_70),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_67_15_LC_26_13_3.C_ON=1'b0;
    defparam shift_srl_67_15_LC_26_13_3.SEQ_MODE=4'b1000;
    defparam shift_srl_67_15_LC_26_13_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_67_15_LC_26_13_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83281),
            .lcout(shift_srl_67Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93335),
            .ce(N__86938),
            .sr(_gnd_net_));
    defparam shift_srl_67_14_LC_26_13_4.C_ON=1'b0;
    defparam shift_srl_67_14_LC_26_13_4.SEQ_MODE=4'b1000;
    defparam shift_srl_67_14_LC_26_13_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_67_14_LC_26_13_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83275),
            .lcout(shift_srl_67Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93335),
            .ce(N__86938),
            .sr(_gnd_net_));
    defparam shift_srl_67_13_LC_26_13_5.C_ON=1'b0;
    defparam shift_srl_67_13_LC_26_13_5.SEQ_MODE=4'b1000;
    defparam shift_srl_67_13_LC_26_13_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_67_13_LC_26_13_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83269),
            .lcout(shift_srl_67Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93335),
            .ce(N__86938),
            .sr(_gnd_net_));
    defparam shift_srl_67_12_LC_26_13_6.C_ON=1'b0;
    defparam shift_srl_67_12_LC_26_13_6.SEQ_MODE=4'b1000;
    defparam shift_srl_67_12_LC_26_13_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_67_12_LC_26_13_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83254),
            .lcout(shift_srl_67Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93335),
            .ce(N__86938),
            .sr(_gnd_net_));
    defparam shift_srl_67_11_LC_26_13_7.C_ON=1'b0;
    defparam shift_srl_67_11_LC_26_13_7.SEQ_MODE=4'b1000;
    defparam shift_srl_67_11_LC_26_13_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_67_11_LC_26_13_7 (
            .in0(N__83263),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_67Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93335),
            .ce(N__86938),
            .sr(_gnd_net_));
    defparam shift_srl_70_4_LC_26_14_0.C_ON=1'b0;
    defparam shift_srl_70_4_LC_26_14_0.SEQ_MODE=4'b1000;
    defparam shift_srl_70_4_LC_26_14_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_70_4_LC_26_14_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83236),
            .lcout(shift_srl_70Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93315),
            .ce(N__85509),
            .sr(_gnd_net_));
    defparam shift_srl_70_1_LC_26_14_1.C_ON=1'b0;
    defparam shift_srl_70_1_LC_26_14_1.SEQ_MODE=4'b1000;
    defparam shift_srl_70_1_LC_26_14_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_70_1_LC_26_14_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85516),
            .lcout(shift_srl_70Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93315),
            .ce(N__85509),
            .sr(_gnd_net_));
    defparam shift_srl_70_2_LC_26_14_2.C_ON=1'b0;
    defparam shift_srl_70_2_LC_26_14_2.SEQ_MODE=4'b1000;
    defparam shift_srl_70_2_LC_26_14_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_70_2_LC_26_14_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83248),
            .lcout(shift_srl_70Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93315),
            .ce(N__85509),
            .sr(_gnd_net_));
    defparam shift_srl_70_3_LC_26_14_3.C_ON=1'b0;
    defparam shift_srl_70_3_LC_26_14_3.SEQ_MODE=4'b1000;
    defparam shift_srl_70_3_LC_26_14_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_70_3_LC_26_14_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83242),
            .lcout(shift_srl_70Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93315),
            .ce(N__85509),
            .sr(_gnd_net_));
    defparam shift_srl_70_5_LC_26_14_4.C_ON=1'b0;
    defparam shift_srl_70_5_LC_26_14_4.SEQ_MODE=4'b1000;
    defparam shift_srl_70_5_LC_26_14_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_70_5_LC_26_14_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83230),
            .lcout(shift_srl_70Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93315),
            .ce(N__85509),
            .sr(_gnd_net_));
    defparam shift_srl_70_8_LC_26_14_5.C_ON=1'b0;
    defparam shift_srl_70_8_LC_26_14_5.SEQ_MODE=4'b1000;
    defparam shift_srl_70_8_LC_26_14_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_70_8_LC_26_14_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83356),
            .lcout(shift_srl_70Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93315),
            .ce(N__85509),
            .sr(_gnd_net_));
    defparam shift_srl_70_6_LC_26_14_6.C_ON=1'b0;
    defparam shift_srl_70_6_LC_26_14_6.SEQ_MODE=4'b1000;
    defparam shift_srl_70_6_LC_26_14_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_70_6_LC_26_14_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83368),
            .lcout(shift_srl_70Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93315),
            .ce(N__85509),
            .sr(_gnd_net_));
    defparam shift_srl_70_7_LC_26_14_7.C_ON=1'b0;
    defparam shift_srl_70_7_LC_26_14_7.SEQ_MODE=4'b1000;
    defparam shift_srl_70_7_LC_26_14_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_70_7_LC_26_14_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83362),
            .lcout(shift_srl_70Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93315),
            .ce(N__85509),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIRS4Q8_15_LC_26_15_0.C_ON=1'b0;
    defparam shift_srl_0_RNIRS4Q8_15_LC_26_15_0.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIRS4Q8_15_LC_26_15_0.LUT_INIT=16'b1100110000000000;
    LogicCell40 shift_srl_0_RNIRS4Q8_15_LC_26_15_0 (
            .in0(_gnd_net_),
            .in1(N__90318),
            .in2(_gnd_net_),
            .in3(N__83609),
            .lcout(clk_en_34),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_34_0_LC_26_15_1.C_ON=1'b0;
    defparam shift_srl_34_0_LC_26_15_1.SEQ_MODE=4'b1000;
    defparam shift_srl_34_0_LC_26_15_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_34_0_LC_26_15_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83339),
            .lcout(shift_srl_34Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93296),
            .ce(N__87120),
            .sr(_gnd_net_));
    defparam shift_srl_34_1_LC_26_15_2.C_ON=1'b0;
    defparam shift_srl_34_1_LC_26_15_2.SEQ_MODE=4'b1000;
    defparam shift_srl_34_1_LC_26_15_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_34_1_LC_26_15_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83305),
            .lcout(shift_srl_34Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93296),
            .ce(N__87120),
            .sr(_gnd_net_));
    defparam shift_srl_34_2_LC_26_15_3.C_ON=1'b0;
    defparam shift_srl_34_2_LC_26_15_3.SEQ_MODE=4'b1000;
    defparam shift_srl_34_2_LC_26_15_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_34_2_LC_26_15_3 (
            .in0(N__83299),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_34Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93296),
            .ce(N__87120),
            .sr(_gnd_net_));
    defparam shift_srl_34_3_LC_26_15_4.C_ON=1'b0;
    defparam shift_srl_34_3_LC_26_15_4.SEQ_MODE=4'b1000;
    defparam shift_srl_34_3_LC_26_15_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_34_3_LC_26_15_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83293),
            .lcout(shift_srl_34Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93296),
            .ce(N__87120),
            .sr(_gnd_net_));
    defparam shift_srl_34_4_LC_26_15_5.C_ON=1'b0;
    defparam shift_srl_34_4_LC_26_15_5.SEQ_MODE=4'b1000;
    defparam shift_srl_34_4_LC_26_15_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_34_4_LC_26_15_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83287),
            .lcout(shift_srl_34Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93296),
            .ce(N__87120),
            .sr(_gnd_net_));
    defparam shift_srl_37_15_LC_26_16_0.C_ON=1'b0;
    defparam shift_srl_37_15_LC_26_16_0.SEQ_MODE=4'b1000;
    defparam shift_srl_37_15_LC_26_16_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_37_15_LC_26_16_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83452),
            .lcout(shift_srl_37Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93282),
            .ce(N__91856),
            .sr(_gnd_net_));
    defparam shift_srl_37_14_LC_26_16_6.C_ON=1'b0;
    defparam shift_srl_37_14_LC_26_16_6.SEQ_MODE=4'b1000;
    defparam shift_srl_37_14_LC_26_16_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_37_14_LC_26_16_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85480),
            .lcout(shift_srl_37Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93282),
            .ce(N__91856),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIK5EK9_15_LC_26_17_0.C_ON=1'b0;
    defparam shift_srl_0_RNIK5EK9_15_LC_26_17_0.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIK5EK9_15_LC_26_17_0.LUT_INIT=16'b1100110000000000;
    LogicCell40 shift_srl_0_RNIK5EK9_15_LC_26_17_0 (
            .in0(_gnd_net_),
            .in1(N__90320),
            .in2(_gnd_net_),
            .in3(N__83526),
            .lcout(clk_en_37),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_37_0_LC_26_17_1.C_ON=1'b0;
    defparam shift_srl_37_0_LC_26_17_1.SEQ_MODE=4'b1000;
    defparam shift_srl_37_0_LC_26_17_1.LUT_INIT=16'b1100110011001100;
    LogicCell40 shift_srl_37_0_LC_26_17_1 (
            .in0(_gnd_net_),
            .in1(N__83433),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_37Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93241),
            .ce(N__91855),
            .sr(_gnd_net_));
    defparam shift_srl_37_1_LC_26_17_2.C_ON=1'b0;
    defparam shift_srl_37_1_LC_26_17_2.SEQ_MODE=4'b1000;
    defparam shift_srl_37_1_LC_26_17_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_37_1_LC_26_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83419),
            .lcout(shift_srl_37Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93241),
            .ce(N__91855),
            .sr(_gnd_net_));
    defparam shift_srl_37_2_LC_26_17_3.C_ON=1'b0;
    defparam shift_srl_37_2_LC_26_17_3.SEQ_MODE=4'b1000;
    defparam shift_srl_37_2_LC_26_17_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_37_2_LC_26_17_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83413),
            .lcout(shift_srl_37Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93241),
            .ce(N__91855),
            .sr(_gnd_net_));
    defparam shift_srl_37_3_LC_26_17_4.C_ON=1'b0;
    defparam shift_srl_37_3_LC_26_17_4.SEQ_MODE=4'b1000;
    defparam shift_srl_37_3_LC_26_17_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_37_3_LC_26_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83407),
            .lcout(shift_srl_37Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93241),
            .ce(N__91855),
            .sr(_gnd_net_));
    defparam shift_srl_37_4_LC_26_17_5.C_ON=1'b0;
    defparam shift_srl_37_4_LC_26_17_5.SEQ_MODE=4'b1000;
    defparam shift_srl_37_4_LC_26_17_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_37_4_LC_26_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83401),
            .lcout(shift_srl_37Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93241),
            .ce(N__91855),
            .sr(_gnd_net_));
    defparam shift_srl_37_5_LC_26_17_6.C_ON=1'b0;
    defparam shift_srl_37_5_LC_26_17_6.SEQ_MODE=4'b1000;
    defparam shift_srl_37_5_LC_26_17_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_37_5_LC_26_17_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83395),
            .lcout(shift_srl_37Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93241),
            .ce(N__91855),
            .sr(_gnd_net_));
    defparam shift_srl_32_RNIFBUO8_15_LC_26_18_0.C_ON=1'b0;
    defparam shift_srl_32_RNIFBUO8_15_LC_26_18_0.SEQ_MODE=4'b0000;
    defparam shift_srl_32_RNIFBUO8_15_LC_26_18_0.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_32_RNIFBUO8_15_LC_26_18_0 (
            .in0(N__85229),
            .in1(N__83583),
            .in2(_gnd_net_),
            .in3(N__87319),
            .lcout(rco_c_32),
            .ltout(rco_c_32_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIANOP8_15_LC_26_18_1.C_ON=1'b0;
    defparam shift_srl_0_RNIANOP8_15_LC_26_18_1.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIANOP8_15_LC_26_18_1.LUT_INIT=16'b1111000000000000;
    LogicCell40 shift_srl_0_RNIANOP8_15_LC_26_18_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__83896),
            .in3(N__90319),
            .lcout(clk_en_33),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_29_RNISHF41_15_LC_26_18_2.C_ON=1'b0;
    defparam shift_srl_29_RNISHF41_15_LC_26_18_2.SEQ_MODE=4'b0000;
    defparam shift_srl_29_RNISHF41_15_LC_26_18_2.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_29_RNISHF41_15_LC_26_18_2 (
            .in0(N__83893),
            .in1(N__83848),
            .in2(_gnd_net_),
            .in3(N__83793),
            .lcout(),
            .ltout(shift_srl_29_RNISHF41Z0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_31_RNIIE682_15_LC_26_18_3.C_ON=1'b0;
    defparam shift_srl_31_RNIIE682_15_LC_26_18_3.SEQ_MODE=4'b0000;
    defparam shift_srl_31_RNIIE682_15_LC_26_18_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_31_RNIIE682_15_LC_26_18_3 (
            .in0(N__83718),
            .in1(N__83680),
            .in2(N__83665),
            .in3(N__83657),
            .lcout(rco_int_0_a2_0_a2_out_4),
            .ltout(rco_int_0_a2_0_a2_out_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_33_RNI0HAP8_15_LC_26_18_4.C_ON=1'b0;
    defparam shift_srl_33_RNI0HAP8_15_LC_26_18_4.SEQ_MODE=4'b0000;
    defparam shift_srl_33_RNI0HAP8_15_LC_26_18_4.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_33_RNI0HAP8_15_LC_26_18_4 (
            .in0(N__85225),
            .in1(N__85555),
            .in2(N__83629),
            .in3(N__87318),
            .lcout(rco_c_33),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_31_RNIV9OC8_15_LC_26_18_5.C_ON=1'b0;
    defparam shift_srl_31_RNIV9OC8_15_LC_26_18_5.SEQ_MODE=4'b0000;
    defparam shift_srl_31_RNIV9OC8_15_LC_26_18_5.LUT_INIT=16'b1100110000000000;
    LogicCell40 shift_srl_31_RNIV9OC8_15_LC_26_18_5 (
            .in0(_gnd_net_),
            .in1(N__83578),
            .in2(_gnd_net_),
            .in3(N__85227),
            .lcout(rco_c_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_35_RNI58L69_15_LC_26_18_6.C_ON=1'b0;
    defparam shift_srl_35_RNI58L69_15_LC_26_18_6.SEQ_MODE=4'b0000;
    defparam shift_srl_35_RNI58L69_15_LC_26_18_6.LUT_INIT=16'b1010000000000000;
    LogicCell40 shift_srl_35_RNI58L69_15_LC_26_18_6 (
            .in0(N__85226),
            .in1(_gnd_net_),
            .in2(N__83584),
            .in3(N__83559),
            .lcout(rco_c_35),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_36_RNIPPJJ9_15_LC_26_18_7.C_ON=1'b0;
    defparam shift_srl_36_RNIPPJJ9_15_LC_26_18_7.SEQ_MODE=4'b0000;
    defparam shift_srl_36_RNIPPJJ9_15_LC_26_18_7.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_36_RNIPPJJ9_15_LC_26_18_7 (
            .in0(N__83582),
            .in1(N__83484),
            .in2(N__83563),
            .in3(N__85228),
            .lcout(rco_c_36),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNI0KF79_15_LC_26_19_0.C_ON=1'b0;
    defparam shift_srl_0_RNI0KF79_15_LC_26_19_0.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNI0KF79_15_LC_26_19_0.LUT_INIT=16'b1100110000000000;
    LogicCell40 shift_srl_0_RNI0KF79_15_LC_26_19_0 (
            .in0(_gnd_net_),
            .in1(N__90309),
            .in2(_gnd_net_),
            .in3(N__83499),
            .lcout(clk_en_36),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_36_0_LC_26_19_1.C_ON=1'b0;
    defparam shift_srl_36_0_LC_26_19_1.SEQ_MODE=4'b1000;
    defparam shift_srl_36_0_LC_26_19_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_36_0_LC_26_19_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83488),
            .lcout(shift_srl_36Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93297),
            .ce(N__90918),
            .sr(_gnd_net_));
    defparam shift_srl_36_1_LC_26_19_2.C_ON=1'b0;
    defparam shift_srl_36_1_LC_26_19_2.SEQ_MODE=4'b1000;
    defparam shift_srl_36_1_LC_26_19_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_36_1_LC_26_19_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84088),
            .lcout(shift_srl_36Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93297),
            .ce(N__90918),
            .sr(_gnd_net_));
    defparam shift_srl_36_2_LC_26_19_3.C_ON=1'b0;
    defparam shift_srl_36_2_LC_26_19_3.SEQ_MODE=4'b1000;
    defparam shift_srl_36_2_LC_26_19_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_36_2_LC_26_19_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84082),
            .lcout(shift_srl_36Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93297),
            .ce(N__90918),
            .sr(_gnd_net_));
    defparam shift_srl_36_3_LC_26_19_4.C_ON=1'b0;
    defparam shift_srl_36_3_LC_26_19_4.SEQ_MODE=4'b1000;
    defparam shift_srl_36_3_LC_26_19_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_36_3_LC_26_19_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84076),
            .lcout(shift_srl_36Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93297),
            .ce(N__90918),
            .sr(_gnd_net_));
    defparam shift_srl_36_4_LC_26_19_5.C_ON=1'b0;
    defparam shift_srl_36_4_LC_26_19_5.SEQ_MODE=4'b1000;
    defparam shift_srl_36_4_LC_26_19_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_36_4_LC_26_19_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84070),
            .lcout(shift_srl_36Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93297),
            .ce(N__90918),
            .sr(_gnd_net_));
    defparam shift_srl_36_5_LC_26_19_6.C_ON=1'b0;
    defparam shift_srl_36_5_LC_26_19_6.SEQ_MODE=4'b1000;
    defparam shift_srl_36_5_LC_26_19_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_36_5_LC_26_19_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84064),
            .lcout(shift_srl_36Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93297),
            .ce(N__90918),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_169_LC_26_20_0.C_ON=1'b0;
    defparam rco_obuf_RNO_169_LC_26_20_0.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_169_LC_26_20_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 rco_obuf_RNO_169_LC_26_20_0 (
            .in0(N__89182),
            .in1(N__87415),
            .in2(N__87712),
            .in3(N__84274),
            .lcout(rco_c_169),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_168_LC_26_20_1.C_ON=1'b0;
    defparam rco_obuf_RNO_168_LC_26_20_1.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_168_LC_26_20_1.LUT_INIT=16'b1000100000000000;
    LogicCell40 rco_obuf_RNO_168_LC_26_20_1 (
            .in0(N__87414),
            .in1(N__89181),
            .in2(_gnd_net_),
            .in3(N__87691),
            .lcout(rco_c_168),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_164_15_LC_26_20_2.C_ON=1'b0;
    defparam shift_srl_164_15_LC_26_20_2.SEQ_MODE=4'b1000;
    defparam shift_srl_164_15_LC_26_20_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_164_15_LC_26_20_2 (
            .in0(N__85738),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_164Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93316),
            .ce(N__87796),
            .sr(_gnd_net_));
    defparam shift_srl_167_RNIUC2T_15_LC_26_20_3.C_ON=1'b0;
    defparam shift_srl_167_RNIUC2T_15_LC_26_20_3.SEQ_MODE=4'b0000;
    defparam shift_srl_167_RNIUC2T_15_LC_26_20_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_167_RNIUC2T_15_LC_26_20_3 (
            .in0(N__84012),
            .in1(N__83964),
            .in2(N__83914),
            .in3(N__87242),
            .lcout(),
            .ltout(shift_srl_167_RNIUC2TZ0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_163_RNI3MR51_15_LC_26_20_4.C_ON=1'b0;
    defparam shift_srl_163_RNI3MR51_15_LC_26_20_4.SEQ_MODE=4'b0000;
    defparam shift_srl_163_RNI3MR51_15_LC_26_20_4.LUT_INIT=16'b1111000010101010;
    LogicCell40 shift_srl_163_RNI3MR51_15_LC_26_20_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__84298),
            .in3(N__87742),
            .lcout(shift_srl_163_RNI3MR51Z0Z_15),
            .ltout(shift_srl_163_RNI3MR51Z0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_170_RNIRM2S1_15_LC_26_20_5.C_ON=1'b0;
    defparam shift_srl_170_RNIRM2S1_15_LC_26_20_5.SEQ_MODE=4'b0000;
    defparam shift_srl_170_RNIRM2S1_15_LC_26_20_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_170_RNIRM2S1_15_LC_26_20_5 (
            .in0(N__84295),
            .in1(N__84273),
            .in2(N__84250),
            .in3(N__89180),
            .lcout(shift_srl_170_RNIRM2S1Z0Z_15),
            .ltout(shift_srl_170_RNIRM2S1Z0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_172_RNI47NL2_15_LC_26_20_6.C_ON=1'b0;
    defparam shift_srl_172_RNI47NL2_15_LC_26_20_6.SEQ_MODE=4'b0000;
    defparam shift_srl_172_RNI47NL2_15_LC_26_20_6.LUT_INIT=16'b1100000000000000;
    LogicCell40 shift_srl_172_RNI47NL2_15_LC_26_20_6 (
            .in0(_gnd_net_),
            .in1(N__88945),
            .in2(N__84247),
            .in3(N__87495),
            .lcout(rco_int_0_a3_0_a2_0_172),
            .ltout(rco_int_0_a3_0_a2_0_172_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIL3KM4_15_LC_26_20_7.C_ON=1'b0;
    defparam shift_srl_0_RNIL3KM4_15_LC_26_20_7.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIL3KM4_15_LC_26_20_7.LUT_INIT=16'b0101111111111111;
    LogicCell40 shift_srl_0_RNIL3KM4_15_LC_26_20_7 (
            .in0(N__90308),
            .in1(_gnd_net_),
            .in2(N__84163),
            .in3(N__87984),
            .lcout(clk_en_0_a3_0_a2cf1_1_176),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_163_10_LC_26_21_0.C_ON=1'b0;
    defparam shift_srl_163_10_LC_26_21_0.SEQ_MODE=4'b1000;
    defparam shift_srl_163_10_LC_26_21_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_163_10_LC_26_21_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84340),
            .lcout(shift_srl_163Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93336),
            .ce(N__85803),
            .sr(_gnd_net_));
    defparam shift_srl_163_11_LC_26_21_1.C_ON=1'b0;
    defparam shift_srl_163_11_LC_26_21_1.SEQ_MODE=4'b1000;
    defparam shift_srl_163_11_LC_26_21_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_163_11_LC_26_21_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84112),
            .lcout(shift_srl_163Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93336),
            .ce(N__85803),
            .sr(_gnd_net_));
    defparam shift_srl_163_12_LC_26_21_2.C_ON=1'b0;
    defparam shift_srl_163_12_LC_26_21_2.SEQ_MODE=4'b1000;
    defparam shift_srl_163_12_LC_26_21_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_163_12_LC_26_21_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84106),
            .lcout(shift_srl_163Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93336),
            .ce(N__85803),
            .sr(_gnd_net_));
    defparam shift_srl_163_13_LC_26_21_3.C_ON=1'b0;
    defparam shift_srl_163_13_LC_26_21_3.SEQ_MODE=4'b1000;
    defparam shift_srl_163_13_LC_26_21_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_163_13_LC_26_21_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84100),
            .lcout(shift_srl_163Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93336),
            .ce(N__85803),
            .sr(_gnd_net_));
    defparam shift_srl_163_14_LC_26_21_4.C_ON=1'b0;
    defparam shift_srl_163_14_LC_26_21_4.SEQ_MODE=4'b1000;
    defparam shift_srl_163_14_LC_26_21_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_163_14_LC_26_21_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84094),
            .lcout(shift_srl_163Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93336),
            .ce(N__85803),
            .sr(_gnd_net_));
    defparam shift_srl_163_15_LC_26_21_5.C_ON=1'b0;
    defparam shift_srl_163_15_LC_26_21_5.SEQ_MODE=4'b1000;
    defparam shift_srl_163_15_LC_26_21_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_163_15_LC_26_21_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84346),
            .lcout(shift_srl_163Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93336),
            .ce(N__85803),
            .sr(_gnd_net_));
    defparam shift_srl_163_9_LC_26_21_6.C_ON=1'b0;
    defparam shift_srl_163_9_LC_26_21_6.SEQ_MODE=4'b1000;
    defparam shift_srl_163_9_LC_26_21_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_163_9_LC_26_21_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84334),
            .lcout(shift_srl_163Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93336),
            .ce(N__85803),
            .sr(_gnd_net_));
    defparam shift_srl_163_8_LC_26_21_7.C_ON=1'b0;
    defparam shift_srl_163_8_LC_26_21_7.SEQ_MODE=4'b1000;
    defparam shift_srl_163_8_LC_26_21_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_163_8_LC_26_21_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85813),
            .lcout(shift_srl_163Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93336),
            .ce(N__85803),
            .sr(_gnd_net_));
    defparam shift_srl_36_10_LC_26_22_0.C_ON=1'b0;
    defparam shift_srl_36_10_LC_26_22_0.SEQ_MODE=4'b1000;
    defparam shift_srl_36_10_LC_26_22_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_36_10_LC_26_22_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84310),
            .lcout(shift_srl_36Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93358),
            .ce(N__90919),
            .sr(_gnd_net_));
    defparam shift_srl_36_11_LC_26_22_1.C_ON=1'b0;
    defparam shift_srl_36_11_LC_26_22_1.SEQ_MODE=4'b1000;
    defparam shift_srl_36_11_LC_26_22_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_36_11_LC_26_22_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84328),
            .lcout(shift_srl_36Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93358),
            .ce(N__90919),
            .sr(_gnd_net_));
    defparam shift_srl_36_12_LC_26_22_2.C_ON=1'b0;
    defparam shift_srl_36_12_LC_26_22_2.SEQ_MODE=4'b1000;
    defparam shift_srl_36_12_LC_26_22_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_36_12_LC_26_22_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84322),
            .lcout(shift_srl_36Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93358),
            .ce(N__90919),
            .sr(_gnd_net_));
    defparam shift_srl_36_13_LC_26_22_3.C_ON=1'b0;
    defparam shift_srl_36_13_LC_26_22_3.SEQ_MODE=4'b1000;
    defparam shift_srl_36_13_LC_26_22_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_36_13_LC_26_22_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84316),
            .lcout(shift_srl_36Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93358),
            .ce(N__90919),
            .sr(_gnd_net_));
    defparam shift_srl_36_9_LC_26_22_5.C_ON=1'b0;
    defparam shift_srl_36_9_LC_26_22_5.SEQ_MODE=4'b1000;
    defparam shift_srl_36_9_LC_26_22_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_36_9_LC_26_22_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84304),
            .lcout(shift_srl_36Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93358),
            .ce(N__90919),
            .sr(_gnd_net_));
    defparam shift_srl_36_8_LC_26_22_6.C_ON=1'b0;
    defparam shift_srl_36_8_LC_26_22_6.SEQ_MODE=4'b1000;
    defparam shift_srl_36_8_LC_26_22_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_36_8_LC_26_22_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84394),
            .lcout(shift_srl_36Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93358),
            .ce(N__90919),
            .sr(_gnd_net_));
    defparam shift_srl_36_7_LC_26_22_7.C_ON=1'b0;
    defparam shift_srl_36_7_LC_26_22_7.SEQ_MODE=4'b1000;
    defparam shift_srl_36_7_LC_26_22_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_36_7_LC_26_22_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84454),
            .lcout(shift_srl_36Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93358),
            .ce(N__90919),
            .sr(_gnd_net_));
    defparam shift_srl_191_10_LC_26_23_0.C_ON=1'b0;
    defparam shift_srl_191_10_LC_26_23_0.SEQ_MODE=4'b1000;
    defparam shift_srl_191_10_LC_26_23_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_191_10_LC_26_23_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84358),
            .lcout(shift_srl_191Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93374),
            .ce(N__86061),
            .sr(_gnd_net_));
    defparam shift_srl_191_11_LC_26_23_1.C_ON=1'b0;
    defparam shift_srl_191_11_LC_26_23_1.SEQ_MODE=4'b1000;
    defparam shift_srl_191_11_LC_26_23_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_191_11_LC_26_23_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84388),
            .lcout(shift_srl_191Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93374),
            .ce(N__86061),
            .sr(_gnd_net_));
    defparam shift_srl_191_12_LC_26_23_2.C_ON=1'b0;
    defparam shift_srl_191_12_LC_26_23_2.SEQ_MODE=4'b1000;
    defparam shift_srl_191_12_LC_26_23_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_191_12_LC_26_23_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84382),
            .lcout(shift_srl_191Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93374),
            .ce(N__86061),
            .sr(_gnd_net_));
    defparam shift_srl_191_13_LC_26_23_3.C_ON=1'b0;
    defparam shift_srl_191_13_LC_26_23_3.SEQ_MODE=4'b1000;
    defparam shift_srl_191_13_LC_26_23_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_191_13_LC_26_23_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84376),
            .lcout(shift_srl_191Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93374),
            .ce(N__86061),
            .sr(_gnd_net_));
    defparam shift_srl_191_14_LC_26_23_4.C_ON=1'b0;
    defparam shift_srl_191_14_LC_26_23_4.SEQ_MODE=4'b1000;
    defparam shift_srl_191_14_LC_26_23_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_191_14_LC_26_23_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84370),
            .lcout(shift_srl_191Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93374),
            .ce(N__86061),
            .sr(_gnd_net_));
    defparam shift_srl_191_15_LC_26_23_5.C_ON=1'b0;
    defparam shift_srl_191_15_LC_26_23_5.SEQ_MODE=4'b1000;
    defparam shift_srl_191_15_LC_26_23_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_191_15_LC_26_23_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84364),
            .lcout(shift_srl_191Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93374),
            .ce(N__86061),
            .sr(_gnd_net_));
    defparam shift_srl_191_9_LC_26_23_6.C_ON=1'b0;
    defparam shift_srl_191_9_LC_26_23_6.SEQ_MODE=4'b1000;
    defparam shift_srl_191_9_LC_26_23_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_191_9_LC_26_23_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84352),
            .lcout(shift_srl_191Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93374),
            .ce(N__86061),
            .sr(_gnd_net_));
    defparam shift_srl_191_8_LC_26_23_7.C_ON=1'b0;
    defparam shift_srl_191_8_LC_26_23_7.SEQ_MODE=4'b1000;
    defparam shift_srl_191_8_LC_26_23_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_191_8_LC_26_23_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86176),
            .lcout(shift_srl_191Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93374),
            .ce(N__86061),
            .sr(_gnd_net_));
    defparam shift_srl_36_6_LC_26_24_7.C_ON=1'b0;
    defparam shift_srl_36_6_LC_26_24_7.SEQ_MODE=4'b1000;
    defparam shift_srl_36_6_LC_26_24_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_36_6_LC_26_24_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84466),
            .lcout(shift_srl_36Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93390),
            .ce(N__90938),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_79_LC_27_1_0.C_ON=1'b0;
    defparam rco_obuf_RNO_79_LC_27_1_0.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_79_LC_27_1_0.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_79_LC_27_1_0 (
            .in0(N__88549),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84541),
            .lcout(rco_c_79),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_81_LC_27_4_3.C_ON=1'b0;
    defparam rco_obuf_RNO_81_LC_27_4_3.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_81_LC_27_4_3.LUT_INIT=16'b1000100000000000;
    LogicCell40 rco_obuf_RNO_81_LC_27_4_3 (
            .in0(N__86347),
            .in1(N__88460),
            .in2(_gnd_net_),
            .in3(N__88545),
            .lcout(N_785),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_81_0_LC_27_5_0.C_ON=1'b0;
    defparam shift_srl_81_0_LC_27_5_0.SEQ_MODE=4'b1000;
    defparam shift_srl_81_0_LC_27_5_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_81_0_LC_27_5_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86334),
            .lcout(shift_srl_81Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93424),
            .ce(N__86283),
            .sr(_gnd_net_));
    defparam shift_srl_81_1_LC_27_5_1.C_ON=1'b0;
    defparam shift_srl_81_1_LC_27_5_1.SEQ_MODE=4'b1000;
    defparam shift_srl_81_1_LC_27_5_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_81_1_LC_27_5_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84424),
            .lcout(shift_srl_81Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93424),
            .ce(N__86283),
            .sr(_gnd_net_));
    defparam shift_srl_81_2_LC_27_5_2.C_ON=1'b0;
    defparam shift_srl_81_2_LC_27_5_2.SEQ_MODE=4'b1000;
    defparam shift_srl_81_2_LC_27_5_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_81_2_LC_27_5_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84418),
            .lcout(shift_srl_81Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93424),
            .ce(N__86283),
            .sr(_gnd_net_));
    defparam shift_srl_81_3_LC_27_5_3.C_ON=1'b0;
    defparam shift_srl_81_3_LC_27_5_3.SEQ_MODE=4'b1000;
    defparam shift_srl_81_3_LC_27_5_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_81_3_LC_27_5_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84412),
            .lcout(shift_srl_81Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93424),
            .ce(N__86283),
            .sr(_gnd_net_));
    defparam shift_srl_81_4_LC_27_5_4.C_ON=1'b0;
    defparam shift_srl_81_4_LC_27_5_4.SEQ_MODE=4'b1000;
    defparam shift_srl_81_4_LC_27_5_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_81_4_LC_27_5_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84406),
            .lcout(shift_srl_81Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93424),
            .ce(N__86283),
            .sr(_gnd_net_));
    defparam shift_srl_81_5_LC_27_5_5.C_ON=1'b0;
    defparam shift_srl_81_5_LC_27_5_5.SEQ_MODE=4'b1000;
    defparam shift_srl_81_5_LC_27_5_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_81_5_LC_27_5_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84400),
            .lcout(shift_srl_81Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93424),
            .ce(N__86283),
            .sr(_gnd_net_));
    defparam shift_srl_81_6_LC_27_5_6.C_ON=1'b0;
    defparam shift_srl_81_6_LC_27_5_6.SEQ_MODE=4'b1000;
    defparam shift_srl_81_6_LC_27_5_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_81_6_LC_27_5_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84553),
            .lcout(shift_srl_81Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93424),
            .ce(N__86283),
            .sr(_gnd_net_));
    defparam shift_srl_81_7_LC_27_5_7.C_ON=1'b0;
    defparam shift_srl_81_7_LC_27_5_7.SEQ_MODE=4'b1000;
    defparam shift_srl_81_7_LC_27_5_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_81_7_LC_27_5_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84547),
            .lcout(shift_srl_81Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93424),
            .ce(N__86283),
            .sr(_gnd_net_));
    defparam shift_srl_79_RNITG241_15_LC_27_6_0.C_ON=1'b0;
    defparam shift_srl_79_RNITG241_15_LC_27_6_0.SEQ_MODE=4'b0000;
    defparam shift_srl_79_RNITG241_15_LC_27_6_0.LUT_INIT=16'b1000100000000000;
    LogicCell40 shift_srl_79_RNITG241_15_LC_27_6_0 (
            .in0(N__86474),
            .in1(N__84504),
            .in2(_gnd_net_),
            .in3(N__88609),
            .lcout(shift_srl_79_RNITG241Z0Z_15),
            .ltout(shift_srl_79_RNITG241Z0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIUOS6K_15_LC_27_6_1.C_ON=1'b0;
    defparam shift_srl_0_RNIUOS6K_15_LC_27_6_1.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIUOS6K_15_LC_27_6_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNIUOS6K_15_LC_27_6_1 (
            .in0(N__86810),
            .in1(N__90728),
            .in2(N__84532),
            .in3(N__89967),
            .lcout(clk_en_80),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIHB9EK_15_LC_27_6_2.C_ON=1'b0;
    defparam shift_srl_0_RNIHB9EK_15_LC_27_6_2.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIHB9EK_15_LC_27_6_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNIHB9EK_15_LC_27_6_2 (
            .in0(N__89968),
            .in1(N__90729),
            .in2(N__88464),
            .in3(N__86809),
            .lcout(N_786),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_78_RNI3734K_15_LC_27_6_4.C_ON=1'b0;
    defparam shift_srl_78_RNI3734K_15_LC_27_6_4.SEQ_MODE=4'b0000;
    defparam shift_srl_78_RNI3734K_15_LC_27_6_4.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_78_RNI3734K_15_LC_27_6_4 (
            .in0(N__88533),
            .in1(N__84505),
            .in2(N__90242),
            .in3(N__88610),
            .lcout(clk_en_79),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_78_LC_27_6_5.C_ON=1'b0;
    defparam rco_obuf_RNO_78_LC_27_6_5.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_78_LC_27_6_5.LUT_INIT=16'b1000100000000000;
    LogicCell40 rco_obuf_RNO_78_LC_27_6_5 (
            .in0(N__84506),
            .in1(N__88611),
            .in2(_gnd_net_),
            .in3(N__88534),
            .lcout(rco_c_78),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_79_0_LC_27_6_6.C_ON=1'b0;
    defparam shift_srl_79_0_LC_27_6_6.SEQ_MODE=4'b1000;
    defparam shift_srl_79_0_LC_27_6_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_79_0_LC_27_6_6 (
            .in0(N__86475),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_79Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93422),
            .ce(N__86426),
            .sr(_gnd_net_));
    defparam shift_srl_79_1_LC_27_6_7.C_ON=1'b0;
    defparam shift_srl_79_1_LC_27_6_7.SEQ_MODE=4'b1000;
    defparam shift_srl_79_1_LC_27_6_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_79_1_LC_27_6_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84514),
            .lcout(shift_srl_79Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93422),
            .ce(N__86426),
            .sr(_gnd_net_));
    defparam shift_srl_80_RNIS8C41_15_LC_27_7_0.C_ON=1'b0;
    defparam shift_srl_80_RNIS8C41_15_LC_27_7_0.SEQ_MODE=4'b0000;
    defparam shift_srl_80_RNIS8C41_15_LC_27_7_0.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_80_RNIS8C41_15_LC_27_7_0 (
            .in0(N__84674),
            .in1(N__86470),
            .in2(N__86338),
            .in3(N__84500),
            .lcout(rco_int_0_a2_0_a2_0_1_83),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_80_15_LC_27_7_1.C_ON=1'b0;
    defparam shift_srl_80_15_LC_27_7_1.SEQ_MODE=4'b1000;
    defparam shift_srl_80_15_LC_27_7_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_80_15_LC_27_7_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84658),
            .lcout(shift_srl_80Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93417),
            .ce(N__84612),
            .sr(_gnd_net_));
    defparam shift_srl_80_14_LC_27_7_2.C_ON=1'b0;
    defparam shift_srl_80_14_LC_27_7_2.SEQ_MODE=4'b1000;
    defparam shift_srl_80_14_LC_27_7_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_80_14_LC_27_7_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84652),
            .lcout(shift_srl_80Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93417),
            .ce(N__84612),
            .sr(_gnd_net_));
    defparam shift_srl_80_13_LC_27_7_3.C_ON=1'b0;
    defparam shift_srl_80_13_LC_27_7_3.SEQ_MODE=4'b1000;
    defparam shift_srl_80_13_LC_27_7_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_80_13_LC_27_7_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84646),
            .lcout(shift_srl_80Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93417),
            .ce(N__84612),
            .sr(_gnd_net_));
    defparam shift_srl_80_12_LC_27_7_4.C_ON=1'b0;
    defparam shift_srl_80_12_LC_27_7_4.SEQ_MODE=4'b1000;
    defparam shift_srl_80_12_LC_27_7_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_80_12_LC_27_7_4 (
            .in0(N__84640),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_80Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93417),
            .ce(N__84612),
            .sr(_gnd_net_));
    defparam shift_srl_80_11_LC_27_7_5.C_ON=1'b0;
    defparam shift_srl_80_11_LC_27_7_5.SEQ_MODE=4'b1000;
    defparam shift_srl_80_11_LC_27_7_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_80_11_LC_27_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84634),
            .lcout(shift_srl_80Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93417),
            .ce(N__84612),
            .sr(_gnd_net_));
    defparam shift_srl_80_10_LC_27_7_6.C_ON=1'b0;
    defparam shift_srl_80_10_LC_27_7_6.SEQ_MODE=4'b1000;
    defparam shift_srl_80_10_LC_27_7_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_80_10_LC_27_7_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84619),
            .lcout(shift_srl_80Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93417),
            .ce(N__84612),
            .sr(_gnd_net_));
    defparam shift_srl_80_9_LC_27_7_7.C_ON=1'b0;
    defparam shift_srl_80_9_LC_27_7_7.SEQ_MODE=4'b1000;
    defparam shift_srl_80_9_LC_27_7_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_80_9_LC_27_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84628),
            .lcout(shift_srl_80Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93417),
            .ce(N__84612),
            .sr(_gnd_net_));
    defparam shift_srl_76_RNIF788_15_LC_27_8_0.C_ON=1'b0;
    defparam shift_srl_76_RNIF788_15_LC_27_8_0.SEQ_MODE=4'b0000;
    defparam shift_srl_76_RNIF788_15_LC_27_8_0.LUT_INIT=16'b1100110000000000;
    LogicCell40 shift_srl_76_RNIF788_15_LC_27_8_0 (
            .in0(_gnd_net_),
            .in1(N__84580),
            .in2(_gnd_net_),
            .in3(N__88390),
            .lcout(shift_srl_76_RNIF788Z0Z_15),
            .ltout(shift_srl_76_RNIF788Z0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIGF2BJ_15_LC_27_8_1.C_ON=1'b0;
    defparam shift_srl_0_RNIGF2BJ_15_LC_27_8_1.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIGF2BJ_15_LC_27_8_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNIGF2BJ_15_LC_27_8_1 (
            .in0(N__86805),
            .in1(N__90238),
            .in2(N__84556),
            .in3(N__90713),
            .lcout(clk_en_77),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNI9PFLJ_15_LC_27_8_2.C_ON=1'b0;
    defparam shift_srl_0_RNI9PFLJ_15_LC_27_8_2.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNI9PFLJ_15_LC_27_8_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNI9PFLJ_15_LC_27_8_2 (
            .in0(N__90714),
            .in1(N__86804),
            .in2(N__90434),
            .in3(N__88605),
            .lcout(clk_en_78),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_75_15_LC_27_8_3.C_ON=1'b0;
    defparam shift_srl_75_15_LC_27_8_3.SEQ_MODE=4'b1000;
    defparam shift_srl_75_15_LC_27_8_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_75_15_LC_27_8_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84718),
            .lcout(shift_srl_75Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93413),
            .ce(N__88700),
            .sr(_gnd_net_));
    defparam shift_srl_75_14_LC_27_8_4.C_ON=1'b0;
    defparam shift_srl_75_14_LC_27_8_4.SEQ_MODE=4'b1000;
    defparam shift_srl_75_14_LC_27_8_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_75_14_LC_27_8_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84712),
            .lcout(shift_srl_75Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93413),
            .ce(N__88700),
            .sr(_gnd_net_));
    defparam shift_srl_75_13_LC_27_8_5.C_ON=1'b0;
    defparam shift_srl_75_13_LC_27_8_5.SEQ_MODE=4'b1000;
    defparam shift_srl_75_13_LC_27_8_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_75_13_LC_27_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84706),
            .lcout(shift_srl_75Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93413),
            .ce(N__88700),
            .sr(_gnd_net_));
    defparam shift_srl_75_12_LC_27_8_6.C_ON=1'b0;
    defparam shift_srl_75_12_LC_27_8_6.SEQ_MODE=4'b1000;
    defparam shift_srl_75_12_LC_27_8_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_75_12_LC_27_8_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84700),
            .lcout(shift_srl_75Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93413),
            .ce(N__88700),
            .sr(_gnd_net_));
    defparam shift_srl_75_11_LC_27_8_7.C_ON=1'b0;
    defparam shift_srl_75_11_LC_27_8_7.SEQ_MODE=4'b1000;
    defparam shift_srl_75_11_LC_27_8_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_75_11_LC_27_8_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88348),
            .lcout(shift_srl_75Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93413),
            .ce(N__88700),
            .sr(_gnd_net_));
    defparam shift_srl_68_0_LC_27_9_0.C_ON=1'b0;
    defparam shift_srl_68_0_LC_27_9_0.SEQ_MODE=4'b1000;
    defparam shift_srl_68_0_LC_27_9_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_68_0_LC_27_9_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86891),
            .lcout(shift_srl_68Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93406),
            .ce(N__86589),
            .sr(_gnd_net_));
    defparam shift_srl_68_1_LC_27_9_1.C_ON=1'b0;
    defparam shift_srl_68_1_LC_27_9_1.SEQ_MODE=4'b1000;
    defparam shift_srl_68_1_LC_27_9_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_68_1_LC_27_9_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84694),
            .lcout(shift_srl_68Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93406),
            .ce(N__86589),
            .sr(_gnd_net_));
    defparam shift_srl_68_2_LC_27_9_2.C_ON=1'b0;
    defparam shift_srl_68_2_LC_27_9_2.SEQ_MODE=4'b1000;
    defparam shift_srl_68_2_LC_27_9_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_68_2_LC_27_9_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84688),
            .lcout(shift_srl_68Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93406),
            .ce(N__86589),
            .sr(_gnd_net_));
    defparam shift_srl_68_3_LC_27_9_3.C_ON=1'b0;
    defparam shift_srl_68_3_LC_27_9_3.SEQ_MODE=4'b1000;
    defparam shift_srl_68_3_LC_27_9_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_68_3_LC_27_9_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84775),
            .lcout(shift_srl_68Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93406),
            .ce(N__86589),
            .sr(_gnd_net_));
    defparam shift_srl_68_4_LC_27_9_4.C_ON=1'b0;
    defparam shift_srl_68_4_LC_27_9_4.SEQ_MODE=4'b1000;
    defparam shift_srl_68_4_LC_27_9_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_68_4_LC_27_9_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84769),
            .lcout(shift_srl_68Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93406),
            .ce(N__86589),
            .sr(_gnd_net_));
    defparam shift_srl_68_5_LC_27_9_5.C_ON=1'b0;
    defparam shift_srl_68_5_LC_27_9_5.SEQ_MODE=4'b1000;
    defparam shift_srl_68_5_LC_27_9_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_68_5_LC_27_9_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84763),
            .lcout(shift_srl_68Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93406),
            .ce(N__86589),
            .sr(_gnd_net_));
    defparam shift_srl_68_6_LC_27_9_6.C_ON=1'b0;
    defparam shift_srl_68_6_LC_27_9_6.SEQ_MODE=4'b1000;
    defparam shift_srl_68_6_LC_27_9_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_68_6_LC_27_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84757),
            .lcout(shift_srl_68Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93406),
            .ce(N__86589),
            .sr(_gnd_net_));
    defparam shift_srl_68_7_LC_27_9_7.C_ON=1'b0;
    defparam shift_srl_68_7_LC_27_9_7.SEQ_MODE=4'b1000;
    defparam shift_srl_68_7_LC_27_9_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_68_7_LC_27_9_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84751),
            .lcout(shift_srl_68Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93406),
            .ce(N__86589),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_70_LC_27_10_0.C_ON=1'b0;
    defparam rco_obuf_RNO_70_LC_27_10_0.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_70_LC_27_10_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 rco_obuf_RNO_70_LC_27_10_0 (
            .in0(N__84828),
            .in1(N__86656),
            .in2(N__90738),
            .in3(N__86698),
            .lcout(rco_c_70),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_71_RNIGP6R_15_LC_27_10_2.C_ON=1'b0;
    defparam shift_srl_71_RNIGP6R_15_LC_27_10_2.SEQ_MODE=4'b0000;
    defparam shift_srl_71_RNIGP6R_15_LC_27_10_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_71_RNIGP6R_15_LC_27_10_2 (
            .in0(N__86719),
            .in1(N__86655),
            .in2(N__84833),
            .in3(N__86697),
            .lcout(shift_srl_71_RNIGP6RZ0Z_15),
            .ltout(shift_srl_71_RNIGP6RZ0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNI2RR5I_15_LC_27_10_3.C_ON=1'b0;
    defparam shift_srl_0_RNI2RR5I_15_LC_27_10_3.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNI2RR5I_15_LC_27_10_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNI2RR5I_15_LC_27_10_3 (
            .in0(N__85020),
            .in1(N__90236),
            .in2(N__84733),
            .in3(N__84865),
            .lcout(clk_en_72),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNI3F1FH_15_LC_27_10_4.C_ON=1'b0;
    defparam shift_srl_0_RNI3F1FH_15_LC_27_10_4.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNI3F1FH_15_LC_27_10_4.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNI3F1FH_15_LC_27_10_4 (
            .in0(N__84866),
            .in1(N__90234),
            .in2(N__84834),
            .in3(N__85021),
            .lcout(clk_en_69),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_48_RNIB5GEF_15_LC_27_10_5.C_ON=1'b0;
    defparam shift_srl_48_RNIB5GEF_15_LC_27_10_5.SEQ_MODE=4'b0000;
    defparam shift_srl_48_RNIB5GEF_15_LC_27_10_5.LUT_INIT=16'b0001000100000000;
    LogicCell40 shift_srl_48_RNIB5GEF_15_LC_27_10_5 (
            .in0(N__85279),
            .in1(N__85266),
            .in2(_gnd_net_),
            .in3(N__85224),
            .lcout(rco_c_59),
            .ltout(rco_c_59_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNI18Q2J_15_LC_27_10_6.C_ON=1'b0;
    defparam shift_srl_0_RNI18Q2J_15_LC_27_10_6.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNI18Q2J_15_LC_27_10_6.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNI18Q2J_15_LC_27_10_6 (
            .in0(N__90235),
            .in1(N__86754),
            .in2(N__85024),
            .in3(N__85018),
            .lcout(clk_en_75),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_67_RNIA6OAH_15_LC_27_10_7.C_ON=1'b0;
    defparam shift_srl_67_RNIA6OAH_15_LC_27_10_7.SEQ_MODE=4'b0000;
    defparam shift_srl_67_RNIA6OAH_15_LC_27_10_7.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_67_RNIA6OAH_15_LC_27_10_7 (
            .in0(N__85019),
            .in1(N__84864),
            .in2(N__86869),
            .in3(N__90237),
            .lcout(clk_en_68),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_70_RNIF9J4I_15_LC_27_11_0.C_ON=1'b0;
    defparam shift_srl_70_RNIF9J4I_15_LC_27_11_0.SEQ_MODE=4'b0000;
    defparam shift_srl_70_RNIF9J4I_15_LC_27_11_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_70_RNIF9J4I_15_LC_27_11_0 (
            .in0(N__86925),
            .in1(N__86696),
            .in2(N__84835),
            .in3(N__86660),
            .lcout(clk_en_71),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_69_15_LC_27_11_1.C_ON=1'b0;
    defparam shift_srl_69_15_LC_27_11_1.SEQ_MODE=4'b1000;
    defparam shift_srl_69_15_LC_27_11_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_69_15_LC_27_11_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84799),
            .lcout(shift_srl_69Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93391),
            .ce(N__85422),
            .sr(_gnd_net_));
    defparam shift_srl_69_14_LC_27_11_2.C_ON=1'b0;
    defparam shift_srl_69_14_LC_27_11_2.SEQ_MODE=4'b1000;
    defparam shift_srl_69_14_LC_27_11_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_69_14_LC_27_11_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84793),
            .lcout(shift_srl_69Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93391),
            .ce(N__85422),
            .sr(_gnd_net_));
    defparam shift_srl_69_13_LC_27_11_3.C_ON=1'b0;
    defparam shift_srl_69_13_LC_27_11_3.SEQ_MODE=4'b1000;
    defparam shift_srl_69_13_LC_27_11_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_69_13_LC_27_11_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84787),
            .lcout(shift_srl_69Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93391),
            .ce(N__85422),
            .sr(_gnd_net_));
    defparam shift_srl_69_12_LC_27_11_4.C_ON=1'b0;
    defparam shift_srl_69_12_LC_27_11_4.SEQ_MODE=4'b1000;
    defparam shift_srl_69_12_LC_27_11_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_69_12_LC_27_11_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84781),
            .lcout(shift_srl_69Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93391),
            .ce(N__85422),
            .sr(_gnd_net_));
    defparam shift_srl_69_11_LC_27_11_5.C_ON=1'b0;
    defparam shift_srl_69_11_LC_27_11_5.SEQ_MODE=4'b1000;
    defparam shift_srl_69_11_LC_27_11_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_69_11_LC_27_11_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85360),
            .lcout(shift_srl_69Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93391),
            .ce(N__85422),
            .sr(_gnd_net_));
    defparam shift_srl_69_10_LC_27_11_6.C_ON=1'b0;
    defparam shift_srl_69_10_LC_27_11_6.SEQ_MODE=4'b1000;
    defparam shift_srl_69_10_LC_27_11_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_69_10_LC_27_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85432),
            .lcout(shift_srl_69Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93391),
            .ce(N__85422),
            .sr(_gnd_net_));
    defparam shift_srl_71_5_LC_27_12_0.C_ON=1'b0;
    defparam shift_srl_71_5_LC_27_12_0.SEQ_MODE=4'b1000;
    defparam shift_srl_71_5_LC_27_12_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_71_5_LC_27_12_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85354),
            .lcout(shift_srl_71Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93375),
            .ce(N__85296),
            .sr(_gnd_net_));
    defparam shift_srl_71_7_LC_27_12_1.C_ON=1'b0;
    defparam shift_srl_71_7_LC_27_12_1.SEQ_MODE=4'b1000;
    defparam shift_srl_71_7_LC_27_12_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_71_7_LC_27_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85342),
            .lcout(shift_srl_71Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93375),
            .ce(N__85296),
            .sr(_gnd_net_));
    defparam shift_srl_71_6_LC_27_12_2.C_ON=1'b0;
    defparam shift_srl_71_6_LC_27_12_2.SEQ_MODE=4'b1000;
    defparam shift_srl_71_6_LC_27_12_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_71_6_LC_27_12_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85348),
            .lcout(shift_srl_71Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93375),
            .ce(N__85296),
            .sr(_gnd_net_));
    defparam shift_srl_71_13_LC_27_12_3.C_ON=1'b0;
    defparam shift_srl_71_13_LC_27_12_3.SEQ_MODE=4'b1000;
    defparam shift_srl_71_13_LC_27_12_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_71_13_LC_27_12_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85318),
            .lcout(shift_srl_71Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93375),
            .ce(N__85296),
            .sr(_gnd_net_));
    defparam shift_srl_71_14_LC_27_12_4.C_ON=1'b0;
    defparam shift_srl_71_14_LC_27_12_4.SEQ_MODE=4'b1000;
    defparam shift_srl_71_14_LC_27_12_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_71_14_LC_27_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85336),
            .lcout(shift_srl_71Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93375),
            .ce(N__85296),
            .sr(_gnd_net_));
    defparam shift_srl_71_15_LC_27_12_5.C_ON=1'b0;
    defparam shift_srl_71_15_LC_27_12_5.SEQ_MODE=4'b1000;
    defparam shift_srl_71_15_LC_27_12_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_71_15_LC_27_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85330),
            .lcout(shift_srl_71Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93375),
            .ce(N__85296),
            .sr(_gnd_net_));
    defparam shift_srl_71_12_LC_27_12_6.C_ON=1'b0;
    defparam shift_srl_71_12_LC_27_12_6.SEQ_MODE=4'b1000;
    defparam shift_srl_71_12_LC_27_12_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_71_12_LC_27_12_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85324),
            .lcout(shift_srl_71Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93375),
            .ce(N__85296),
            .sr(_gnd_net_));
    defparam shift_srl_71_8_LC_27_12_7.C_ON=1'b0;
    defparam shift_srl_71_8_LC_27_12_7.SEQ_MODE=4'b1000;
    defparam shift_srl_71_8_LC_27_12_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_71_8_LC_27_12_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85312),
            .lcout(shift_srl_71Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93375),
            .ce(N__85296),
            .sr(_gnd_net_));
    defparam shift_srl_69_8_LC_27_13_0.C_ON=1'b0;
    defparam shift_srl_69_8_LC_27_13_0.SEQ_MODE=4'b1000;
    defparam shift_srl_69_8_LC_27_13_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_69_8_LC_27_13_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85444),
            .lcout(shift_srl_69Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93359),
            .ce(N__85423),
            .sr(_gnd_net_));
    defparam shift_srl_69_7_LC_27_13_2.C_ON=1'b0;
    defparam shift_srl_69_7_LC_27_13_2.SEQ_MODE=4'b1000;
    defparam shift_srl_69_7_LC_27_13_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_69_7_LC_27_13_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85456),
            .lcout(shift_srl_69Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93359),
            .ce(N__85423),
            .sr(_gnd_net_));
    defparam shift_srl_69_9_LC_27_13_4.C_ON=1'b0;
    defparam shift_srl_69_9_LC_27_13_4.SEQ_MODE=4'b1000;
    defparam shift_srl_69_9_LC_27_13_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_69_9_LC_27_13_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85438),
            .lcout(shift_srl_69Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93359),
            .ce(N__85423),
            .sr(_gnd_net_));
    defparam shift_srl_70_10_LC_27_14_0.C_ON=1'b0;
    defparam shift_srl_70_10_LC_27_14_0.SEQ_MODE=4'b1000;
    defparam shift_srl_70_10_LC_27_14_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_70_10_LC_27_14_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85522),
            .lcout(shift_srl_70Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93337),
            .ce(N__85510),
            .sr(_gnd_net_));
    defparam shift_srl_70_11_LC_27_14_1.C_ON=1'b0;
    defparam shift_srl_70_11_LC_27_14_1.SEQ_MODE=4'b1000;
    defparam shift_srl_70_11_LC_27_14_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_70_11_LC_27_14_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85390),
            .lcout(shift_srl_70Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93337),
            .ce(N__85510),
            .sr(_gnd_net_));
    defparam shift_srl_70_12_LC_27_14_2.C_ON=1'b0;
    defparam shift_srl_70_12_LC_27_14_2.SEQ_MODE=4'b1000;
    defparam shift_srl_70_12_LC_27_14_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_70_12_LC_27_14_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85384),
            .lcout(shift_srl_70Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93337),
            .ce(N__85510),
            .sr(_gnd_net_));
    defparam shift_srl_70_13_LC_27_14_3.C_ON=1'b0;
    defparam shift_srl_70_13_LC_27_14_3.SEQ_MODE=4'b1000;
    defparam shift_srl_70_13_LC_27_14_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_70_13_LC_27_14_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85378),
            .lcout(shift_srl_70Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93337),
            .ce(N__85510),
            .sr(_gnd_net_));
    defparam shift_srl_70_14_LC_27_14_4.C_ON=1'b0;
    defparam shift_srl_70_14_LC_27_14_4.SEQ_MODE=4'b1000;
    defparam shift_srl_70_14_LC_27_14_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_70_14_LC_27_14_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85372),
            .lcout(shift_srl_70Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93337),
            .ce(N__85510),
            .sr(_gnd_net_));
    defparam shift_srl_70_15_LC_27_14_5.C_ON=1'b0;
    defparam shift_srl_70_15_LC_27_14_5.SEQ_MODE=4'b1000;
    defparam shift_srl_70_15_LC_27_14_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_70_15_LC_27_14_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85366),
            .lcout(shift_srl_70Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93337),
            .ce(N__85510),
            .sr(_gnd_net_));
    defparam shift_srl_70_9_LC_27_14_6.C_ON=1'b0;
    defparam shift_srl_70_9_LC_27_14_6.SEQ_MODE=4'b1000;
    defparam shift_srl_70_9_LC_27_14_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_70_9_LC_27_14_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85528),
            .lcout(shift_srl_70Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93337),
            .ce(N__85510),
            .sr(_gnd_net_));
    defparam shift_srl_70_0_LC_27_14_7.C_ON=1'b0;
    defparam shift_srl_70_0_LC_27_14_7.SEQ_MODE=4'b1000;
    defparam shift_srl_70_0_LC_27_14_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_70_0_LC_27_14_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86694),
            .lcout(shift_srl_70Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93337),
            .ce(N__85510),
            .sr(_gnd_net_));
    defparam shift_srl_34_5_LC_27_15_1.C_ON=1'b0;
    defparam shift_srl_34_5_LC_27_15_1.SEQ_MODE=4'b1000;
    defparam shift_srl_34_5_LC_27_15_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_34_5_LC_27_15_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85498),
            .lcout(shift_srl_34Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93317),
            .ce(N__87121),
            .sr(_gnd_net_));
    defparam shift_srl_34_6_LC_27_15_5.C_ON=1'b0;
    defparam shift_srl_34_6_LC_27_15_5.SEQ_MODE=4'b1000;
    defparam shift_srl_34_6_LC_27_15_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_34_6_LC_27_15_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85492),
            .lcout(shift_srl_34Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93317),
            .ce(N__87121),
            .sr(_gnd_net_));
    defparam shift_srl_37_10_LC_27_17_0.C_ON=1'b0;
    defparam shift_srl_37_10_LC_27_17_0.SEQ_MODE=4'b1000;
    defparam shift_srl_37_10_LC_27_17_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_37_10_LC_27_17_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85462),
            .lcout(shift_srl_37Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93263),
            .ce(N__91857),
            .sr(_gnd_net_));
    defparam shift_srl_37_7_LC_27_17_1.C_ON=1'b0;
    defparam shift_srl_37_7_LC_27_17_1.SEQ_MODE=4'b1000;
    defparam shift_srl_37_7_LC_27_17_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_37_7_LC_27_17_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85468),
            .lcout(shift_srl_37Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93263),
            .ce(N__91857),
            .sr(_gnd_net_));
    defparam shift_srl_37_12_LC_27_17_2.C_ON=1'b0;
    defparam shift_srl_37_12_LC_27_17_2.SEQ_MODE=4'b1000;
    defparam shift_srl_37_12_LC_27_17_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_37_12_LC_27_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__93436),
            .lcout(shift_srl_37Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93263),
            .ce(N__91857),
            .sr(_gnd_net_));
    defparam shift_srl_37_13_LC_27_17_3.C_ON=1'b0;
    defparam shift_srl_37_13_LC_27_17_3.SEQ_MODE=4'b1000;
    defparam shift_srl_37_13_LC_27_17_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_37_13_LC_27_17_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85486),
            .lcout(shift_srl_37Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93263),
            .ce(N__91857),
            .sr(_gnd_net_));
    defparam shift_srl_37_6_LC_27_17_5.C_ON=1'b0;
    defparam shift_srl_37_6_LC_27_17_5.SEQ_MODE=4'b1000;
    defparam shift_srl_37_6_LC_27_17_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_37_6_LC_27_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85474),
            .lcout(shift_srl_37Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93263),
            .ce(N__91857),
            .sr(_gnd_net_));
    defparam shift_srl_37_9_LC_27_17_6.C_ON=1'b0;
    defparam shift_srl_37_9_LC_27_17_6.SEQ_MODE=4'b1000;
    defparam shift_srl_37_9_LC_27_17_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_37_9_LC_27_17_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85621),
            .lcout(shift_srl_37Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93263),
            .ce(N__91857),
            .sr(_gnd_net_));
    defparam shift_srl_37_8_LC_27_17_7.C_ON=1'b0;
    defparam shift_srl_37_8_LC_27_17_7.SEQ_MODE=4'b1000;
    defparam shift_srl_37_8_LC_27_17_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_37_8_LC_27_17_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85627),
            .lcout(shift_srl_37Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93263),
            .ce(N__91857),
            .sr(_gnd_net_));
    defparam shift_srl_33_0_LC_27_18_0.C_ON=1'b0;
    defparam shift_srl_33_0_LC_27_18_0.SEQ_MODE=4'b1000;
    defparam shift_srl_33_0_LC_27_18_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_33_0_LC_27_18_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85556),
            .lcout(shift_srl_33Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93298),
            .ce(N__85644),
            .sr(_gnd_net_));
    defparam shift_srl_33_1_LC_27_18_1.C_ON=1'b0;
    defparam shift_srl_33_1_LC_27_18_1.SEQ_MODE=4'b1000;
    defparam shift_srl_33_1_LC_27_18_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_33_1_LC_27_18_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85615),
            .lcout(shift_srl_33Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93298),
            .ce(N__85644),
            .sr(_gnd_net_));
    defparam shift_srl_33_2_LC_27_18_2.C_ON=1'b0;
    defparam shift_srl_33_2_LC_27_18_2.SEQ_MODE=4'b1000;
    defparam shift_srl_33_2_LC_27_18_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_33_2_LC_27_18_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85609),
            .lcout(shift_srl_33Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93298),
            .ce(N__85644),
            .sr(_gnd_net_));
    defparam shift_srl_33_3_LC_27_18_3.C_ON=1'b0;
    defparam shift_srl_33_3_LC_27_18_3.SEQ_MODE=4'b1000;
    defparam shift_srl_33_3_LC_27_18_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_33_3_LC_27_18_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85603),
            .lcout(shift_srl_33Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93298),
            .ce(N__85644),
            .sr(_gnd_net_));
    defparam shift_srl_33_4_LC_27_18_4.C_ON=1'b0;
    defparam shift_srl_33_4_LC_27_18_4.SEQ_MODE=4'b1000;
    defparam shift_srl_33_4_LC_27_18_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_33_4_LC_27_18_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85597),
            .lcout(shift_srl_33Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93298),
            .ce(N__85644),
            .sr(_gnd_net_));
    defparam shift_srl_33_13_LC_27_18_5.C_ON=1'b0;
    defparam shift_srl_33_13_LC_27_18_5.SEQ_MODE=4'b1000;
    defparam shift_srl_33_13_LC_27_18_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_33_13_LC_27_18_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85690),
            .lcout(shift_srl_33Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93298),
            .ce(N__85644),
            .sr(_gnd_net_));
    defparam shift_srl_33_14_LC_27_18_6.C_ON=1'b0;
    defparam shift_srl_33_14_LC_27_18_6.SEQ_MODE=4'b1000;
    defparam shift_srl_33_14_LC_27_18_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_33_14_LC_27_18_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85591),
            .lcout(shift_srl_33Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93298),
            .ce(N__85644),
            .sr(_gnd_net_));
    defparam shift_srl_33_15_LC_27_18_7.C_ON=1'b0;
    defparam shift_srl_33_15_LC_27_18_7.SEQ_MODE=4'b1000;
    defparam shift_srl_33_15_LC_27_18_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_33_15_LC_27_18_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85585),
            .lcout(shift_srl_33Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93298),
            .ce(N__85644),
            .sr(_gnd_net_));
    defparam shift_srl_33_10_LC_27_19_0.C_ON=1'b0;
    defparam shift_srl_33_10_LC_27_19_0.SEQ_MODE=4'b1000;
    defparam shift_srl_33_10_LC_27_19_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_33_10_LC_27_19_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85666),
            .lcout(shift_srl_33Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93318),
            .ce(N__85648),
            .sr(_gnd_net_));
    defparam shift_srl_33_11_LC_27_19_1.C_ON=1'b0;
    defparam shift_srl_33_11_LC_27_19_1.SEQ_MODE=4'b1000;
    defparam shift_srl_33_11_LC_27_19_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_33_11_LC_27_19_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85702),
            .lcout(shift_srl_33Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93318),
            .ce(N__85648),
            .sr(_gnd_net_));
    defparam shift_srl_33_12_LC_27_19_2.C_ON=1'b0;
    defparam shift_srl_33_12_LC_27_19_2.SEQ_MODE=4'b1000;
    defparam shift_srl_33_12_LC_27_19_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_33_12_LC_27_19_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85696),
            .lcout(shift_srl_33Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93318),
            .ce(N__85648),
            .sr(_gnd_net_));
    defparam shift_srl_33_5_LC_27_19_3.C_ON=1'b0;
    defparam shift_srl_33_5_LC_27_19_3.SEQ_MODE=4'b1000;
    defparam shift_srl_33_5_LC_27_19_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_33_5_LC_27_19_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85684),
            .lcout(shift_srl_33Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93318),
            .ce(N__85648),
            .sr(_gnd_net_));
    defparam shift_srl_33_6_LC_27_19_4.C_ON=1'b0;
    defparam shift_srl_33_6_LC_27_19_4.SEQ_MODE=4'b1000;
    defparam shift_srl_33_6_LC_27_19_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_33_6_LC_27_19_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85678),
            .lcout(shift_srl_33Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93318),
            .ce(N__85648),
            .sr(_gnd_net_));
    defparam shift_srl_33_7_LC_27_19_5.C_ON=1'b0;
    defparam shift_srl_33_7_LC_27_19_5.SEQ_MODE=4'b1000;
    defparam shift_srl_33_7_LC_27_19_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_33_7_LC_27_19_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85672),
            .lcout(shift_srl_33Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93318),
            .ce(N__85648),
            .sr(_gnd_net_));
    defparam shift_srl_33_9_LC_27_19_6.C_ON=1'b0;
    defparam shift_srl_33_9_LC_27_19_6.SEQ_MODE=4'b1000;
    defparam shift_srl_33_9_LC_27_19_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_33_9_LC_27_19_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85654),
            .lcout(shift_srl_33Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93318),
            .ce(N__85648),
            .sr(_gnd_net_));
    defparam shift_srl_33_8_LC_27_19_7.C_ON=1'b0;
    defparam shift_srl_33_8_LC_27_19_7.SEQ_MODE=4'b1000;
    defparam shift_srl_33_8_LC_27_19_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_33_8_LC_27_19_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85660),
            .lcout(shift_srl_33Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93318),
            .ce(N__85648),
            .sr(_gnd_net_));
    defparam shift_srl_164_10_LC_27_20_0.C_ON=1'b0;
    defparam shift_srl_164_10_LC_27_20_0.SEQ_MODE=4'b1000;
    defparam shift_srl_164_10_LC_27_20_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_164_10_LC_27_20_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85726),
            .lcout(shift_srl_164Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93338),
            .ce(N__87785),
            .sr(_gnd_net_));
    defparam shift_srl_164_8_LC_27_20_1.C_ON=1'b0;
    defparam shift_srl_164_8_LC_27_20_1.SEQ_MODE=4'b1000;
    defparam shift_srl_164_8_LC_27_20_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_164_8_LC_27_20_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85714),
            .lcout(shift_srl_164Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93338),
            .ce(N__87785),
            .sr(_gnd_net_));
    defparam shift_srl_164_11_LC_27_20_2.C_ON=1'b0;
    defparam shift_srl_164_11_LC_27_20_2.SEQ_MODE=4'b1000;
    defparam shift_srl_164_11_LC_27_20_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_164_11_LC_27_20_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85750),
            .lcout(shift_srl_164Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93338),
            .ce(N__87785),
            .sr(_gnd_net_));
    defparam shift_srl_164_13_LC_27_20_3.C_ON=1'b0;
    defparam shift_srl_164_13_LC_27_20_3.SEQ_MODE=4'b1000;
    defparam shift_srl_164_13_LC_27_20_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_164_13_LC_27_20_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87514),
            .lcout(shift_srl_164Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93338),
            .ce(N__87785),
            .sr(_gnd_net_));
    defparam shift_srl_164_14_LC_27_20_4.C_ON=1'b0;
    defparam shift_srl_164_14_LC_27_20_4.SEQ_MODE=4'b1000;
    defparam shift_srl_164_14_LC_27_20_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_164_14_LC_27_20_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85744),
            .lcout(shift_srl_164Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93338),
            .ce(N__87785),
            .sr(_gnd_net_));
    defparam shift_srl_164_9_LC_27_20_5.C_ON=1'b0;
    defparam shift_srl_164_9_LC_27_20_5.SEQ_MODE=4'b1000;
    defparam shift_srl_164_9_LC_27_20_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_164_9_LC_27_20_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85732),
            .lcout(shift_srl_164Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93338),
            .ce(N__87785),
            .sr(_gnd_net_));
    defparam shift_srl_164_6_LC_27_20_6.C_ON=1'b0;
    defparam shift_srl_164_6_LC_27_20_6.SEQ_MODE=4'b1000;
    defparam shift_srl_164_6_LC_27_20_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_164_6_LC_27_20_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87526),
            .lcout(shift_srl_164Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93338),
            .ce(N__87785),
            .sr(_gnd_net_));
    defparam shift_srl_164_7_LC_27_20_7.C_ON=1'b0;
    defparam shift_srl_164_7_LC_27_20_7.SEQ_MODE=4'b1000;
    defparam shift_srl_164_7_LC_27_20_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_164_7_LC_27_20_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85720),
            .lcout(shift_srl_164Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93338),
            .ce(N__87785),
            .sr(_gnd_net_));
    defparam shift_srl_163_0_LC_27_21_0.C_ON=1'b0;
    defparam shift_srl_163_0_LC_27_21_0.SEQ_MODE=4'b1000;
    defparam shift_srl_163_0_LC_27_21_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_163_0_LC_27_21_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87749),
            .lcout(shift_srl_163Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93360),
            .ce(N__85807),
            .sr(_gnd_net_));
    defparam shift_srl_163_1_LC_27_21_1.C_ON=1'b0;
    defparam shift_srl_163_1_LC_27_21_1.SEQ_MODE=4'b1000;
    defparam shift_srl_163_1_LC_27_21_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_163_1_LC_27_21_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85708),
            .lcout(shift_srl_163Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93360),
            .ce(N__85807),
            .sr(_gnd_net_));
    defparam shift_srl_163_2_LC_27_21_2.C_ON=1'b0;
    defparam shift_srl_163_2_LC_27_21_2.SEQ_MODE=4'b1000;
    defparam shift_srl_163_2_LC_27_21_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_163_2_LC_27_21_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85849),
            .lcout(shift_srl_163Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93360),
            .ce(N__85807),
            .sr(_gnd_net_));
    defparam shift_srl_163_3_LC_27_21_3.C_ON=1'b0;
    defparam shift_srl_163_3_LC_27_21_3.SEQ_MODE=4'b1000;
    defparam shift_srl_163_3_LC_27_21_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_163_3_LC_27_21_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85843),
            .lcout(shift_srl_163Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93360),
            .ce(N__85807),
            .sr(_gnd_net_));
    defparam shift_srl_163_4_LC_27_21_4.C_ON=1'b0;
    defparam shift_srl_163_4_LC_27_21_4.SEQ_MODE=4'b1000;
    defparam shift_srl_163_4_LC_27_21_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_163_4_LC_27_21_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85837),
            .lcout(shift_srl_163Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93360),
            .ce(N__85807),
            .sr(_gnd_net_));
    defparam shift_srl_163_5_LC_27_21_5.C_ON=1'b0;
    defparam shift_srl_163_5_LC_27_21_5.SEQ_MODE=4'b1000;
    defparam shift_srl_163_5_LC_27_21_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_163_5_LC_27_21_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85831),
            .lcout(shift_srl_163Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93360),
            .ce(N__85807),
            .sr(_gnd_net_));
    defparam shift_srl_163_6_LC_27_21_6.C_ON=1'b0;
    defparam shift_srl_163_6_LC_27_21_6.SEQ_MODE=4'b1000;
    defparam shift_srl_163_6_LC_27_21_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_163_6_LC_27_21_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85825),
            .lcout(shift_srl_163Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93360),
            .ce(N__85807),
            .sr(_gnd_net_));
    defparam shift_srl_163_7_LC_27_21_7.C_ON=1'b0;
    defparam shift_srl_163_7_LC_27_21_7.SEQ_MODE=4'b1000;
    defparam shift_srl_163_7_LC_27_21_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_163_7_LC_27_21_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85819),
            .lcout(shift_srl_163Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93360),
            .ce(N__85807),
            .sr(_gnd_net_));
    defparam shift_srl_191_0_LC_27_22_0.C_ON=1'b0;
    defparam shift_srl_191_0_LC_27_22_0.SEQ_MODE=4'b1000;
    defparam shift_srl_191_0_LC_27_22_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_191_0_LC_27_22_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85776),
            .lcout(shift_srl_191Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93376),
            .ce(N__86062),
            .sr(_gnd_net_));
    defparam shift_srl_191_1_LC_27_22_1.C_ON=1'b0;
    defparam shift_srl_191_1_LC_27_22_1.SEQ_MODE=4'b1000;
    defparam shift_srl_191_1_LC_27_22_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_191_1_LC_27_22_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85762),
            .lcout(shift_srl_191Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93376),
            .ce(N__86062),
            .sr(_gnd_net_));
    defparam shift_srl_191_2_LC_27_22_2.C_ON=1'b0;
    defparam shift_srl_191_2_LC_27_22_2.SEQ_MODE=4'b1000;
    defparam shift_srl_191_2_LC_27_22_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_191_2_LC_27_22_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85756),
            .lcout(shift_srl_191Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93376),
            .ce(N__86062),
            .sr(_gnd_net_));
    defparam shift_srl_191_3_LC_27_22_3.C_ON=1'b0;
    defparam shift_srl_191_3_LC_27_22_3.SEQ_MODE=4'b1000;
    defparam shift_srl_191_3_LC_27_22_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_191_3_LC_27_22_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86206),
            .lcout(shift_srl_191Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93376),
            .ce(N__86062),
            .sr(_gnd_net_));
    defparam shift_srl_191_4_LC_27_22_4.C_ON=1'b0;
    defparam shift_srl_191_4_LC_27_22_4.SEQ_MODE=4'b1000;
    defparam shift_srl_191_4_LC_27_22_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_191_4_LC_27_22_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86200),
            .lcout(shift_srl_191Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93376),
            .ce(N__86062),
            .sr(_gnd_net_));
    defparam shift_srl_191_5_LC_27_22_5.C_ON=1'b0;
    defparam shift_srl_191_5_LC_27_22_5.SEQ_MODE=4'b1000;
    defparam shift_srl_191_5_LC_27_22_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_191_5_LC_27_22_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86194),
            .lcout(shift_srl_191Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93376),
            .ce(N__86062),
            .sr(_gnd_net_));
    defparam shift_srl_191_6_LC_27_22_6.C_ON=1'b0;
    defparam shift_srl_191_6_LC_27_22_6.SEQ_MODE=4'b1000;
    defparam shift_srl_191_6_LC_27_22_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_191_6_LC_27_22_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86188),
            .lcout(shift_srl_191Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93376),
            .ce(N__86062),
            .sr(_gnd_net_));
    defparam shift_srl_191_7_LC_27_22_7.C_ON=1'b0;
    defparam shift_srl_191_7_LC_27_22_7.SEQ_MODE=4'b1000;
    defparam shift_srl_191_7_LC_27_22_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_191_7_LC_27_22_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86182),
            .lcout(shift_srl_191Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93376),
            .ce(N__86062),
            .sr(_gnd_net_));
    defparam shift_srl_187_RNI6LJV_0_15_LC_27_23_1.C_ON=1'b0;
    defparam shift_srl_187_RNI6LJV_0_15_LC_27_23_1.SEQ_MODE=4'b0000;
    defparam shift_srl_187_RNI6LJV_0_15_LC_27_23_1.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_187_RNI6LJV_0_15_LC_27_23_1 (
            .in0(N__91821),
            .in1(N__91767),
            .in2(N__86170),
            .in3(N__91682),
            .lcout(),
            .ltout(clk_en_0_a3_0_a2_0_sx_190_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_189_RNIV7I81_15_LC_27_23_2.C_ON=1'b0;
    defparam shift_srl_189_RNIV7I81_15_LC_27_23_2.SEQ_MODE=4'b0000;
    defparam shift_srl_189_RNIV7I81_15_LC_27_23_2.LUT_INIT=16'b0000110000000000;
    LogicCell40 shift_srl_189_RNIV7I81_15_LC_27_23_2 (
            .in0(_gnd_net_),
            .in1(N__86140),
            .in2(N__86107),
            .in3(N__86104),
            .lcout(N_4175),
            .ltout(N_4175_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_190_RNIISOTF1_15_LC_27_23_3.C_ON=1'b0;
    defparam shift_srl_190_RNIISOTF1_15_LC_27_23_3.SEQ_MODE=4'b0000;
    defparam shift_srl_190_RNIISOTF1_15_LC_27_23_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_190_RNIISOTF1_15_LC_27_23_3 (
            .in0(N__90454),
            .in1(N__91606),
            .in2(N__86065),
            .in3(N__91493),
            .lcout(clk_en_191),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIDGJIF1_15_LC_27_23_5.C_ON=1'b0;
    defparam shift_srl_0_RNIDGJIF1_15_LC_27_23_5.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIDGJIF1_15_LC_27_23_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNIDGJIF1_15_LC_27_23_5 (
            .in0(N__90453),
            .in1(N__86050),
            .in2(N__91565),
            .in3(N__85984),
            .lcout(clk_en_190),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_79_2_LC_28_5_0.C_ON=1'b0;
    defparam shift_srl_79_2_LC_28_5_0.SEQ_MODE=4'b1000;
    defparam shift_srl_79_2_LC_28_5_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_79_2_LC_28_5_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86254),
            .lcout(shift_srl_79Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93426),
            .ce(N__86427),
            .sr(_gnd_net_));
    defparam shift_srl_79_3_LC_28_5_1.C_ON=1'b0;
    defparam shift_srl_79_3_LC_28_5_1.SEQ_MODE=4'b1000;
    defparam shift_srl_79_3_LC_28_5_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_79_3_LC_28_5_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86248),
            .lcout(shift_srl_79Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93426),
            .ce(N__86427),
            .sr(_gnd_net_));
    defparam shift_srl_79_4_LC_28_5_2.C_ON=1'b0;
    defparam shift_srl_79_4_LC_28_5_2.SEQ_MODE=4'b1000;
    defparam shift_srl_79_4_LC_28_5_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_79_4_LC_28_5_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86242),
            .lcout(shift_srl_79Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93426),
            .ce(N__86427),
            .sr(_gnd_net_));
    defparam shift_srl_79_5_LC_28_5_3.C_ON=1'b0;
    defparam shift_srl_79_5_LC_28_5_3.SEQ_MODE=4'b1000;
    defparam shift_srl_79_5_LC_28_5_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_79_5_LC_28_5_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86236),
            .lcout(shift_srl_79Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93426),
            .ce(N__86427),
            .sr(_gnd_net_));
    defparam shift_srl_79_6_LC_28_5_4.C_ON=1'b0;
    defparam shift_srl_79_6_LC_28_5_4.SEQ_MODE=4'b1000;
    defparam shift_srl_79_6_LC_28_5_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_79_6_LC_28_5_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86230),
            .lcout(shift_srl_79Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93426),
            .ce(N__86427),
            .sr(_gnd_net_));
    defparam shift_srl_79_7_LC_28_5_5.C_ON=1'b0;
    defparam shift_srl_79_7_LC_28_5_5.SEQ_MODE=4'b1000;
    defparam shift_srl_79_7_LC_28_5_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_79_7_LC_28_5_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86224),
            .lcout(shift_srl_79Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93426),
            .ce(N__86427),
            .sr(_gnd_net_));
    defparam shift_srl_81_10_LC_28_6_0.C_ON=1'b0;
    defparam shift_srl_81_10_LC_28_6_0.SEQ_MODE=4'b1000;
    defparam shift_srl_81_10_LC_28_6_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_81_10_LC_28_6_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86302),
            .lcout(shift_srl_81Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93425),
            .ce(N__86284),
            .sr(_gnd_net_));
    defparam shift_srl_81_11_LC_28_6_1.C_ON=1'b0;
    defparam shift_srl_81_11_LC_28_6_1.SEQ_MODE=4'b1000;
    defparam shift_srl_81_11_LC_28_6_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_81_11_LC_28_6_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86218),
            .lcout(shift_srl_81Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93425),
            .ce(N__86284),
            .sr(_gnd_net_));
    defparam shift_srl_81_12_LC_28_6_2.C_ON=1'b0;
    defparam shift_srl_81_12_LC_28_6_2.SEQ_MODE=4'b1000;
    defparam shift_srl_81_12_LC_28_6_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_81_12_LC_28_6_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86212),
            .lcout(shift_srl_81Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93425),
            .ce(N__86284),
            .sr(_gnd_net_));
    defparam shift_srl_81_13_LC_28_6_3.C_ON=1'b0;
    defparam shift_srl_81_13_LC_28_6_3.SEQ_MODE=4'b1000;
    defparam shift_srl_81_13_LC_28_6_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_81_13_LC_28_6_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86371),
            .lcout(shift_srl_81Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93425),
            .ce(N__86284),
            .sr(_gnd_net_));
    defparam shift_srl_81_14_LC_28_6_4.C_ON=1'b0;
    defparam shift_srl_81_14_LC_28_6_4.SEQ_MODE=4'b1000;
    defparam shift_srl_81_14_LC_28_6_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_81_14_LC_28_6_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86365),
            .lcout(shift_srl_81Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93425),
            .ce(N__86284),
            .sr(_gnd_net_));
    defparam shift_srl_81_15_LC_28_6_5.C_ON=1'b0;
    defparam shift_srl_81_15_LC_28_6_5.SEQ_MODE=4'b1000;
    defparam shift_srl_81_15_LC_28_6_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_81_15_LC_28_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86359),
            .lcout(shift_srl_81Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93425),
            .ce(N__86284),
            .sr(_gnd_net_));
    defparam shift_srl_81_9_LC_28_6_6.C_ON=1'b0;
    defparam shift_srl_81_9_LC_28_6_6.SEQ_MODE=4'b1000;
    defparam shift_srl_81_9_LC_28_6_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_81_9_LC_28_6_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86290),
            .lcout(shift_srl_81Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93425),
            .ce(N__86284),
            .sr(_gnd_net_));
    defparam shift_srl_81_8_LC_28_6_7.C_ON=1'b0;
    defparam shift_srl_81_8_LC_28_6_7.SEQ_MODE=4'b1000;
    defparam shift_srl_81_8_LC_28_6_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_81_8_LC_28_6_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86296),
            .lcout(shift_srl_81Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93425),
            .ce(N__86284),
            .sr(_gnd_net_));
    defparam shift_srl_79_10_LC_28_7_0.C_ON=1'b0;
    defparam shift_srl_79_10_LC_28_7_0.SEQ_MODE=4'b1000;
    defparam shift_srl_79_10_LC_28_7_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_79_10_LC_28_7_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86452),
            .lcout(shift_srl_79Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93423),
            .ce(N__86431),
            .sr(_gnd_net_));
    defparam shift_srl_79_11_LC_28_7_1.C_ON=1'b0;
    defparam shift_srl_79_11_LC_28_7_1.SEQ_MODE=4'b1000;
    defparam shift_srl_79_11_LC_28_7_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_79_11_LC_28_7_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86272),
            .lcout(shift_srl_79Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93423),
            .ce(N__86431),
            .sr(_gnd_net_));
    defparam shift_srl_79_12_LC_28_7_2.C_ON=1'b0;
    defparam shift_srl_79_12_LC_28_7_2.SEQ_MODE=4'b1000;
    defparam shift_srl_79_12_LC_28_7_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_79_12_LC_28_7_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86266),
            .lcout(shift_srl_79Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93423),
            .ce(N__86431),
            .sr(_gnd_net_));
    defparam shift_srl_79_13_LC_28_7_3.C_ON=1'b0;
    defparam shift_srl_79_13_LC_28_7_3.SEQ_MODE=4'b1000;
    defparam shift_srl_79_13_LC_28_7_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_79_13_LC_28_7_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86260),
            .lcout(shift_srl_79Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93423),
            .ce(N__86431),
            .sr(_gnd_net_));
    defparam shift_srl_79_14_LC_28_7_4.C_ON=1'b0;
    defparam shift_srl_79_14_LC_28_7_4.SEQ_MODE=4'b1000;
    defparam shift_srl_79_14_LC_28_7_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_79_14_LC_28_7_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86488),
            .lcout(shift_srl_79Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93423),
            .ce(N__86431),
            .sr(_gnd_net_));
    defparam shift_srl_79_15_LC_28_7_5.C_ON=1'b0;
    defparam shift_srl_79_15_LC_28_7_5.SEQ_MODE=4'b1000;
    defparam shift_srl_79_15_LC_28_7_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_79_15_LC_28_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86482),
            .lcout(shift_srl_79Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93423),
            .ce(N__86431),
            .sr(_gnd_net_));
    defparam shift_srl_79_9_LC_28_7_6.C_ON=1'b0;
    defparam shift_srl_79_9_LC_28_7_6.SEQ_MODE=4'b1000;
    defparam shift_srl_79_9_LC_28_7_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_79_9_LC_28_7_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86437),
            .lcout(shift_srl_79Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93423),
            .ce(N__86431),
            .sr(_gnd_net_));
    defparam shift_srl_79_8_LC_28_7_7.C_ON=1'b0;
    defparam shift_srl_79_8_LC_28_7_7.SEQ_MODE=4'b1000;
    defparam shift_srl_79_8_LC_28_7_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_79_8_LC_28_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86446),
            .lcout(shift_srl_79Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93423),
            .ce(N__86431),
            .sr(_gnd_net_));
    defparam shift_srl_77_10_LC_28_8_0.C_ON=1'b0;
    defparam shift_srl_77_10_LC_28_8_0.SEQ_MODE=4'b1000;
    defparam shift_srl_77_10_LC_28_8_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_77_10_LC_28_8_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86530),
            .lcout(shift_srl_77Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93418),
            .ce(N__88203),
            .sr(_gnd_net_));
    defparam shift_srl_77_11_LC_28_8_1.C_ON=1'b0;
    defparam shift_srl_77_11_LC_28_8_1.SEQ_MODE=4'b1000;
    defparam shift_srl_77_11_LC_28_8_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_77_11_LC_28_8_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86395),
            .lcout(shift_srl_77Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93418),
            .ce(N__88203),
            .sr(_gnd_net_));
    defparam shift_srl_77_12_LC_28_8_2.C_ON=1'b0;
    defparam shift_srl_77_12_LC_28_8_2.SEQ_MODE=4'b1000;
    defparam shift_srl_77_12_LC_28_8_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_77_12_LC_28_8_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86389),
            .lcout(shift_srl_77Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93418),
            .ce(N__88203),
            .sr(_gnd_net_));
    defparam shift_srl_77_13_LC_28_8_3.C_ON=1'b0;
    defparam shift_srl_77_13_LC_28_8_3.SEQ_MODE=4'b1000;
    defparam shift_srl_77_13_LC_28_8_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_77_13_LC_28_8_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86383),
            .lcout(shift_srl_77Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93418),
            .ce(N__88203),
            .sr(_gnd_net_));
    defparam shift_srl_77_14_LC_28_8_4.C_ON=1'b0;
    defparam shift_srl_77_14_LC_28_8_4.SEQ_MODE=4'b1000;
    defparam shift_srl_77_14_LC_28_8_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_77_14_LC_28_8_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86377),
            .lcout(shift_srl_77Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93418),
            .ce(N__88203),
            .sr(_gnd_net_));
    defparam shift_srl_77_15_LC_28_8_5.C_ON=1'b0;
    defparam shift_srl_77_15_LC_28_8_5.SEQ_MODE=4'b1000;
    defparam shift_srl_77_15_LC_28_8_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_77_15_LC_28_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86536),
            .lcout(shift_srl_77Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93418),
            .ce(N__88203),
            .sr(_gnd_net_));
    defparam shift_srl_77_9_LC_28_8_6.C_ON=1'b0;
    defparam shift_srl_77_9_LC_28_8_6.SEQ_MODE=4'b1000;
    defparam shift_srl_77_9_LC_28_8_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_77_9_LC_28_8_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86524),
            .lcout(shift_srl_77Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93418),
            .ce(N__88203),
            .sr(_gnd_net_));
    defparam shift_srl_77_8_LC_28_8_7.C_ON=1'b0;
    defparam shift_srl_77_8_LC_28_8_7.SEQ_MODE=4'b1000;
    defparam shift_srl_77_8_LC_28_8_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_77_8_LC_28_8_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88219),
            .lcout(shift_srl_77Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93418),
            .ce(N__88203),
            .sr(_gnd_net_));
    defparam shift_srl_68_10_LC_28_9_0.C_ON=1'b0;
    defparam shift_srl_68_10_LC_28_9_0.SEQ_MODE=4'b1000;
    defparam shift_srl_68_10_LC_28_9_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_68_10_LC_28_9_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86608),
            .lcout(shift_srl_68Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93414),
            .ce(N__86590),
            .sr(_gnd_net_));
    defparam shift_srl_68_11_LC_28_9_1.C_ON=1'b0;
    defparam shift_srl_68_11_LC_28_9_1.SEQ_MODE=4'b1000;
    defparam shift_srl_68_11_LC_28_9_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_68_11_LC_28_9_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86518),
            .lcout(shift_srl_68Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93414),
            .ce(N__86590),
            .sr(_gnd_net_));
    defparam shift_srl_68_12_LC_28_9_2.C_ON=1'b0;
    defparam shift_srl_68_12_LC_28_9_2.SEQ_MODE=4'b1000;
    defparam shift_srl_68_12_LC_28_9_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_68_12_LC_28_9_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86512),
            .lcout(shift_srl_68Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93414),
            .ce(N__86590),
            .sr(_gnd_net_));
    defparam shift_srl_68_13_LC_28_9_3.C_ON=1'b0;
    defparam shift_srl_68_13_LC_28_9_3.SEQ_MODE=4'b1000;
    defparam shift_srl_68_13_LC_28_9_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_68_13_LC_28_9_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86506),
            .lcout(shift_srl_68Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93414),
            .ce(N__86590),
            .sr(_gnd_net_));
    defparam shift_srl_68_14_LC_28_9_4.C_ON=1'b0;
    defparam shift_srl_68_14_LC_28_9_4.SEQ_MODE=4'b1000;
    defparam shift_srl_68_14_LC_28_9_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_68_14_LC_28_9_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86500),
            .lcout(shift_srl_68Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93414),
            .ce(N__86590),
            .sr(_gnd_net_));
    defparam shift_srl_68_15_LC_28_9_5.C_ON=1'b0;
    defparam shift_srl_68_15_LC_28_9_5.SEQ_MODE=4'b1000;
    defparam shift_srl_68_15_LC_28_9_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_68_15_LC_28_9_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86494),
            .lcout(shift_srl_68Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93414),
            .ce(N__86590),
            .sr(_gnd_net_));
    defparam shift_srl_68_9_LC_28_9_6.C_ON=1'b0;
    defparam shift_srl_68_9_LC_28_9_6.SEQ_MODE=4'b1000;
    defparam shift_srl_68_9_LC_28_9_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_68_9_LC_28_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86596),
            .lcout(shift_srl_68Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93414),
            .ce(N__86590),
            .sr(_gnd_net_));
    defparam shift_srl_68_8_LC_28_9_7.C_ON=1'b0;
    defparam shift_srl_68_8_LC_28_9_7.SEQ_MODE=4'b1000;
    defparam shift_srl_68_8_LC_28_9_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_68_8_LC_28_9_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86602),
            .lcout(shift_srl_68Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93414),
            .ce(N__86590),
            .sr(_gnd_net_));
    defparam shift_srl_72_0_LC_28_10_0.C_ON=1'b0;
    defparam shift_srl_72_0_LC_28_10_0.SEQ_MODE=4'b1000;
    defparam shift_srl_72_0_LC_28_10_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_72_0_LC_28_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__90834),
            .lcout(shift_srl_72Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93407),
            .ce(N__87002),
            .sr(_gnd_net_));
    defparam shift_srl_72_1_LC_28_10_1.C_ON=1'b0;
    defparam shift_srl_72_1_LC_28_10_1.SEQ_MODE=4'b1000;
    defparam shift_srl_72_1_LC_28_10_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_72_1_LC_28_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86572),
            .lcout(shift_srl_72Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93407),
            .ce(N__87002),
            .sr(_gnd_net_));
    defparam shift_srl_72_2_LC_28_10_2.C_ON=1'b0;
    defparam shift_srl_72_2_LC_28_10_2.SEQ_MODE=4'b1000;
    defparam shift_srl_72_2_LC_28_10_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_72_2_LC_28_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86566),
            .lcout(shift_srl_72Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93407),
            .ce(N__87002),
            .sr(_gnd_net_));
    defparam shift_srl_72_3_LC_28_10_3.C_ON=1'b0;
    defparam shift_srl_72_3_LC_28_10_3.SEQ_MODE=4'b1000;
    defparam shift_srl_72_3_LC_28_10_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_72_3_LC_28_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86560),
            .lcout(shift_srl_72Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93407),
            .ce(N__87002),
            .sr(_gnd_net_));
    defparam shift_srl_72_4_LC_28_10_4.C_ON=1'b0;
    defparam shift_srl_72_4_LC_28_10_4.SEQ_MODE=4'b1000;
    defparam shift_srl_72_4_LC_28_10_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_72_4_LC_28_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86554),
            .lcout(shift_srl_72Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93407),
            .ce(N__87002),
            .sr(_gnd_net_));
    defparam shift_srl_72_5_LC_28_10_5.C_ON=1'b0;
    defparam shift_srl_72_5_LC_28_10_5.SEQ_MODE=4'b1000;
    defparam shift_srl_72_5_LC_28_10_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_72_5_LC_28_10_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86548),
            .lcout(shift_srl_72Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93407),
            .ce(N__87002),
            .sr(_gnd_net_));
    defparam shift_srl_72_6_LC_28_10_6.C_ON=1'b0;
    defparam shift_srl_72_6_LC_28_10_6.SEQ_MODE=4'b1000;
    defparam shift_srl_72_6_LC_28_10_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_72_6_LC_28_10_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86542),
            .lcout(shift_srl_72Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93407),
            .ce(N__87002),
            .sr(_gnd_net_));
    defparam shift_srl_72_7_LC_28_10_7.C_ON=1'b0;
    defparam shift_srl_72_7_LC_28_10_7.SEQ_MODE=4'b1000;
    defparam shift_srl_72_7_LC_28_10_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_72_7_LC_28_10_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86944),
            .lcout(shift_srl_72Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93407),
            .ce(N__87002),
            .sr(_gnd_net_));
    defparam shift_srl_73_RNIBAVKI_15_LC_28_11_3.C_ON=1'b0;
    defparam shift_srl_73_RNIBAVKI_15_LC_28_11_3.SEQ_MODE=4'b0000;
    defparam shift_srl_73_RNIBAVKI_15_LC_28_11_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_73_RNIBAVKI_15_LC_28_11_3 (
            .in0(N__90827),
            .in1(N__90883),
            .in2(N__90766),
            .in3(N__86926),
            .lcout(clk_en_74),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_72_15_LC_28_11_4.C_ON=1'b0;
    defparam shift_srl_72_15_LC_28_11_4.SEQ_MODE=4'b1000;
    defparam shift_srl_72_15_LC_28_11_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_72_15_LC_28_11_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87037),
            .lcout(shift_srl_72Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93398),
            .ce(N__87003),
            .sr(_gnd_net_));
    defparam shift_srl_74_RNIS4SR_15_LC_28_11_5.C_ON=1'b0;
    defparam shift_srl_74_RNIS4SR_15_LC_28_11_5.SEQ_MODE=4'b0000;
    defparam shift_srl_74_RNIS4SR_15_LC_28_11_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_74_RNIS4SR_15_LC_28_11_5 (
            .in0(N__90882),
            .in1(N__86892),
            .in2(N__86868),
            .in3(N__88911),
            .lcout(),
            .ltout(shift_srl_74_RNIS4SRZ0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_71_RNIF65O1_15_LC_28_11_6.C_ON=1'b0;
    defparam shift_srl_71_RNIF65O1_15_LC_28_11_6.SEQ_MODE=4'b0000;
    defparam shift_srl_71_RNIF65O1_15_LC_28_11_6.LUT_INIT=16'b1010101011110000;
    LogicCell40 shift_srl_71_RNIF65O1_15_LC_28_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__86824),
            .in3(N__86626),
            .lcout(rco_int_0_a3_0_a2_0_74),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_71_RNIJ19S_15_LC_28_11_7.C_ON=1'b0;
    defparam shift_srl_71_RNIJ19S_15_LC_28_11_7.SEQ_MODE=4'b0000;
    defparam shift_srl_71_RNIJ19S_15_LC_28_11_7.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_srl_71_RNIJ19S_15_LC_28_11_7 (
            .in0(N__86714),
            .in1(N__86695),
            .in2(N__90838),
            .in3(N__86654),
            .lcout(rco_int_0_a3_0_a2_0_1_74),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_72_10_LC_28_12_0.C_ON=1'b0;
    defparam shift_srl_72_10_LC_28_12_0.SEQ_MODE=4'b1000;
    defparam shift_srl_72_10_LC_28_12_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_72_10_LC_28_12_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87031),
            .lcout(shift_srl_72Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93392),
            .ce(N__87010),
            .sr(_gnd_net_));
    defparam shift_srl_72_11_LC_28_12_1.C_ON=1'b0;
    defparam shift_srl_72_11_LC_28_12_1.SEQ_MODE=4'b1000;
    defparam shift_srl_72_11_LC_28_12_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_72_11_LC_28_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86620),
            .lcout(shift_srl_72Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93392),
            .ce(N__87010),
            .sr(_gnd_net_));
    defparam shift_srl_72_12_LC_28_12_2.C_ON=1'b0;
    defparam shift_srl_72_12_LC_28_12_2.SEQ_MODE=4'b1000;
    defparam shift_srl_72_12_LC_28_12_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_72_12_LC_28_12_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86614),
            .lcout(shift_srl_72Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93392),
            .ce(N__87010),
            .sr(_gnd_net_));
    defparam shift_srl_72_13_LC_28_12_3.C_ON=1'b0;
    defparam shift_srl_72_13_LC_28_12_3.SEQ_MODE=4'b1000;
    defparam shift_srl_72_13_LC_28_12_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_72_13_LC_28_12_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87049),
            .lcout(shift_srl_72Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93392),
            .ce(N__87010),
            .sr(_gnd_net_));
    defparam shift_srl_72_14_LC_28_12_4.C_ON=1'b0;
    defparam shift_srl_72_14_LC_28_12_4.SEQ_MODE=4'b1000;
    defparam shift_srl_72_14_LC_28_12_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_72_14_LC_28_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87043),
            .lcout(shift_srl_72Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93392),
            .ce(N__87010),
            .sr(_gnd_net_));
    defparam shift_srl_72_9_LC_28_12_5.C_ON=1'b0;
    defparam shift_srl_72_9_LC_28_12_5.SEQ_MODE=4'b1000;
    defparam shift_srl_72_9_LC_28_12_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_72_9_LC_28_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87016),
            .lcout(shift_srl_72Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93392),
            .ce(N__87010),
            .sr(_gnd_net_));
    defparam shift_srl_72_8_LC_28_12_6.C_ON=1'b0;
    defparam shift_srl_72_8_LC_28_12_6.SEQ_MODE=4'b1000;
    defparam shift_srl_72_8_LC_28_12_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_72_8_LC_28_12_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87025),
            .lcout(shift_srl_72Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93392),
            .ce(N__87010),
            .sr(_gnd_net_));
    defparam shift_srl_34_7_LC_28_13_5.C_ON=1'b0;
    defparam shift_srl_34_7_LC_28_13_5.SEQ_MODE=4'b1000;
    defparam shift_srl_34_7_LC_28_13_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_34_7_LC_28_13_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86986),
            .lcout(shift_srl_34Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93377),
            .ce(N__87135),
            .sr(_gnd_net_));
    defparam shift_srl_54_5_LC_28_14_0.C_ON=1'b0;
    defparam shift_srl_54_5_LC_28_14_0.SEQ_MODE=4'b1000;
    defparam shift_srl_54_5_LC_28_14_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_54_5_LC_28_14_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86977),
            .lcout(shift_srl_54Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93361),
            .ce(N__87186),
            .sr(_gnd_net_));
    defparam shift_srl_54_6_LC_28_14_1.C_ON=1'b0;
    defparam shift_srl_54_6_LC_28_14_1.SEQ_MODE=4'b1000;
    defparam shift_srl_54_6_LC_28_14_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_54_6_LC_28_14_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86962),
            .lcout(shift_srl_54Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93361),
            .ce(N__87186),
            .sr(_gnd_net_));
    defparam shift_srl_54_7_LC_28_14_2.C_ON=1'b0;
    defparam shift_srl_54_7_LC_28_14_2.SEQ_MODE=4'b1000;
    defparam shift_srl_54_7_LC_28_14_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_54_7_LC_28_14_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86956),
            .lcout(shift_srl_54Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93361),
            .ce(N__87186),
            .sr(_gnd_net_));
    defparam shift_srl_54_8_LC_28_14_3.C_ON=1'b0;
    defparam shift_srl_54_8_LC_28_14_3.SEQ_MODE=4'b1000;
    defparam shift_srl_54_8_LC_28_14_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_54_8_LC_28_14_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86950),
            .lcout(shift_srl_54Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93361),
            .ce(N__87186),
            .sr(_gnd_net_));
    defparam shift_srl_54_9_LC_28_14_4.C_ON=1'b0;
    defparam shift_srl_54_9_LC_28_14_4.SEQ_MODE=4'b1000;
    defparam shift_srl_54_9_LC_28_14_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_54_9_LC_28_14_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87208),
            .lcout(shift_srl_54Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93361),
            .ce(N__87186),
            .sr(_gnd_net_));
    defparam shift_srl_34_8_LC_28_15_1.C_ON=1'b0;
    defparam shift_srl_34_8_LC_28_15_1.SEQ_MODE=4'b1000;
    defparam shift_srl_34_8_LC_28_15_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_34_8_LC_28_15_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87154),
            .lcout(shift_srl_34Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93339),
            .ce(N__87136),
            .sr(_gnd_net_));
    defparam shift_srl_32_10_LC_28_17_0.C_ON=1'b0;
    defparam shift_srl_32_10_LC_28_17_0.SEQ_MODE=4'b1000;
    defparam shift_srl_32_10_LC_28_17_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_32_10_LC_28_17_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87055),
            .lcout(shift_srl_32Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93283),
            .ce(N__88834),
            .sr(_gnd_net_));
    defparam shift_srl_32_11_LC_28_17_1.C_ON=1'b0;
    defparam shift_srl_32_11_LC_28_17_1.SEQ_MODE=4'b1000;
    defparam shift_srl_32_11_LC_28_17_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_32_11_LC_28_17_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87085),
            .lcout(shift_srl_32Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93283),
            .ce(N__88834),
            .sr(_gnd_net_));
    defparam shift_srl_32_12_LC_28_17_2.C_ON=1'b0;
    defparam shift_srl_32_12_LC_28_17_2.SEQ_MODE=4'b1000;
    defparam shift_srl_32_12_LC_28_17_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_32_12_LC_28_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87079),
            .lcout(shift_srl_32Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93283),
            .ce(N__88834),
            .sr(_gnd_net_));
    defparam shift_srl_32_13_LC_28_17_3.C_ON=1'b0;
    defparam shift_srl_32_13_LC_28_17_3.SEQ_MODE=4'b1000;
    defparam shift_srl_32_13_LC_28_17_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_32_13_LC_28_17_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87073),
            .lcout(shift_srl_32Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93283),
            .ce(N__88834),
            .sr(_gnd_net_));
    defparam shift_srl_32_14_LC_28_17_4.C_ON=1'b0;
    defparam shift_srl_32_14_LC_28_17_4.SEQ_MODE=4'b1000;
    defparam shift_srl_32_14_LC_28_17_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_32_14_LC_28_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87067),
            .lcout(shift_srl_32Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93283),
            .ce(N__88834),
            .sr(_gnd_net_));
    defparam shift_srl_32_15_LC_28_17_5.C_ON=1'b0;
    defparam shift_srl_32_15_LC_28_17_5.SEQ_MODE=4'b1000;
    defparam shift_srl_32_15_LC_28_17_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_32_15_LC_28_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87061),
            .lcout(shift_srl_32Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93283),
            .ce(N__88834),
            .sr(_gnd_net_));
    defparam shift_srl_32_9_LC_28_17_6.C_ON=1'b0;
    defparam shift_srl_32_9_LC_28_17_6.SEQ_MODE=4'b1000;
    defparam shift_srl_32_9_LC_28_17_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_32_9_LC_28_17_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87373),
            .lcout(shift_srl_32Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93283),
            .ce(N__88834),
            .sr(_gnd_net_));
    defparam shift_srl_32_8_LC_28_17_7.C_ON=1'b0;
    defparam shift_srl_32_8_LC_28_17_7.SEQ_MODE=4'b1000;
    defparam shift_srl_32_8_LC_28_17_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_32_8_LC_28_17_7 (
            .in0(N__88870),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_32Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93283),
            .ce(N__88834),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIQLID8_15_LC_28_18_0.C_ON=1'b0;
    defparam shift_srl_0_RNIQLID8_15_LC_28_18_0.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIQLID8_15_LC_28_18_0.LUT_INIT=16'b1100110000000000;
    LogicCell40 shift_srl_0_RNIQLID8_15_LC_28_18_0 (
            .in0(_gnd_net_),
            .in1(N__90133),
            .in2(_gnd_net_),
            .in3(N__87347),
            .lcout(clk_en_32),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_32_0_LC_28_18_1.C_ON=1'b0;
    defparam shift_srl_32_0_LC_28_18_1.SEQ_MODE=4'b1000;
    defparam shift_srl_32_0_LC_28_18_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_32_0_LC_28_18_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87298),
            .lcout(shift_srl_32Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93319),
            .ce(N__88825),
            .sr(_gnd_net_));
    defparam shift_srl_32_1_LC_28_18_2.C_ON=1'b0;
    defparam shift_srl_32_1_LC_28_18_2.SEQ_MODE=4'b1000;
    defparam shift_srl_32_1_LC_28_18_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_32_1_LC_28_18_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87268),
            .lcout(shift_srl_32Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93319),
            .ce(N__88825),
            .sr(_gnd_net_));
    defparam shift_srl_32_2_LC_28_18_3.C_ON=1'b0;
    defparam shift_srl_32_2_LC_28_18_3.SEQ_MODE=4'b1000;
    defparam shift_srl_32_2_LC_28_18_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_32_2_LC_28_18_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87262),
            .lcout(shift_srl_32Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93319),
            .ce(N__88825),
            .sr(_gnd_net_));
    defparam shift_srl_164_0_LC_28_19_0.C_ON=1'b0;
    defparam shift_srl_164_0_LC_28_19_0.SEQ_MODE=4'b1000;
    defparam shift_srl_164_0_LC_28_19_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_164_0_LC_28_19_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87256),
            .lcout(shift_srl_164Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93340),
            .ce(N__87795),
            .sr(_gnd_net_));
    defparam shift_srl_164_1_LC_28_19_1.C_ON=1'b0;
    defparam shift_srl_164_1_LC_28_19_1.SEQ_MODE=4'b1000;
    defparam shift_srl_164_1_LC_28_19_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_164_1_LC_28_19_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87226),
            .lcout(shift_srl_164Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93340),
            .ce(N__87795),
            .sr(_gnd_net_));
    defparam shift_srl_164_2_LC_28_19_2.C_ON=1'b0;
    defparam shift_srl_164_2_LC_28_19_2.SEQ_MODE=4'b1000;
    defparam shift_srl_164_2_LC_28_19_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_164_2_LC_28_19_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87220),
            .lcout(shift_srl_164Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93340),
            .ce(N__87795),
            .sr(_gnd_net_));
    defparam shift_srl_164_3_LC_28_19_3.C_ON=1'b0;
    defparam shift_srl_164_3_LC_28_19_3.SEQ_MODE=4'b1000;
    defparam shift_srl_164_3_LC_28_19_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_164_3_LC_28_19_3 (
            .in0(N__87214),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_164Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93340),
            .ce(N__87795),
            .sr(_gnd_net_));
    defparam shift_srl_164_4_LC_28_19_4.C_ON=1'b0;
    defparam shift_srl_164_4_LC_28_19_4.SEQ_MODE=4'b1000;
    defparam shift_srl_164_4_LC_28_19_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_164_4_LC_28_19_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87538),
            .lcout(shift_srl_164Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93340),
            .ce(N__87795),
            .sr(_gnd_net_));
    defparam shift_srl_164_5_LC_28_19_5.C_ON=1'b0;
    defparam shift_srl_164_5_LC_28_19_5.SEQ_MODE=4'b1000;
    defparam shift_srl_164_5_LC_28_19_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_164_5_LC_28_19_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87532),
            .lcout(shift_srl_164Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93340),
            .ce(N__87795),
            .sr(_gnd_net_));
    defparam shift_srl_164_12_LC_28_19_7.C_ON=1'b0;
    defparam shift_srl_164_12_LC_28_19_7.SEQ_MODE=4'b1000;
    defparam shift_srl_164_12_LC_28_19_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_164_12_LC_28_19_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87520),
            .lcout(shift_srl_164Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93340),
            .ce(N__87795),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_171_LC_28_20_0.C_ON=1'b0;
    defparam rco_obuf_RNO_171_LC_28_20_0.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_171_LC_28_20_0.LUT_INIT=16'b1000100010001000;
    LogicCell40 rco_obuf_RNO_171_LC_28_20_0 (
            .in0(N__87719),
            .in1(N__87475),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(rco_c_171),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_171_RNIVSP62_15_LC_28_20_1.C_ON=1'b0;
    defparam shift_srl_171_RNIVSP62_15_LC_28_20_1.SEQ_MODE=4'b0000;
    defparam shift_srl_171_RNIVSP62_15_LC_28_20_1.LUT_INIT=16'b1100110000000000;
    LogicCell40 shift_srl_171_RNIVSP62_15_LC_28_20_1 (
            .in0(_gnd_net_),
            .in1(N__87496),
            .in2(_gnd_net_),
            .in3(N__87461),
            .lcout(shift_srl_171_RNIVSP62Z0Z_15),
            .ltout(shift_srl_171_RNIVSP62Z0Z_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIKHP0B1_15_LC_28_20_2.C_ON=1'b0;
    defparam shift_srl_0_RNIKHP0B1_15_LC_28_20_2.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIKHP0B1_15_LC_28_20_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNIKHP0B1_15_LC_28_20_2 (
            .in0(N__88010),
            .in1(N__90472),
            .in2(N__87469),
            .in3(N__87875),
            .lcout(clk_en_172),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_170_LC_28_20_3.C_ON=1'b0;
    defparam rco_obuf_RNO_170_LC_28_20_3.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_170_LC_28_20_3.LUT_INIT=16'b1100110000000000;
    LogicCell40 rco_obuf_RNO_170_LC_28_20_3 (
            .in0(_gnd_net_),
            .in1(N__87718),
            .in2(_gnd_net_),
            .in3(N__87462),
            .lcout(rco_c_170),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_0_RNIOARV91_15_LC_28_20_4.C_ON=1'b0;
    defparam shift_srl_0_RNIOARV91_15_LC_28_20_4.SEQ_MODE=4'b0000;
    defparam shift_srl_0_RNIOARV91_15_LC_28_20_4.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_0_RNIOARV91_15_LC_28_20_4 (
            .in0(N__88011),
            .in1(N__90471),
            .in2(N__87425),
            .in3(N__87874),
            .lcout(clk_en_168),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_167_LC_28_20_5.C_ON=1'b0;
    defparam rco_obuf_RNO_167_LC_28_20_5.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_167_LC_28_20_5.LUT_INIT=16'b1100110000000000;
    LogicCell40 rco_obuf_RNO_167_LC_28_20_5 (
            .in0(_gnd_net_),
            .in1(N__87717),
            .in2(_gnd_net_),
            .in3(N__87419),
            .lcout(rco_c_167),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_163_RNIQTO291_15_LC_28_20_6.C_ON=1'b0;
    defparam shift_srl_163_RNIQTO291_15_LC_28_20_6.SEQ_MODE=4'b0000;
    defparam shift_srl_163_RNIQTO291_15_LC_28_20_6.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_163_RNIQTO291_15_LC_28_20_6 (
            .in0(N__88009),
            .in1(N__87761),
            .in2(N__90550),
            .in3(N__87873),
            .lcout(clk_en_164),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_163_LC_28_20_7.C_ON=1'b0;
    defparam rco_obuf_RNO_163_LC_28_20_7.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_163_LC_28_20_7.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_163_LC_28_20_7 (
            .in0(N__87762),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87716),
            .lcout(rco_c_163),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_168_0_LC_28_21_0.C_ON=1'b0;
    defparam shift_srl_168_0_LC_28_21_0.SEQ_MODE=4'b1000;
    defparam shift_srl_168_0_LC_28_21_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_168_0_LC_28_21_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__89170),
            .lcout(shift_srl_168Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93378),
            .ce(N__89105),
            .sr(_gnd_net_));
    defparam shift_srl_168_1_LC_28_21_1.C_ON=1'b0;
    defparam shift_srl_168_1_LC_28_21_1.SEQ_MODE=4'b1000;
    defparam shift_srl_168_1_LC_28_21_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_168_1_LC_28_21_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87574),
            .lcout(shift_srl_168Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93378),
            .ce(N__89105),
            .sr(_gnd_net_));
    defparam shift_srl_168_2_LC_28_21_2.C_ON=1'b0;
    defparam shift_srl_168_2_LC_28_21_2.SEQ_MODE=4'b1000;
    defparam shift_srl_168_2_LC_28_21_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_168_2_LC_28_21_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87568),
            .lcout(shift_srl_168Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93378),
            .ce(N__89105),
            .sr(_gnd_net_));
    defparam shift_srl_168_3_LC_28_21_3.C_ON=1'b0;
    defparam shift_srl_168_3_LC_28_21_3.SEQ_MODE=4'b1000;
    defparam shift_srl_168_3_LC_28_21_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_168_3_LC_28_21_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87562),
            .lcout(shift_srl_168Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93378),
            .ce(N__89105),
            .sr(_gnd_net_));
    defparam shift_srl_168_4_LC_28_21_4.C_ON=1'b0;
    defparam shift_srl_168_4_LC_28_21_4.SEQ_MODE=4'b1000;
    defparam shift_srl_168_4_LC_28_21_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_168_4_LC_28_21_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87556),
            .lcout(shift_srl_168Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93378),
            .ce(N__89105),
            .sr(_gnd_net_));
    defparam shift_srl_168_5_LC_28_21_5.C_ON=1'b0;
    defparam shift_srl_168_5_LC_28_21_5.SEQ_MODE=4'b1000;
    defparam shift_srl_168_5_LC_28_21_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_168_5_LC_28_21_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87550),
            .lcout(shift_srl_168Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93378),
            .ce(N__89105),
            .sr(_gnd_net_));
    defparam shift_srl_168_6_LC_28_21_6.C_ON=1'b0;
    defparam shift_srl_168_6_LC_28_21_6.SEQ_MODE=4'b1000;
    defparam shift_srl_168_6_LC_28_21_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_168_6_LC_28_21_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87544),
            .lcout(shift_srl_168Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93378),
            .ce(N__89105),
            .sr(_gnd_net_));
    defparam shift_srl_168_7_LC_28_21_7.C_ON=1'b0;
    defparam shift_srl_168_7_LC_28_21_7.SEQ_MODE=4'b1000;
    defparam shift_srl_168_7_LC_28_21_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_168_7_LC_28_21_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88054),
            .lcout(shift_srl_168Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93378),
            .ce(N__89105),
            .sr(_gnd_net_));
    defparam shift_srl_190_10_LC_28_22_0.C_ON=1'b0;
    defparam shift_srl_190_10_LC_28_22_0.SEQ_MODE=4'b1000;
    defparam shift_srl_190_10_LC_28_22_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_190_10_LC_28_22_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88048),
            .lcout(shift_srl_190Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93393),
            .ce(N__88132),
            .sr(_gnd_net_));
    defparam shift_srl_190_9_LC_28_22_1.C_ON=1'b0;
    defparam shift_srl_190_9_LC_28_22_1.SEQ_MODE=4'b1000;
    defparam shift_srl_190_9_LC_28_22_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_190_9_LC_28_22_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88186),
            .lcout(shift_srl_190Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93393),
            .ce(N__88132),
            .sr(_gnd_net_));
    defparam shift_srl_190_5_LC_28_22_2.C_ON=1'b0;
    defparam shift_srl_190_5_LC_28_22_2.SEQ_MODE=4'b1000;
    defparam shift_srl_190_5_LC_28_22_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_190_5_LC_28_22_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88036),
            .lcout(shift_srl_190Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93393),
            .ce(N__88132),
            .sr(_gnd_net_));
    defparam shift_srl_190_3_LC_28_22_3.C_ON=1'b0;
    defparam shift_srl_190_3_LC_28_22_3.SEQ_MODE=4'b1000;
    defparam shift_srl_190_3_LC_28_22_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_190_3_LC_28_22_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88150),
            .lcout(shift_srl_190Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93393),
            .ce(N__88132),
            .sr(_gnd_net_));
    defparam shift_srl_190_4_LC_28_22_4.C_ON=1'b0;
    defparam shift_srl_190_4_LC_28_22_4.SEQ_MODE=4'b1000;
    defparam shift_srl_190_4_LC_28_22_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_190_4_LC_28_22_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88042),
            .lcout(shift_srl_190Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93393),
            .ce(N__88132),
            .sr(_gnd_net_));
    defparam shift_srl_190_11_LC_28_22_5.C_ON=1'b0;
    defparam shift_srl_190_11_LC_28_22_5.SEQ_MODE=4'b1000;
    defparam shift_srl_190_11_LC_28_22_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_190_11_LC_28_22_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88030),
            .lcout(shift_srl_190Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93393),
            .ce(N__88132),
            .sr(_gnd_net_));
    defparam shift_srl_190_6_LC_28_22_6.C_ON=1'b0;
    defparam shift_srl_190_6_LC_28_22_6.SEQ_MODE=4'b1000;
    defparam shift_srl_190_6_LC_28_22_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_190_6_LC_28_22_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88024),
            .lcout(shift_srl_190Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93393),
            .ce(N__88132),
            .sr(_gnd_net_));
    defparam shift_srl_190_12_LC_28_22_7.C_ON=1'b0;
    defparam shift_srl_190_12_LC_28_22_7.SEQ_MODE=4'b1000;
    defparam shift_srl_190_12_LC_28_22_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_190_12_LC_28_22_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88018),
            .lcout(shift_srl_190Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93393),
            .ce(N__88132),
            .sr(_gnd_net_));
    defparam shift_srl_190_14_LC_28_23_0.C_ON=1'b0;
    defparam shift_srl_190_14_LC_28_23_0.SEQ_MODE=4'b1000;
    defparam shift_srl_190_14_LC_28_23_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_190_14_LC_28_23_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88162),
            .lcout(shift_srl_190Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93399),
            .ce(N__88128),
            .sr(_gnd_net_));
    defparam shift_srl_190_8_LC_28_23_1.C_ON=1'b0;
    defparam shift_srl_190_8_LC_28_23_1.SEQ_MODE=4'b1000;
    defparam shift_srl_190_8_LC_28_23_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_190_8_LC_28_23_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88174),
            .lcout(shift_srl_190Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93399),
            .ce(N__88128),
            .sr(_gnd_net_));
    defparam shift_srl_190_7_LC_28_23_2.C_ON=1'b0;
    defparam shift_srl_190_7_LC_28_23_2.SEQ_MODE=4'b1000;
    defparam shift_srl_190_7_LC_28_23_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_190_7_LC_28_23_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88180),
            .lcout(shift_srl_190Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93399),
            .ce(N__88128),
            .sr(_gnd_net_));
    defparam shift_srl_190_13_LC_28_23_3.C_ON=1'b0;
    defparam shift_srl_190_13_LC_28_23_3.SEQ_MODE=4'b1000;
    defparam shift_srl_190_13_LC_28_23_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_190_13_LC_28_23_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88168),
            .lcout(shift_srl_190Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93399),
            .ce(N__88128),
            .sr(_gnd_net_));
    defparam shift_srl_190_0_LC_28_23_4.C_ON=1'b0;
    defparam shift_srl_190_0_LC_28_23_4.SEQ_MODE=4'b1000;
    defparam shift_srl_190_0_LC_28_23_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_190_0_LC_28_23_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__91607),
            .lcout(shift_srl_190Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93399),
            .ce(N__88128),
            .sr(_gnd_net_));
    defparam shift_srl_190_15_LC_28_23_5.C_ON=1'b0;
    defparam shift_srl_190_15_LC_28_23_5.SEQ_MODE=4'b1000;
    defparam shift_srl_190_15_LC_28_23_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_190_15_LC_28_23_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88156),
            .lcout(shift_srl_190Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93399),
            .ce(N__88128),
            .sr(_gnd_net_));
    defparam shift_srl_190_2_LC_28_23_6.C_ON=1'b0;
    defparam shift_srl_190_2_LC_28_23_6.SEQ_MODE=4'b1000;
    defparam shift_srl_190_2_LC_28_23_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_190_2_LC_28_23_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88138),
            .lcout(shift_srl_190Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93399),
            .ce(N__88128),
            .sr(_gnd_net_));
    defparam shift_srl_190_1_LC_28_23_7.C_ON=1'b0;
    defparam shift_srl_190_1_LC_28_23_7.SEQ_MODE=4'b1000;
    defparam shift_srl_190_1_LC_28_23_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_190_1_LC_28_23_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88144),
            .lcout(shift_srl_190Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93399),
            .ce(N__88128),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_139_LC_28_24_6.C_ON=1'b0;
    defparam rco_obuf_RNO_139_LC_28_24_6.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_139_LC_28_24_6.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_139_LC_28_24_6 (
            .in0(N__91112),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88114),
            .lcout(rco_c_139),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_50_LC_29_2_3.C_ON=1'b0;
    defparam rco_obuf_RNO_50_LC_29_2_3.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_50_LC_29_2_3.LUT_INIT=16'b1100110000000000;
    LogicCell40 rco_obuf_RNO_50_LC_29_2_3 (
            .in0(_gnd_net_),
            .in1(N__88336),
            .in2(_gnd_net_),
            .in3(N__93615),
            .lcout(rco_c_50),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_77_0_LC_29_5_0.C_ON=1'b0;
    defparam shift_srl_77_0_LC_29_5_0.SEQ_MODE=4'b1000;
    defparam shift_srl_77_0_LC_29_5_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_77_0_LC_29_5_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88279),
            .lcout(shift_srl_77Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93427),
            .ce(N__88207),
            .sr(_gnd_net_));
    defparam shift_srl_77_1_LC_29_5_1.C_ON=1'b0;
    defparam shift_srl_77_1_LC_29_5_1.SEQ_MODE=4'b1000;
    defparam shift_srl_77_1_LC_29_5_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_77_1_LC_29_5_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88261),
            .lcout(shift_srl_77Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93427),
            .ce(N__88207),
            .sr(_gnd_net_));
    defparam shift_srl_77_2_LC_29_5_2.C_ON=1'b0;
    defparam shift_srl_77_2_LC_29_5_2.SEQ_MODE=4'b1000;
    defparam shift_srl_77_2_LC_29_5_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_77_2_LC_29_5_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88255),
            .lcout(shift_srl_77Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93427),
            .ce(N__88207),
            .sr(_gnd_net_));
    defparam shift_srl_77_3_LC_29_5_3.C_ON=1'b0;
    defparam shift_srl_77_3_LC_29_5_3.SEQ_MODE=4'b1000;
    defparam shift_srl_77_3_LC_29_5_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_77_3_LC_29_5_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88249),
            .lcout(shift_srl_77Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93427),
            .ce(N__88207),
            .sr(_gnd_net_));
    defparam shift_srl_77_4_LC_29_5_4.C_ON=1'b0;
    defparam shift_srl_77_4_LC_29_5_4.SEQ_MODE=4'b1000;
    defparam shift_srl_77_4_LC_29_5_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_77_4_LC_29_5_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88243),
            .lcout(shift_srl_77Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93427),
            .ce(N__88207),
            .sr(_gnd_net_));
    defparam shift_srl_77_5_LC_29_5_5.C_ON=1'b0;
    defparam shift_srl_77_5_LC_29_5_5.SEQ_MODE=4'b1000;
    defparam shift_srl_77_5_LC_29_5_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_77_5_LC_29_5_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88237),
            .lcout(shift_srl_77Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93427),
            .ce(N__88207),
            .sr(_gnd_net_));
    defparam shift_srl_77_6_LC_29_5_6.C_ON=1'b0;
    defparam shift_srl_77_6_LC_29_5_6.SEQ_MODE=4'b1000;
    defparam shift_srl_77_6_LC_29_5_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_77_6_LC_29_5_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88231),
            .lcout(shift_srl_77Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93427),
            .ce(N__88207),
            .sr(_gnd_net_));
    defparam shift_srl_77_7_LC_29_5_7.C_ON=1'b0;
    defparam shift_srl_77_7_LC_29_5_7.SEQ_MODE=4'b1000;
    defparam shift_srl_77_7_LC_29_5_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_77_7_LC_29_5_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88225),
            .lcout(shift_srl_77Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93427),
            .ce(N__88207),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_75_LC_29_9_0.C_ON=1'b0;
    defparam rco_obuf_RNO_75_LC_29_9_0.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_75_LC_29_9_0.LUT_INIT=16'b1100110000000000;
    LogicCell40 rco_obuf_RNO_75_LC_29_9_0 (
            .in0(_gnd_net_),
            .in1(N__88541),
            .in2(_gnd_net_),
            .in3(N__88405),
            .lcout(rco_c_75),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_76_LC_29_9_1.C_ON=1'b0;
    defparam rco_obuf_RNO_76_LC_29_9_1.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_76_LC_29_9_1.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_76_LC_29_9_1 (
            .in0(N__88542),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88639),
            .lcout(rco_c_76),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_77_LC_29_9_2.C_ON=1'b0;
    defparam rco_obuf_RNO_77_LC_29_9_2.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_77_LC_29_9_2.LUT_INIT=16'b1100110000000000;
    LogicCell40 rco_obuf_RNO_77_LC_29_9_2 (
            .in0(_gnd_net_),
            .in1(N__88543),
            .in2(_gnd_net_),
            .in3(N__88615),
            .lcout(rco_c_77),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_80_LC_29_9_3.C_ON=1'b0;
    defparam rco_obuf_RNO_80_LC_29_9_3.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_80_LC_29_9_3.LUT_INIT=16'b1000100010001000;
    LogicCell40 rco_obuf_RNO_80_LC_29_9_3 (
            .in0(N__88544),
            .in1(N__88465),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(rco_c_80),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_75_0_LC_29_9_4.C_ON=1'b0;
    defparam shift_srl_75_0_LC_29_9_4.SEQ_MODE=4'b1000;
    defparam shift_srl_75_0_LC_29_9_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_75_0_LC_29_9_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88404),
            .lcout(shift_srl_75Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93419),
            .ce(N__88702),
            .sr(_gnd_net_));
    defparam shift_srl_75_1_LC_29_9_5.C_ON=1'b0;
    defparam shift_srl_75_1_LC_29_9_5.SEQ_MODE=4'b1000;
    defparam shift_srl_75_1_LC_29_9_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_75_1_LC_29_9_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88366),
            .lcout(shift_srl_75Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93419),
            .ce(N__88702),
            .sr(_gnd_net_));
    defparam shift_srl_75_2_LC_29_9_6.C_ON=1'b0;
    defparam shift_srl_75_2_LC_29_9_6.SEQ_MODE=4'b1000;
    defparam shift_srl_75_2_LC_29_9_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_75_2_LC_29_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88360),
            .lcout(shift_srl_75Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93419),
            .ce(N__88702),
            .sr(_gnd_net_));
    defparam shift_srl_75_3_LC_29_9_7.C_ON=1'b0;
    defparam shift_srl_75_3_LC_29_9_7.SEQ_MODE=4'b1000;
    defparam shift_srl_75_3_LC_29_9_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_75_3_LC_29_9_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88354),
            .lcout(shift_srl_75Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93419),
            .ce(N__88702),
            .sr(_gnd_net_));
    defparam shift_srl_75_10_LC_29_10_0.C_ON=1'b0;
    defparam shift_srl_75_10_LC_29_10_0.SEQ_MODE=4'b1000;
    defparam shift_srl_75_10_LC_29_10_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_75_10_LC_29_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88744),
            .lcout(shift_srl_75Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93415),
            .ce(N__88701),
            .sr(_gnd_net_));
    defparam shift_srl_75_9_LC_29_10_1.C_ON=1'b0;
    defparam shift_srl_75_9_LC_29_10_1.SEQ_MODE=4'b1000;
    defparam shift_srl_75_9_LC_29_10_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_75_9_LC_29_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88738),
            .lcout(shift_srl_75Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93415),
            .ce(N__88701),
            .sr(_gnd_net_));
    defparam shift_srl_75_8_LC_29_10_2.C_ON=1'b0;
    defparam shift_srl_75_8_LC_29_10_2.SEQ_MODE=4'b1000;
    defparam shift_srl_75_8_LC_29_10_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_75_8_LC_29_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88732),
            .lcout(shift_srl_75Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93415),
            .ce(N__88701),
            .sr(_gnd_net_));
    defparam shift_srl_75_7_LC_29_10_3.C_ON=1'b0;
    defparam shift_srl_75_7_LC_29_10_3.SEQ_MODE=4'b1000;
    defparam shift_srl_75_7_LC_29_10_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_75_7_LC_29_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88726),
            .lcout(shift_srl_75Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93415),
            .ce(N__88701),
            .sr(_gnd_net_));
    defparam shift_srl_75_6_LC_29_10_4.C_ON=1'b0;
    defparam shift_srl_75_6_LC_29_10_4.SEQ_MODE=4'b1000;
    defparam shift_srl_75_6_LC_29_10_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_75_6_LC_29_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88720),
            .lcout(shift_srl_75Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93415),
            .ce(N__88701),
            .sr(_gnd_net_));
    defparam shift_srl_75_5_LC_29_10_5.C_ON=1'b0;
    defparam shift_srl_75_5_LC_29_10_5.SEQ_MODE=4'b1000;
    defparam shift_srl_75_5_LC_29_10_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_75_5_LC_29_10_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88708),
            .lcout(shift_srl_75Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93415),
            .ce(N__88701),
            .sr(_gnd_net_));
    defparam shift_srl_75_4_LC_29_10_6.C_ON=1'b0;
    defparam shift_srl_75_4_LC_29_10_6.SEQ_MODE=4'b1000;
    defparam shift_srl_75_4_LC_29_10_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_75_4_LC_29_10_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88714),
            .lcout(shift_srl_75Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93415),
            .ce(N__88701),
            .sr(_gnd_net_));
    defparam shift_srl_74_0_LC_29_11_0.C_ON=1'b0;
    defparam shift_srl_74_0_LC_29_11_0.SEQ_MODE=4'b1000;
    defparam shift_srl_74_0_LC_29_11_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_74_0_LC_29_11_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88912),
            .lcout(shift_srl_74Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93408),
            .ce(N__88881),
            .sr(_gnd_net_));
    defparam shift_srl_74_1_LC_29_11_1.C_ON=1'b0;
    defparam shift_srl_74_1_LC_29_11_1.SEQ_MODE=4'b1000;
    defparam shift_srl_74_1_LC_29_11_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_74_1_LC_29_11_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88666),
            .lcout(shift_srl_74Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93408),
            .ce(N__88881),
            .sr(_gnd_net_));
    defparam shift_srl_74_2_LC_29_11_2.C_ON=1'b0;
    defparam shift_srl_74_2_LC_29_11_2.SEQ_MODE=4'b1000;
    defparam shift_srl_74_2_LC_29_11_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_74_2_LC_29_11_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88660),
            .lcout(shift_srl_74Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93408),
            .ce(N__88881),
            .sr(_gnd_net_));
    defparam shift_srl_74_3_LC_29_11_3.C_ON=1'b0;
    defparam shift_srl_74_3_LC_29_11_3.SEQ_MODE=4'b1000;
    defparam shift_srl_74_3_LC_29_11_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_74_3_LC_29_11_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88792),
            .lcout(shift_srl_74Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93408),
            .ce(N__88881),
            .sr(_gnd_net_));
    defparam shift_srl_74_4_LC_29_11_4.C_ON=1'b0;
    defparam shift_srl_74_4_LC_29_11_4.SEQ_MODE=4'b1000;
    defparam shift_srl_74_4_LC_29_11_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_74_4_LC_29_11_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88786),
            .lcout(shift_srl_74Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93408),
            .ce(N__88881),
            .sr(_gnd_net_));
    defparam shift_srl_74_5_LC_29_11_5.C_ON=1'b0;
    defparam shift_srl_74_5_LC_29_11_5.SEQ_MODE=4'b1000;
    defparam shift_srl_74_5_LC_29_11_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_74_5_LC_29_11_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88780),
            .lcout(shift_srl_74Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93408),
            .ce(N__88881),
            .sr(_gnd_net_));
    defparam shift_srl_74_6_LC_29_11_6.C_ON=1'b0;
    defparam shift_srl_74_6_LC_29_11_6.SEQ_MODE=4'b1000;
    defparam shift_srl_74_6_LC_29_11_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_74_6_LC_29_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88774),
            .lcout(shift_srl_74Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93408),
            .ce(N__88881),
            .sr(_gnd_net_));
    defparam shift_srl_74_7_LC_29_11_7.C_ON=1'b0;
    defparam shift_srl_74_7_LC_29_11_7.SEQ_MODE=4'b1000;
    defparam shift_srl_74_7_LC_29_11_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_74_7_LC_29_11_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88768),
            .lcout(shift_srl_74Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93408),
            .ce(N__88881),
            .sr(_gnd_net_));
    defparam shift_srl_74_10_LC_29_12_0.C_ON=1'b0;
    defparam shift_srl_74_10_LC_29_12_0.SEQ_MODE=4'b1000;
    defparam shift_srl_74_10_LC_29_12_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_74_10_LC_29_12_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88900),
            .lcout(shift_srl_74Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93400),
            .ce(N__88882),
            .sr(_gnd_net_));
    defparam shift_srl_74_11_LC_29_12_1.C_ON=1'b0;
    defparam shift_srl_74_11_LC_29_12_1.SEQ_MODE=4'b1000;
    defparam shift_srl_74_11_LC_29_12_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_74_11_LC_29_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88762),
            .lcout(shift_srl_74Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93400),
            .ce(N__88882),
            .sr(_gnd_net_));
    defparam shift_srl_74_12_LC_29_12_2.C_ON=1'b0;
    defparam shift_srl_74_12_LC_29_12_2.SEQ_MODE=4'b1000;
    defparam shift_srl_74_12_LC_29_12_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_74_12_LC_29_12_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88756),
            .lcout(shift_srl_74Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93400),
            .ce(N__88882),
            .sr(_gnd_net_));
    defparam shift_srl_74_13_LC_29_12_3.C_ON=1'b0;
    defparam shift_srl_74_13_LC_29_12_3.SEQ_MODE=4'b1000;
    defparam shift_srl_74_13_LC_29_12_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_74_13_LC_29_12_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88750),
            .lcout(shift_srl_74Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93400),
            .ce(N__88882),
            .sr(_gnd_net_));
    defparam shift_srl_74_14_LC_29_12_4.C_ON=1'b0;
    defparam shift_srl_74_14_LC_29_12_4.SEQ_MODE=4'b1000;
    defparam shift_srl_74_14_LC_29_12_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_74_14_LC_29_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88924),
            .lcout(shift_srl_74Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93400),
            .ce(N__88882),
            .sr(_gnd_net_));
    defparam shift_srl_74_15_LC_29_12_5.C_ON=1'b0;
    defparam shift_srl_74_15_LC_29_12_5.SEQ_MODE=4'b1000;
    defparam shift_srl_74_15_LC_29_12_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_74_15_LC_29_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88918),
            .lcout(shift_srl_74Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93400),
            .ce(N__88882),
            .sr(_gnd_net_));
    defparam shift_srl_74_9_LC_29_12_6.C_ON=1'b0;
    defparam shift_srl_74_9_LC_29_12_6.SEQ_MODE=4'b1000;
    defparam shift_srl_74_9_LC_29_12_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_74_9_LC_29_12_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88888),
            .lcout(shift_srl_74Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93400),
            .ce(N__88882),
            .sr(_gnd_net_));
    defparam shift_srl_74_8_LC_29_12_7.C_ON=1'b0;
    defparam shift_srl_74_8_LC_29_12_7.SEQ_MODE=4'b1000;
    defparam shift_srl_74_8_LC_29_12_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_74_8_LC_29_12_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88894),
            .lcout(shift_srl_74Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93400),
            .ce(N__88882),
            .sr(_gnd_net_));
    defparam shift_srl_32_7_LC_29_17_0.C_ON=1'b0;
    defparam shift_srl_32_7_LC_29_17_0.SEQ_MODE=4'b1000;
    defparam shift_srl_32_7_LC_29_17_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_32_7_LC_29_17_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88864),
            .lcout(shift_srl_32Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93299),
            .ce(N__88833),
            .sr(_gnd_net_));
    defparam shift_srl_32_6_LC_29_17_1.C_ON=1'b0;
    defparam shift_srl_32_6_LC_29_17_1.SEQ_MODE=4'b1000;
    defparam shift_srl_32_6_LC_29_17_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_32_6_LC_29_17_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88852),
            .lcout(shift_srl_32Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93299),
            .ce(N__88833),
            .sr(_gnd_net_));
    defparam shift_srl_32_4_LC_29_17_4.C_ON=1'b0;
    defparam shift_srl_32_4_LC_29_17_4.SEQ_MODE=4'b1000;
    defparam shift_srl_32_4_LC_29_17_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_32_4_LC_29_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88840),
            .lcout(shift_srl_32Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93299),
            .ce(N__88833),
            .sr(_gnd_net_));
    defparam shift_srl_32_5_LC_29_17_6.C_ON=1'b0;
    defparam shift_srl_32_5_LC_29_17_6.SEQ_MODE=4'b1000;
    defparam shift_srl_32_5_LC_29_17_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_32_5_LC_29_17_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88858),
            .lcout(shift_srl_32Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93299),
            .ce(N__88833),
            .sr(_gnd_net_));
    defparam shift_srl_32_3_LC_29_18_5.C_ON=1'b0;
    defparam shift_srl_32_3_LC_29_18_5.SEQ_MODE=4'b1000;
    defparam shift_srl_32_3_LC_29_18_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_32_3_LC_29_18_5 (
            .in0(N__88846),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_32Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93341),
            .ce(N__88832),
            .sr(_gnd_net_));
    defparam shift_srl_172_10_LC_29_19_0.C_ON=1'b0;
    defparam shift_srl_172_10_LC_29_19_0.SEQ_MODE=4'b1000;
    defparam shift_srl_172_10_LC_29_19_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_172_10_LC_29_19_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88957),
            .lcout(shift_srl_172Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93362),
            .ce(N__89005),
            .sr(_gnd_net_));
    defparam shift_srl_172_11_LC_29_19_1.C_ON=1'b0;
    defparam shift_srl_172_11_LC_29_19_1.SEQ_MODE=4'b1000;
    defparam shift_srl_172_11_LC_29_19_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_172_11_LC_29_19_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88987),
            .lcout(shift_srl_172Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93362),
            .ce(N__89005),
            .sr(_gnd_net_));
    defparam shift_srl_172_12_LC_29_19_2.C_ON=1'b0;
    defparam shift_srl_172_12_LC_29_19_2.SEQ_MODE=4'b1000;
    defparam shift_srl_172_12_LC_29_19_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_172_12_LC_29_19_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88981),
            .lcout(shift_srl_172Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93362),
            .ce(N__89005),
            .sr(_gnd_net_));
    defparam shift_srl_172_13_LC_29_19_3.C_ON=1'b0;
    defparam shift_srl_172_13_LC_29_19_3.SEQ_MODE=4'b1000;
    defparam shift_srl_172_13_LC_29_19_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_172_13_LC_29_19_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88975),
            .lcout(shift_srl_172Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93362),
            .ce(N__89005),
            .sr(_gnd_net_));
    defparam shift_srl_172_14_LC_29_19_4.C_ON=1'b0;
    defparam shift_srl_172_14_LC_29_19_4.SEQ_MODE=4'b1000;
    defparam shift_srl_172_14_LC_29_19_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_172_14_LC_29_19_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88969),
            .lcout(shift_srl_172Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93362),
            .ce(N__89005),
            .sr(_gnd_net_));
    defparam shift_srl_172_15_LC_29_19_5.C_ON=1'b0;
    defparam shift_srl_172_15_LC_29_19_5.SEQ_MODE=4'b1000;
    defparam shift_srl_172_15_LC_29_19_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_172_15_LC_29_19_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88963),
            .lcout(shift_srl_172Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93362),
            .ce(N__89005),
            .sr(_gnd_net_));
    defparam shift_srl_172_9_LC_29_19_6.C_ON=1'b0;
    defparam shift_srl_172_9_LC_29_19_6.SEQ_MODE=4'b1000;
    defparam shift_srl_172_9_LC_29_19_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_172_9_LC_29_19_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88951),
            .lcout(shift_srl_172Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93362),
            .ce(N__89005),
            .sr(_gnd_net_));
    defparam shift_srl_172_8_LC_29_19_7.C_ON=1'b0;
    defparam shift_srl_172_8_LC_29_19_7.SEQ_MODE=4'b1000;
    defparam shift_srl_172_8_LC_29_19_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_172_8_LC_29_19_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__89011),
            .lcout(shift_srl_172Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93362),
            .ce(N__89005),
            .sr(_gnd_net_));
    defparam shift_srl_172_0_LC_29_20_0.C_ON=1'b0;
    defparam shift_srl_172_0_LC_29_20_0.SEQ_MODE=4'b1000;
    defparam shift_srl_172_0_LC_29_20_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_172_0_LC_29_20_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88938),
            .lcout(shift_srl_172Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93379),
            .ce(N__89004),
            .sr(_gnd_net_));
    defparam shift_srl_172_1_LC_29_20_1.C_ON=1'b0;
    defparam shift_srl_172_1_LC_29_20_1.SEQ_MODE=4'b1000;
    defparam shift_srl_172_1_LC_29_20_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_172_1_LC_29_20_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__89053),
            .lcout(shift_srl_172Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93379),
            .ce(N__89004),
            .sr(_gnd_net_));
    defparam shift_srl_172_2_LC_29_20_2.C_ON=1'b0;
    defparam shift_srl_172_2_LC_29_20_2.SEQ_MODE=4'b1000;
    defparam shift_srl_172_2_LC_29_20_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_172_2_LC_29_20_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__89047),
            .lcout(shift_srl_172Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93379),
            .ce(N__89004),
            .sr(_gnd_net_));
    defparam shift_srl_172_3_LC_29_20_3.C_ON=1'b0;
    defparam shift_srl_172_3_LC_29_20_3.SEQ_MODE=4'b1000;
    defparam shift_srl_172_3_LC_29_20_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_172_3_LC_29_20_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__89041),
            .lcout(shift_srl_172Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93379),
            .ce(N__89004),
            .sr(_gnd_net_));
    defparam shift_srl_172_4_LC_29_20_4.C_ON=1'b0;
    defparam shift_srl_172_4_LC_29_20_4.SEQ_MODE=4'b1000;
    defparam shift_srl_172_4_LC_29_20_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_172_4_LC_29_20_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__89035),
            .lcout(shift_srl_172Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93379),
            .ce(N__89004),
            .sr(_gnd_net_));
    defparam shift_srl_172_5_LC_29_20_5.C_ON=1'b0;
    defparam shift_srl_172_5_LC_29_20_5.SEQ_MODE=4'b1000;
    defparam shift_srl_172_5_LC_29_20_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_172_5_LC_29_20_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__89029),
            .lcout(shift_srl_172Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93379),
            .ce(N__89004),
            .sr(_gnd_net_));
    defparam shift_srl_172_6_LC_29_20_6.C_ON=1'b0;
    defparam shift_srl_172_6_LC_29_20_6.SEQ_MODE=4'b1000;
    defparam shift_srl_172_6_LC_29_20_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_172_6_LC_29_20_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__89023),
            .lcout(shift_srl_172Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93379),
            .ce(N__89004),
            .sr(_gnd_net_));
    defparam shift_srl_172_7_LC_29_20_7.C_ON=1'b0;
    defparam shift_srl_172_7_LC_29_20_7.SEQ_MODE=4'b1000;
    defparam shift_srl_172_7_LC_29_20_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_172_7_LC_29_20_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__89017),
            .lcout(shift_srl_172Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93379),
            .ce(N__89004),
            .sr(_gnd_net_));
    defparam shift_srl_168_13_LC_29_21_0.C_ON=1'b0;
    defparam shift_srl_168_13_LC_29_21_0.SEQ_MODE=4'b1000;
    defparam shift_srl_168_13_LC_29_21_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_168_13_LC_29_21_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__89146),
            .lcout(shift_srl_168Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93394),
            .ce(N__89106),
            .sr(_gnd_net_));
    defparam shift_srl_168_9_LC_29_21_3.C_ON=1'b0;
    defparam shift_srl_168_9_LC_29_21_3.SEQ_MODE=4'b1000;
    defparam shift_srl_168_9_LC_29_21_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_168_9_LC_29_21_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__89134),
            .lcout(shift_srl_168Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93394),
            .ce(N__89106),
            .sr(_gnd_net_));
    defparam shift_srl_168_14_LC_29_21_4.C_ON=1'b0;
    defparam shift_srl_168_14_LC_29_21_4.SEQ_MODE=4'b1000;
    defparam shift_srl_168_14_LC_29_21_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_168_14_LC_29_21_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88993),
            .lcout(shift_srl_168Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93394),
            .ce(N__89106),
            .sr(_gnd_net_));
    defparam shift_srl_168_15_LC_29_21_5.C_ON=1'b0;
    defparam shift_srl_168_15_LC_29_21_5.SEQ_MODE=4'b1000;
    defparam shift_srl_168_15_LC_29_21_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_168_15_LC_29_21_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__89188),
            .lcout(shift_srl_168Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93394),
            .ce(N__89106),
            .sr(_gnd_net_));
    defparam shift_srl_168_12_LC_29_21_6.C_ON=1'b0;
    defparam shift_srl_168_12_LC_29_21_6.SEQ_MODE=4'b1000;
    defparam shift_srl_168_12_LC_29_21_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_168_12_LC_29_21_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__89116),
            .lcout(shift_srl_168Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93394),
            .ce(N__89106),
            .sr(_gnd_net_));
    defparam shift_srl_168_8_LC_29_21_7.C_ON=1'b0;
    defparam shift_srl_168_8_LC_29_21_7.SEQ_MODE=4'b1000;
    defparam shift_srl_168_8_LC_29_21_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_168_8_LC_29_21_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__89140),
            .lcout(shift_srl_168Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93394),
            .ce(N__89106),
            .sr(_gnd_net_));
    defparam shift_srl_168_10_LC_29_22_3.C_ON=1'b0;
    defparam shift_srl_168_10_LC_29_22_3.SEQ_MODE=4'b1000;
    defparam shift_srl_168_10_LC_29_22_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_srl_168_10_LC_29_22_3 (
            .in0(N__89128),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_srl_168Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93401),
            .ce(N__89104),
            .sr(_gnd_net_));
    defparam shift_srl_168_11_LC_29_23_2.C_ON=1'b0;
    defparam shift_srl_168_11_LC_29_23_2.SEQ_MODE=4'b1000;
    defparam shift_srl_168_11_LC_29_23_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_168_11_LC_29_23_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__89122),
            .lcout(shift_srl_168Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93409),
            .ce(N__89107),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_72_LC_30_9_0.C_ON=1'b0;
    defparam rco_obuf_RNO_72_LC_30_9_0.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_72_LC_30_9_0.LUT_INIT=16'b1000100000000000;
    LogicCell40 rco_obuf_RNO_72_LC_30_9_0 (
            .in0(N__90786),
            .in1(N__90734),
            .in2(_gnd_net_),
            .in3(N__90847),
            .lcout(rco_c_72),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_73_10_LC_30_10_0.C_ON=1'b0;
    defparam shift_srl_73_10_LC_30_10_0.SEQ_MODE=4'b1000;
    defparam shift_srl_73_10_LC_30_10_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_73_10_LC_30_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__90598),
            .lcout(shift_srl_73Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93420),
            .ce(N__90997),
            .sr(_gnd_net_));
    defparam shift_srl_73_11_LC_30_10_1.C_ON=1'b0;
    defparam shift_srl_73_11_LC_30_10_1.SEQ_MODE=4'b1000;
    defparam shift_srl_73_11_LC_30_10_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_73_11_LC_30_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__89059),
            .lcout(shift_srl_73Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93420),
            .ce(N__90997),
            .sr(_gnd_net_));
    defparam shift_srl_73_12_LC_30_10_2.C_ON=1'b0;
    defparam shift_srl_73_12_LC_30_10_2.SEQ_MODE=4'b1000;
    defparam shift_srl_73_12_LC_30_10_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_73_12_LC_30_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__90622),
            .lcout(shift_srl_73Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93420),
            .ce(N__90997),
            .sr(_gnd_net_));
    defparam shift_srl_73_13_LC_30_10_3.C_ON=1'b0;
    defparam shift_srl_73_13_LC_30_10_3.SEQ_MODE=4'b1000;
    defparam shift_srl_73_13_LC_30_10_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_73_13_LC_30_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__90616),
            .lcout(shift_srl_73Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93420),
            .ce(N__90997),
            .sr(_gnd_net_));
    defparam shift_srl_73_14_LC_30_10_4.C_ON=1'b0;
    defparam shift_srl_73_14_LC_30_10_4.SEQ_MODE=4'b1000;
    defparam shift_srl_73_14_LC_30_10_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_73_14_LC_30_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__90610),
            .lcout(shift_srl_73Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93420),
            .ce(N__90997),
            .sr(_gnd_net_));
    defparam shift_srl_73_15_LC_30_10_5.C_ON=1'b0;
    defparam shift_srl_73_15_LC_30_10_5.SEQ_MODE=4'b1000;
    defparam shift_srl_73_15_LC_30_10_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_73_15_LC_30_10_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__90604),
            .lcout(shift_srl_73Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93420),
            .ce(N__90997),
            .sr(_gnd_net_));
    defparam shift_srl_73_9_LC_30_10_6.C_ON=1'b0;
    defparam shift_srl_73_9_LC_30_10_6.SEQ_MODE=4'b1000;
    defparam shift_srl_73_9_LC_30_10_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_73_9_LC_30_10_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__90592),
            .lcout(shift_srl_73Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93420),
            .ce(N__90997),
            .sr(_gnd_net_));
    defparam shift_srl_73_8_LC_30_10_7.C_ON=1'b0;
    defparam shift_srl_73_8_LC_30_10_7.SEQ_MODE=4'b1000;
    defparam shift_srl_73_8_LC_30_10_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_73_8_LC_30_10_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__91006),
            .lcout(shift_srl_73Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93420),
            .ce(N__90997),
            .sr(_gnd_net_));
    defparam shift_srl_72_RNIMGABI_15_LC_30_11_6.C_ON=1'b0;
    defparam shift_srl_72_RNIMGABI_15_LC_30_11_6.SEQ_MODE=4'b0000;
    defparam shift_srl_72_RNIMGABI_15_LC_30_11_6.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_srl_72_RNIMGABI_15_LC_30_11_6 (
            .in0(N__90292),
            .in1(N__90693),
            .in2(N__90785),
            .in3(N__90839),
            .lcout(clk_en_73),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_73_0_LC_30_12_0.C_ON=1'b0;
    defparam shift_srl_73_0_LC_30_12_0.SEQ_MODE=4'b1000;
    defparam shift_srl_73_0_LC_30_12_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_73_0_LC_30_12_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__90875),
            .lcout(shift_srl_73Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93410),
            .ce(N__90996),
            .sr(_gnd_net_));
    defparam shift_srl_73_1_LC_30_12_1.C_ON=1'b0;
    defparam shift_srl_73_1_LC_30_12_1.SEQ_MODE=4'b1000;
    defparam shift_srl_73_1_LC_30_12_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_73_1_LC_30_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__89200),
            .lcout(shift_srl_73Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93410),
            .ce(N__90996),
            .sr(_gnd_net_));
    defparam shift_srl_73_2_LC_30_12_2.C_ON=1'b0;
    defparam shift_srl_73_2_LC_30_12_2.SEQ_MODE=4'b1000;
    defparam shift_srl_73_2_LC_30_12_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_73_2_LC_30_12_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__89194),
            .lcout(shift_srl_73Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93410),
            .ce(N__90996),
            .sr(_gnd_net_));
    defparam shift_srl_73_3_LC_30_12_3.C_ON=1'b0;
    defparam shift_srl_73_3_LC_30_12_3.SEQ_MODE=4'b1000;
    defparam shift_srl_73_3_LC_30_12_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_73_3_LC_30_12_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__91036),
            .lcout(shift_srl_73Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93410),
            .ce(N__90996),
            .sr(_gnd_net_));
    defparam shift_srl_73_4_LC_30_12_4.C_ON=1'b0;
    defparam shift_srl_73_4_LC_30_12_4.SEQ_MODE=4'b1000;
    defparam shift_srl_73_4_LC_30_12_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_73_4_LC_30_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__91030),
            .lcout(shift_srl_73Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93410),
            .ce(N__90996),
            .sr(_gnd_net_));
    defparam shift_srl_73_5_LC_30_12_5.C_ON=1'b0;
    defparam shift_srl_73_5_LC_30_12_5.SEQ_MODE=4'b1000;
    defparam shift_srl_73_5_LC_30_12_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_73_5_LC_30_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__91024),
            .lcout(shift_srl_73Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93410),
            .ce(N__90996),
            .sr(_gnd_net_));
    defparam shift_srl_73_6_LC_30_12_6.C_ON=1'b0;
    defparam shift_srl_73_6_LC_30_12_6.SEQ_MODE=4'b1000;
    defparam shift_srl_73_6_LC_30_12_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_73_6_LC_30_12_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__91018),
            .lcout(shift_srl_73Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93410),
            .ce(N__90996),
            .sr(_gnd_net_));
    defparam shift_srl_73_7_LC_30_12_7.C_ON=1'b0;
    defparam shift_srl_73_7_LC_30_12_7.SEQ_MODE=4'b1000;
    defparam shift_srl_73_7_LC_30_12_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_73_7_LC_30_12_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__91012),
            .lcout(shift_srl_73Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93410),
            .ce(N__90996),
            .sr(_gnd_net_));
    defparam shift_srl_36_14_LC_30_21_2.C_ON=1'b0;
    defparam shift_srl_36_14_LC_30_21_2.SEQ_MODE=4'b1000;
    defparam shift_srl_36_14_LC_30_21_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_36_14_LC_30_21_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__90976),
            .lcout(shift_srl_36Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93402),
            .ce(N__90943),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_73_LC_31_9_1.C_ON=1'b0;
    defparam rco_obuf_RNO_73_LC_31_9_1.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_73_LC_31_9_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 rco_obuf_RNO_73_LC_31_9_1 (
            .in0(N__90869),
            .in1(N__90787),
            .in2(N__90739),
            .in3(N__90846),
            .lcout(rco_c_73),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_71_LC_31_10_2.C_ON=1'b0;
    defparam rco_obuf_RNO_71_LC_31_10_2.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_71_LC_31_10_2.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_71_LC_31_10_2 (
            .in0(N__90775),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__90733),
            .lcout(rco_c_71),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_srl_37_11_LC_31_17_0.C_ON=1'b0;
    defparam shift_srl_37_11_LC_31_17_0.SEQ_MODE=4'b1000;
    defparam shift_srl_37_11_LC_31_17_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_srl_37_11_LC_31_17_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__93445),
            .lcout(shift_srl_37Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93342),
            .ce(N__91858),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_186_LC_31_21_4.C_ON=1'b0;
    defparam rco_obuf_RNO_186_LC_31_21_4.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_186_LC_31_21_4.LUT_INIT=16'b1000000000000000;
    LogicCell40 rco_obuf_RNO_186_LC_31_21_4 (
            .in0(N__91699),
            .in1(N__91825),
            .in2(N__91768),
            .in3(N__91539),
            .lcout(rco_c_186),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_185_LC_31_22_5.C_ON=1'b0;
    defparam rco_obuf_RNO_185_LC_31_22_5.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_185_LC_31_22_5.LUT_INIT=16'b1000100000000000;
    LogicCell40 rco_obuf_RNO_185_LC_31_22_5 (
            .in0(N__91763),
            .in1(N__91698),
            .in2(_gnd_net_),
            .in3(N__91537),
            .lcout(rco_c_185),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_190_LC_31_22_7.C_ON=1'b0;
    defparam rco_obuf_RNO_190_LC_31_22_7.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_190_LC_31_22_7.LUT_INIT=16'b1000100000000000;
    LogicCell40 rco_obuf_RNO_190_LC_31_22_7 (
            .in0(N__91612),
            .in1(N__91570),
            .in2(_gnd_net_),
            .in3(N__91538),
            .lcout(rco_c_190),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_189_LC_31_23_1.C_ON=1'b0;
    defparam rco_obuf_RNO_189_LC_31_23_1.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_189_LC_31_23_1.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_189_LC_31_23_1 (
            .in0(N__91566),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__91527),
            .lcout(rco_c_189),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_129_LC_31_24_3.C_ON=1'b0;
    defparam rco_obuf_RNO_129_LC_31_24_3.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_129_LC_31_24_3.LUT_INIT=16'b1100110000000000;
    LogicCell40 rco_obuf_RNO_129_LC_31_24_3 (
            .in0(_gnd_net_),
            .in1(N__91306),
            .in2(_gnd_net_),
            .in3(N__91387),
            .lcout(rco_c_129),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_128_LC_31_25_1.C_ON=1'b0;
    defparam rco_obuf_RNO_128_LC_31_25_1.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_128_LC_31_25_1.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_128_LC_31_25_1 (
            .in0(N__91325),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__91276),
            .lcout(rco_c_128),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_140_LC_31_27_7.C_ON=1'b0;
    defparam rco_obuf_RNO_140_LC_31_27_7.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_140_LC_31_27_7.LUT_INIT=16'b1010101000000000;
    LogicCell40 rco_obuf_RNO_140_LC_31_27_7 (
            .in0(N__91162),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__91113),
            .lcout(N_125_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rco_obuf_RNO_49_LC_32_7_2.C_ON=1'b0;
    defparam rco_obuf_RNO_49_LC_32_7_2.SEQ_MODE=4'b0000;
    defparam rco_obuf_RNO_49_LC_32_7_2.LUT_INIT=16'b1100110000000000;
    LogicCell40 rco_obuf_RNO_49_LC_32_7_2 (
            .in0(_gnd_net_),
            .in1(N__93603),
            .in2(_gnd_net_),
            .in3(N__93499),
            .lcout(rco_c_49),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // big_counter
