module pudc_and2(
    input a,
    input b,
    output o
);

assign o = a & b;

endmodule