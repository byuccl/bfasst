// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 12 2017 08:25:46

// File Generated:     Jan 24 2019 13:19:30

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "bcd_adder" view "INTERFACE"

module bcd_adder (
    sum_o,
    a_i,
    b_i,
    cout_o,
    clk_i,
    cin_i);

    output [15:0] sum_o;
    input [15:0] a_i;
    input [15:0] b_i;
    output cout_o;
    input clk_i;
    input cin_i;

    wire N__3728;
    wire N__3727;
    wire N__3726;
    wire N__3717;
    wire N__3716;
    wire N__3715;
    wire N__3708;
    wire N__3707;
    wire N__3706;
    wire N__3699;
    wire N__3698;
    wire N__3697;
    wire N__3690;
    wire N__3689;
    wire N__3688;
    wire N__3681;
    wire N__3680;
    wire N__3679;
    wire N__3672;
    wire N__3671;
    wire N__3670;
    wire N__3663;
    wire N__3662;
    wire N__3661;
    wire N__3654;
    wire N__3653;
    wire N__3652;
    wire N__3645;
    wire N__3644;
    wire N__3643;
    wire N__3636;
    wire N__3635;
    wire N__3634;
    wire N__3627;
    wire N__3626;
    wire N__3625;
    wire N__3618;
    wire N__3617;
    wire N__3616;
    wire N__3609;
    wire N__3608;
    wire N__3607;
    wire N__3600;
    wire N__3599;
    wire N__3598;
    wire N__3591;
    wire N__3590;
    wire N__3589;
    wire N__3582;
    wire N__3581;
    wire N__3580;
    wire N__3573;
    wire N__3572;
    wire N__3571;
    wire N__3564;
    wire N__3563;
    wire N__3562;
    wire N__3555;
    wire N__3554;
    wire N__3553;
    wire N__3546;
    wire N__3545;
    wire N__3544;
    wire N__3537;
    wire N__3536;
    wire N__3535;
    wire N__3528;
    wire N__3527;
    wire N__3526;
    wire N__3519;
    wire N__3518;
    wire N__3517;
    wire N__3510;
    wire N__3509;
    wire N__3508;
    wire N__3501;
    wire N__3500;
    wire N__3499;
    wire N__3492;
    wire N__3491;
    wire N__3490;
    wire N__3483;
    wire N__3482;
    wire N__3481;
    wire N__3474;
    wire N__3473;
    wire N__3472;
    wire N__3465;
    wire N__3464;
    wire N__3463;
    wire N__3456;
    wire N__3455;
    wire N__3454;
    wire N__3447;
    wire N__3446;
    wire N__3445;
    wire N__3438;
    wire N__3437;
    wire N__3436;
    wire N__3429;
    wire N__3428;
    wire N__3427;
    wire N__3420;
    wire N__3419;
    wire N__3418;
    wire N__3411;
    wire N__3410;
    wire N__3409;
    wire N__3402;
    wire N__3401;
    wire N__3400;
    wire N__3393;
    wire N__3392;
    wire N__3391;
    wire N__3384;
    wire N__3383;
    wire N__3382;
    wire N__3375;
    wire N__3374;
    wire N__3373;
    wire N__3366;
    wire N__3365;
    wire N__3364;
    wire N__3357;
    wire N__3356;
    wire N__3355;
    wire N__3348;
    wire N__3347;
    wire N__3346;
    wire N__3339;
    wire N__3338;
    wire N__3337;
    wire N__3330;
    wire N__3329;
    wire N__3328;
    wire N__3321;
    wire N__3320;
    wire N__3319;
    wire N__3312;
    wire N__3311;
    wire N__3310;
    wire N__3303;
    wire N__3302;
    wire N__3301;
    wire N__3294;
    wire N__3293;
    wire N__3292;
    wire N__3285;
    wire N__3284;
    wire N__3283;
    wire N__3276;
    wire N__3275;
    wire N__3274;
    wire N__3257;
    wire N__3254;
    wire N__3251;
    wire N__3248;
    wire N__3245;
    wire N__3242;
    wire N__3241;
    wire N__3240;
    wire N__3235;
    wire N__3232;
    wire N__3227;
    wire N__3224;
    wire N__3221;
    wire N__3218;
    wire N__3215;
    wire N__3212;
    wire N__3211;
    wire N__3208;
    wire N__3205;
    wire N__3200;
    wire N__3197;
    wire N__3194;
    wire N__3191;
    wire N__3188;
    wire N__3185;
    wire N__3182;
    wire N__3179;
    wire N__3176;
    wire N__3173;
    wire N__3170;
    wire N__3167;
    wire N__3164;
    wire N__3163;
    wire N__3158;
    wire N__3155;
    wire N__3154;
    wire N__3153;
    wire N__3152;
    wire N__3151;
    wire N__3150;
    wire N__3149;
    wire N__3148;
    wire N__3147;
    wire N__3146;
    wire N__3145;
    wire N__3144;
    wire N__3119;
    wire N__3116;
    wire N__3113;
    wire N__3110;
    wire N__3107;
    wire N__3104;
    wire N__3101;
    wire N__3098;
    wire N__3095;
    wire N__3092;
    wire N__3089;
    wire N__3086;
    wire N__3083;
    wire N__3080;
    wire N__3077;
    wire N__3074;
    wire N__3071;
    wire N__3068;
    wire N__3065;
    wire N__3062;
    wire N__3061;
    wire N__3060;
    wire N__3057;
    wire N__3052;
    wire N__3049;
    wire N__3046;
    wire N__3043;
    wire N__3038;
    wire N__3035;
    wire N__3032;
    wire N__3029;
    wire N__3026;
    wire N__3023;
    wire N__3020;
    wire N__3017;
    wire N__3014;
    wire N__3013;
    wire N__3010;
    wire N__3007;
    wire N__3004;
    wire N__3001;
    wire N__2996;
    wire N__2995;
    wire N__2992;
    wire N__2989;
    wire N__2986;
    wire N__2983;
    wire N__2978;
    wire N__2975;
    wire N__2972;
    wire N__2969;
    wire N__2966;
    wire N__2965;
    wire N__2962;
    wire N__2959;
    wire N__2954;
    wire N__2951;
    wire N__2948;
    wire N__2945;
    wire N__2944;
    wire N__2941;
    wire N__2938;
    wire N__2935;
    wire N__2930;
    wire N__2927;
    wire N__2924;
    wire N__2921;
    wire N__2920;
    wire N__2919;
    wire N__2916;
    wire N__2913;
    wire N__2910;
    wire N__2907;
    wire N__2902;
    wire N__2897;
    wire N__2894;
    wire N__2891;
    wire N__2888;
    wire N__2885;
    wire N__2882;
    wire N__2879;
    wire N__2876;
    wire N__2875;
    wire N__2874;
    wire N__2871;
    wire N__2866;
    wire N__2861;
    wire N__2860;
    wire N__2859;
    wire N__2856;
    wire N__2853;
    wire N__2850;
    wire N__2847;
    wire N__2840;
    wire N__2837;
    wire N__2836;
    wire N__2833;
    wire N__2830;
    wire N__2825;
    wire N__2822;
    wire N__2819;
    wire N__2816;
    wire N__2813;
    wire N__2810;
    wire N__2807;
    wire N__2804;
    wire N__2801;
    wire N__2798;
    wire N__2797;
    wire N__2794;
    wire N__2793;
    wire N__2790;
    wire N__2787;
    wire N__2784;
    wire N__2781;
    wire N__2774;
    wire N__2771;
    wire N__2770;
    wire N__2769;
    wire N__2766;
    wire N__2763;
    wire N__2760;
    wire N__2753;
    wire N__2752;
    wire N__2751;
    wire N__2748;
    wire N__2745;
    wire N__2742;
    wire N__2735;
    wire N__2732;
    wire N__2729;
    wire N__2726;
    wire N__2723;
    wire N__2720;
    wire N__2717;
    wire N__2714;
    wire N__2713;
    wire N__2710;
    wire N__2707;
    wire N__2702;
    wire N__2699;
    wire N__2696;
    wire N__2693;
    wire N__2690;
    wire N__2687;
    wire N__2684;
    wire N__2681;
    wire N__2678;
    wire N__2677;
    wire N__2676;
    wire N__2669;
    wire N__2666;
    wire N__2663;
    wire N__2660;
    wire N__2657;
    wire N__2654;
    wire N__2651;
    wire N__2648;
    wire N__2645;
    wire N__2644;
    wire N__2641;
    wire N__2638;
    wire N__2635;
    wire N__2630;
    wire N__2627;
    wire N__2624;
    wire N__2621;
    wire N__2618;
    wire N__2615;
    wire N__2614;
    wire N__2613;
    wire N__2610;
    wire N__2607;
    wire N__2604;
    wire N__2597;
    wire N__2594;
    wire N__2591;
    wire N__2588;
    wire N__2585;
    wire N__2584;
    wire N__2583;
    wire N__2580;
    wire N__2577;
    wire N__2574;
    wire N__2567;
    wire N__2564;
    wire N__2563;
    wire N__2560;
    wire N__2557;
    wire N__2552;
    wire N__2549;
    wire N__2548;
    wire N__2545;
    wire N__2542;
    wire N__2539;
    wire N__2534;
    wire N__2531;
    wire N__2528;
    wire N__2525;
    wire N__2522;
    wire N__2519;
    wire N__2516;
    wire N__2515;
    wire N__2514;
    wire N__2511;
    wire N__2506;
    wire N__2505;
    wire N__2502;
    wire N__2499;
    wire N__2496;
    wire N__2493;
    wire N__2486;
    wire N__2485;
    wire N__2482;
    wire N__2481;
    wire N__2478;
    wire N__2473;
    wire N__2472;
    wire N__2469;
    wire N__2466;
    wire N__2463;
    wire N__2460;
    wire N__2453;
    wire N__2452;
    wire N__2451;
    wire N__2450;
    wire N__2447;
    wire N__2440;
    wire N__2435;
    wire N__2432;
    wire N__2429;
    wire N__2426;
    wire N__2423;
    wire N__2422;
    wire N__2419;
    wire N__2416;
    wire N__2413;
    wire N__2408;
    wire N__2405;
    wire N__2402;
    wire N__2399;
    wire N__2396;
    wire N__2395;
    wire N__2392;
    wire N__2389;
    wire N__2386;
    wire N__2383;
    wire N__2380;
    wire N__2377;
    wire N__2372;
    wire N__2369;
    wire N__2366;
    wire N__2363;
    wire N__2360;
    wire N__2357;
    wire N__2354;
    wire N__2351;
    wire N__2348;
    wire N__2345;
    wire N__2342;
    wire N__2339;
    wire N__2336;
    wire N__2333;
    wire N__2330;
    wire N__2327;
    wire N__2324;
    wire N__2321;
    wire N__2318;
    wire N__2315;
    wire N__2314;
    wire N__2311;
    wire N__2310;
    wire N__2307;
    wire N__2304;
    wire N__2299;
    wire N__2294;
    wire N__2291;
    wire N__2288;
    wire N__2285;
    wire N__2282;
    wire N__2281;
    wire N__2276;
    wire N__2273;
    wire N__2270;
    wire N__2267;
    wire N__2264;
    wire N__2261;
    wire N__2258;
    wire N__2255;
    wire N__2252;
    wire N__2251;
    wire N__2250;
    wire N__2247;
    wire N__2244;
    wire N__2241;
    wire N__2238;
    wire N__2231;
    wire N__2230;
    wire N__2229;
    wire N__2222;
    wire N__2219;
    wire N__2216;
    wire N__2213;
    wire N__2210;
    wire N__2207;
    wire N__2204;
    wire N__2201;
    wire N__2198;
    wire N__2195;
    wire N__2192;
    wire N__2189;
    wire N__2186;
    wire N__2183;
    wire N__2180;
    wire N__2177;
    wire N__2174;
    wire N__2171;
    wire N__2168;
    wire N__2165;
    wire N__2162;
    wire N__2159;
    wire N__2156;
    wire N__2153;
    wire N__2150;
    wire N__2147;
    wire N__2144;
    wire N__2141;
    wire N__2138;
    wire N__2135;
    wire N__2132;
    wire N__2129;
    wire N__2126;
    wire N__2123;
    wire N__2120;
    wire N__2117;
    wire N__2114;
    wire N__2111;
    wire N__2108;
    wire N__2105;
    wire N__2104;
    wire N__2101;
    wire N__2098;
    wire N__2093;
    wire N__2090;
    wire N__2087;
    wire N__2084;
    wire N__2081;
    wire N__2078;
    wire N__2075;
    wire N__2072;
    wire N__2069;
    wire N__2066;
    wire N__2063;
    wire N__2060;
    wire N__2057;
    wire N__2054;
    wire N__2051;
    wire N__2048;
    wire N__2045;
    wire N__2042;
    wire N__2039;
    wire N__2038;
    wire N__2033;
    wire N__2030;
    wire N__2027;
    wire N__2024;
    wire N__2021;
    wire N__2018;
    wire N__2015;
    wire N__2012;
    wire N__2009;
    wire N__2006;
    wire N__2003;
    wire N__2000;
    wire N__1997;
    wire N__1994;
    wire N__1991;
    wire N__1988;
    wire N__1985;
    wire N__1982;
    wire N__1979;
    wire N__1976;
    wire N__1973;
    wire N__1970;
    wire N__1967;
    wire N__1964;
    wire N__1961;
    wire N__1958;
    wire N__1955;
    wire N__1952;
    wire N__1949;
    wire N__1946;
    wire N__1943;
    wire N__1940;
    wire N__1937;
    wire N__1934;
    wire N__1931;
    wire N__1928;
    wire N__1925;
    wire N__1922;
    wire N__1919;
    wire N__1916;
    wire N__1913;
    wire N__1910;
    wire N__1907;
    wire N__1904;
    wire N__1901;
    wire N__1898;
    wire N__1895;
    wire N__1892;
    wire N__1889;
    wire N__1886;
    wire N__1883;
    wire N__1880;
    wire N__1877;
    wire N__1874;
    wire N__1871;
    wire N__1868;
    wire N__1865;
    wire N__1862;
    wire N__1859;
    wire N__1856;
    wire N__1853;
    wire N__1850;
    wire N__1847;
    wire N__1844;
    wire N__1841;
    wire N__1838;
    wire N__1835;
    wire N__1832;
    wire N__1829;
    wire N__1826;
    wire N__1825;
    wire N__1824;
    wire N__1817;
    wire N__1814;
    wire N__1813;
    wire N__1808;
    wire N__1805;
    wire N__1802;
    wire N__1799;
    wire N__1796;
    wire N__1793;
    wire N__1790;
    wire N__1787;
    wire N__1784;
    wire N__1781;
    wire N__1778;
    wire N__1775;
    wire N__1772;
    wire N__1769;
    wire N__1766;
    wire N__1763;
    wire N__1760;
    wire N__1757;
    wire N__1754;
    wire N__1751;
    wire N__1748;
    wire N__1745;
    wire N__1742;
    wire N__1739;
    wire N__1736;
    wire N__1733;
    wire N__1730;
    wire N__1727;
    wire N__1724;
    wire N__1721;
    wire N__1718;
    wire N__1715;
    wire N__1712;
    wire N__1709;
    wire N__1706;
    wire N__1703;
    wire N__1700;
    wire N__1697;
    wire N__1694;
    wire N__1691;
    wire N__1688;
    wire N__1685;
    wire N__1682;
    wire N__1679;
    wire N__1676;
    wire N__1673;
    wire N__1670;
    wire N__1667;
    wire N__1664;
    wire N__1661;
    wire N__1658;
    wire N__1655;
    wire N__1652;
    wire N__1649;
    wire N__1646;
    wire N__1643;
    wire N__1640;
    wire N__1637;
    wire N__1634;
    wire N__1631;
    wire N__1628;
    wire VCCG0;
    wire GNDG0;
    wire a_i_c_15;
    wire b_i_c_4;
    wire a_i_c_14;
    wire b_i_c_14;
    wire b_i_c_0;
    wire b_i_c_13;
    wire a_i_c_9;
    wire b_i_c_15;
    wire sum_o_c_12;
    wire sum_o_c_9;
    wire a_i_c_5;
    wire b_rZ0Z_15;
    wire un68_sum_v_cascade_;
    wire sum_o_c_11;
    wire b_rZ0Z_13;
    wire b_rZ0Z_14;
    wire sum_o_c_10;
    wire sum_o_c_13;
    wire a_i_c_1;
    wire sum_o_c_5;
    wire a_i_c_6;
    wire a_i_c_8;
    wire sum_o_c_14;
    wire sum_o_c_8;
    wire b_i_c_3;
    wire b_rZ0Z_3;
    wire cout_o_c;
    wire b_i_c_8;
    wire b_i_c_2;
    wire b_rZ0Z_2;
    wire a_i_c_11;
    wire a_i_c_12;
    wire b_i_c_12;
    wire b_i_c_11;
    wire b_rZ0Z_11;
    wire m4_0;
    wire b_i_c_10;
    wire cin_i_c;
    wire sum_o_c_3;
    wire sum_o_c_1;
    wire sum_o_c_4;
    wire un13_sum_v;
    wire un13_sum_v_cascade_;
    wire sum_o_c_2;
    wire a_i_c_0;
    wire cin_rZ0;
    wire bfn_2_16_0_;
    wire b_rZ0Z_0;
    wire a_rZ0Z_0;
    wire sum_o_c_0;
    wire un5_sum_v_cry_0_c_THRU_CO;
    wire a_rZ0Z_1;
    wire b_r_i_1;
    wire b_r_sbtinv_RNIB4UQZ0Z_1;
    wire un5_sum_v_cry_0;
    wire b_r_RNILOR9Z0Z_2;
    wire un5_sum_v_cry_1_c_RNIHJLZ0Z01;
    wire un5_sum_v_cry_1;
    wire b_r_RNIKF8BZ0Z_3;
    wire sum_r_RNO_0Z0Z_3;
    wire un5_sum_v_cry_2;
    wire b_rZ0Z_4;
    wire un5_sum_v_cry_3_c_RNIVN8OZ0;
    wire un5_sum_v_cry_3;
    wire a_rZ0Z_5;
    wire un5_sum_v_cry_4;
    wire un5_sum_v_cry_5;
    wire un5_sum_v_cry_6;
    wire bfn_2_17_0_;
    wire un5_sum_v_cry_7;
    wire a_rZ0Z_9;
    wire b_r_sbtinv_RNI357RZ0Z_9;
    wire un5_sum_v_cry_8;
    wire un5_sum_v_cry_9_c_RNIEOBIZ0Z1;
    wire un5_sum_v_cry_9;
    wire a_rZ0Z_11;
    wire b_r_RNI95R61Z0Z_11;
    wire sum_r_RNO_0Z0Z_11;
    wire un5_sum_v_cry_10;
    wire a_rZ0Z_12;
    wire b_rZ0Z_12;
    wire un5_sum_v_cry_11_c_RNICJ0TZ0;
    wire un5_sum_v_cry_11;
    wire b_r_i_13;
    wire un5_sum_v_cry_12;
    wire a_rZ0Z_14;
    wire b_r_RNIEIE51Z0Z_14;
    wire un5_sum_v_cry_13;
    wire un5_sum_v_cry_14;
    wire a_rZ0Z_15;
    wire b_r_RNI0TDJ1Z0Z_15;
    wire bfn_2_18_0_;
    wire un5_sum_v_cry_15;
    wire un5_sum_v_cry_15_THRU_CO;
    wire un5_sum_v_cry_12_c_RNI45JOZ0;
    wire un5_sum_v_cry_13_c_RNIG5IKZ0Z1;
    wire un5_sum_v_cry_15_THRU_CO_cascade_;
    wire sum_r_RNO_0Z0Z_15;
    wire sum_o_c_15;
    wire a_rZ0Z_8;
    wire b_rZ0Z_8;
    wire un5_sum_v_cry_7_c_RNIB8DOZ0;
    wire un40_sum_v_cascade_;
    wire sum_o_c_6;
    wire b_rZ0Z_10;
    wire b_r_RNIRUROZ0Z_10;
    wire b_i_c_1;
    wire b_rZ0Z_1;
    wire b_r_i_9;
    wire a_i_c_10;
    wire a_rZ0Z_10;
    wire b_i_c_9;
    wire b_rZ0Z_9;
    wire a_i_c_7;
    wire a_i_c_13;
    wire a_rZ0Z_13;
    wire a_i_c_4;
    wire a_rZ0Z_4;
    wire b_r_i_5;
    wire a_i_c_2;
    wire a_rZ0Z_2;
    wire a_rZ0Z_7;
    wire b_r_RNI409BZ0Z_7;
    wire a_rZ0Z_6;
    wire b_r_RNI15S9Z0Z_6;
    wire un5_sum_v_cry_5_c_RNI5CQZ0Z01;
    wire sum_r_RNO_0Z0Z_7;
    wire b_r_sbtinv_RNINK2RZ0Z_5;
    wire un40_sum_v;
    wire sum_o_c_7;
    wire b_i_c_5;
    wire b_rZ0Z_5;
    wire a_i_c_3;
    wire a_rZ0Z_3;
    wire b_i_c_7;
    wire b_rZ0Z_7;
    wire b_i_c_6;
    wire b_rZ0Z_6;
    wire clk_i_c_g;
    wire _gnd_net_;

    PRE_IO_GBUF clk_i_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__3726),
            .GLOBALBUFFEROUTPUT(clk_i_c_g));
    IO_PAD clk_i_ibuf_gb_io_iopad (
            .OE(N__3728),
            .DIN(N__3727),
            .DOUT(N__3726),
            .PACKAGEPIN(clk_i));
    defparam clk_i_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam clk_i_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_i_ibuf_gb_io_preio (
            .PADOEN(N__3728),
            .PADOUT(N__3727),
            .PADIN(N__3726),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD a_i_ibuf_0_iopad (
            .OE(N__3717),
            .DIN(N__3716),
            .DOUT(N__3715),
            .PACKAGEPIN(a_i[0]));
    defparam a_i_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam a_i_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO a_i_ibuf_0_preio (
            .PADOEN(N__3717),
            .PADOUT(N__3716),
            .PADIN(N__3715),
            .CLOCKENABLE(),
            .DIN0(a_i_c_0),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD a_i_ibuf_1_iopad (
            .OE(N__3708),
            .DIN(N__3707),
            .DOUT(N__3706),
            .PACKAGEPIN(a_i[1]));
    defparam a_i_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam a_i_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO a_i_ibuf_1_preio (
            .PADOEN(N__3708),
            .PADOUT(N__3707),
            .PADIN(N__3706),
            .CLOCKENABLE(),
            .DIN0(a_i_c_1),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD a_i_ibuf_10_iopad (
            .OE(N__3699),
            .DIN(N__3698),
            .DOUT(N__3697),
            .PACKAGEPIN(a_i[10]));
    defparam a_i_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam a_i_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO a_i_ibuf_10_preio (
            .PADOEN(N__3699),
            .PADOUT(N__3698),
            .PADIN(N__3697),
            .CLOCKENABLE(),
            .DIN0(a_i_c_10),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD a_i_ibuf_11_iopad (
            .OE(N__3690),
            .DIN(N__3689),
            .DOUT(N__3688),
            .PACKAGEPIN(a_i[11]));
    defparam a_i_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam a_i_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO a_i_ibuf_11_preio (
            .PADOEN(N__3690),
            .PADOUT(N__3689),
            .PADIN(N__3688),
            .CLOCKENABLE(),
            .DIN0(a_i_c_11),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD a_i_ibuf_12_iopad (
            .OE(N__3681),
            .DIN(N__3680),
            .DOUT(N__3679),
            .PACKAGEPIN(a_i[12]));
    defparam a_i_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam a_i_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO a_i_ibuf_12_preio (
            .PADOEN(N__3681),
            .PADOUT(N__3680),
            .PADIN(N__3679),
            .CLOCKENABLE(),
            .DIN0(a_i_c_12),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD a_i_ibuf_13_iopad (
            .OE(N__3672),
            .DIN(N__3671),
            .DOUT(N__3670),
            .PACKAGEPIN(a_i[13]));
    defparam a_i_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam a_i_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO a_i_ibuf_13_preio (
            .PADOEN(N__3672),
            .PADOUT(N__3671),
            .PADIN(N__3670),
            .CLOCKENABLE(),
            .DIN0(a_i_c_13),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD a_i_ibuf_14_iopad (
            .OE(N__3663),
            .DIN(N__3662),
            .DOUT(N__3661),
            .PACKAGEPIN(a_i[14]));
    defparam a_i_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam a_i_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO a_i_ibuf_14_preio (
            .PADOEN(N__3663),
            .PADOUT(N__3662),
            .PADIN(N__3661),
            .CLOCKENABLE(),
            .DIN0(a_i_c_14),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD a_i_ibuf_15_iopad (
            .OE(N__3654),
            .DIN(N__3653),
            .DOUT(N__3652),
            .PACKAGEPIN(a_i[15]));
    defparam a_i_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam a_i_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO a_i_ibuf_15_preio (
            .PADOEN(N__3654),
            .PADOUT(N__3653),
            .PADIN(N__3652),
            .CLOCKENABLE(),
            .DIN0(a_i_c_15),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD a_i_ibuf_2_iopad (
            .OE(N__3645),
            .DIN(N__3644),
            .DOUT(N__3643),
            .PACKAGEPIN(a_i[2]));
    defparam a_i_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam a_i_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO a_i_ibuf_2_preio (
            .PADOEN(N__3645),
            .PADOUT(N__3644),
            .PADIN(N__3643),
            .CLOCKENABLE(),
            .DIN0(a_i_c_2),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD a_i_ibuf_3_iopad (
            .OE(N__3636),
            .DIN(N__3635),
            .DOUT(N__3634),
            .PACKAGEPIN(a_i[3]));
    defparam a_i_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam a_i_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO a_i_ibuf_3_preio (
            .PADOEN(N__3636),
            .PADOUT(N__3635),
            .PADIN(N__3634),
            .CLOCKENABLE(),
            .DIN0(a_i_c_3),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD a_i_ibuf_4_iopad (
            .OE(N__3627),
            .DIN(N__3626),
            .DOUT(N__3625),
            .PACKAGEPIN(a_i[4]));
    defparam a_i_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam a_i_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO a_i_ibuf_4_preio (
            .PADOEN(N__3627),
            .PADOUT(N__3626),
            .PADIN(N__3625),
            .CLOCKENABLE(),
            .DIN0(a_i_c_4),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD a_i_ibuf_5_iopad (
            .OE(N__3618),
            .DIN(N__3617),
            .DOUT(N__3616),
            .PACKAGEPIN(a_i[5]));
    defparam a_i_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam a_i_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO a_i_ibuf_5_preio (
            .PADOEN(N__3618),
            .PADOUT(N__3617),
            .PADIN(N__3616),
            .CLOCKENABLE(),
            .DIN0(a_i_c_5),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD a_i_ibuf_6_iopad (
            .OE(N__3609),
            .DIN(N__3608),
            .DOUT(N__3607),
            .PACKAGEPIN(a_i[6]));
    defparam a_i_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam a_i_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO a_i_ibuf_6_preio (
            .PADOEN(N__3609),
            .PADOUT(N__3608),
            .PADIN(N__3607),
            .CLOCKENABLE(),
            .DIN0(a_i_c_6),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD a_i_ibuf_7_iopad (
            .OE(N__3600),
            .DIN(N__3599),
            .DOUT(N__3598),
            .PACKAGEPIN(a_i[7]));
    defparam a_i_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam a_i_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO a_i_ibuf_7_preio (
            .PADOEN(N__3600),
            .PADOUT(N__3599),
            .PADIN(N__3598),
            .CLOCKENABLE(),
            .DIN0(a_i_c_7),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD a_i_ibuf_8_iopad (
            .OE(N__3591),
            .DIN(N__3590),
            .DOUT(N__3589),
            .PACKAGEPIN(a_i[8]));
    defparam a_i_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam a_i_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO a_i_ibuf_8_preio (
            .PADOEN(N__3591),
            .PADOUT(N__3590),
            .PADIN(N__3589),
            .CLOCKENABLE(),
            .DIN0(a_i_c_8),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD a_i_ibuf_9_iopad (
            .OE(N__3582),
            .DIN(N__3581),
            .DOUT(N__3580),
            .PACKAGEPIN(a_i[9]));
    defparam a_i_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam a_i_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO a_i_ibuf_9_preio (
            .PADOEN(N__3582),
            .PADOUT(N__3581),
            .PADIN(N__3580),
            .CLOCKENABLE(),
            .DIN0(a_i_c_9),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD b_i_ibuf_0_iopad (
            .OE(N__3573),
            .DIN(N__3572),
            .DOUT(N__3571),
            .PACKAGEPIN(b_i[0]));
    defparam b_i_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam b_i_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO b_i_ibuf_0_preio (
            .PADOEN(N__3573),
            .PADOUT(N__3572),
            .PADIN(N__3571),
            .CLOCKENABLE(),
            .DIN0(b_i_c_0),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD b_i_ibuf_1_iopad (
            .OE(N__3564),
            .DIN(N__3563),
            .DOUT(N__3562),
            .PACKAGEPIN(b_i[1]));
    defparam b_i_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam b_i_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO b_i_ibuf_1_preio (
            .PADOEN(N__3564),
            .PADOUT(N__3563),
            .PADIN(N__3562),
            .CLOCKENABLE(),
            .DIN0(b_i_c_1),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD b_i_ibuf_10_iopad (
            .OE(N__3555),
            .DIN(N__3554),
            .DOUT(N__3553),
            .PACKAGEPIN(b_i[10]));
    defparam b_i_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam b_i_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO b_i_ibuf_10_preio (
            .PADOEN(N__3555),
            .PADOUT(N__3554),
            .PADIN(N__3553),
            .CLOCKENABLE(),
            .DIN0(b_i_c_10),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD b_i_ibuf_11_iopad (
            .OE(N__3546),
            .DIN(N__3545),
            .DOUT(N__3544),
            .PACKAGEPIN(b_i[11]));
    defparam b_i_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam b_i_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO b_i_ibuf_11_preio (
            .PADOEN(N__3546),
            .PADOUT(N__3545),
            .PADIN(N__3544),
            .CLOCKENABLE(),
            .DIN0(b_i_c_11),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD b_i_ibuf_12_iopad (
            .OE(N__3537),
            .DIN(N__3536),
            .DOUT(N__3535),
            .PACKAGEPIN(b_i[12]));
    defparam b_i_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam b_i_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO b_i_ibuf_12_preio (
            .PADOEN(N__3537),
            .PADOUT(N__3536),
            .PADIN(N__3535),
            .CLOCKENABLE(),
            .DIN0(b_i_c_12),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD b_i_ibuf_13_iopad (
            .OE(N__3528),
            .DIN(N__3527),
            .DOUT(N__3526),
            .PACKAGEPIN(b_i[13]));
    defparam b_i_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam b_i_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO b_i_ibuf_13_preio (
            .PADOEN(N__3528),
            .PADOUT(N__3527),
            .PADIN(N__3526),
            .CLOCKENABLE(),
            .DIN0(b_i_c_13),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD b_i_ibuf_14_iopad (
            .OE(N__3519),
            .DIN(N__3518),
            .DOUT(N__3517),
            .PACKAGEPIN(b_i[14]));
    defparam b_i_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam b_i_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO b_i_ibuf_14_preio (
            .PADOEN(N__3519),
            .PADOUT(N__3518),
            .PADIN(N__3517),
            .CLOCKENABLE(),
            .DIN0(b_i_c_14),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD b_i_ibuf_15_iopad (
            .OE(N__3510),
            .DIN(N__3509),
            .DOUT(N__3508),
            .PACKAGEPIN(b_i[15]));
    defparam b_i_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam b_i_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO b_i_ibuf_15_preio (
            .PADOEN(N__3510),
            .PADOUT(N__3509),
            .PADIN(N__3508),
            .CLOCKENABLE(),
            .DIN0(b_i_c_15),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD b_i_ibuf_2_iopad (
            .OE(N__3501),
            .DIN(N__3500),
            .DOUT(N__3499),
            .PACKAGEPIN(b_i[2]));
    defparam b_i_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam b_i_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO b_i_ibuf_2_preio (
            .PADOEN(N__3501),
            .PADOUT(N__3500),
            .PADIN(N__3499),
            .CLOCKENABLE(),
            .DIN0(b_i_c_2),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD b_i_ibuf_3_iopad (
            .OE(N__3492),
            .DIN(N__3491),
            .DOUT(N__3490),
            .PACKAGEPIN(b_i[3]));
    defparam b_i_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam b_i_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO b_i_ibuf_3_preio (
            .PADOEN(N__3492),
            .PADOUT(N__3491),
            .PADIN(N__3490),
            .CLOCKENABLE(),
            .DIN0(b_i_c_3),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD b_i_ibuf_4_iopad (
            .OE(N__3483),
            .DIN(N__3482),
            .DOUT(N__3481),
            .PACKAGEPIN(b_i[4]));
    defparam b_i_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam b_i_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO b_i_ibuf_4_preio (
            .PADOEN(N__3483),
            .PADOUT(N__3482),
            .PADIN(N__3481),
            .CLOCKENABLE(),
            .DIN0(b_i_c_4),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD b_i_ibuf_5_iopad (
            .OE(N__3474),
            .DIN(N__3473),
            .DOUT(N__3472),
            .PACKAGEPIN(b_i[5]));
    defparam b_i_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam b_i_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO b_i_ibuf_5_preio (
            .PADOEN(N__3474),
            .PADOUT(N__3473),
            .PADIN(N__3472),
            .CLOCKENABLE(),
            .DIN0(b_i_c_5),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD b_i_ibuf_6_iopad (
            .OE(N__3465),
            .DIN(N__3464),
            .DOUT(N__3463),
            .PACKAGEPIN(b_i[6]));
    defparam b_i_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam b_i_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO b_i_ibuf_6_preio (
            .PADOEN(N__3465),
            .PADOUT(N__3464),
            .PADIN(N__3463),
            .CLOCKENABLE(),
            .DIN0(b_i_c_6),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD b_i_ibuf_7_iopad (
            .OE(N__3456),
            .DIN(N__3455),
            .DOUT(N__3454),
            .PACKAGEPIN(b_i[7]));
    defparam b_i_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam b_i_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO b_i_ibuf_7_preio (
            .PADOEN(N__3456),
            .PADOUT(N__3455),
            .PADIN(N__3454),
            .CLOCKENABLE(),
            .DIN0(b_i_c_7),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD b_i_ibuf_8_iopad (
            .OE(N__3447),
            .DIN(N__3446),
            .DOUT(N__3445),
            .PACKAGEPIN(b_i[8]));
    defparam b_i_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam b_i_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO b_i_ibuf_8_preio (
            .PADOEN(N__3447),
            .PADOUT(N__3446),
            .PADIN(N__3445),
            .CLOCKENABLE(),
            .DIN0(b_i_c_8),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD b_i_ibuf_9_iopad (
            .OE(N__3438),
            .DIN(N__3437),
            .DOUT(N__3436),
            .PACKAGEPIN(b_i[9]));
    defparam b_i_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam b_i_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO b_i_ibuf_9_preio (
            .PADOEN(N__3438),
            .PADOUT(N__3437),
            .PADIN(N__3436),
            .CLOCKENABLE(),
            .DIN0(b_i_c_9),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD cin_i_ibuf_iopad (
            .OE(N__3429),
            .DIN(N__3428),
            .DOUT(N__3427),
            .PACKAGEPIN(cin_i));
    defparam cin_i_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam cin_i_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO cin_i_ibuf_preio (
            .PADOEN(N__3429),
            .PADOUT(N__3428),
            .PADIN(N__3427),
            .CLOCKENABLE(),
            .DIN0(cin_i_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD cout_o_obuf_iopad (
            .OE(N__3420),
            .DIN(N__3419),
            .DOUT(N__3418),
            .PACKAGEPIN(cout_o));
    defparam cout_o_obuf_preio.NEG_TRIGGER=1'b0;
    defparam cout_o_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO cout_o_obuf_preio (
            .PADOEN(N__3420),
            .PADOUT(N__3419),
            .PADIN(N__3418),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__2084),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD sum_o_obuf_0_iopad (
            .OE(N__3411),
            .DIN(N__3410),
            .DOUT(N__3409),
            .PACKAGEPIN(sum_o[0]));
    defparam sum_o_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam sum_o_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO sum_o_obuf_0_preio (
            .PADOEN(N__3411),
            .PADOUT(N__3410),
            .PADIN(N__3409),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__2348),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD sum_o_obuf_1_iopad (
            .OE(N__3402),
            .DIN(N__3401),
            .DOUT(N__3400),
            .PACKAGEPIN(sum_o[1]));
    defparam sum_o_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam sum_o_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO sum_o_obuf_1_preio (
            .PADOEN(N__3402),
            .PADOUT(N__3401),
            .PADIN(N__3400),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__2171),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD sum_o_obuf_10_iopad (
            .OE(N__3393),
            .DIN(N__3392),
            .DOUT(N__3391),
            .PACKAGEPIN(sum_o[10]));
    defparam sum_o_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam sum_o_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO sum_o_obuf_10_preio (
            .PADOEN(N__3393),
            .PADOUT(N__3392),
            .PADIN(N__3391),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__1805),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD sum_o_obuf_11_iopad (
            .OE(N__3384),
            .DIN(N__3383),
            .DOUT(N__3382),
            .PACKAGEPIN(sum_o[11]));
    defparam sum_o_obuf_11_preio.NEG_TRIGGER=1'b0;
    defparam sum_o_obuf_11_preio.PIN_TYPE=6'b011001;
    PRE_IO sum_o_obuf_11_preio (
            .PADOEN(N__3384),
            .PADOUT(N__3383),
            .PADIN(N__3382),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__1844),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD sum_o_obuf_12_iopad (
            .OE(N__3375),
            .DIN(N__3374),
            .DOUT(N__3373),
            .PACKAGEPIN(sum_o[12]));
    defparam sum_o_obuf_12_preio.NEG_TRIGGER=1'b0;
    defparam sum_o_obuf_12_preio.PIN_TYPE=6'b011001;
    PRE_IO sum_o_obuf_12_preio (
            .PADOEN(N__3375),
            .PADOUT(N__3374),
            .PADIN(N__3373),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__1670),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD sum_o_obuf_13_iopad (
            .OE(N__3366),
            .DIN(N__3365),
            .DOUT(N__3364),
            .PACKAGEPIN(sum_o[13]));
    defparam sum_o_obuf_13_preio.NEG_TRIGGER=1'b0;
    defparam sum_o_obuf_13_preio.PIN_TYPE=6'b011001;
    PRE_IO sum_o_obuf_13_preio (
            .PADOEN(N__3366),
            .PADOUT(N__3365),
            .PADIN(N__3364),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__1790),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD sum_o_obuf_14_iopad (
            .OE(N__3357),
            .DIN(N__3356),
            .DOUT(N__3355),
            .PACKAGEPIN(sum_o[14]));
    defparam sum_o_obuf_14_preio.NEG_TRIGGER=1'b0;
    defparam sum_o_obuf_14_preio.PIN_TYPE=6'b011001;
    PRE_IO sum_o_obuf_14_preio (
            .PADOEN(N__3357),
            .PADOUT(N__3356),
            .PADIN(N__3355),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__1898),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD sum_o_obuf_15_iopad (
            .OE(N__3348),
            .DIN(N__3347),
            .DOUT(N__3346),
            .PACKAGEPIN(sum_o[15]));
    defparam sum_o_obuf_15_preio.NEG_TRIGGER=1'b0;
    defparam sum_o_obuf_15_preio.PIN_TYPE=6'b011001;
    PRE_IO sum_o_obuf_15_preio (
            .PADOEN(N__3348),
            .PADOUT(N__3347),
            .PADIN(N__3346),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__2816),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD sum_o_obuf_2_iopad (
            .OE(N__3339),
            .DIN(N__3338),
            .DOUT(N__3337),
            .PACKAGEPIN(sum_o[2]));
    defparam sum_o_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam sum_o_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO sum_o_obuf_2_preio (
            .PADOEN(N__3339),
            .PADOUT(N__3338),
            .PADIN(N__3337),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__2135),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD sum_o_obuf_3_iopad (
            .OE(N__3330),
            .DIN(N__3329),
            .DOUT(N__3328),
            .PACKAGEPIN(sum_o[3]));
    defparam sum_o_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam sum_o_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO sum_o_obuf_3_preio (
            .PADOEN(N__3330),
            .PADOUT(N__3329),
            .PADIN(N__3328),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__2183),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD sum_o_obuf_4_iopad (
            .OE(N__3321),
            .DIN(N__3320),
            .DOUT(N__3319),
            .PACKAGEPIN(sum_o[4]));
    defparam sum_o_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam sum_o_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO sum_o_obuf_4_preio (
            .PADOEN(N__3321),
            .PADOUT(N__3320),
            .PADIN(N__3319),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__2156),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD sum_o_obuf_5_iopad (
            .OE(N__3312),
            .DIN(N__3311),
            .DOUT(N__3310),
            .PACKAGEPIN(sum_o[5]));
    defparam sum_o_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam sum_o_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO sum_o_obuf_5_preio (
            .PADOEN(N__3312),
            .PADOUT(N__3311),
            .PADIN(N__3310),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__1931),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD sum_o_obuf_6_iopad (
            .OE(N__3303),
            .DIN(N__3302),
            .DOUT(N__3301),
            .PACKAGEPIN(sum_o[6]));
    defparam sum_o_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam sum_o_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO sum_o_obuf_6_preio (
            .PADOEN(N__3303),
            .PADOUT(N__3302),
            .PADIN(N__3301),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__2732),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD sum_o_obuf_7_iopad (
            .OE(N__3294),
            .DIN(N__3293),
            .DOUT(N__3292),
            .PACKAGEPIN(sum_o[7]));
    defparam sum_o_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam sum_o_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO sum_o_obuf_7_preio (
            .PADOEN(N__3294),
            .PADOUT(N__3293),
            .PADIN(N__3292),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__2891),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD sum_o_obuf_8_iopad (
            .OE(N__3285),
            .DIN(N__3284),
            .DOUT(N__3283),
            .PACKAGEPIN(sum_o[8]));
    defparam sum_o_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam sum_o_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO sum_o_obuf_8_preio (
            .PADOEN(N__3285),
            .PADOUT(N__3284),
            .PADIN(N__3283),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__1892),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD sum_o_obuf_9_iopad (
            .OE(N__3276),
            .DIN(N__3275),
            .DOUT(N__3274),
            .PACKAGEPIN(sum_o[9]));
    defparam sum_o_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam sum_o_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO sum_o_obuf_9_preio (
            .PADOEN(N__3276),
            .PADOUT(N__3275),
            .PADIN(N__3274),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__1655),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    InMux I__683 (
            .O(N__3257),
            .I(N__3254));
    LocalMux I__682 (
            .O(N__3254),
            .I(N__3251));
    Span4Mux_v I__681 (
            .O(N__3251),
            .I(N__3248));
    Span4Mux_v I__680 (
            .O(N__3248),
            .I(N__3245));
    Odrv4 I__679 (
            .O(N__3245),
            .I(b_i_c_5));
    InMux I__678 (
            .O(N__3242),
            .I(N__3235));
    InMux I__677 (
            .O(N__3241),
            .I(N__3235));
    InMux I__676 (
            .O(N__3240),
            .I(N__3232));
    LocalMux I__675 (
            .O(N__3235),
            .I(b_rZ0Z_5));
    LocalMux I__674 (
            .O(N__3232),
            .I(b_rZ0Z_5));
    InMux I__673 (
            .O(N__3227),
            .I(N__3224));
    LocalMux I__672 (
            .O(N__3224),
            .I(N__3221));
    Span12Mux_v I__671 (
            .O(N__3221),
            .I(N__3218));
    Odrv12 I__670 (
            .O(N__3218),
            .I(a_i_c_3));
    InMux I__669 (
            .O(N__3215),
            .I(N__3212));
    LocalMux I__668 (
            .O(N__3212),
            .I(N__3208));
    InMux I__667 (
            .O(N__3211),
            .I(N__3205));
    Odrv4 I__666 (
            .O(N__3208),
            .I(a_rZ0Z_3));
    LocalMux I__665 (
            .O(N__3205),
            .I(a_rZ0Z_3));
    InMux I__664 (
            .O(N__3200),
            .I(N__3197));
    LocalMux I__663 (
            .O(N__3197),
            .I(N__3194));
    IoSpan4Mux I__662 (
            .O(N__3194),
            .I(N__3191));
    Odrv4 I__661 (
            .O(N__3191),
            .I(b_i_c_7));
    InMux I__660 (
            .O(N__3188),
            .I(N__3185));
    LocalMux I__659 (
            .O(N__3185),
            .I(b_rZ0Z_7));
    InMux I__658 (
            .O(N__3182),
            .I(N__3179));
    LocalMux I__657 (
            .O(N__3179),
            .I(N__3176));
    Span4Mux_h I__656 (
            .O(N__3176),
            .I(N__3173));
    Span4Mux_v I__655 (
            .O(N__3173),
            .I(N__3170));
    Odrv4 I__654 (
            .O(N__3170),
            .I(b_i_c_6));
    CascadeMux I__653 (
            .O(N__3167),
            .I(N__3164));
    InMux I__652 (
            .O(N__3164),
            .I(N__3158));
    InMux I__651 (
            .O(N__3163),
            .I(N__3158));
    LocalMux I__650 (
            .O(N__3158),
            .I(b_rZ0Z_6));
    ClkMux I__649 (
            .O(N__3155),
            .I(N__3119));
    ClkMux I__648 (
            .O(N__3154),
            .I(N__3119));
    ClkMux I__647 (
            .O(N__3153),
            .I(N__3119));
    ClkMux I__646 (
            .O(N__3152),
            .I(N__3119));
    ClkMux I__645 (
            .O(N__3151),
            .I(N__3119));
    ClkMux I__644 (
            .O(N__3150),
            .I(N__3119));
    ClkMux I__643 (
            .O(N__3149),
            .I(N__3119));
    ClkMux I__642 (
            .O(N__3148),
            .I(N__3119));
    ClkMux I__641 (
            .O(N__3147),
            .I(N__3119));
    ClkMux I__640 (
            .O(N__3146),
            .I(N__3119));
    ClkMux I__639 (
            .O(N__3145),
            .I(N__3119));
    ClkMux I__638 (
            .O(N__3144),
            .I(N__3119));
    GlobalMux I__637 (
            .O(N__3119),
            .I(N__3116));
    gio2CtrlBuf I__636 (
            .O(N__3116),
            .I(clk_i_c_g));
    InMux I__635 (
            .O(N__3113),
            .I(N__3110));
    LocalMux I__634 (
            .O(N__3110),
            .I(N__3107));
    Span12Mux_v I__633 (
            .O(N__3107),
            .I(N__3104));
    Odrv12 I__632 (
            .O(N__3104),
            .I(a_i_c_7));
    InMux I__631 (
            .O(N__3101),
            .I(N__3098));
    LocalMux I__630 (
            .O(N__3098),
            .I(N__3095));
    Span4Mux_v I__629 (
            .O(N__3095),
            .I(N__3092));
    Odrv4 I__628 (
            .O(N__3092),
            .I(a_i_c_13));
    CascadeMux I__627 (
            .O(N__3089),
            .I(N__3086));
    InMux I__626 (
            .O(N__3086),
            .I(N__3083));
    LocalMux I__625 (
            .O(N__3083),
            .I(N__3080));
    Odrv4 I__624 (
            .O(N__3080),
            .I(a_rZ0Z_13));
    InMux I__623 (
            .O(N__3077),
            .I(N__3074));
    LocalMux I__622 (
            .O(N__3074),
            .I(N__3071));
    Span12Mux_h I__621 (
            .O(N__3071),
            .I(N__3068));
    Span12Mux_v I__620 (
            .O(N__3068),
            .I(N__3065));
    Odrv12 I__619 (
            .O(N__3065),
            .I(a_i_c_4));
    InMux I__618 (
            .O(N__3062),
            .I(N__3057));
    InMux I__617 (
            .O(N__3061),
            .I(N__3052));
    InMux I__616 (
            .O(N__3060),
            .I(N__3052));
    LocalMux I__615 (
            .O(N__3057),
            .I(N__3049));
    LocalMux I__614 (
            .O(N__3052),
            .I(N__3046));
    Span4Mux_h I__613 (
            .O(N__3049),
            .I(N__3043));
    Odrv12 I__612 (
            .O(N__3046),
            .I(a_rZ0Z_4));
    Odrv4 I__611 (
            .O(N__3043),
            .I(a_rZ0Z_4));
    CascadeMux I__610 (
            .O(N__3038),
            .I(N__3035));
    InMux I__609 (
            .O(N__3035),
            .I(N__3032));
    LocalMux I__608 (
            .O(N__3032),
            .I(b_r_i_5));
    InMux I__607 (
            .O(N__3029),
            .I(N__3026));
    LocalMux I__606 (
            .O(N__3026),
            .I(N__3023));
    Sp12to4 I__605 (
            .O(N__3023),
            .I(N__3020));
    Span12Mux_v I__604 (
            .O(N__3020),
            .I(N__3017));
    Odrv12 I__603 (
            .O(N__3017),
            .I(a_i_c_2));
    InMux I__602 (
            .O(N__3014),
            .I(N__3010));
    InMux I__601 (
            .O(N__3013),
            .I(N__3007));
    LocalMux I__600 (
            .O(N__3010),
            .I(N__3004));
    LocalMux I__599 (
            .O(N__3007),
            .I(N__3001));
    Odrv4 I__598 (
            .O(N__3004),
            .I(a_rZ0Z_2));
    Odrv4 I__597 (
            .O(N__3001),
            .I(a_rZ0Z_2));
    InMux I__596 (
            .O(N__2996),
            .I(N__2992));
    InMux I__595 (
            .O(N__2995),
            .I(N__2989));
    LocalMux I__594 (
            .O(N__2992),
            .I(N__2986));
    LocalMux I__593 (
            .O(N__2989),
            .I(N__2983));
    Odrv4 I__592 (
            .O(N__2986),
            .I(a_rZ0Z_7));
    Odrv4 I__591 (
            .O(N__2983),
            .I(a_rZ0Z_7));
    CascadeMux I__590 (
            .O(N__2978),
            .I(N__2975));
    InMux I__589 (
            .O(N__2975),
            .I(N__2972));
    LocalMux I__588 (
            .O(N__2972),
            .I(b_r_RNI409BZ0Z_7));
    InMux I__587 (
            .O(N__2969),
            .I(N__2966));
    LocalMux I__586 (
            .O(N__2966),
            .I(N__2962));
    InMux I__585 (
            .O(N__2965),
            .I(N__2959));
    Odrv4 I__584 (
            .O(N__2962),
            .I(a_rZ0Z_6));
    LocalMux I__583 (
            .O(N__2959),
            .I(a_rZ0Z_6));
    CascadeMux I__582 (
            .O(N__2954),
            .I(N__2951));
    InMux I__581 (
            .O(N__2951),
            .I(N__2948));
    LocalMux I__580 (
            .O(N__2948),
            .I(b_r_RNI15S9Z0Z_6));
    InMux I__579 (
            .O(N__2945),
            .I(N__2941));
    InMux I__578 (
            .O(N__2944),
            .I(N__2938));
    LocalMux I__577 (
            .O(N__2941),
            .I(N__2935));
    LocalMux I__576 (
            .O(N__2938),
            .I(un5_sum_v_cry_5_c_RNI5CQZ0Z01));
    Odrv4 I__575 (
            .O(N__2935),
            .I(un5_sum_v_cry_5_c_RNI5CQZ0Z01));
    InMux I__574 (
            .O(N__2930),
            .I(N__2927));
    LocalMux I__573 (
            .O(N__2927),
            .I(sum_r_RNO_0Z0Z_7));
    CascadeMux I__572 (
            .O(N__2924),
            .I(N__2921));
    InMux I__571 (
            .O(N__2921),
            .I(N__2916));
    InMux I__570 (
            .O(N__2920),
            .I(N__2913));
    InMux I__569 (
            .O(N__2919),
            .I(N__2910));
    LocalMux I__568 (
            .O(N__2916),
            .I(N__2907));
    LocalMux I__567 (
            .O(N__2913),
            .I(N__2902));
    LocalMux I__566 (
            .O(N__2910),
            .I(N__2902));
    Odrv4 I__565 (
            .O(N__2907),
            .I(b_r_sbtinv_RNINK2RZ0Z_5));
    Odrv4 I__564 (
            .O(N__2902),
            .I(b_r_sbtinv_RNINK2RZ0Z_5));
    InMux I__563 (
            .O(N__2897),
            .I(N__2894));
    LocalMux I__562 (
            .O(N__2894),
            .I(un40_sum_v));
    IoInMux I__561 (
            .O(N__2891),
            .I(N__2888));
    LocalMux I__560 (
            .O(N__2888),
            .I(N__2885));
    Span4Mux_s2_h I__559 (
            .O(N__2885),
            .I(N__2882));
    Odrv4 I__558 (
            .O(N__2882),
            .I(sum_o_c_7));
    InMux I__557 (
            .O(N__2879),
            .I(un5_sum_v_cry_15));
    InMux I__556 (
            .O(N__2876),
            .I(N__2871));
    InMux I__555 (
            .O(N__2875),
            .I(N__2866));
    InMux I__554 (
            .O(N__2874),
            .I(N__2866));
    LocalMux I__553 (
            .O(N__2871),
            .I(un5_sum_v_cry_15_THRU_CO));
    LocalMux I__552 (
            .O(N__2866),
            .I(un5_sum_v_cry_15_THRU_CO));
    CascadeMux I__551 (
            .O(N__2861),
            .I(N__2856));
    InMux I__550 (
            .O(N__2860),
            .I(N__2853));
    InMux I__549 (
            .O(N__2859),
            .I(N__2850));
    InMux I__548 (
            .O(N__2856),
            .I(N__2847));
    LocalMux I__547 (
            .O(N__2853),
            .I(un5_sum_v_cry_12_c_RNI45JOZ0));
    LocalMux I__546 (
            .O(N__2850),
            .I(un5_sum_v_cry_12_c_RNI45JOZ0));
    LocalMux I__545 (
            .O(N__2847),
            .I(un5_sum_v_cry_12_c_RNI45JOZ0));
    CascadeMux I__544 (
            .O(N__2840),
            .I(N__2837));
    InMux I__543 (
            .O(N__2837),
            .I(N__2833));
    InMux I__542 (
            .O(N__2836),
            .I(N__2830));
    LocalMux I__541 (
            .O(N__2833),
            .I(un5_sum_v_cry_13_c_RNIG5IKZ0Z1));
    LocalMux I__540 (
            .O(N__2830),
            .I(un5_sum_v_cry_13_c_RNIG5IKZ0Z1));
    CascadeMux I__539 (
            .O(N__2825),
            .I(un5_sum_v_cry_15_THRU_CO_cascade_));
    InMux I__538 (
            .O(N__2822),
            .I(N__2819));
    LocalMux I__537 (
            .O(N__2819),
            .I(sum_r_RNO_0Z0Z_15));
    IoInMux I__536 (
            .O(N__2816),
            .I(N__2813));
    LocalMux I__535 (
            .O(N__2813),
            .I(N__2810));
    IoSpan4Mux I__534 (
            .O(N__2810),
            .I(N__2807));
    Span4Mux_s1_h I__533 (
            .O(N__2807),
            .I(N__2804));
    Span4Mux_v I__532 (
            .O(N__2804),
            .I(N__2801));
    Odrv4 I__531 (
            .O(N__2801),
            .I(sum_o_c_15));
    CascadeMux I__530 (
            .O(N__2798),
            .I(N__2794));
    CascadeMux I__529 (
            .O(N__2797),
            .I(N__2790));
    InMux I__528 (
            .O(N__2794),
            .I(N__2787));
    InMux I__527 (
            .O(N__2793),
            .I(N__2784));
    InMux I__526 (
            .O(N__2790),
            .I(N__2781));
    LocalMux I__525 (
            .O(N__2787),
            .I(N__2774));
    LocalMux I__524 (
            .O(N__2784),
            .I(N__2774));
    LocalMux I__523 (
            .O(N__2781),
            .I(N__2774));
    Odrv4 I__522 (
            .O(N__2774),
            .I(a_rZ0Z_8));
    InMux I__521 (
            .O(N__2771),
            .I(N__2766));
    InMux I__520 (
            .O(N__2770),
            .I(N__2763));
    InMux I__519 (
            .O(N__2769),
            .I(N__2760));
    LocalMux I__518 (
            .O(N__2766),
            .I(b_rZ0Z_8));
    LocalMux I__517 (
            .O(N__2763),
            .I(b_rZ0Z_8));
    LocalMux I__516 (
            .O(N__2760),
            .I(b_rZ0Z_8));
    InMux I__515 (
            .O(N__2753),
            .I(N__2748));
    InMux I__514 (
            .O(N__2752),
            .I(N__2745));
    InMux I__513 (
            .O(N__2751),
            .I(N__2742));
    LocalMux I__512 (
            .O(N__2748),
            .I(un5_sum_v_cry_7_c_RNIB8DOZ0));
    LocalMux I__511 (
            .O(N__2745),
            .I(un5_sum_v_cry_7_c_RNIB8DOZ0));
    LocalMux I__510 (
            .O(N__2742),
            .I(un5_sum_v_cry_7_c_RNIB8DOZ0));
    CascadeMux I__509 (
            .O(N__2735),
            .I(un40_sum_v_cascade_));
    IoInMux I__508 (
            .O(N__2732),
            .I(N__2729));
    LocalMux I__507 (
            .O(N__2729),
            .I(N__2726));
    Span4Mux_s1_h I__506 (
            .O(N__2726),
            .I(N__2723));
    Odrv4 I__505 (
            .O(N__2723),
            .I(sum_o_c_6));
    CascadeMux I__504 (
            .O(N__2720),
            .I(N__2717));
    InMux I__503 (
            .O(N__2717),
            .I(N__2714));
    LocalMux I__502 (
            .O(N__2714),
            .I(N__2710));
    InMux I__501 (
            .O(N__2713),
            .I(N__2707));
    Odrv4 I__500 (
            .O(N__2710),
            .I(b_rZ0Z_10));
    LocalMux I__499 (
            .O(N__2707),
            .I(b_rZ0Z_10));
    CascadeMux I__498 (
            .O(N__2702),
            .I(N__2699));
    InMux I__497 (
            .O(N__2699),
            .I(N__2696));
    LocalMux I__496 (
            .O(N__2696),
            .I(b_r_RNIRUROZ0Z_10));
    InMux I__495 (
            .O(N__2693),
            .I(N__2690));
    LocalMux I__494 (
            .O(N__2690),
            .I(N__2687));
    Sp12to4 I__493 (
            .O(N__2687),
            .I(N__2684));
    Span12Mux_v I__492 (
            .O(N__2684),
            .I(N__2681));
    Odrv12 I__491 (
            .O(N__2681),
            .I(b_i_c_1));
    InMux I__490 (
            .O(N__2678),
            .I(N__2669));
    InMux I__489 (
            .O(N__2677),
            .I(N__2669));
    InMux I__488 (
            .O(N__2676),
            .I(N__2669));
    LocalMux I__487 (
            .O(N__2669),
            .I(b_rZ0Z_1));
    CascadeMux I__486 (
            .O(N__2666),
            .I(N__2663));
    InMux I__485 (
            .O(N__2663),
            .I(N__2660));
    LocalMux I__484 (
            .O(N__2660),
            .I(b_r_i_9));
    InMux I__483 (
            .O(N__2657),
            .I(N__2654));
    LocalMux I__482 (
            .O(N__2654),
            .I(N__2651));
    Span12Mux_v I__481 (
            .O(N__2651),
            .I(N__2648));
    Odrv12 I__480 (
            .O(N__2648),
            .I(a_i_c_10));
    InMux I__479 (
            .O(N__2645),
            .I(N__2641));
    InMux I__478 (
            .O(N__2644),
            .I(N__2638));
    LocalMux I__477 (
            .O(N__2641),
            .I(N__2635));
    LocalMux I__476 (
            .O(N__2638),
            .I(a_rZ0Z_10));
    Odrv4 I__475 (
            .O(N__2635),
            .I(a_rZ0Z_10));
    InMux I__474 (
            .O(N__2630),
            .I(N__2627));
    LocalMux I__473 (
            .O(N__2627),
            .I(N__2624));
    IoSpan4Mux I__472 (
            .O(N__2624),
            .I(N__2621));
    IoSpan4Mux I__471 (
            .O(N__2621),
            .I(N__2618));
    Odrv4 I__470 (
            .O(N__2618),
            .I(b_i_c_9));
    InMux I__469 (
            .O(N__2615),
            .I(N__2610));
    InMux I__468 (
            .O(N__2614),
            .I(N__2607));
    InMux I__467 (
            .O(N__2613),
            .I(N__2604));
    LocalMux I__466 (
            .O(N__2610),
            .I(b_rZ0Z_9));
    LocalMux I__465 (
            .O(N__2607),
            .I(b_rZ0Z_9));
    LocalMux I__464 (
            .O(N__2604),
            .I(b_rZ0Z_9));
    InMux I__463 (
            .O(N__2597),
            .I(N__2594));
    LocalMux I__462 (
            .O(N__2594),
            .I(N__2591));
    Span4Mux_h I__461 (
            .O(N__2591),
            .I(N__2588));
    Odrv4 I__460 (
            .O(N__2588),
            .I(a_rZ0Z_9));
    InMux I__459 (
            .O(N__2585),
            .I(N__2580));
    InMux I__458 (
            .O(N__2584),
            .I(N__2577));
    InMux I__457 (
            .O(N__2583),
            .I(N__2574));
    LocalMux I__456 (
            .O(N__2580),
            .I(b_r_sbtinv_RNI357RZ0Z_9));
    LocalMux I__455 (
            .O(N__2577),
            .I(b_r_sbtinv_RNI357RZ0Z_9));
    LocalMux I__454 (
            .O(N__2574),
            .I(b_r_sbtinv_RNI357RZ0Z_9));
    InMux I__453 (
            .O(N__2567),
            .I(un5_sum_v_cry_8));
    InMux I__452 (
            .O(N__2564),
            .I(N__2560));
    InMux I__451 (
            .O(N__2563),
            .I(N__2557));
    LocalMux I__450 (
            .O(N__2560),
            .I(un5_sum_v_cry_9_c_RNIEOBIZ0Z1));
    LocalMux I__449 (
            .O(N__2557),
            .I(un5_sum_v_cry_9_c_RNIEOBIZ0Z1));
    InMux I__448 (
            .O(N__2552),
            .I(un5_sum_v_cry_9));
    InMux I__447 (
            .O(N__2549),
            .I(N__2545));
    InMux I__446 (
            .O(N__2548),
            .I(N__2542));
    LocalMux I__445 (
            .O(N__2545),
            .I(N__2539));
    LocalMux I__444 (
            .O(N__2542),
            .I(a_rZ0Z_11));
    Odrv4 I__443 (
            .O(N__2539),
            .I(a_rZ0Z_11));
    CascadeMux I__442 (
            .O(N__2534),
            .I(N__2531));
    InMux I__441 (
            .O(N__2531),
            .I(N__2528));
    LocalMux I__440 (
            .O(N__2528),
            .I(b_r_RNI95R61Z0Z_11));
    InMux I__439 (
            .O(N__2525),
            .I(N__2522));
    LocalMux I__438 (
            .O(N__2522),
            .I(sum_r_RNO_0Z0Z_11));
    InMux I__437 (
            .O(N__2519),
            .I(un5_sum_v_cry_10));
    InMux I__436 (
            .O(N__2516),
            .I(N__2511));
    InMux I__435 (
            .O(N__2515),
            .I(N__2506));
    InMux I__434 (
            .O(N__2514),
            .I(N__2506));
    LocalMux I__433 (
            .O(N__2511),
            .I(N__2502));
    LocalMux I__432 (
            .O(N__2506),
            .I(N__2499));
    InMux I__431 (
            .O(N__2505),
            .I(N__2496));
    Span4Mux_h I__430 (
            .O(N__2502),
            .I(N__2493));
    Odrv4 I__429 (
            .O(N__2499),
            .I(a_rZ0Z_12));
    LocalMux I__428 (
            .O(N__2496),
            .I(a_rZ0Z_12));
    Odrv4 I__427 (
            .O(N__2493),
            .I(a_rZ0Z_12));
    CascadeMux I__426 (
            .O(N__2486),
            .I(N__2482));
    CascadeMux I__425 (
            .O(N__2485),
            .I(N__2478));
    InMux I__424 (
            .O(N__2482),
            .I(N__2473));
    InMux I__423 (
            .O(N__2481),
            .I(N__2473));
    InMux I__422 (
            .O(N__2478),
            .I(N__2469));
    LocalMux I__421 (
            .O(N__2473),
            .I(N__2466));
    InMux I__420 (
            .O(N__2472),
            .I(N__2463));
    LocalMux I__419 (
            .O(N__2469),
            .I(N__2460));
    Odrv4 I__418 (
            .O(N__2466),
            .I(b_rZ0Z_12));
    LocalMux I__417 (
            .O(N__2463),
            .I(b_rZ0Z_12));
    Odrv4 I__416 (
            .O(N__2460),
            .I(b_rZ0Z_12));
    InMux I__415 (
            .O(N__2453),
            .I(N__2447));
    InMux I__414 (
            .O(N__2452),
            .I(N__2440));
    InMux I__413 (
            .O(N__2451),
            .I(N__2440));
    InMux I__412 (
            .O(N__2450),
            .I(N__2440));
    LocalMux I__411 (
            .O(N__2447),
            .I(un5_sum_v_cry_11_c_RNICJ0TZ0));
    LocalMux I__410 (
            .O(N__2440),
            .I(un5_sum_v_cry_11_c_RNICJ0TZ0));
    InMux I__409 (
            .O(N__2435),
            .I(un5_sum_v_cry_11));
    InMux I__408 (
            .O(N__2432),
            .I(N__2429));
    LocalMux I__407 (
            .O(N__2429),
            .I(b_r_i_13));
    InMux I__406 (
            .O(N__2426),
            .I(un5_sum_v_cry_12));
    InMux I__405 (
            .O(N__2423),
            .I(N__2419));
    InMux I__404 (
            .O(N__2422),
            .I(N__2416));
    LocalMux I__403 (
            .O(N__2419),
            .I(N__2413));
    LocalMux I__402 (
            .O(N__2416),
            .I(a_rZ0Z_14));
    Odrv4 I__401 (
            .O(N__2413),
            .I(a_rZ0Z_14));
    CascadeMux I__400 (
            .O(N__2408),
            .I(N__2405));
    InMux I__399 (
            .O(N__2405),
            .I(N__2402));
    LocalMux I__398 (
            .O(N__2402),
            .I(b_r_RNIEIE51Z0Z_14));
    InMux I__397 (
            .O(N__2399),
            .I(un5_sum_v_cry_13));
    CascadeMux I__396 (
            .O(N__2396),
            .I(N__2392));
    InMux I__395 (
            .O(N__2395),
            .I(N__2389));
    InMux I__394 (
            .O(N__2392),
            .I(N__2386));
    LocalMux I__393 (
            .O(N__2389),
            .I(N__2383));
    LocalMux I__392 (
            .O(N__2386),
            .I(N__2380));
    Span4Mux_v I__391 (
            .O(N__2383),
            .I(N__2377));
    Odrv4 I__390 (
            .O(N__2380),
            .I(a_rZ0Z_15));
    Odrv4 I__389 (
            .O(N__2377),
            .I(a_rZ0Z_15));
    CascadeMux I__388 (
            .O(N__2372),
            .I(N__2369));
    InMux I__387 (
            .O(N__2369),
            .I(N__2366));
    LocalMux I__386 (
            .O(N__2366),
            .I(N__2363));
    Odrv4 I__385 (
            .O(N__2363),
            .I(b_r_RNI0TDJ1Z0Z_15));
    InMux I__384 (
            .O(N__2360),
            .I(bfn_2_18_0_));
    CascadeMux I__383 (
            .O(N__2357),
            .I(N__2354));
    InMux I__382 (
            .O(N__2354),
            .I(N__2351));
    LocalMux I__381 (
            .O(N__2351),
            .I(a_rZ0Z_0));
    IoInMux I__380 (
            .O(N__2348),
            .I(N__2345));
    LocalMux I__379 (
            .O(N__2345),
            .I(N__2342));
    Span4Mux_s1_h I__378 (
            .O(N__2342),
            .I(N__2339));
    Span4Mux_v I__377 (
            .O(N__2339),
            .I(N__2336));
    Odrv4 I__376 (
            .O(N__2336),
            .I(sum_o_c_0));
    InMux I__375 (
            .O(N__2333),
            .I(un5_sum_v_cry_0_c_THRU_CO));
    InMux I__374 (
            .O(N__2330),
            .I(N__2327));
    LocalMux I__373 (
            .O(N__2327),
            .I(a_rZ0Z_1));
    CascadeMux I__372 (
            .O(N__2324),
            .I(N__2321));
    InMux I__371 (
            .O(N__2321),
            .I(N__2318));
    LocalMux I__370 (
            .O(N__2318),
            .I(b_r_i_1));
    CascadeMux I__369 (
            .O(N__2315),
            .I(N__2311));
    CascadeMux I__368 (
            .O(N__2314),
            .I(N__2307));
    InMux I__367 (
            .O(N__2311),
            .I(N__2304));
    InMux I__366 (
            .O(N__2310),
            .I(N__2299));
    InMux I__365 (
            .O(N__2307),
            .I(N__2299));
    LocalMux I__364 (
            .O(N__2304),
            .I(b_r_sbtinv_RNIB4UQZ0Z_1));
    LocalMux I__363 (
            .O(N__2299),
            .I(b_r_sbtinv_RNIB4UQZ0Z_1));
    InMux I__362 (
            .O(N__2294),
            .I(un5_sum_v_cry_0));
    CascadeMux I__361 (
            .O(N__2291),
            .I(N__2288));
    InMux I__360 (
            .O(N__2288),
            .I(N__2285));
    LocalMux I__359 (
            .O(N__2285),
            .I(b_r_RNILOR9Z0Z_2));
    InMux I__358 (
            .O(N__2282),
            .I(N__2276));
    InMux I__357 (
            .O(N__2281),
            .I(N__2276));
    LocalMux I__356 (
            .O(N__2276),
            .I(un5_sum_v_cry_1_c_RNIHJLZ0Z01));
    InMux I__355 (
            .O(N__2273),
            .I(un5_sum_v_cry_1));
    CascadeMux I__354 (
            .O(N__2270),
            .I(N__2267));
    InMux I__353 (
            .O(N__2267),
            .I(N__2264));
    LocalMux I__352 (
            .O(N__2264),
            .I(b_r_RNIKF8BZ0Z_3));
    InMux I__351 (
            .O(N__2261),
            .I(N__2258));
    LocalMux I__350 (
            .O(N__2258),
            .I(sum_r_RNO_0Z0Z_3));
    InMux I__349 (
            .O(N__2255),
            .I(un5_sum_v_cry_2));
    CascadeMux I__348 (
            .O(N__2252),
            .I(N__2247));
    InMux I__347 (
            .O(N__2251),
            .I(N__2244));
    InMux I__346 (
            .O(N__2250),
            .I(N__2241));
    InMux I__345 (
            .O(N__2247),
            .I(N__2238));
    LocalMux I__344 (
            .O(N__2244),
            .I(b_rZ0Z_4));
    LocalMux I__343 (
            .O(N__2241),
            .I(b_rZ0Z_4));
    LocalMux I__342 (
            .O(N__2238),
            .I(b_rZ0Z_4));
    InMux I__341 (
            .O(N__2231),
            .I(N__2222));
    InMux I__340 (
            .O(N__2230),
            .I(N__2222));
    InMux I__339 (
            .O(N__2229),
            .I(N__2222));
    LocalMux I__338 (
            .O(N__2222),
            .I(un5_sum_v_cry_3_c_RNIVN8OZ0));
    InMux I__337 (
            .O(N__2219),
            .I(un5_sum_v_cry_3));
    InMux I__336 (
            .O(N__2216),
            .I(N__2213));
    LocalMux I__335 (
            .O(N__2213),
            .I(a_rZ0Z_5));
    InMux I__334 (
            .O(N__2210),
            .I(un5_sum_v_cry_4));
    InMux I__333 (
            .O(N__2207),
            .I(un5_sum_v_cry_5));
    InMux I__332 (
            .O(N__2204),
            .I(bfn_2_17_0_));
    InMux I__331 (
            .O(N__2201),
            .I(un5_sum_v_cry_7));
    InMux I__330 (
            .O(N__2198),
            .I(N__2195));
    LocalMux I__329 (
            .O(N__2195),
            .I(N__2192));
    Span12Mux_h I__328 (
            .O(N__2192),
            .I(N__2189));
    Span12Mux_v I__327 (
            .O(N__2189),
            .I(N__2186));
    Odrv12 I__326 (
            .O(N__2186),
            .I(cin_i_c));
    IoInMux I__325 (
            .O(N__2183),
            .I(N__2180));
    LocalMux I__324 (
            .O(N__2180),
            .I(N__2177));
    Span4Mux_s1_h I__323 (
            .O(N__2177),
            .I(N__2174));
    Odrv4 I__322 (
            .O(N__2174),
            .I(sum_o_c_3));
    IoInMux I__321 (
            .O(N__2171),
            .I(N__2168));
    LocalMux I__320 (
            .O(N__2168),
            .I(N__2165));
    Span4Mux_s1_h I__319 (
            .O(N__2165),
            .I(N__2162));
    Sp12to4 I__318 (
            .O(N__2162),
            .I(N__2159));
    Odrv12 I__317 (
            .O(N__2159),
            .I(sum_o_c_1));
    IoInMux I__316 (
            .O(N__2156),
            .I(N__2153));
    LocalMux I__315 (
            .O(N__2153),
            .I(N__2150));
    Span4Mux_s1_h I__314 (
            .O(N__2150),
            .I(N__2147));
    Odrv4 I__313 (
            .O(N__2147),
            .I(sum_o_c_4));
    InMux I__312 (
            .O(N__2144),
            .I(N__2141));
    LocalMux I__311 (
            .O(N__2141),
            .I(un13_sum_v));
    CascadeMux I__310 (
            .O(N__2138),
            .I(un13_sum_v_cascade_));
    IoInMux I__309 (
            .O(N__2135),
            .I(N__2132));
    LocalMux I__308 (
            .O(N__2132),
            .I(N__2129));
    Span4Mux_s0_h I__307 (
            .O(N__2129),
            .I(N__2126));
    Span4Mux_v I__306 (
            .O(N__2126),
            .I(N__2123));
    Odrv4 I__305 (
            .O(N__2123),
            .I(sum_o_c_2));
    InMux I__304 (
            .O(N__2120),
            .I(N__2117));
    LocalMux I__303 (
            .O(N__2117),
            .I(N__2114));
    Span12Mux_v I__302 (
            .O(N__2114),
            .I(N__2111));
    Odrv12 I__301 (
            .O(N__2111),
            .I(a_i_c_0));
    CascadeMux I__300 (
            .O(N__2108),
            .I(N__2105));
    InMux I__299 (
            .O(N__2105),
            .I(N__2101));
    InMux I__298 (
            .O(N__2104),
            .I(N__2098));
    LocalMux I__297 (
            .O(N__2101),
            .I(cin_rZ0));
    LocalMux I__296 (
            .O(N__2098),
            .I(cin_rZ0));
    InMux I__295 (
            .O(N__2093),
            .I(N__2090));
    LocalMux I__294 (
            .O(N__2090),
            .I(N__2087));
    Odrv4 I__293 (
            .O(N__2087),
            .I(b_rZ0Z_0));
    IoInMux I__292 (
            .O(N__2084),
            .I(N__2081));
    LocalMux I__291 (
            .O(N__2081),
            .I(N__2078));
    Span4Mux_s0_h I__290 (
            .O(N__2078),
            .I(N__2075));
    Span4Mux_v I__289 (
            .O(N__2075),
            .I(N__2072));
    Span4Mux_v I__288 (
            .O(N__2072),
            .I(N__2069));
    Span4Mux_v I__287 (
            .O(N__2069),
            .I(N__2066));
    Odrv4 I__286 (
            .O(N__2066),
            .I(cout_o_c));
    InMux I__285 (
            .O(N__2063),
            .I(N__2060));
    LocalMux I__284 (
            .O(N__2060),
            .I(b_i_c_8));
    InMux I__283 (
            .O(N__2057),
            .I(N__2054));
    LocalMux I__282 (
            .O(N__2054),
            .I(N__2051));
    Sp12to4 I__281 (
            .O(N__2051),
            .I(N__2048));
    Span12Mux_v I__280 (
            .O(N__2048),
            .I(N__2045));
    Odrv12 I__279 (
            .O(N__2045),
            .I(b_i_c_2));
    CascadeMux I__278 (
            .O(N__2042),
            .I(N__2039));
    InMux I__277 (
            .O(N__2039),
            .I(N__2033));
    InMux I__276 (
            .O(N__2038),
            .I(N__2033));
    LocalMux I__275 (
            .O(N__2033),
            .I(b_rZ0Z_2));
    InMux I__274 (
            .O(N__2030),
            .I(N__2027));
    LocalMux I__273 (
            .O(N__2027),
            .I(N__2024));
    Span4Mux_v I__272 (
            .O(N__2024),
            .I(N__2021));
    Span4Mux_v I__271 (
            .O(N__2021),
            .I(N__2018));
    Span4Mux_v I__270 (
            .O(N__2018),
            .I(N__2015));
    Odrv4 I__269 (
            .O(N__2015),
            .I(a_i_c_11));
    InMux I__268 (
            .O(N__2012),
            .I(N__2009));
    LocalMux I__267 (
            .O(N__2009),
            .I(N__2006));
    IoSpan4Mux I__266 (
            .O(N__2006),
            .I(N__2003));
    IoSpan4Mux I__265 (
            .O(N__2003),
            .I(N__2000));
    Odrv4 I__264 (
            .O(N__2000),
            .I(a_i_c_12));
    InMux I__263 (
            .O(N__1997),
            .I(N__1994));
    LocalMux I__262 (
            .O(N__1994),
            .I(N__1991));
    Span4Mux_v I__261 (
            .O(N__1991),
            .I(N__1988));
    Span4Mux_v I__260 (
            .O(N__1988),
            .I(N__1985));
    Odrv4 I__259 (
            .O(N__1985),
            .I(b_i_c_12));
    InMux I__258 (
            .O(N__1982),
            .I(N__1979));
    LocalMux I__257 (
            .O(N__1979),
            .I(N__1976));
    Span4Mux_v I__256 (
            .O(N__1976),
            .I(N__1973));
    Span4Mux_v I__255 (
            .O(N__1973),
            .I(N__1970));
    Span4Mux_v I__254 (
            .O(N__1970),
            .I(N__1967));
    Odrv4 I__253 (
            .O(N__1967),
            .I(b_i_c_11));
    InMux I__252 (
            .O(N__1964),
            .I(N__1961));
    LocalMux I__251 (
            .O(N__1961),
            .I(b_rZ0Z_11));
    CascadeMux I__250 (
            .O(N__1958),
            .I(N__1955));
    InMux I__249 (
            .O(N__1955),
            .I(N__1952));
    LocalMux I__248 (
            .O(N__1952),
            .I(N__1949));
    Odrv4 I__247 (
            .O(N__1949),
            .I(m4_0));
    InMux I__246 (
            .O(N__1946),
            .I(N__1943));
    LocalMux I__245 (
            .O(N__1943),
            .I(N__1940));
    Sp12to4 I__244 (
            .O(N__1940),
            .I(N__1937));
    Span12Mux_v I__243 (
            .O(N__1937),
            .I(N__1934));
    Odrv12 I__242 (
            .O(N__1934),
            .I(b_i_c_10));
    IoInMux I__241 (
            .O(N__1931),
            .I(N__1928));
    LocalMux I__240 (
            .O(N__1928),
            .I(N__1925));
    IoSpan4Mux I__239 (
            .O(N__1925),
            .I(N__1922));
    Odrv4 I__238 (
            .O(N__1922),
            .I(sum_o_c_5));
    InMux I__237 (
            .O(N__1919),
            .I(N__1916));
    LocalMux I__236 (
            .O(N__1916),
            .I(N__1913));
    IoSpan4Mux I__235 (
            .O(N__1913),
            .I(N__1910));
    IoSpan4Mux I__234 (
            .O(N__1910),
            .I(N__1907));
    Odrv4 I__233 (
            .O(N__1907),
            .I(a_i_c_6));
    InMux I__232 (
            .O(N__1904),
            .I(N__1901));
    LocalMux I__231 (
            .O(N__1901),
            .I(a_i_c_8));
    IoInMux I__230 (
            .O(N__1898),
            .I(N__1895));
    LocalMux I__229 (
            .O(N__1895),
            .I(sum_o_c_14));
    IoInMux I__228 (
            .O(N__1892),
            .I(N__1889));
    LocalMux I__227 (
            .O(N__1889),
            .I(N__1886));
    Span4Mux_s0_h I__226 (
            .O(N__1886),
            .I(N__1883));
    Odrv4 I__225 (
            .O(N__1883),
            .I(sum_o_c_8));
    InMux I__224 (
            .O(N__1880),
            .I(N__1877));
    LocalMux I__223 (
            .O(N__1877),
            .I(N__1874));
    Sp12to4 I__222 (
            .O(N__1874),
            .I(N__1871));
    Span12Mux_v I__221 (
            .O(N__1871),
            .I(N__1868));
    Odrv12 I__220 (
            .O(N__1868),
            .I(b_i_c_3));
    InMux I__219 (
            .O(N__1865),
            .I(N__1862));
    LocalMux I__218 (
            .O(N__1862),
            .I(b_rZ0Z_3));
    InMux I__217 (
            .O(N__1859),
            .I(N__1856));
    LocalMux I__216 (
            .O(N__1856),
            .I(a_i_c_5));
    InMux I__215 (
            .O(N__1853),
            .I(N__1850));
    LocalMux I__214 (
            .O(N__1850),
            .I(b_rZ0Z_15));
    CascadeMux I__213 (
            .O(N__1847),
            .I(un68_sum_v_cascade_));
    IoInMux I__212 (
            .O(N__1844),
            .I(N__1841));
    LocalMux I__211 (
            .O(N__1841),
            .I(N__1838));
    Span4Mux_s0_h I__210 (
            .O(N__1838),
            .I(N__1835));
    Span4Mux_v I__209 (
            .O(N__1835),
            .I(N__1832));
    Span4Mux_v I__208 (
            .O(N__1832),
            .I(N__1829));
    Odrv4 I__207 (
            .O(N__1829),
            .I(sum_o_c_11));
    InMux I__206 (
            .O(N__1826),
            .I(N__1817));
    InMux I__205 (
            .O(N__1825),
            .I(N__1817));
    InMux I__204 (
            .O(N__1824),
            .I(N__1817));
    LocalMux I__203 (
            .O(N__1817),
            .I(b_rZ0Z_13));
    InMux I__202 (
            .O(N__1814),
            .I(N__1808));
    InMux I__201 (
            .O(N__1813),
            .I(N__1808));
    LocalMux I__200 (
            .O(N__1808),
            .I(b_rZ0Z_14));
    IoInMux I__199 (
            .O(N__1805),
            .I(N__1802));
    LocalMux I__198 (
            .O(N__1802),
            .I(N__1799));
    Span4Mux_s0_h I__197 (
            .O(N__1799),
            .I(N__1796));
    Sp12to4 I__196 (
            .O(N__1796),
            .I(N__1793));
    Odrv12 I__195 (
            .O(N__1793),
            .I(sum_o_c_10));
    IoInMux I__194 (
            .O(N__1790),
            .I(N__1787));
    LocalMux I__193 (
            .O(N__1787),
            .I(N__1784));
    Span4Mux_s0_h I__192 (
            .O(N__1784),
            .I(N__1781));
    Sp12to4 I__191 (
            .O(N__1781),
            .I(N__1778));
    Odrv12 I__190 (
            .O(N__1778),
            .I(sum_o_c_13));
    InMux I__189 (
            .O(N__1775),
            .I(N__1772));
    LocalMux I__188 (
            .O(N__1772),
            .I(a_i_c_1));
    InMux I__187 (
            .O(N__1769),
            .I(N__1766));
    LocalMux I__186 (
            .O(N__1766),
            .I(N__1763));
    Span4Mux_s3_h I__185 (
            .O(N__1763),
            .I(N__1760));
    Span4Mux_v I__184 (
            .O(N__1760),
            .I(N__1757));
    Sp12to4 I__183 (
            .O(N__1757),
            .I(N__1754));
    Span12Mux_v I__182 (
            .O(N__1754),
            .I(N__1751));
    Odrv12 I__181 (
            .O(N__1751),
            .I(b_i_c_4));
    InMux I__180 (
            .O(N__1748),
            .I(N__1745));
    LocalMux I__179 (
            .O(N__1745),
            .I(N__1742));
    Span12Mux_s3_h I__178 (
            .O(N__1742),
            .I(N__1739));
    Span12Mux_v I__177 (
            .O(N__1739),
            .I(N__1736));
    Odrv12 I__176 (
            .O(N__1736),
            .I(a_i_c_14));
    InMux I__175 (
            .O(N__1733),
            .I(N__1730));
    LocalMux I__174 (
            .O(N__1730),
            .I(N__1727));
    Sp12to4 I__173 (
            .O(N__1727),
            .I(N__1724));
    Span12Mux_v I__172 (
            .O(N__1724),
            .I(N__1721));
    Odrv12 I__171 (
            .O(N__1721),
            .I(b_i_c_14));
    InMux I__170 (
            .O(N__1718),
            .I(N__1715));
    LocalMux I__169 (
            .O(N__1715),
            .I(b_i_c_0));
    InMux I__168 (
            .O(N__1712),
            .I(N__1709));
    LocalMux I__167 (
            .O(N__1709),
            .I(N__1706));
    Span4Mux_v I__166 (
            .O(N__1706),
            .I(N__1703));
    Span4Mux_v I__165 (
            .O(N__1703),
            .I(N__1700));
    Span4Mux_v I__164 (
            .O(N__1700),
            .I(N__1697));
    Odrv4 I__163 (
            .O(N__1697),
            .I(b_i_c_13));
    InMux I__162 (
            .O(N__1694),
            .I(N__1691));
    LocalMux I__161 (
            .O(N__1691),
            .I(a_i_c_9));
    InMux I__160 (
            .O(N__1688),
            .I(N__1685));
    LocalMux I__159 (
            .O(N__1685),
            .I(N__1682));
    Span4Mux_v I__158 (
            .O(N__1682),
            .I(N__1679));
    Span4Mux_v I__157 (
            .O(N__1679),
            .I(N__1676));
    Span4Mux_v I__156 (
            .O(N__1676),
            .I(N__1673));
    Odrv4 I__155 (
            .O(N__1673),
            .I(b_i_c_15));
    IoInMux I__154 (
            .O(N__1670),
            .I(N__1667));
    LocalMux I__153 (
            .O(N__1667),
            .I(N__1664));
    Span4Mux_s0_h I__152 (
            .O(N__1664),
            .I(N__1661));
    Sp12to4 I__151 (
            .O(N__1661),
            .I(N__1658));
    Odrv12 I__150 (
            .O(N__1658),
            .I(sum_o_c_12));
    IoInMux I__149 (
            .O(N__1655),
            .I(N__1652));
    LocalMux I__148 (
            .O(N__1652),
            .I(N__1649));
    IoSpan4Mux I__147 (
            .O(N__1649),
            .I(N__1646));
    IoSpan4Mux I__146 (
            .O(N__1646),
            .I(N__1643));
    Odrv4 I__145 (
            .O(N__1643),
            .I(sum_o_c_9));
    InMux I__144 (
            .O(N__1640),
            .I(N__1637));
    LocalMux I__143 (
            .O(N__1637),
            .I(N__1634));
    Sp12to4 I__142 (
            .O(N__1634),
            .I(N__1631));
    Span12Mux_v I__141 (
            .O(N__1631),
            .I(N__1628));
    Odrv12 I__140 (
            .O(N__1628),
            .I(a_i_c_15));
    defparam IN_MUX_bfv_2_16_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_16_0_));
    defparam IN_MUX_bfv_2_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_17_0_ (
            .carryinitin(un5_sum_v_cry_6),
            .carryinitout(bfn_2_17_0_));
    defparam IN_MUX_bfv_2_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_18_0_ (
            .carryinitin(un5_sum_v_cry_14),
            .carryinitout(bfn_2_18_0_));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam a_r_15_LC_1_14_7.C_ON=1'b0;
    defparam a_r_15_LC_1_14_7.SEQ_MODE=4'b1000;
    defparam a_r_15_LC_1_14_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 a_r_15_LC_1_14_7 (
            .in0(N__1640),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(a_rZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3152),
            .ce(),
            .sr(_gnd_net_));
    defparam b_r_4_LC_1_15_0.C_ON=1'b0;
    defparam b_r_4_LC_1_15_0.SEQ_MODE=4'b1000;
    defparam b_r_4_LC_1_15_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 b_r_4_LC_1_15_0 (
            .in0(N__1769),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(b_rZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3148),
            .ce(),
            .sr(_gnd_net_));
    defparam a_r_14_LC_1_15_1.C_ON=1'b0;
    defparam a_r_14_LC_1_15_1.SEQ_MODE=4'b1000;
    defparam a_r_14_LC_1_15_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 a_r_14_LC_1_15_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1748),
            .lcout(a_rZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3148),
            .ce(),
            .sr(_gnd_net_));
    defparam b_r_14_LC_1_15_2.C_ON=1'b0;
    defparam b_r_14_LC_1_15_2.SEQ_MODE=4'b1000;
    defparam b_r_14_LC_1_15_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 b_r_14_LC_1_15_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1733),
            .lcout(b_rZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3148),
            .ce(),
            .sr(_gnd_net_));
    defparam b_r_0_LC_1_15_4.C_ON=1'b0;
    defparam b_r_0_LC_1_15_4.SEQ_MODE=4'b1000;
    defparam b_r_0_LC_1_15_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 b_r_0_LC_1_15_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1718),
            .lcout(b_rZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3148),
            .ce(),
            .sr(_gnd_net_));
    defparam b_r_13_LC_1_15_5.C_ON=1'b0;
    defparam b_r_13_LC_1_15_5.SEQ_MODE=4'b1000;
    defparam b_r_13_LC_1_15_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 b_r_13_LC_1_15_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1712),
            .lcout(b_rZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3148),
            .ce(),
            .sr(_gnd_net_));
    defparam a_r_9_LC_1_15_6.C_ON=1'b0;
    defparam a_r_9_LC_1_15_6.SEQ_MODE=4'b1000;
    defparam a_r_9_LC_1_15_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 a_r_9_LC_1_15_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1694),
            .lcout(a_rZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3148),
            .ce(),
            .sr(_gnd_net_));
    defparam b_r_15_LC_1_15_7.C_ON=1'b0;
    defparam b_r_15_LC_1_15_7.SEQ_MODE=4'b1000;
    defparam b_r_15_LC_1_15_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 b_r_15_LC_1_15_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1688),
            .lcout(b_rZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3148),
            .ce(),
            .sr(_gnd_net_));
    defparam sum_r_12_LC_1_16_0.C_ON=1'b0;
    defparam sum_r_12_LC_1_16_0.SEQ_MODE=4'b1000;
    defparam sum_r_12_LC_1_16_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sum_r_12_LC_1_16_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2452),
            .lcout(sum_o_c_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3145),
            .ce(),
            .sr(_gnd_net_));
    defparam sum_r_9_LC_1_16_1.C_ON=1'b0;
    defparam sum_r_9_LC_1_16_1.SEQ_MODE=4'b1000;
    defparam sum_r_9_LC_1_16_1.LUT_INIT=16'b1001011001101001;
    LogicCell40 sum_r_9_LC_1_16_1 (
            .in0(N__2451),
            .in1(N__2515),
            .in2(N__2486),
            .in3(N__2585),
            .lcout(sum_o_c_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3145),
            .ce(),
            .sr(_gnd_net_));
    defparam a_r_5_LC_1_16_2.C_ON=1'b0;
    defparam a_r_5_LC_1_16_2.SEQ_MODE=4'b1000;
    defparam a_r_5_LC_1_16_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 a_r_5_LC_1_16_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1859),
            .lcout(a_rZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3145),
            .ce(),
            .sr(_gnd_net_));
    defparam b_r_RNI0TDJ1_15_LC_1_16_3.C_ON=1'b0;
    defparam b_r_RNI0TDJ1_15_LC_1_16_3.SEQ_MODE=4'b0000;
    defparam b_r_RNI0TDJ1_15_LC_1_16_3.LUT_INIT=16'b1111111111101110;
    LogicCell40 b_r_RNI0TDJ1_15_LC_1_16_3 (
            .in0(N__1826),
            .in1(N__1853),
            .in2(N__2396),
            .in3(N__1814),
            .lcout(b_r_RNI0TDJ1Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sum_r_RNO_1_11_LC_1_16_4.C_ON=1'b0;
    defparam sum_r_RNO_1_11_LC_1_16_4.SEQ_MODE=4'b0000;
    defparam sum_r_RNO_1_11_LC_1_16_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 sum_r_RNO_1_11_LC_1_16_4 (
            .in0(N__2514),
            .in1(N__2481),
            .in2(_gnd_net_),
            .in3(N__2450),
            .lcout(),
            .ltout(un68_sum_v_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sum_r_11_LC_1_16_5.C_ON=1'b0;
    defparam sum_r_11_LC_1_16_5.SEQ_MODE=4'b1000;
    defparam sum_r_11_LC_1_16_5.LUT_INIT=16'b1111100000000000;
    LogicCell40 sum_r_11_LC_1_16_5 (
            .in0(N__2584),
            .in1(N__2564),
            .in2(N__1847),
            .in3(N__2525),
            .lcout(sum_o_c_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3145),
            .ce(),
            .sr(_gnd_net_));
    defparam b_r_sbtinv_13_LC_1_16_6.C_ON=1'b0;
    defparam b_r_sbtinv_13_LC_1_16_6.SEQ_MODE=4'b0000;
    defparam b_r_sbtinv_13_LC_1_16_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 b_r_sbtinv_13_LC_1_16_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1824),
            .lcout(b_r_i_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam b_r_RNIEIE51_14_LC_1_16_7.C_ON=1'b0;
    defparam b_r_RNIEIE51_14_LC_1_16_7.SEQ_MODE=4'b0000;
    defparam b_r_RNIEIE51_14_LC_1_16_7.LUT_INIT=16'b1010101001010101;
    LogicCell40 b_r_RNIEIE51_14_LC_1_16_7 (
            .in0(N__1825),
            .in1(N__2422),
            .in2(_gnd_net_),
            .in3(N__1813),
            .lcout(b_r_RNIEIE51Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sum_r_10_LC_1_17_0.C_ON=1'b0;
    defparam sum_r_10_LC_1_17_0.SEQ_MODE=4'b1000;
    defparam sum_r_10_LC_1_17_0.LUT_INIT=16'b0110110011000110;
    LogicCell40 sum_r_10_LC_1_17_0 (
            .in0(N__2583),
            .in1(N__2563),
            .in2(N__1958),
            .in3(N__2453),
            .lcout(sum_o_c_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3144),
            .ce(),
            .sr(_gnd_net_));
    defparam sum_r_13_LC_1_17_1.C_ON=1'b0;
    defparam sum_r_13_LC_1_17_1.SEQ_MODE=4'b1000;
    defparam sum_r_13_LC_1_17_1.LUT_INIT=16'b1010010110100101;
    LogicCell40 sum_r_13_LC_1_17_1 (
            .in0(N__2876),
            .in1(_gnd_net_),
            .in2(N__2861),
            .in3(_gnd_net_),
            .lcout(sum_o_c_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3144),
            .ce(),
            .sr(_gnd_net_));
    defparam a_r_1_LC_1_17_2.C_ON=1'b0;
    defparam a_r_1_LC_1_17_2.SEQ_MODE=4'b1000;
    defparam a_r_1_LC_1_17_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 a_r_1_LC_1_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1775),
            .lcout(a_rZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3144),
            .ce(),
            .sr(_gnd_net_));
    defparam b_r_RNILOR9_2_LC_1_17_3.C_ON=1'b0;
    defparam b_r_RNILOR9_2_LC_1_17_3.SEQ_MODE=4'b0000;
    defparam b_r_RNILOR9_2_LC_1_17_3.LUT_INIT=16'b1100110000110011;
    LogicCell40 b_r_RNILOR9_2_LC_1_17_3 (
            .in0(N__3014),
            .in1(N__2677),
            .in2(_gnd_net_),
            .in3(N__2038),
            .lcout(b_r_RNILOR9Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam b_r_RNIKF8B_3_LC_1_17_4.C_ON=1'b0;
    defparam b_r_RNIKF8B_3_LC_1_17_4.SEQ_MODE=4'b0000;
    defparam b_r_RNIKF8B_3_LC_1_17_4.LUT_INIT=16'b1111111111111010;
    LogicCell40 b_r_RNIKF8B_3_LC_1_17_4 (
            .in0(N__2678),
            .in1(N__3215),
            .in2(N__2042),
            .in3(N__1865),
            .lcout(b_r_RNIKF8BZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sum_r_5_LC_1_17_5.C_ON=1'b0;
    defparam sum_r_5_LC_1_17_5.SEQ_MODE=4'b1000;
    defparam sum_r_5_LC_1_17_5.LUT_INIT=16'b1001011001101001;
    LogicCell40 sum_r_5_LC_1_17_5 (
            .in0(N__2771),
            .in1(N__2920),
            .in2(N__2798),
            .in3(N__2752),
            .lcout(sum_o_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3144),
            .ce(),
            .sr(_gnd_net_));
    defparam a_r_6_LC_1_17_6.C_ON=1'b0;
    defparam a_r_6_LC_1_17_6.SEQ_MODE=4'b1000;
    defparam a_r_6_LC_1_17_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 a_r_6_LC_1_17_6 (
            .in0(N__1919),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(a_rZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3144),
            .ce(),
            .sr(_gnd_net_));
    defparam b_r_sbtinv_1_LC_1_17_7.C_ON=1'b0;
    defparam b_r_sbtinv_1_LC_1_17_7.SEQ_MODE=4'b0000;
    defparam b_r_sbtinv_1_LC_1_17_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 b_r_sbtinv_1_LC_1_17_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2676),
            .lcout(b_r_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam a_r_8_LC_1_18_0.C_ON=1'b0;
    defparam a_r_8_LC_1_18_0.SEQ_MODE=4'b1000;
    defparam a_r_8_LC_1_18_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 a_r_8_LC_1_18_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1904),
            .lcout(a_rZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3146),
            .ce(),
            .sr(_gnd_net_));
    defparam sum_r_14_LC_1_18_1.C_ON=1'b0;
    defparam sum_r_14_LC_1_18_1.SEQ_MODE=4'b1000;
    defparam sum_r_14_LC_1_18_1.LUT_INIT=16'b1010010111110000;
    LogicCell40 sum_r_14_LC_1_18_1 (
            .in0(N__2875),
            .in1(_gnd_net_),
            .in2(N__2840),
            .in3(N__2860),
            .lcout(sum_o_c_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3146),
            .ce(),
            .sr(_gnd_net_));
    defparam sum_r_8_LC_1_18_2.C_ON=1'b0;
    defparam sum_r_8_LC_1_18_2.SEQ_MODE=4'b1000;
    defparam sum_r_8_LC_1_18_2.LUT_INIT=16'b1100110011001100;
    LogicCell40 sum_r_8_LC_1_18_2 (
            .in0(_gnd_net_),
            .in1(N__2753),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sum_o_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3146),
            .ce(),
            .sr(_gnd_net_));
    defparam b_r_3_LC_1_18_3.C_ON=1'b0;
    defparam b_r_3_LC_1_18_3.SEQ_MODE=4'b1000;
    defparam b_r_3_LC_1_18_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 b_r_3_LC_1_18_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1880),
            .lcout(b_rZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3146),
            .ce(),
            .sr(_gnd_net_));
    defparam cout_r_LC_1_18_4.C_ON=1'b0;
    defparam cout_r_LC_1_18_4.SEQ_MODE=4'b1000;
    defparam cout_r_LC_1_18_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 cout_r_LC_1_18_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2874),
            .lcout(cout_o_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3146),
            .ce(),
            .sr(_gnd_net_));
    defparam b_r_8_LC_1_18_5.C_ON=1'b0;
    defparam b_r_8_LC_1_18_5.SEQ_MODE=4'b1000;
    defparam b_r_8_LC_1_18_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 b_r_8_LC_1_18_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2063),
            .lcout(b_rZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3146),
            .ce(),
            .sr(_gnd_net_));
    defparam b_r_2_LC_1_18_6.C_ON=1'b0;
    defparam b_r_2_LC_1_18_6.SEQ_MODE=4'b1000;
    defparam b_r_2_LC_1_18_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 b_r_2_LC_1_18_6 (
            .in0(N__2057),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(b_rZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3146),
            .ce(),
            .sr(_gnd_net_));
    defparam b_r_RNI95R61_11_LC_1_18_7.C_ON=1'b0;
    defparam b_r_RNI95R61_11_LC_1_18_7.SEQ_MODE=4'b0000;
    defparam b_r_RNI95R61_11_LC_1_18_7.LUT_INIT=16'b1111111111111100;
    LogicCell40 b_r_RNI95R61_11_LC_1_18_7 (
            .in0(N__2548),
            .in1(N__2615),
            .in2(N__2720),
            .in3(N__1964),
            .lcout(b_r_RNI95R61Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam a_r_11_LC_1_19_0.C_ON=1'b0;
    defparam a_r_11_LC_1_19_0.SEQ_MODE=4'b1000;
    defparam a_r_11_LC_1_19_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 a_r_11_LC_1_19_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2030),
            .lcout(a_rZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3149),
            .ce(),
            .sr(_gnd_net_));
    defparam a_r_12_LC_1_19_1.C_ON=1'b0;
    defparam a_r_12_LC_1_19_1.SEQ_MODE=4'b1000;
    defparam a_r_12_LC_1_19_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 a_r_12_LC_1_19_1 (
            .in0(N__2012),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(a_rZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3149),
            .ce(),
            .sr(_gnd_net_));
    defparam b_r_12_LC_1_19_2.C_ON=1'b0;
    defparam b_r_12_LC_1_19_2.SEQ_MODE=4'b1000;
    defparam b_r_12_LC_1_19_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 b_r_12_LC_1_19_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1997),
            .lcout(b_rZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3149),
            .ce(),
            .sr(_gnd_net_));
    defparam b_r_11_LC_1_19_3.C_ON=1'b0;
    defparam b_r_11_LC_1_19_3.SEQ_MODE=4'b1000;
    defparam b_r_11_LC_1_19_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 b_r_11_LC_1_19_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1982),
            .lcout(b_rZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3149),
            .ce(),
            .sr(_gnd_net_));
    defparam sum_r_RNO_0_10_LC_1_19_4.C_ON=1'b0;
    defparam sum_r_RNO_0_10_LC_1_19_4.SEQ_MODE=4'b0000;
    defparam sum_r_RNO_0_10_LC_1_19_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 sum_r_RNO_0_10_LC_1_19_4 (
            .in0(_gnd_net_),
            .in1(N__2505),
            .in2(_gnd_net_),
            .in3(N__2472),
            .lcout(m4_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam b_r_10_LC_1_19_7.C_ON=1'b0;
    defparam b_r_10_LC_1_19_7.SEQ_MODE=4'b1000;
    defparam b_r_10_LC_1_19_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 b_r_10_LC_1_19_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1946),
            .lcout(b_rZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3149),
            .ce(),
            .sr(_gnd_net_));
    defparam cin_r_LC_2_15_0.C_ON=1'b0;
    defparam cin_r_LC_2_15_0.SEQ_MODE=4'b1000;
    defparam cin_r_LC_2_15_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 cin_r_LC_2_15_0 (
            .in0(N__2198),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(cin_rZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3153),
            .ce(),
            .sr(_gnd_net_));
    defparam sum_r_3_LC_2_15_1.C_ON=1'b0;
    defparam sum_r_3_LC_2_15_1.SEQ_MODE=4'b1000;
    defparam sum_r_3_LC_2_15_1.LUT_INIT=16'b1100110010000000;
    LogicCell40 sum_r_3_LC_2_15_1 (
            .in0(N__2282),
            .in1(N__2261),
            .in2(N__2315),
            .in3(N__2144),
            .lcout(sum_o_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3153),
            .ce(),
            .sr(_gnd_net_));
    defparam sum_r_1_LC_2_15_2.C_ON=1'b0;
    defparam sum_r_1_LC_2_15_2.SEQ_MODE=4'b1000;
    defparam sum_r_1_LC_2_15_2.LUT_INIT=16'b1001011001101001;
    LogicCell40 sum_r_1_LC_2_15_2 (
            .in0(N__2230),
            .in1(N__3061),
            .in2(N__2314),
            .in3(N__2251),
            .lcout(sum_o_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3153),
            .ce(),
            .sr(_gnd_net_));
    defparam sum_r_4_LC_2_15_3.C_ON=1'b0;
    defparam sum_r_4_LC_2_15_3.SEQ_MODE=4'b1000;
    defparam sum_r_4_LC_2_15_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sum_r_4_LC_2_15_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2231),
            .lcout(sum_o_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3153),
            .ce(),
            .sr(_gnd_net_));
    defparam b_r_RNIS0O01_4_LC_2_15_5.C_ON=1'b0;
    defparam b_r_RNIS0O01_4_LC_2_15_5.SEQ_MODE=4'b0000;
    defparam b_r_RNIS0O01_4_LC_2_15_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 b_r_RNIS0O01_4_LC_2_15_5 (
            .in0(N__3060),
            .in1(N__2250),
            .in2(_gnd_net_),
            .in3(N__2229),
            .lcout(un13_sum_v),
            .ltout(un13_sum_v_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sum_r_2_LC_2_15_6.C_ON=1'b0;
    defparam sum_r_2_LC_2_15_6.SEQ_MODE=4'b1000;
    defparam sum_r_2_LC_2_15_6.LUT_INIT=16'b1111010100001010;
    LogicCell40 sum_r_2_LC_2_15_6 (
            .in0(N__2310),
            .in1(_gnd_net_),
            .in2(N__2138),
            .in3(N__2281),
            .lcout(sum_o_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3153),
            .ce(),
            .sr(_gnd_net_));
    defparam a_r_0_LC_2_15_7.C_ON=1'b0;
    defparam a_r_0_LC_2_15_7.SEQ_MODE=4'b1000;
    defparam a_r_0_LC_2_15_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 a_r_0_LC_2_15_7 (
            .in0(N__2120),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(a_rZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3153),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sum_v_cry_0_c_THRU_CRY_0_LC_2_16_0.C_ON=1'b1;
    defparam un5_sum_v_cry_0_c_THRU_CRY_0_LC_2_16_0.SEQ_MODE=4'b0000;
    defparam un5_sum_v_cry_0_c_THRU_CRY_0_LC_2_16_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un5_sum_v_cry_0_c_THRU_CRY_0_LC_2_16_0 (
            .in0(_gnd_net_),
            .in1(N__2104),
            .in2(N__2108),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_16_0_),
            .carryout(un5_sum_v_cry_0_c_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sum_r_0_LC_2_16_1.C_ON=1'b1;
    defparam sum_r_0_LC_2_16_1.SEQ_MODE=4'b1000;
    defparam sum_r_0_LC_2_16_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 sum_r_0_LC_2_16_1 (
            .in0(_gnd_net_),
            .in1(N__2093),
            .in2(N__2357),
            .in3(N__2333),
            .lcout(sum_o_c_0),
            .ltout(),
            .carryin(un5_sum_v_cry_0_c_THRU_CO),
            .carryout(un5_sum_v_cry_0),
            .clk(N__3150),
            .ce(),
            .sr(_gnd_net_));
    defparam b_r_sbtinv_RNIB4UQ_1_LC_2_16_2.C_ON=1'b1;
    defparam b_r_sbtinv_RNIB4UQ_1_LC_2_16_2.SEQ_MODE=4'b0000;
    defparam b_r_sbtinv_RNIB4UQ_1_LC_2_16_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 b_r_sbtinv_RNIB4UQ_1_LC_2_16_2 (
            .in0(_gnd_net_),
            .in1(N__2330),
            .in2(N__2324),
            .in3(N__2294),
            .lcout(b_r_sbtinv_RNIB4UQZ0Z_1),
            .ltout(),
            .carryin(un5_sum_v_cry_0),
            .carryout(un5_sum_v_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sum_v_cry_1_c_RNIHJL01_LC_2_16_3.C_ON=1'b1;
    defparam un5_sum_v_cry_1_c_RNIHJL01_LC_2_16_3.SEQ_MODE=4'b0000;
    defparam un5_sum_v_cry_1_c_RNIHJL01_LC_2_16_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_sum_v_cry_1_c_RNIHJL01_LC_2_16_3 (
            .in0(_gnd_net_),
            .in1(N__3013),
            .in2(N__2291),
            .in3(N__2273),
            .lcout(un5_sum_v_cry_1_c_RNIHJLZ0Z01),
            .ltout(),
            .carryin(un5_sum_v_cry_1),
            .carryout(un5_sum_v_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sum_r_RNO_0_3_LC_2_16_4.C_ON=1'b1;
    defparam sum_r_RNO_0_3_LC_2_16_4.SEQ_MODE=4'b0000;
    defparam sum_r_RNO_0_3_LC_2_16_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 sum_r_RNO_0_3_LC_2_16_4 (
            .in0(_gnd_net_),
            .in1(N__3211),
            .in2(N__2270),
            .in3(N__2255),
            .lcout(sum_r_RNO_0Z0Z_3),
            .ltout(),
            .carryin(un5_sum_v_cry_2),
            .carryout(un5_sum_v_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sum_v_cry_3_c_RNIVN8O_LC_2_16_5.C_ON=1'b1;
    defparam un5_sum_v_cry_3_c_RNIVN8O_LC_2_16_5.SEQ_MODE=4'b0000;
    defparam un5_sum_v_cry_3_c_RNIVN8O_LC_2_16_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_sum_v_cry_3_c_RNIVN8O_LC_2_16_5 (
            .in0(_gnd_net_),
            .in1(N__3062),
            .in2(N__2252),
            .in3(N__2219),
            .lcout(un5_sum_v_cry_3_c_RNIVN8OZ0),
            .ltout(),
            .carryin(un5_sum_v_cry_3),
            .carryout(un5_sum_v_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam b_r_sbtinv_RNINK2R_5_LC_2_16_6.C_ON=1'b1;
    defparam b_r_sbtinv_RNINK2R_5_LC_2_16_6.SEQ_MODE=4'b0000;
    defparam b_r_sbtinv_RNINK2R_5_LC_2_16_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 b_r_sbtinv_RNINK2R_5_LC_2_16_6 (
            .in0(_gnd_net_),
            .in1(N__2216),
            .in2(N__3038),
            .in3(N__2210),
            .lcout(b_r_sbtinv_RNINK2RZ0Z_5),
            .ltout(),
            .carryin(un5_sum_v_cry_4),
            .carryout(un5_sum_v_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sum_v_cry_5_c_RNI5CQ01_LC_2_16_7.C_ON=1'b1;
    defparam un5_sum_v_cry_5_c_RNI5CQ01_LC_2_16_7.SEQ_MODE=4'b0000;
    defparam un5_sum_v_cry_5_c_RNI5CQ01_LC_2_16_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_sum_v_cry_5_c_RNI5CQ01_LC_2_16_7 (
            .in0(_gnd_net_),
            .in1(N__2965),
            .in2(N__2954),
            .in3(N__2207),
            .lcout(un5_sum_v_cry_5_c_RNI5CQZ0Z01),
            .ltout(),
            .carryin(un5_sum_v_cry_5),
            .carryout(un5_sum_v_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sum_r_RNO_0_7_LC_2_17_0.C_ON=1'b1;
    defparam sum_r_RNO_0_7_LC_2_17_0.SEQ_MODE=4'b0000;
    defparam sum_r_RNO_0_7_LC_2_17_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 sum_r_RNO_0_7_LC_2_17_0 (
            .in0(_gnd_net_),
            .in1(N__2995),
            .in2(N__2978),
            .in3(N__2204),
            .lcout(sum_r_RNO_0Z0Z_7),
            .ltout(),
            .carryin(bfn_2_17_0_),
            .carryout(un5_sum_v_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sum_v_cry_7_c_RNIB8DO_LC_2_17_1.C_ON=1'b1;
    defparam un5_sum_v_cry_7_c_RNIB8DO_LC_2_17_1.SEQ_MODE=4'b0000;
    defparam un5_sum_v_cry_7_c_RNIB8DO_LC_2_17_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_sum_v_cry_7_c_RNIB8DO_LC_2_17_1 (
            .in0(_gnd_net_),
            .in1(N__2769),
            .in2(N__2797),
            .in3(N__2201),
            .lcout(un5_sum_v_cry_7_c_RNIB8DOZ0),
            .ltout(),
            .carryin(un5_sum_v_cry_7),
            .carryout(un5_sum_v_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam b_r_sbtinv_RNI357R_9_LC_2_17_2.C_ON=1'b1;
    defparam b_r_sbtinv_RNI357R_9_LC_2_17_2.SEQ_MODE=4'b0000;
    defparam b_r_sbtinv_RNI357R_9_LC_2_17_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 b_r_sbtinv_RNI357R_9_LC_2_17_2 (
            .in0(_gnd_net_),
            .in1(N__2597),
            .in2(N__2666),
            .in3(N__2567),
            .lcout(b_r_sbtinv_RNI357RZ0Z_9),
            .ltout(),
            .carryin(un5_sum_v_cry_8),
            .carryout(un5_sum_v_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sum_v_cry_9_c_RNIEOBI1_LC_2_17_3.C_ON=1'b1;
    defparam un5_sum_v_cry_9_c_RNIEOBI1_LC_2_17_3.SEQ_MODE=4'b0000;
    defparam un5_sum_v_cry_9_c_RNIEOBI1_LC_2_17_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_sum_v_cry_9_c_RNIEOBI1_LC_2_17_3 (
            .in0(_gnd_net_),
            .in1(N__2645),
            .in2(N__2702),
            .in3(N__2552),
            .lcout(un5_sum_v_cry_9_c_RNIEOBIZ0Z1),
            .ltout(),
            .carryin(un5_sum_v_cry_9),
            .carryout(un5_sum_v_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sum_r_RNO_0_11_LC_2_17_4.C_ON=1'b1;
    defparam sum_r_RNO_0_11_LC_2_17_4.SEQ_MODE=4'b0000;
    defparam sum_r_RNO_0_11_LC_2_17_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 sum_r_RNO_0_11_LC_2_17_4 (
            .in0(_gnd_net_),
            .in1(N__2549),
            .in2(N__2534),
            .in3(N__2519),
            .lcout(sum_r_RNO_0Z0Z_11),
            .ltout(),
            .carryin(un5_sum_v_cry_10),
            .carryout(un5_sum_v_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sum_v_cry_11_c_RNICJ0T_LC_2_17_5.C_ON=1'b1;
    defparam un5_sum_v_cry_11_c_RNICJ0T_LC_2_17_5.SEQ_MODE=4'b0000;
    defparam un5_sum_v_cry_11_c_RNICJ0T_LC_2_17_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_sum_v_cry_11_c_RNICJ0T_LC_2_17_5 (
            .in0(_gnd_net_),
            .in1(N__2516),
            .in2(N__2485),
            .in3(N__2435),
            .lcout(un5_sum_v_cry_11_c_RNICJ0TZ0),
            .ltout(),
            .carryin(un5_sum_v_cry_11),
            .carryout(un5_sum_v_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sum_v_cry_12_c_RNI45JO_LC_2_17_6.C_ON=1'b1;
    defparam un5_sum_v_cry_12_c_RNI45JO_LC_2_17_6.SEQ_MODE=4'b0000;
    defparam un5_sum_v_cry_12_c_RNI45JO_LC_2_17_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_sum_v_cry_12_c_RNI45JO_LC_2_17_6 (
            .in0(_gnd_net_),
            .in1(N__2432),
            .in2(N__3089),
            .in3(N__2426),
            .lcout(un5_sum_v_cry_12_c_RNI45JOZ0),
            .ltout(),
            .carryin(un5_sum_v_cry_12),
            .carryout(un5_sum_v_cry_13),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sum_v_cry_13_c_RNIG5IK1_LC_2_17_7.C_ON=1'b1;
    defparam un5_sum_v_cry_13_c_RNIG5IK1_LC_2_17_7.SEQ_MODE=4'b0000;
    defparam un5_sum_v_cry_13_c_RNIG5IK1_LC_2_17_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_sum_v_cry_13_c_RNIG5IK1_LC_2_17_7 (
            .in0(_gnd_net_),
            .in1(N__2423),
            .in2(N__2408),
            .in3(N__2399),
            .lcout(un5_sum_v_cry_13_c_RNIG5IKZ0Z1),
            .ltout(),
            .carryin(un5_sum_v_cry_13),
            .carryout(un5_sum_v_cry_14),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sum_r_RNO_0_15_LC_2_18_0.C_ON=1'b1;
    defparam sum_r_RNO_0_15_LC_2_18_0.SEQ_MODE=4'b0000;
    defparam sum_r_RNO_0_15_LC_2_18_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 sum_r_RNO_0_15_LC_2_18_0 (
            .in0(_gnd_net_),
            .in1(N__2395),
            .in2(N__2372),
            .in3(N__2360),
            .lcout(sum_r_RNO_0Z0Z_15),
            .ltout(),
            .carryin(bfn_2_18_0_),
            .carryout(un5_sum_v_cry_15),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sum_v_cry_15_THRU_LUT4_0_LC_2_18_1.C_ON=1'b0;
    defparam un5_sum_v_cry_15_THRU_LUT4_0_LC_2_18_1.SEQ_MODE=4'b0000;
    defparam un5_sum_v_cry_15_THRU_LUT4_0_LC_2_18_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 un5_sum_v_cry_15_THRU_LUT4_0_LC_2_18_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2879),
            .lcout(un5_sum_v_cry_15_THRU_CO),
            .ltout(un5_sum_v_cry_15_THRU_CO_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sum_r_15_LC_2_18_2.C_ON=1'b0;
    defparam sum_r_15_LC_2_18_2.SEQ_MODE=4'b1000;
    defparam sum_r_15_LC_2_18_2.LUT_INIT=16'b1111100000000000;
    LogicCell40 sum_r_15_LC_2_18_2 (
            .in0(N__2859),
            .in1(N__2836),
            .in2(N__2825),
            .in3(N__2822),
            .lcout(sum_o_c_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3151),
            .ce(),
            .sr(_gnd_net_));
    defparam b_r_RNIGPS01_8_LC_2_18_3.C_ON=1'b0;
    defparam b_r_RNIGPS01_8_LC_2_18_3.SEQ_MODE=4'b0000;
    defparam b_r_RNIGPS01_8_LC_2_18_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 b_r_RNIGPS01_8_LC_2_18_3 (
            .in0(N__2793),
            .in1(N__2770),
            .in2(_gnd_net_),
            .in3(N__2751),
            .lcout(un40_sum_v),
            .ltout(un40_sum_v_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sum_r_6_LC_2_18_4.C_ON=1'b0;
    defparam sum_r_6_LC_2_18_4.SEQ_MODE=4'b1000;
    defparam sum_r_6_LC_2_18_4.LUT_INIT=16'b1111001100001100;
    LogicCell40 sum_r_6_LC_2_18_4 (
            .in0(_gnd_net_),
            .in1(N__2919),
            .in2(N__2735),
            .in3(N__2945),
            .lcout(sum_o_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3151),
            .ce(),
            .sr(_gnd_net_));
    defparam b_r_RNIRURO_10_LC_2_18_5.C_ON=1'b0;
    defparam b_r_RNIRURO_10_LC_2_18_5.SEQ_MODE=4'b0000;
    defparam b_r_RNIRURO_10_LC_2_18_5.LUT_INIT=16'b1010101001010101;
    LogicCell40 b_r_RNIRURO_10_LC_2_18_5 (
            .in0(N__2614),
            .in1(N__2644),
            .in2(_gnd_net_),
            .in3(N__2713),
            .lcout(b_r_RNIRUROZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam b_r_1_LC_2_18_6.C_ON=1'b0;
    defparam b_r_1_LC_2_18_6.SEQ_MODE=4'b1000;
    defparam b_r_1_LC_2_18_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 b_r_1_LC_2_18_6 (
            .in0(N__2693),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(b_rZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3151),
            .ce(),
            .sr(_gnd_net_));
    defparam b_r_sbtinv_9_LC_2_18_7.C_ON=1'b0;
    defparam b_r_sbtinv_9_LC_2_18_7.SEQ_MODE=4'b0000;
    defparam b_r_sbtinv_9_LC_2_18_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 b_r_sbtinv_9_LC_2_18_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2613),
            .lcout(b_r_i_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam a_r_10_LC_2_19_0.C_ON=1'b0;
    defparam a_r_10_LC_2_19_0.SEQ_MODE=4'b1000;
    defparam a_r_10_LC_2_19_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 a_r_10_LC_2_19_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2657),
            .lcout(a_rZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3154),
            .ce(),
            .sr(_gnd_net_));
    defparam b_r_9_LC_2_19_2.C_ON=1'b0;
    defparam b_r_9_LC_2_19_2.SEQ_MODE=4'b1000;
    defparam b_r_9_LC_2_19_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 b_r_9_LC_2_19_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2630),
            .lcout(b_rZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3154),
            .ce(),
            .sr(_gnd_net_));
    defparam a_r_7_LC_2_19_4.C_ON=1'b0;
    defparam a_r_7_LC_2_19_4.SEQ_MODE=4'b1000;
    defparam a_r_7_LC_2_19_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 a_r_7_LC_2_19_4 (
            .in0(N__3113),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(a_rZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3154),
            .ce(),
            .sr(_gnd_net_));
    defparam a_r_13_LC_2_19_5.C_ON=1'b0;
    defparam a_r_13_LC_2_19_5.SEQ_MODE=4'b1000;
    defparam a_r_13_LC_2_19_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 a_r_13_LC_2_19_5 (
            .in0(N__3101),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(a_rZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3154),
            .ce(),
            .sr(_gnd_net_));
    defparam a_r_4_LC_2_19_7.C_ON=1'b0;
    defparam a_r_4_LC_2_19_7.SEQ_MODE=4'b1000;
    defparam a_r_4_LC_2_19_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 a_r_4_LC_2_19_7 (
            .in0(N__3077),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(a_rZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3154),
            .ce(),
            .sr(_gnd_net_));
    defparam b_r_sbtinv_5_LC_3_16_0.C_ON=1'b0;
    defparam b_r_sbtinv_5_LC_3_16_0.SEQ_MODE=4'b0000;
    defparam b_r_sbtinv_5_LC_3_16_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 b_r_sbtinv_5_LC_3_16_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3240),
            .lcout(b_r_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam a_r_2_LC_3_17_0.C_ON=1'b0;
    defparam a_r_2_LC_3_17_0.SEQ_MODE=4'b1000;
    defparam a_r_2_LC_3_17_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 a_r_2_LC_3_17_0 (
            .in0(N__3029),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(a_rZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3147),
            .ce(),
            .sr(_gnd_net_));
    defparam b_r_RNI409B_7_LC_3_17_3.C_ON=1'b0;
    defparam b_r_RNI409B_7_LC_3_17_3.SEQ_MODE=4'b0000;
    defparam b_r_RNI409B_7_LC_3_17_3.LUT_INIT=16'b1111111111111010;
    LogicCell40 b_r_RNI409B_7_LC_3_17_3 (
            .in0(N__3242),
            .in1(N__2996),
            .in2(N__3167),
            .in3(N__3188),
            .lcout(b_r_RNI409BZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam b_r_RNI15S9_6_LC_3_17_4.C_ON=1'b0;
    defparam b_r_RNI15S9_6_LC_3_17_4.SEQ_MODE=4'b0000;
    defparam b_r_RNI15S9_6_LC_3_17_4.LUT_INIT=16'b1100110000110011;
    LogicCell40 b_r_RNI15S9_6_LC_3_17_4 (
            .in0(N__2969),
            .in1(N__3241),
            .in2(_gnd_net_),
            .in3(N__3163),
            .lcout(b_r_RNI15S9Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sum_r_7_LC_3_17_5.C_ON=1'b0;
    defparam sum_r_7_LC_3_17_5.SEQ_MODE=4'b1000;
    defparam sum_r_7_LC_3_17_5.LUT_INIT=16'b1100110010000000;
    LogicCell40 sum_r_7_LC_3_17_5 (
            .in0(N__2944),
            .in1(N__2930),
            .in2(N__2924),
            .in3(N__2897),
            .lcout(sum_o_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3147),
            .ce(),
            .sr(_gnd_net_));
    defparam b_r_5_LC_3_17_6.C_ON=1'b0;
    defparam b_r_5_LC_3_17_6.SEQ_MODE=4'b1000;
    defparam b_r_5_LC_3_17_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 b_r_5_LC_3_17_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3257),
            .lcout(b_rZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3147),
            .ce(),
            .sr(_gnd_net_));
    defparam a_r_3_LC_3_17_7.C_ON=1'b0;
    defparam a_r_3_LC_3_17_7.SEQ_MODE=4'b1000;
    defparam a_r_3_LC_3_17_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 a_r_3_LC_3_17_7 (
            .in0(N__3227),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(a_rZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3147),
            .ce(),
            .sr(_gnd_net_));
    defparam b_r_7_LC_3_18_3.C_ON=1'b0;
    defparam b_r_7_LC_3_18_3.SEQ_MODE=4'b1000;
    defparam b_r_7_LC_3_18_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 b_r_7_LC_3_18_3 (
            .in0(N__3200),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(b_rZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3155),
            .ce(),
            .sr(_gnd_net_));
    defparam b_r_6_LC_3_18_5.C_ON=1'b0;
    defparam b_r_6_LC_3_18_5.SEQ_MODE=4'b1000;
    defparam b_r_6_LC_3_18_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 b_r_6_LC_3_18_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3182),
            .lcout(b_rZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3155),
            .ce(),
            .sr(_gnd_net_));
endmodule // bcd_adder
