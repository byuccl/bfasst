
 module ucsb_152_tap_fir(clk, In_X, Out_Y); 

 input clk;
 input [11:0] In_X; 
 output [28 :0] Out_Y; 

 reg [11:0] x0 ;

 wire [14:0] x1 ;
 wire [17:0] x5 ;
 wire [22:0] x16 ;
 wire [22:0] x102 ;
 wire [22:0] y53 ;
 wire [22:0] y97 ;
 wire [22:0] x16_1_1 ;
 wire [22:0] y11 ;
 wire [22:0] x16_2_1 ;
 wire [22:0] y139 ;
 wire [21:0] x47 ;
 wire [21:0] x47_0_1 ;
 wire [22:0] y9 ;
 wire [21:0] x47_1_1 ;
 wire [22:0] y141 ;
 wire [22:0] x48 ;
 wire [22:0] x48_0_1 ;
 wire [22:0] y18 ;
 wire [22:0] x48_1_1 ;
 wire [22:0] y132 ;
 wire [22:0] x49 ;
 wire [22:0] x103 ;
 wire [23:0] y57 ;
 wire [23:0] y93 ;
 wire [23:0] x50 ;
 wire [23:0] x50_0_1 ;
 wire [23:0] y59 ;
 wire [23:0] x50_1_1 ;
 wire [23:0] y91 ;
 wire [21:0] x62 ;
 wire [21:0] x62_0_1 ;
 wire [22:0] y50 ;
 wire [21:0] x62_1_1 ;
 wire [22:0] y100 ;
 wire [24:0] x73 ;
 wire [24:0] x73_0_1 ;
 wire [24:0] y54 ;
 wire [24:0] x73_1_1 ;
 wire [24:0] y96 ;
 wire [17:0] x6 ;
 wire [21:0] x51 ;
 wire [21:0] x51_0_1 ;
 wire [21:0] y7 ;
 wire [21:0] x51_1_1 ;
 wire [21:0] y143 ;
 wire [22:0] x52 ;
 wire [22:0] x52_0_1 ;
 wire [23:0] y39 ;
 wire [22:0] x52_1_1 ;
 wire [23:0] y111 ;
 wire [23:0] x53 ;
 wire [23:0] x53_0_1 ;
 wire [23:0] y41 ;
 wire [23:0] x53_1_1 ;
 wire [23:0] y109 ;
 wire [23:0] x63 ;
 wire [23:0] x92 ;
 wire [23:0] y19 ;
 wire [23:0] y131 ;
 wire [21:0] x64 ;
 wire [21:0] x64_0_1 ;
 wire [21:0] y33 ;
 wire [21:0] x64_1_1 ;
 wire [21:0] y117 ;
 wire [23:0] x75 ;
 wire [23:0] x98 ;
 wire [23:0] y38 ;
 wire [19:0] x77 ;
 wire [19:0] x77_0_1 ;
 wire [23:0] y66 ;
 wire [19:0] x84 ;
 wire [19:0] x84_0_1 ;
 wire [23:0] y84 ;
 wire [23:0] x86 ;
 wire [23:0] x109 ;
 wire [23:0] y112 ;
 wire [18:0] x8 ;
 wire [22:0] x17 ;
 wire [22:0] x99 ;
 wire [22:0] y43 ;
 wire [22:0] y107 ;
 wire [22:0] x17_1_1 ;
 wire [22:0] y17 ;
 wire [22:0] x17_2_1 ;
 wire [22:0] y133 ;
 wire [22:0] x55 ;
 wire [22:0] x89 ;
 wire [22:0] y5 ;
 wire [22:0] y145 ;
 wire [24:0] x74 ;
 wire [24:0] x74_0_1 ;
 wire [24:0] y8 ;
 wire [21:0] x76 ;
 wire [21:0] x76_0_1 ;
 wire [21:0] y46 ;
 wire [21:0] x85 ;
 wire [21:0] x85_0_1 ;
 wire [21:0] y104 ;
 wire [24:0] x87 ;
 wire [24:0] x87_0_1 ;
 wire [24:0] y142 ;
 wire [18:0] x8_6_1 ;
 wire [18:0] x8_6_2 ;
 wire [22:0] y45 ;
 wire [18:0] x8_7_1 ;
 wire [18:0] x8_7_2 ;
 wire [22:0] y105 ;
 wire [22:0] x9 ;
 wire [23:0] x65 ;
 wire [23:0] x65_0_1 ;
 wire [23:0] y37 ;
 wire [23:0] x65_1_1 ;
 wire [23:0] y113 ;
 wire [23:0] x66 ;
 wire [23:0] x66_0_1 ;
 wire [23:0] y63 ;
 wire [23:0] x66_1_1 ;
 wire [23:0] y87 ;
 wire [22:0] x9_2_1 ;
 wire [22:0] x9_2_2 ;
 wire [22:0] y49 ;
 wire [22:0] x9_3_1 ;
 wire [22:0] x9_3_2 ;
 wire [22:0] y101 ;
 wire [18:0] x12 ;
 wire [24:0] x68 ;
 wire [24:0] x68_0_1 ;
 wire [24:0] y1 ;
 wire [24:0] x68_1_1 ;
 wire [24:0] y149 ;
 wire [18:0] x12_1_1 ;
 wire [18:0] x12_1_2 ;
 wire [21:0] y24 ;
 wire [18:0] x12_2_1 ;
 wire [18:0] x12_2_2 ;
 wire [21:0] y126 ;
 wire [20:0] x15 ;
 wire [20:0] x104 ;
 wire [20:0] x104_0_1 ;
 wire [22:0] y61 ;
 wire [20:0] x104_1_1 ;
 wire [22:0] y89 ;
 wire [20:0] x15_1_1 ;
 wire [20:0] x15_1_2 ;
 wire [21:0] y26 ;
 wire [20:0] x15_2_1 ;
 wire [20:0] x15_2_2 ;
 wire [21:0] y124 ;
 wire [23:0] x18 ;
 wire [23:0] x105 ;
 wire [24:0] y62 ;
 wire [24:0] y88 ;
 wire [23:0] x18_1_1 ;
 wire [23:0] y52 ;
 wire [23:0] x18_2_1 ;
 wire [23:0] y98 ;
 wire [17:0] x21 ;
 wire [23:0] x72 ;
 wire [23:0] x72_0_1 ;
 wire [24:0] y3 ;
 wire [23:0] x72_1_1 ;
 wire [24:0] y147 ;
 wire [19:0] x22 ;
 wire [19:0] x22_0_1 ;
 wire [19:0] x22_0_2 ;
 wire [22:0] y40 ;
 wire [19:0] x22_1_1 ;
 wire [19:0] x22_1_2 ;
 wire [22:0] y110 ;
 wire [19:0] x23 ;
 wire [19:0] x91 ;
 wire [19:0] x91_0_1 ;
 wire [22:0] y15 ;
 wire [19:0] x91_1_1 ;
 wire [22:0] y135 ;
 wire [20:0] x24 ;
 wire [20:0] x24_0_1 ;
 wire [20:0] x24_0_2 ;
 wire [21:0] y22 ;
 wire [20:0] x24_1_1 ;
 wire [20:0] x24_1_2 ;
 wire [21:0] y128 ;
 wire [21:0] x25 ;
 wire [22:0] x70 ;
 wire [22:0] x70_0_1 ;
 wire [22:0] y48 ;
 wire [22:0] x70_1_1 ;
 wire [22:0] y102 ;
 wire [19:0] x34 ;
 wire [24:0] x57 ;
 wire [24:0] x57_0_1 ;
 wire [26:0] y68 ;
 wire [24:0] x57_1_1 ;
 wire [26:0] y82 ;
 wire [21:0] x35 ;
 wire [21:0] x101 ;
 wire [21:0] x101_0_1 ;
 wire [22:0] y51 ;
 wire [21:0] x101_1_1 ;
 wire [22:0] y99 ;
 wire [21:0] x36 ;
 wire [21:0] x36_0_1 ;
 wire [21:0] x36_0_2 ;
 wire [22:0] y13 ;
 wire [21:0] x36_1_1 ;
 wire [21:0] x36_1_2 ;
 wire [22:0] y137 ;
 wire [21:0] x37 ;
 wire [21:0] x37_0_1 ;
 wire [21:0] x37_0_2 ;
 wire [21:0] y27 ;
 wire [21:0] x37_1_1 ;
 wire [21:0] x37_1_2 ;
 wire [21:0] y123 ;
 wire [20:0] x38 ;
 wire [20:0] x38_0_1 ;
 wire [20:0] x38_0_2 ;
 wire [21:0] y29 ;
 wire [20:0] x38_1_1 ;
 wire [20:0] x38_1_2 ;
 wire [21:0] y121 ;
 wire [22:0] x39 ;
 wire [22:0] x39_0_1 ;
 wire [22:0] x39_0_2 ;
 wire [27:0] y74 ;
 wire [22:0] x39_1_1 ;
 wire [22:0] x39_1_2 ;
 wire [27:0] y76 ;
 wire [21:0] x40 ;
 wire [21:0] x40_0_1 ;
 wire [21:0] x40_0_2 ;
 wire [21:0] y14 ;
 wire [21:0] x40_1_1 ;
 wire [21:0] x40_1_2 ;
 wire [21:0] y136 ;
 wire [21:0] x41 ;
 wire [21:0] x41_0_1 ;
 wire [21:0] x41_0_2 ;
 wire [21:0] y34 ;
 wire [21:0] x41_1_1 ;
 wire [21:0] x41_1_2 ;
 wire [21:0] y116 ;
 wire [21:0] x42 ;
 wire [21:0] x42_0_1 ;
 wire [21:0] x42_0_2 ;
 wire [22:0] y55 ;
 wire [21:0] x42_1_1 ;
 wire [21:0] x42_1_2 ;
 wire [22:0] y95 ;
 wire [21:0] x43 ;
 wire [21:0] x43_0_1 ;
 wire [21:0] x43_0_2 ;
 wire [21:0] y20 ;
 wire [21:0] x43_1_1 ;
 wire [21:0] x43_1_2 ;
 wire [21:0] y130 ;
 wire [22:0] x44 ;
 wire [22:0] x100 ;
 wire [22:0] x100_0_1 ;
 wire [22:0] y47 ;
 wire [22:0] x100_1_1 ;
 wire [22:0] y103 ;
 wire [24:0] x45 ;
 wire [24:0] x45_0_1 ;
 wire [24:0] x45_0_2 ;
 wire [24:0] y64 ;
 wire [24:0] x45_1_1 ;
 wire [24:0] x45_1_2 ;
 wire [24:0] y86 ;
 wire [20:0] x46 ;
 wire [20:0] x107 ;
 wire [20:0] x107_0_1 ;
 wire [22:0] y73 ;
 wire [20:0] x107_1_1 ;
 wire [22:0] y77 ;
 wire [22:0] x54 ;
 wire [22:0] x54_0_1 ;
 wire [22:0] x54_0_2 ;
 wire [22:0] y12 ;
 wire [22:0] x54_1_1 ;
 wire [22:0] x54_1_2 ;
 wire [22:0] y138 ;
 wire [24:0] x56 ;
 wire [24:0] x56_0_1 ;
 wire [24:0] y4 ;
 wire [24:0] x56_1_1 ;
 wire [24:0] y146 ;
 wire [14:0] x2 ;
 wire [17:0] x10 ;
 wire [17:0] x10_1_1 ;
 wire [17:0] x10_1_2 ;
 wire [21:0] y35 ;
 wire [17:0] x10_2_1 ;
 wire [17:0] x10_2_2 ;
 wire [21:0] y115 ;
 wire [17:0] x11 ;
 wire [22:0] x67 ;
 wire [22:0] x67_0_1 ;
 wire [22:0] y65 ;
 wire [22:0] x67_1_1 ;
 wire [22:0] y85 ;
 wire [23:0] x71 ;
 wire [23:0] x71_0_1 ;
 wire [26:0] y72 ;
 wire [23:0] x71_1_1 ;
 wire [26:0] y78 ;
 wire [21:0] x78 ;
 wire [21:0] x78_0_1 ;
 wire [22:0] y67 ;
 wire [22:0] x79 ;
 wire [22:0] x106 ;
 wire [22:0] y69 ;
 wire [21:0] x80 ;
 wire [21:0] x80_0_1 ;
 wire [22:0] y71 ;
 wire [21:0] x81 ;
 wire [21:0] x81_0_1 ;
 wire [22:0] y79 ;
 wire [22:0] x82 ;
 wire [22:0] x108 ;
 wire [22:0] y81 ;
 wire [21:0] x83 ;
 wire [21:0] x83_0_1 ;
 wire [22:0] y83 ;
 wire [17:0] x11_8_1 ;
 wire [17:0] x11_8_2 ;
 wire [21:0] y42 ;
 wire [17:0] x11_9_1 ;
 wire [17:0] x11_9_2 ;
 wire [21:0] y108 ;
 wire [19:0] x13 ;
 wire [19:0] x13_1_1 ;
 wire [19:0] x13_1_2 ;
 wire [20:0] y0 ;
 wire [19:0] x13_2_1 ;
 wire [19:0] x13_2_2 ;
 wire [20:0] y150 ;
 wire [18:0] x26 ;
 wire [18:0] x26_0_1 ;
 wire [18:0] x26_0_2 ;
 wire [21:0] y23 ;
 wire [18:0] x26_1_1 ;
 wire [18:0] x26_1_2 ;
 wire [21:0] y127 ;
 wire [19:0] x27 ;
 wire [19:0] x94 ;
 wire [19:0] x94_0_1 ;
 wire [21:0] y25 ;
 wire [19:0] x94_1_1 ;
 wire [21:0] y125 ;
 wire [20:0] x58 ;
 wire [20:0] x93 ;
 wire [20:0] x93_0_1 ;
 wire [21:0] y21 ;
 wire [20:0] x93_1_1 ;
 wire [21:0] y129 ;
 wire [23:0] x59 ;
 wire [23:0] x59_0_1 ;
 wire [23:0] x59_0_2 ;
 wire [23:0] y60 ;
 wire [23:0] x59_1_1 ;
 wire [23:0] x59_1_2 ;
 wire [23:0] y90 ;
 wire [24:0] x60 ;
 wire [24:0] x88 ;
 wire [24:0] x88_0_1 ;
 wire [24:0] y2 ;
 wire [24:0] x88_1_1 ;
 wire [24:0] y148 ;
 wire [21:0] x61 ;
 wire [21:0] x61_0_1 ;
 wire [21:0] x61_0_2 ;
 wire [21:0] y31 ;
 wire [21:0] x61_1_1 ;
 wire [21:0] x61_1_2 ;
 wire [21:0] y119 ;
 wire [23:0] x69 ;
 wire [23:0] x69_0_1 ;
 wire [23:0] x69_0_2 ;
 wire [23:0] y6 ;
 wire [23:0] x69_1_1 ;
 wire [23:0] x69_1_2 ;
 wire [23:0] y144 ;
 wire [14:0] x97 ;
 wire [14:0] x97_0_1 ;
 wire [14:0] x97_0_2 ;
 wire [20:0] y36 ;
 wire [14:0] x97_1_1 ;
 wire [14:0] x97_1_2 ;
 wire [20:0] y114 ;
 wire [15:0] x3 ;
 wire [19:0] x28 ;
 wire [19:0] x28_0_1 ;
 wire [19:0] x28_0_2 ;
 wire [20:0] y16 ;
 wire [19:0] x28_1_1 ;
 wire [19:0] x28_1_2 ;
 wire [20:0] y134 ;
 wire [20:0] x29 ;
 wire [20:0] x96 ;
 wire [20:0] x96_0_1 ;
 wire [20:0] y32 ;
 wire [20:0] x96_1_1 ;
 wire [20:0] y118 ;
 wire [19:0] x30 ;
 wire [19:0] x30_0_1 ;
 wire [19:0] x30_0_2 ;
 wire [22:0] y58 ;
 wire [19:0] x30_1_1 ;
 wire [19:0] x30_1_2 ;
 wire [22:0] y92 ;
 wire [15:0] x4 ;
 wire [20:0] x31 ;
 wire [20:0] x95 ;
 wire [20:0] x95_0_1 ;
 wire [21:0] y28 ;
 wire [20:0] x95_1_1 ;
 wire [21:0] y122 ;
 wire [19:0] x32 ;
 wire [19:0] x32_0_1 ;
 wire [19:0] x32_0_2 ;
 wire [20:0] y30 ;
 wire [19:0] x32_1_1 ;
 wire [19:0] x32_1_2 ;
 wire [20:0] y120 ;
 wire [16:0] x7 ;
 wire [22:0] x14 ;
 wire [22:0] x14_0_1 ;
 wire [22:0] x14_0_2 ;
 wire [22:0] y44 ;
 wire [22:0] x14_1_1 ;
 wire [22:0] x14_1_2 ;
 wire [23:0] y56 ;
 wire [22:0] x14_2_1 ;
 wire [22:0] x14_2_2 ;
 wire [23:0] y94 ;
 wire [22:0] x14_3_1 ;
 wire [22:0] x14_3_2 ;
 wire [22:0] y106 ;
 wire [24:0] x33 ;
 wire [24:0] x33_0_1 ;
 wire [24:0] x33_0_2 ;
 wire [24:0] y70 ;
 wire [24:0] x33_1_1 ;
 wire [24:0] x33_1_2 ;
 wire [24:0] y80 ;
 wire [19:0] x19 ;
 wire [19:0] x90 ;
 wire [19:0] x90_0_1 ;
 wire [19:0] x90_0_2 ;
 wire [21:0] y10 ;
 wire [19:0] x90_1_1 ;
 wire [19:0] x90_1_2 ;
 wire [21:0] y140 ;
 wire [22:0] x20 ;
 wire [11:0] x74_36_1 ;
 wire [11:0] x74_36_2 ;
 wire [11:0] x75_37_1 ;
 wire [11:0] x75_37_2 ;
 wire [11:0] x76_38_1 ;
 wire [11:0] x76_38_2 ;
 wire [11:0] x77_39_1 ;
 wire [11:0] x77_39_2 ;
 wire [11:0] x78_40_1 ;
 wire [11:0] x78_40_2 ;
 wire [11:0] x79_41_1 ;
 wire [11:0] x79_41_2 ;
 wire [11:0] x80_42_1 ;
 wire [11:0] x80_42_2 ;
 wire [11:0] x81_43_1 ;
 wire [11:0] x81_43_2 ;
 wire [11:0] x82_44_1 ;
 wire [11:0] x82_44_2 ;
 wire [11:0] x83_45_1 ;
 wire [11:0] x83_45_2 ;
 wire [11:0] x84_46_1 ;
 wire [11:0] x84_46_2 ;
 wire [11:0] x85_47_1 ;
 wire [11:0] x85_47_2 ;
 wire [11:0] x86_48_1 ;
 wire [11:0] x86_48_2 ;
 wire [11:0] x87_49_1 ;
 wire [11:0] x87_49_2 ;
 wire [11:0] x0_50_1 ;
 wire [11:0] x0_50_2 ;
 wire [11:0] x0_50_3 ;
 wire [11:0] x0_50_4 ;
 wire [26:0] y75 ;
 wire [20:0] x110 ;
 wire [25:0] x111 ;
 wire [25:0] x111_1 ;
 wire [26:0] x112 ;
 wire [26:0] x112_1 ;
 wire [27:0] x113 ;
 wire [27:0] x113_1 ;
 wire [28:0] x114 ;
 wire [28:0] x114_1 ;
 wire [28:0] x115 ;
 wire [28:0] x115_1 ;
 wire [28:0] x116 ;
 wire [28:0] x116_1 ;
 wire [28:0] x117 ;
 wire [28:0] x117_1 ;
 wire [28:0] x118 ;
 wire [28:0] x118_1 ;
 wire [28:0] x119 ;
 wire [28:0] x119_1 ;
 wire [28:0] x120 ;
 wire [28:0] x120_1 ;
 wire [28:0] x121 ;
 wire [28:0] x121_1 ;
 wire [28:0] x122 ;
 wire [28:0] x122_1 ;
 wire [28:0] x123 ;
 wire [28:0] x123_1 ;
 wire [28:0] x124 ;
 wire [28:0] x124_1 ;
 wire [28:0] x125 ;
 wire [28:0] x125_1 ;
 wire [28:0] x126 ;
 wire [28:0] x126_1 ;
 wire [28:0] x127 ;
 wire [28:0] x127_1 ;
 wire [28:0] x128 ;
 wire [28:0] x128_1 ;
 wire [28:0] x129 ;
 wire [28:0] x129_1 ;
 wire [28:0] x130 ;
 wire [28:0] x130_1 ;
 wire [28:0] x131 ;
 wire [28:0] x131_1 ;
 wire [28:0] x132 ;
 wire [28:0] x132_1 ;
 wire [28:0] x133 ;
 wire [28:0] x133_1 ;
 wire [28:0] x134 ;
 wire [28:0] x134_1 ;
 wire [28:0] x135 ;
 wire [28:0] x135_1 ;
 wire [28:0] x136 ;
 wire [28:0] x136_1 ;
 wire [28:0] x137 ;
 wire [28:0] x137_1 ;
 wire [28:0] x138 ;
 wire [28:0] x138_1 ;
 wire [28:0] x139 ;
 wire [28:0] x139_1 ;
 wire [28:0] x140 ;
 wire [28:0] x140_1 ;
 wire [28:0] x141 ;
 wire [28:0] x141_1 ;
 wire [28:0] x142 ;
 wire [28:0] x142_1 ;
 wire [28:0] x143 ;
 wire [28:0] x143_1 ;
 wire [28:0] x144 ;
 wire [28:0] x144_1 ;
 wire [28:0] x145 ;
 wire [28:0] x145_1 ;
 wire [28:0] x146 ;
 wire [28:0] x146_1 ;
 wire [28:0] x147 ;
 wire [28:0] x147_1 ;
 wire [28:0] x148 ;
 wire [28:0] x148_1 ;
 wire [28:0] x149 ;
 wire [28:0] x149_1 ;
 wire [28:0] x150 ;
 wire [28:0] x150_1 ;
 wire [28:0] x151 ;
 wire [28:0] x151_1 ;
 wire [28:0] x152 ;
 wire [28:0] x152_1 ;
 wire [28:0] x153 ;
 wire [28:0] x153_1 ;
 wire [28:0] x154 ;
 wire [28:0] x154_1 ;
 wire [28:0] x155 ;
 wire [28:0] x155_1 ;
 wire [28:0] x156 ;
 wire [28:0] x156_1 ;
 wire [28:0] x157 ;
 wire [28:0] x157_1 ;
 wire [28:0] x158 ;
 wire [28:0] x158_1 ;
 wire [28:0] x159 ;
 wire [28:0] x159_1 ;
 wire [28:0] x160 ;
 wire [28:0] x160_1 ;
 wire [28:0] x161 ;
 wire [28:0] x161_1 ;
 wire [28:0] x162 ;
 wire [28:0] x162_1 ;
 wire [28:0] x163 ;
 wire [28:0] x163_1 ;
 wire [28:0] x164 ;
 wire [28:0] x164_1 ;
 wire [28:0] x165 ;
 wire [28:0] x165_1 ;
 wire [28:0] x166 ;
 wire [28:0] x166_1 ;
 wire [28:0] x167 ;
 wire [28:0] x167_1 ;
 wire [28:0] x168 ;
 wire [28:0] x168_1 ;
 wire [28:0] x169 ;
 wire [28:0] x169_1 ;
 wire [28:0] x170 ;
 wire [28:0] x170_1 ;
 wire [28:0] x171 ;
 wire [28:0] x171_1 ;
 wire [28:0] x172 ;
 wire [28:0] x172_1 ;
 wire [28:0] x173 ;
 wire [28:0] x173_1 ;
 wire [28:0] x174 ;
 wire [28:0] x174_1 ;
 wire [28:0] x175 ;
 wire [28:0] x175_1 ;
 wire [28:0] x176 ;
 wire [28:0] x176_1 ;
 wire [28:0] x177 ;
 wire [28:0] x177_1 ;
 wire [28:0] x178 ;
 wire [28:0] x178_1 ;
 wire [28:0] x179 ;
 wire [28:0] x179_1 ;
 wire [28:0] x180 ;
 wire [28:0] x180_1 ;
 wire [28:0] x181 ;
 wire [28:0] x181_1 ;
 wire [28:0] x182 ;
 wire [28:0] x182_1 ;
 wire [28:0] x183 ;
 wire [28:0] x183_1 ;
 wire [28:0] x184 ;
 wire [28:0] x184_1 ;
 wire [28:0] x185 ;
 wire [28:0] x185_1 ;
 wire [28:0] x186 ;
 wire [28:0] x186_1 ;
 wire [28:0] x187 ;
 wire [28:0] x187_1 ;
 wire [28:0] x188 ;
 wire [28:0] x188_1 ;
 wire [28:0] x189 ;
 wire [28:0] x189_1 ;
 wire [28:0] x190 ;
 wire [28:0] x190_1 ;
 wire [28:0] x191 ;
 wire [28:0] x191_1 ;
 wire [28:0] x192 ;
 wire [28:0] x192_1 ;
 wire [28:0] x193 ;
 wire [28:0] x193_1 ;
 wire [28:0] x194 ;
 wire [28:0] x194_1 ;
 wire [28:0] x195 ;
 wire [28:0] x195_1 ;
 wire [28:0] x196 ;
 wire [28:0] x196_1 ;
 wire [28:0] x197 ;
 wire [28:0] x197_1 ;
 wire [28:0] x198 ;
 wire [28:0] x198_1 ;
 wire [28:0] x199 ;
 wire [28:0] x199_1 ;
 wire [28:0] x200 ;
 wire [28:0] x200_1 ;
 wire [28:0] x201 ;
 wire [28:0] x201_1 ;
 wire [28:0] x202 ;
 wire [28:0] x202_1 ;
 wire [28:0] x203 ;
 wire [28:0] x203_1 ;
 wire [28:0] x204 ;
 wire [28:0] x204_1 ;
 wire [28:0] x205 ;
 wire [28:0] x205_1 ;
 wire [28:0] x206 ;
 wire [28:0] x206_1 ;
 wire [28:0] x207 ;
 wire [28:0] x207_1 ;
 wire [28:0] x208 ;
 wire [28:0] x208_1 ;
 wire [28:0] x209 ;
 wire [28:0] x209_1 ;
 wire [28:0] x210 ;
 wire [28:0] x210_1 ;
 wire [28:0] x211 ;
 wire [28:0] x211_1 ;
 wire [28:0] x212 ;
 wire [28:0] x212_1 ;
 wire [28:0] x213 ;
 wire [28:0] x213_1 ;
 wire [28:0] x214 ;
 wire [28:0] x214_1 ;
 wire [28:0] x215 ;
 wire [28:0] x215_1 ;
 wire [28:0] x216 ;
 wire [28:0] x216_1 ;
 wire [28:0] x217 ;
 wire [28:0] x217_1 ;
 wire [28:0] x218 ;
 wire [28:0] x218_1 ;
 wire [28:0] x219 ;
 wire [28:0] x219_1 ;
 wire [28:0] x220 ;
 wire [28:0] x220_1 ;
 wire [28:0] x221 ;
 wire [28:0] x221_1 ;
 wire [28:0] x222 ;
 wire [28:0] x222_1 ;
 wire [28:0] x223 ;
 wire [28:0] x223_1 ;
 wire [28:0] x224 ;
 wire [28:0] x224_1 ;
 wire [28:0] x225 ;
 wire [28:0] x225_1 ;
 wire [28:0] x226 ;
 wire [28:0] x226_1 ;
 wire [28:0] x227 ;
 wire [28:0] x227_1 ;
 wire [28:0] x228 ;
 wire [28:0] x228_1 ;
 wire [28:0] x229 ;
 wire [28:0] x229_1 ;
 wire [28:0] x230 ;
 wire [28:0] x230_1 ;
 wire [28:0] x231 ;
 wire [28:0] x231_1 ;
 wire [28:0] x232 ;
 wire [28:0] x232_1 ;
 wire [28:0] x233 ;
 wire [28:0] x233_1 ;
 wire [28:0] x234 ;
 wire [28:0] x234_1 ;
 wire [28:0] x235 ;
 wire [28:0] x235_1 ;
 wire [28:0] x236 ;
 wire [28:0] x236_1 ;
 wire [28:0] x237 ;
 wire [28:0] x237_1 ;
 wire [28:0] x238 ;
 wire [28:0] x238_1 ;
 wire [28:0] x239 ;
 wire [28:0] x239_1 ;
 wire [28:0] x240 ;
 wire [28:0] x240_1 ;
 wire [28:0] x241 ;
 wire [28:0] x241_1 ;
 wire [28:0] x242 ;
 wire [28:0] x242_1 ;
 wire [28:0] x243 ;
 wire [28:0] x243_1 ;
 wire [28:0] x244 ;
 wire [28:0] x244_1 ;
 wire [28:0] x245 ;
 wire [28:0] x245_1 ;
 wire [28:0] x246 ;
 wire [28:0] x246_1 ;
 wire [28:0] x247 ;
 wire [28:0] x247_1 ;
 wire [28:0] x248 ;
 wire [28:0] x248_1 ;
 wire [28:0] x249 ;
 wire [28:0] x249_1 ;
 wire [28:0] x250 ;
 wire [28:0] x250_1 ;
 wire [28:0] x251 ;
 wire [28:0] x251_1 ;
 wire [28:0] x252 ;
 wire [28:0] x252_1 ;
 wire [28:0] x253 ;
 wire [28:0] x253_1 ;
 wire [28:0] x254 ;
 wire [28:0] x254_1 ;
 wire [28:0] x255 ;
 wire [28:0] x255_1 ;
 wire [28:0] x256 ;
 wire [28:0] x256_1 ;
 wire [28:0] x257 ;
 wire [28:0] x257_1 ;
 wire [28:0] x258 ;
 wire [28:0] x258_1 ;
 wire [28:0] x259 ;
 wire [28:0] x259_1 ;
 wire [28:0] Out_Y_wire ;
 reg [28:0] Out_Y;


 always @(posedge clk) 
 begin
 x0 <= In_X; 
 end 


 always @(posedge clk) 
 begin
 Out_Y = Out_Y_wire;
 end


 Subtractor14Bit Sub0(clk, {x0[11],x0[11], x0[11: 0] },  { x0[11: 0], 2'b0 },x1); 


 Subtractor17Bit Sub1(clk, {x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] },  { x1[14: 0], 2'b0 },x5); 


 Subtractor22Bit Sub2(clk, {x5[17],x5[17],x5[17],x5[17], x5[17: 0] },  { x1[14: 0], 7'b0 },x16); 

 Negator23Bit Neg0(clk, x16, x102 );
 Register23Bit Reg0 (clk,x102, y53 );
 Register23Bit Reg1 (clk,x102, y97 );
 Register23Bit Reg2 (clk,x16, x16_1_1 );
 Register23Bit Reg3 (clk,x16_1_1, y11 );
 Register23Bit Reg4 (clk,x16, x16_2_1 );
 Register23Bit Reg5 (clk,x16_2_1, y139 );

 Adder21Bit Adder0(clk,  { x1[14: 0], 6'b0 }, {x5[17],x5[17],x5[17], x5[17: 0]  }, x47); 

 Register22Bit Reg6 (clk,x47, x47_0_1 );
 Register23Bit Reg7 (clk, {x47_0_1, 1'b0}, y9 );
 Register22Bit Reg8 (clk,x47, x47_1_1 );
 Register23Bit Reg9 (clk, {x47_1_1, 1'b0}, y141 );

 Subtractor22Bit Sub3(clk, { x5[17: 0], 4'b0 }, {x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0] }, x48); 

 Register23Bit Reg10 (clk,x48, x48_0_1 );
 Register23Bit Reg11 (clk,x48_0_1, y18 );
 Register23Bit Reg12 (clk,x48, x48_1_1 );
 Register23Bit Reg13 (clk,x48_1_1, y132 );

 Adder22Bit Adder1(clk,  {x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0] },  { x5[17: 0], 4'b0 },x49); 

 Negator23Bit Neg1(clk, x49, x103 );
 Register24Bit Reg14 (clk, {x103, 1'b0}, y57 );
 Register24Bit Reg15 (clk, {x103, 1'b0}, y93 );

 Adder23Bit Adder2(clk,  {x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0] },  { x5[17: 0], 5'b0 },x50); 

 Register24Bit Reg16 (clk,x50, x50_0_1 );
 Register24Bit Reg17 (clk,x50_0_1, y59 );
 Register24Bit Reg18 (clk,x50, x50_1_1 );
 Register24Bit Reg19 (clk,x50_1_1, y91 );

 Adder17Bit Adder3(clk,  {x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] },  { x1[14: 0], 2'b0 },x6); 


 Subtractor21Bit Sub4(clk, {x6[17],x6[17],x6[17], x6[17: 0] },  { x1[14: 0], 6'b0 },x51); 

 Register22Bit Reg20 (clk,x51, x51_0_1 );
 Register22Bit Reg21 (clk,x51_0_1, y7 );
 Register22Bit Reg22 (clk,x51, x51_1_1 );
 Register22Bit Reg23 (clk,x51_1_1, y143 );

 Subtractor22Bit Sub5(clk, {x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0] },  { x6[17: 0], 4'b0 },x52); 

 Register23Bit Reg24 (clk,x52, x52_0_1 );
 Register24Bit Reg25 (clk, {x52_0_1, 1'b0}, y39 );
 Register23Bit Reg26 (clk,x52, x52_1_1 );
 Register24Bit Reg27 (clk, {x52_1_1, 1'b0}, y111 );

 Adder23Bit Adder4(clk,  {x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0] },  { x6[17: 0], 5'b0 },x53); 

 Register24Bit Reg28 (clk,x53, x53_0_1 );
 Register24Bit Reg29 (clk,x53_0_1, y41 );
 Register24Bit Reg30 (clk,x53, x53_1_1 );
 Register24Bit Reg31 (clk,x53_1_1, y109 );

 Subtractor24Bit Sub6(clk, { x5[17: 0], 6'b0 }, {x6[17],x6[17],x6[17],x6[17],x6[17],x6[17], x6[17: 0] }, x73); 

 Register25Bit Reg32 (clk,x73, x73_0_1 );
 Register25Bit Reg33 (clk,x73_0_1, y54 );
 Register25Bit Reg34 (clk,x73, x73_1_1 );
 Register25Bit Reg35 (clk,x73_1_1, y96 );

 Adder18Bit Adder5(clk,  {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] },  { x1[14: 0], 3'b0 },x8); 


 Subtractor22Bit Sub7(clk, { x1[14: 0], 7'b0 }, {x8[18],x8[18],x8[18], x8[18: 0] }, x17); 

 Negator23Bit Neg2(clk, x17, x99 );
 Register23Bit Reg36 (clk,x99, y43 );
 Register23Bit Reg37 (clk,x99, y107 );
 Register23Bit Reg38 (clk,x17, x17_1_1 );
 Register23Bit Reg39 (clk,x17_1_1, y17 );
 Register23Bit Reg40 (clk,x17, x17_2_1 );
 Register23Bit Reg41 (clk,x17_2_1, y133 );

 Adder22Bit Adder6(clk,  { x1[14: 0], 7'b0 }, {x8[18],x8[18],x8[18], x8[18: 0]  }, x55); 

 Negator23Bit Neg3(clk, x55, x89 );
 Register23Bit Reg42 (clk,x89, y5 );
 Register23Bit Reg43 (clk,x89, y145 );
 Register19Bit Reg44 (clk,x8, x8_6_1 );
 Register19Bit Reg45 (clk,x8_6_1, x8_6_2 );
 Register23Bit Reg46 (clk, {x8_6_2, 4'b0}, y45 );
 Register19Bit Reg47 (clk,x8, x8_7_1 );
 Register19Bit Reg48 (clk,x8_7_1, x8_7_2 );
 Register23Bit Reg49 (clk, {x8_7_2, 4'b0}, y105 );

 Adder22Bit Adder7(clk,  {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] },  { x1[14: 0], 7'b0 },x9); 

 Register23Bit Reg50 (clk,x9, x9_2_1 );
 Register23Bit Reg51 (clk,x9_2_1, x9_2_2 );
 Register23Bit Reg52 (clk,x9_2_2, y49 );
 Register23Bit Reg53 (clk,x9, x9_3_1 );
 Register23Bit Reg54 (clk,x9_3_1, x9_3_2 );
 Register23Bit Reg55 (clk,x9_3_2, y101 );

 Subtractor18Bit Sub8(clk, { x1[14: 0], 3'b0 }, {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] }, x12); 

 Register19Bit Reg56 (clk,x12, x12_1_1 );
 Register19Bit Reg57 (clk,x12_1_1, x12_1_2 );
 Register22Bit Reg58 (clk, {x12_1_2, 3'b0}, y24 );
 Register19Bit Reg59 (clk,x12, x12_2_1 );
 Register19Bit Reg60 (clk,x12_2_1, x12_2_2 );
 Register22Bit Reg61 (clk, {x12_2_2, 3'b0}, y126 );

 Subtractor17Bit Sub9(clk, {x1[14],x1[14], x1[14: 0] },  { x0[11: 0], 5'b0 },x21); 


 Subtractor19Bit Sub10(clk, { x1[14: 0], 4'b0 }, {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] }, x22); 

 Register20Bit Reg62 (clk,x22, x22_0_1 );
 Register20Bit Reg63 (clk,x22_0_1, x22_0_2 );
 Register23Bit Reg64 (clk, {x22_0_2, 3'b0}, y40 );
 Register20Bit Reg65 (clk,x22, x22_1_1 );
 Register20Bit Reg66 (clk,x22_1_1, x22_1_2 );
 Register23Bit Reg67 (clk, {x22_1_2, 3'b0}, y110 );

 Adder19Bit Adder8(clk,  {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] },  { x1[14: 0], 4'b0 },x23); 

 Negator20Bit Neg4(clk, x23, x91 );
 Register20Bit Reg68 (clk,x91, x91_0_1 );
 Register23Bit Reg69 (clk, {x91_0_1, 3'b0}, y15 );
 Register20Bit Reg70 (clk,x91, x91_1_1 );
 Register23Bit Reg71 (clk, {x91_1_1, 3'b0}, y135 );

 Subtractor20Bit Sub11(clk, {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] },  { x1[14: 0], 5'b0 },x24); 

 Register21Bit Reg72 (clk,x24, x24_0_1 );
 Register21Bit Reg73 (clk,x24_0_1, x24_0_2 );
 Register22Bit Reg74 (clk, {x24_0_2, 1'b0}, y22 );
 Register21Bit Reg75 (clk,x24, x24_1_1 );
 Register21Bit Reg76 (clk,x24_1_1, x24_1_2 );
 Register22Bit Reg77 (clk, {x24_1_2, 1'b0}, y128 );

 Subtractor21Bit Sub12(clk, {x1[14],x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0] },  { x0[11: 0], 9'b0 },x25); 


 Subtractor19Bit Sub13(clk, {x1[14],x1[14],x1[14],x1[14], x1[14: 0] },  { x1[14: 0], 4'b0 },x34); 


 Subtractor24Bit Sub14(clk, {x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0] },  { x34[19: 0], 4'b0 },x57); 

 Register25Bit Reg78 (clk,x57, x57_0_1 );
 Register27Bit Reg79 (clk, {x57_0_1, 2'b0}, y68 );
 Register25Bit Reg80 (clk,x57, x57_1_1 );
 Register27Bit Reg81 (clk, {x57_1_1, 2'b0}, y82 );

 Adder21Bit Adder9(clk,  {x1[14],x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0] },  { x1[14: 0], 6'b0 },x35); 

 Negator22Bit Neg5(clk, x35, x101 );
 Register22Bit Reg82 (clk,x101, x101_0_1 );
 Register23Bit Reg83 (clk, {x101_0_1, 1'b0}, y51 );
 Register22Bit Reg84 (clk,x101, x101_1_1 );
 Register23Bit Reg85 (clk, {x101_1_1, 1'b0}, y99 );

 Adder14Bit Adder10(clk,  {x0[11],x0[11], x0[11: 0] },  { x0[11: 0], 2'b0 },x2); 


 Adder17Bit Adder11(clk,  {x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] },  { x2[14: 0], 2'b0 },x10); 


 Adder23Bit Adder12(clk,  { x1[14: 0], 8'b0 }, {x10[17],x10[17],x10[17],x10[17],x10[17], x10[17: 0]  }, x18); 

 Negator24Bit Neg6(clk, x18, x105 );
 Register25Bit Reg86 (clk, {x105, 1'b0}, y62 );
 Register25Bit Reg87 (clk, {x105, 1'b0}, y88 );
 Register24Bit Reg88 (clk,x18, x18_1_1 );
 Register24Bit Reg89 (clk,x18_1_1, y52 );
 Register24Bit Reg90 (clk,x18, x18_2_1 );
 Register24Bit Reg91 (clk,x18_2_1, y98 );
 Register18Bit Reg92 (clk,x10, x10_1_1 );
 Register18Bit Reg93 (clk,x10_1_1, x10_1_2 );
 Register22Bit Reg94 (clk, {x10_1_2, 4'b0}, y35 );
 Register18Bit Reg95 (clk,x10, x10_2_1 );
 Register18Bit Reg96 (clk,x10_2_1, x10_2_2 );
 Register22Bit Reg97 (clk, {x10_2_2, 4'b0}, y115 );

 Subtractor17Bit Sub15(clk, { x0[11: 0], 5'b0 }, {x2[14],x2[14], x2[14: 0] }, x11); 


 Subtractor22Bit Sub16(clk, {x2[14],x2[14],x2[14],x2[14],x2[14],x2[14],x2[14], x2[14: 0] },  { x11[17: 0], 4'b0 },x67); 

 Register23Bit Reg98 (clk,x67, x67_0_1 );
 Register23Bit Reg99 (clk,x67_0_1, y65 );
 Register23Bit Reg100 (clk,x67, x67_1_1 );
 Register23Bit Reg101 (clk,x67_1_1, y85 );
 Register18Bit Reg102 (clk,x11, x11_8_1 );
 Register18Bit Reg103 (clk,x11_8_1, x11_8_2 );
 Register22Bit Reg104 (clk, {x11_8_2, 4'b0}, y42 );
 Register18Bit Reg105 (clk,x11, x11_9_1 );
 Register18Bit Reg106 (clk,x11_9_1, x11_9_2 );
 Register22Bit Reg107 (clk, {x11_9_2, 4'b0}, y108 );

 Subtractor19Bit Sub17(clk, {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] },  { x2[14: 0], 4'b0 },x13); 


 Subtractor24Bit Sub18(clk, { x13[19: 0], 4'b0 }, {x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0] }, x56); 

 Register25Bit Reg108 (clk,x56, x56_0_1 );
 Register25Bit Reg109 (clk,x56_0_1, y4 );
 Register25Bit Reg110 (clk,x56, x56_1_1 );
 Register25Bit Reg111 (clk,x56_1_1, y146 );
 Register20Bit Reg112 (clk,x13, x13_1_1 );
 Register20Bit Reg113 (clk,x13_1_1, x13_1_2 );
 Register21Bit Reg114 (clk, {x13_1_2, 1'b0}, y0 );
 Register20Bit Reg115 (clk,x13, x13_2_1 );
 Register20Bit Reg116 (clk,x13_2_1, x13_2_2 );
 Register21Bit Reg117 (clk, {x13_2_2, 1'b0}, y150 );

 Adder18Bit Adder13(clk,  {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] },  { x2[14: 0], 3'b0 },x26); 

 Register19Bit Reg118 (clk,x26, x26_0_1 );
 Register19Bit Reg119 (clk,x26_0_1, x26_0_2 );
 Register22Bit Reg120 (clk, {x26_0_2, 3'b0}, y23 );
 Register19Bit Reg121 (clk,x26, x26_1_1 );
 Register19Bit Reg122 (clk,x26_1_1, x26_1_2 );
 Register22Bit Reg123 (clk, {x26_1_2, 3'b0}, y127 );

 Adder19Bit Adder14(clk,  {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] },  { x2[14: 0], 4'b0 },x27); 

 Negator20Bit Neg7(clk, x27, x94 );
 Register20Bit Reg124 (clk,x94, x94_0_1 );
 Register22Bit Reg125 (clk, {x94_0_1, 2'b0}, y25 );
 Register20Bit Reg126 (clk,x94, x94_1_1 );
 Register22Bit Reg127 (clk, {x94_1_1, 2'b0}, y125 );

 Subtractor21Bit Sub19(clk, { x1[14: 0], 6'b0 }, {x2[14],x2[14],x2[14],x2[14],x2[14],x2[14], x2[14: 0] }, x36); 

 Register22Bit Reg128 (clk,x36, x36_0_1 );
 Register22Bit Reg129 (clk,x36_0_1, x36_0_2 );
 Register23Bit Reg130 (clk, {x36_0_2, 1'b0}, y13 );
 Register22Bit Reg131 (clk,x36, x36_1_1 );
 Register22Bit Reg132 (clk,x36_1_1, x36_1_2 );
 Register23Bit Reg133 (clk, {x36_1_2, 1'b0}, y137 );

 Subtractor21Bit Sub20(clk, { x2[14: 0], 6'b0 }, {x1[14],x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0] }, x37); 

 Register22Bit Reg134 (clk,x37, x37_0_1 );
 Register22Bit Reg135 (clk,x37_0_1, x37_0_2 );
 Register22Bit Reg136 (clk,x37_0_2, y27 );
 Register22Bit Reg137 (clk,x37, x37_1_1 );
 Register22Bit Reg138 (clk,x37_1_1, x37_1_2 );
 Register22Bit Reg139 (clk,x37_1_2, y123 );

 Subtractor20Bit Sub21(clk, {x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0] },  { x2[14: 0], 5'b0 },x38); 

 Register21Bit Reg140 (clk,x38, x38_0_1 );
 Register21Bit Reg141 (clk,x38_0_1, x38_0_2 );
 Register22Bit Reg142 (clk, {x38_0_2, 1'b0}, y29 );
 Register21Bit Reg143 (clk,x38, x38_1_1 );
 Register21Bit Reg144 (clk,x38_1_1, x38_1_2 );
 Register22Bit Reg145 (clk, {x38_1_2, 1'b0}, y121 );

 Subtractor22Bit Sub22(clk, { x2[14: 0], 7'b0 }, {x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0] }, x39); 

 Register23Bit Reg146 (clk,x39, x39_0_1 );
 Register23Bit Reg147 (clk,x39_0_1, x39_0_2 );
 Register28Bit Reg148 (clk, {x39_0_2, 5'b0}, y74 );
 Register23Bit Reg149 (clk,x39, x39_1_1 );
 Register23Bit Reg150 (clk,x39_1_1, x39_1_2 );
 Register28Bit Reg151 (clk, {x39_1_2, 5'b0}, y76 );

 Adder21Bit Adder15(clk,  { x2[14: 0], 6'b0 }, {x5[17],x5[17],x5[17], x5[17: 0]  }, x62); 

 Register22Bit Reg152 (clk,x62, x62_0_1 );
 Register23Bit Reg153 (clk, {x62_0_1, 1'b0}, y50 );
 Register22Bit Reg154 (clk,x62, x62_1_1 );
 Register23Bit Reg155 (clk, {x62_1_1, 1'b0}, y100 );

 Adder23Bit Adder16(clk,  {x2[14],x2[14],x2[14],x2[14],x2[14],x2[14],x2[14],x2[14], x2[14: 0] },  { x6[17: 0], 5'b0 },x63); 

 Negator24Bit Neg8(clk, x63, x92 );
 Register24Bit Reg156 (clk,x92, y19 );
 Register24Bit Reg157 (clk,x92, y131 );

 Subtractor21Bit Sub23(clk, {x6[17],x6[17],x6[17], x6[17: 0] },  { x2[14: 0], 6'b0 },x64); 

 Register22Bit Reg158 (clk,x64, x64_0_1 );
 Register22Bit Reg159 (clk,x64_0_1, y33 );
 Register22Bit Reg160 (clk,x64, x64_1_1 );
 Register22Bit Reg161 (clk,x64_1_1, y117 );

 Adder23Bit Adder17(clk,  {x2[14],x2[14],x2[14],x2[14],x2[14], x2[14: 0], 3'b0 }, { x9[22: 0]  }, x65); 

 Register24Bit Reg162 (clk,x65, x65_0_1 );
 Register24Bit Reg163 (clk,x65_0_1, y37 );
 Register24Bit Reg164 (clk,x65, x65_1_1 );
 Register24Bit Reg165 (clk,x65_1_1, y113 );

 Subtractor23Bit Sub24(clk, {x2[14],x2[14],x2[14],x2[14],x2[14], x2[14: 0], 3'b0 }, { x9[22: 0] }, x66); 

 Register24Bit Reg166 (clk,x66, x66_0_1 );
 Register24Bit Reg167 (clk,x66_0_1, y63 );
 Register24Bit Reg168 (clk,x66, x66_1_1 );
 Register24Bit Reg169 (clk,x66_1_1, y87 );

 Subtractor24Bit Sub25(clk, { x12[18: 0], 5'b0 }, {x2[14],x2[14],x2[14],x2[14],x2[14],x2[14],x2[14],x2[14],x2[14], x2[14: 0] }, x68); 

 Register25Bit Reg170 (clk,x68, x68_0_1 );
 Register25Bit Reg171 (clk,x68_0_1, y1 );
 Register25Bit Reg172 (clk,x68, x68_1_1 );
 Register25Bit Reg173 (clk,x68_1_1, y149 );

 Subtractor22Bit Sub26(clk, { x25[21: 0] },  {x2[14],x2[14],x2[14], x2[14: 0], 4'b0 },x70); 

 Register23Bit Reg174 (clk,x70, x70_0_1 );
 Register23Bit Reg175 (clk,x70_0_1, y48 );
 Register23Bit Reg176 (clk,x70, x70_1_1 );
 Register23Bit Reg177 (clk,x70_1_1, y102 );
 Negator15Bit Neg9(clk, x2, x97 );
 Register15Bit Reg178 (clk,x97, x97_0_1 );
 Register15Bit Reg179 (clk,x97_0_1, x97_0_2 );
 Register21Bit Reg180 (clk, {x97_0_2, 6'b0}, y36 );
 Register15Bit Reg181 (clk,x97, x97_1_1 );
 Register15Bit Reg182 (clk,x97_1_1, x97_1_2 );
 Register21Bit Reg183 (clk, {x97_1_2, 6'b0}, y114 );

 Adder15Bit Adder18(clk,  {x0[11],x0[11],x0[11], x0[11: 0] },  { x0[11: 0], 3'b0 },x3); 


 Subtractor20Bit Sub27(clk, {x3[15],x3[15],x3[15],x3[15], x3[15: 0] },  { x1[14: 0], 5'b0 },x15); 

 Negator21Bit Neg10(clk, x15, x104 );
 Register21Bit Reg184 (clk,x104, x104_0_1 );
 Register23Bit Reg185 (clk, {x104_0_1, 2'b0}, y61 );
 Register21Bit Reg186 (clk,x104, x104_1_1 );
 Register23Bit Reg187 (clk, {x104_1_1, 2'b0}, y89 );
 Register21Bit Reg188 (clk,x15, x15_1_1 );
 Register21Bit Reg189 (clk,x15_1_1, x15_1_2 );
 Register22Bit Reg190 (clk, {x15_1_2, 1'b0}, y26 );
 Register21Bit Reg191 (clk,x15, x15_2_1 );
 Register21Bit Reg192 (clk,x15_2_1, x15_2_2 );
 Register22Bit Reg193 (clk, {x15_2_2, 1'b0}, y124 );

 Subtractor19Bit Sub28(clk, {x3[15],x3[15],x3[15], x3[15: 0] },  { x0[11: 0], 7'b0 },x28); 

 Register20Bit Reg194 (clk,x28, x28_0_1 );
 Register20Bit Reg195 (clk,x28_0_1, x28_0_2 );
 Register21Bit Reg196 (clk, {x28_0_2, 1'b0}, y16 );
 Register20Bit Reg197 (clk,x28, x28_1_1 );
 Register20Bit Reg198 (clk,x28_1_1, x28_1_2 );
 Register21Bit Reg199 (clk, {x28_1_2, 1'b0}, y134 );

 Adder20Bit Adder19(clk,  { x0[11: 0], 8'b0 }, {x3[15],x3[15],x3[15],x3[15], x3[15: 0]  }, x29); 

 Negator21Bit Neg11(clk, x29, x96 );
 Register21Bit Reg200 (clk,x96, x96_0_1 );
 Register21Bit Reg201 (clk,x96_0_1, y32 );
 Register21Bit Reg202 (clk,x96, x96_1_1 );
 Register21Bit Reg203 (clk,x96_1_1, y118 );

 Adder19Bit Adder20(clk,  { x0[11: 0], 7'b0 }, {x3[15],x3[15],x3[15], x3[15: 0]  }, x30); 

 Register20Bit Reg204 (clk,x30, x30_0_1 );
 Register20Bit Reg205 (clk,x30_0_1, x30_0_2 );
 Register23Bit Reg206 (clk, {x30_0_2, 3'b0}, y58 );
 Register20Bit Reg207 (clk,x30, x30_1_1 );
 Register20Bit Reg208 (clk,x30_1_1, x30_1_2 );
 Register23Bit Reg209 (clk, {x30_1_2, 3'b0}, y92 );

 Adder21Bit Adder21(clk,  {x1[14],x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0] },  { x3[15: 0], 5'b0 },x40); 

 Register22Bit Reg210 (clk,x40, x40_0_1 );
 Register22Bit Reg211 (clk,x40_0_1, x40_0_2 );
 Register22Bit Reg212 (clk,x40_0_2, y14 );
 Register22Bit Reg213 (clk,x40, x40_1_1 );
 Register22Bit Reg214 (clk,x40_1_1, x40_1_2 );
 Register22Bit Reg215 (clk,x40_1_2, y136 );

 Subtractor21Bit Sub29(clk, { x3[15: 0], 5'b0 }, {x1[14],x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0] }, x41); 

 Register22Bit Reg216 (clk,x41, x41_0_1 );
 Register22Bit Reg217 (clk,x41_0_1, x41_0_2 );
 Register22Bit Reg218 (clk,x41_0_2, y34 );
 Register22Bit Reg219 (clk,x41, x41_1_1 );
 Register22Bit Reg220 (clk,x41_1_1, x41_1_2 );
 Register22Bit Reg221 (clk,x41_1_2, y116 );

 Subtractor21Bit Sub30(clk, {x3[15],x3[15],x3[15],x3[15],x3[15], x3[15: 0] },  { x1[14: 0], 6'b0 },x42); 

 Register22Bit Reg222 (clk,x42, x42_0_1 );
 Register22Bit Reg223 (clk,x42_0_1, x42_0_2 );
 Register23Bit Reg224 (clk, {x42_0_2, 1'b0}, y55 );
 Register22Bit Reg225 (clk,x42, x42_1_1 );
 Register22Bit Reg226 (clk,x42_1_1, x42_1_2 );
 Register23Bit Reg227 (clk, {x42_1_2, 1'b0}, y95 );

 Adder20Bit Adder22(clk,  { x2[14: 0], 5'b0 }, {x3[15],x3[15],x3[15],x3[15], x3[15: 0]  }, x58); 

 Negator21Bit Neg12(clk, x58, x93 );
 Register21Bit Reg228 (clk,x93, x93_0_1 );
 Register22Bit Reg229 (clk, {x93_0_1, 1'b0}, y21 );
 Register21Bit Reg230 (clk,x93, x93_1_1 );
 Register22Bit Reg231 (clk, {x93_1_1, 1'b0}, y129 );

 Subtractor23Bit Sub31(clk, {x3[15],x3[15],x3[15],x3[15],x3[15],x3[15],x3[15], x3[15: 0] },  { x2[14: 0], 8'b0 },x59); 

 Register24Bit Reg232 (clk,x59, x59_0_1 );
 Register24Bit Reg233 (clk,x59_0_1, x59_0_2 );
 Register24Bit Reg234 (clk,x59_0_2, y60 );
 Register24Bit Reg235 (clk,x59, x59_1_1 );
 Register24Bit Reg236 (clk,x59_1_1, x59_1_2 );
 Register24Bit Reg237 (clk,x59_1_2, y90 );

 Subtractor23Bit Sub32(clk, {x3[15],x3[15],x3[15],x3[15],x3[15],x3[15],x3[15], x3[15: 0] },  { x11[17: 0], 5'b0 },x71); 

 Register24Bit Reg238 (clk,x71, x71_0_1 );
 Register27Bit Reg239 (clk, {x71_0_1, 3'b0}, y72 );
 Register24Bit Reg240 (clk,x71, x71_1_1 );
 Register27Bit Reg241 (clk, {x71_1_1, 3'b0}, y78 );

 Adder23Bit Adder23(clk,  {x3[15],x3[15],x3[15],x3[15],x3[15],x3[15],x3[15], x3[15: 0] },  { x21[17: 0], 5'b0 },x72); 

 Register24Bit Reg242 (clk,x72, x72_0_1 );
 Register25Bit Reg243 (clk, {x72_0_1, 1'b0}, y3 );
 Register24Bit Reg244 (clk,x72, x72_1_1 );
 Register25Bit Reg245 (clk, {x72_1_1, 1'b0}, y147 );

 Subtractor15Bit Sub33(clk, { x0[11: 0], 3'b0 }, {x0[11],x0[11],x0[11], x0[11: 0] }, x4); 


 Adder20Bit Adder24(clk,  {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] },  { x4[15: 0], 4'b0 },x31); 

 Negator21Bit Neg13(clk, x31, x95 );
 Register21Bit Reg246 (clk,x95, x95_0_1 );
 Register22Bit Reg247 (clk, {x95_0_1, 1'b0}, y28 );
 Register21Bit Reg248 (clk,x95, x95_1_1 );
 Register22Bit Reg249 (clk, {x95_1_1, 1'b0}, y122 );

 Subtractor19Bit Sub34(clk, { x0[11: 0], 7'b0 }, {x4[15],x4[15],x4[15], x4[15: 0] }, x32); 

 Register20Bit Reg250 (clk,x32, x32_0_1 );
 Register20Bit Reg251 (clk,x32_0_1, x32_0_2 );
 Register21Bit Reg252 (clk, {x32_0_2, 1'b0}, y30 );
 Register20Bit Reg253 (clk,x32, x32_1_1 );
 Register20Bit Reg254 (clk,x32_1_1, x32_1_2 );
 Register21Bit Reg255 (clk, {x32_1_2, 1'b0}, y120 );

 Subtractor21Bit Sub35(clk, { x1[14: 0], 6'b0 }, {x4[15],x4[15],x4[15],x4[15],x4[15], x4[15: 0] }, x43); 

 Register22Bit Reg256 (clk,x43, x43_0_1 );
 Register22Bit Reg257 (clk,x43_0_1, x43_0_2 );
 Register22Bit Reg258 (clk,x43_0_2, y20 );
 Register22Bit Reg259 (clk,x43, x43_1_1 );
 Register22Bit Reg260 (clk,x43_1_1, x43_1_2 );
 Register22Bit Reg261 (clk,x43_1_2, y130 );

 Adder22Bit Adder25(clk,  { x1[14: 0], 7'b0 }, {x4[15],x4[15],x4[15],x4[15],x4[15],x4[15], x4[15: 0]  }, x44); 

 Negator23Bit Neg14(clk, x44, x100 );
 Register23Bit Reg262 (clk,x100, x100_0_1 );
 Register23Bit Reg263 (clk,x100_0_1, y47 );
 Register23Bit Reg264 (clk,x100, x100_1_1 );
 Register23Bit Reg265 (clk,x100_1_1, y103 );

 Subtractor24Bit Sub36(clk, {x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0] },  { x4[15: 0], 8'b0 },x45); 

 Register25Bit Reg266 (clk,x45, x45_0_1 );
 Register25Bit Reg267 (clk,x45_0_1, x45_0_2 );
 Register25Bit Reg268 (clk,x45_0_2, y64 );
 Register25Bit Reg269 (clk,x45, x45_1_1 );
 Register25Bit Reg270 (clk,x45_1_1, x45_1_2 );
 Register25Bit Reg271 (clk,x45_1_2, y86 );

 Adder20Bit Adder26(clk,  {x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0] },  { x4[15: 0], 4'b0 },x46); 

 Negator21Bit Neg15(clk, x46, x107 );
 Register21Bit Reg272 (clk,x107, x107_0_1 );
 Register23Bit Reg273 (clk, {x107_0_1, 2'b0}, y73 );
 Register21Bit Reg274 (clk,x107, x107_1_1 );
 Register23Bit Reg275 (clk, {x107_1_1, 2'b0}, y77 );

 Adder24Bit Adder27(clk,  {x2[14],x2[14],x2[14],x2[14],x2[14],x2[14],x2[14],x2[14],x2[14], x2[14: 0] },  { x4[15: 0], 8'b0 },x60); 

 Negator25Bit Neg16(clk, x60, x88 );
 Register25Bit Reg276 (clk,x88, x88_0_1 );
 Register25Bit Reg277 (clk,x88_0_1, y2 );
 Register25Bit Reg278 (clk,x88, x88_1_1 );
 Register25Bit Reg279 (clk,x88_1_1, y148 );

 Adder21Bit Adder28(clk,  { x2[14: 0], 6'b0 }, {x4[15],x4[15],x4[15],x4[15],x4[15], x4[15: 0]  }, x61); 

 Register22Bit Reg280 (clk,x61, x61_0_1 );
 Register22Bit Reg281 (clk,x61_0_1, x61_0_2 );
 Register22Bit Reg282 (clk,x61_0_2, y31 );
 Register22Bit Reg283 (clk,x61, x61_1_1 );
 Register22Bit Reg284 (clk,x61_1_1, x61_1_2 );
 Register22Bit Reg285 (clk,x61_1_2, y119 );

 Subtractor16Bit Sub37(clk, {x0[11],x0[11],x0[11],x0[11], x0[11: 0] },  { x0[11: 0], 4'b0 },x7); 


 Adder22Bit Adder29(clk,  {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] },  { x7[16: 0], 5'b0 },x14); 

 Register23Bit Reg286 (clk,x14, x14_0_1 );
 Register23Bit Reg287 (clk,x14_0_1, x14_0_2 );
 Register23Bit Reg288 (clk,x14_0_2, y44 );
 Register23Bit Reg289 (clk,x14, x14_1_1 );
 Register23Bit Reg290 (clk,x14_1_1, x14_1_2 );
 Register24Bit Reg291 (clk, {x14_1_2, 1'b0}, y56 );
 Register23Bit Reg292 (clk,x14, x14_2_1 );
 Register23Bit Reg293 (clk,x14_2_1, x14_2_2 );
 Register24Bit Reg294 (clk, {x14_2_2, 1'b0}, y94 );
 Register23Bit Reg295 (clk,x14, x14_3_1 );
 Register23Bit Reg296 (clk,x14_3_1, x14_3_2 );
 Register23Bit Reg297 (clk,x14_3_2, y106 );

 Adder24Bit Adder30(clk,  { x0[11: 0], 12'b0 }, {x7[16],x7[16],x7[16],x7[16],x7[16],x7[16],x7[16], x7[16: 0]  }, x33); 

 Register25Bit Reg298 (clk,x33, x33_0_1 );
 Register25Bit Reg299 (clk,x33_0_1, x33_0_2 );
 Register25Bit Reg300 (clk,x33_0_2, y70 );
 Register25Bit Reg301 (clk,x33, x33_1_1 );
 Register25Bit Reg302 (clk,x33_1_1, x33_1_2 );
 Register25Bit Reg303 (clk,x33_1_2, y80 );

 Subtractor22Bit Sub38(clk, { x1[14: 0], 7'b0 }, {x7[16],x7[16],x7[16],x7[16],x7[16], x7[16: 0] }, x54); 

 Register23Bit Reg304 (clk,x54, x54_0_1 );
 Register23Bit Reg305 (clk,x54_0_1, x54_0_2 );
 Register23Bit Reg306 (clk,x54_0_2, y12 );
 Register23Bit Reg307 (clk,x54, x54_1_1 );
 Register23Bit Reg308 (clk,x54_1_1, x54_1_2 );
 Register23Bit Reg309 (clk,x54_1_2, y138 );

 Subtractor19Bit Sub39(clk, {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] },  { x0[11: 0], 7'b0 },x19); 

 Negator20Bit Neg17(clk, x19, x90 );
 Register20Bit Reg310 (clk,x90, x90_0_1 );
 Register20Bit Reg311 (clk,x90_0_1, x90_0_2 );
 Register22Bit Reg312 (clk, {x90_0_2, 2'b0}, y10 );
 Register20Bit Reg313 (clk,x90, x90_1_1 );
 Register20Bit Reg314 (clk,x90_1_1, x90_1_2 );
 Register22Bit Reg315 (clk, {x90_1_2, 2'b0}, y140 );

 Subtractor22Bit Sub40(clk, {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] },  { x0[11: 0], 10'b0 },x20); 


 Subtractor23Bit Sub41(clk, {x2[14],x2[14],x2[14],x2[14],x2[14], x2[14: 0], 3'b0 }, { x20[22: 0] }, x69); 

 Register24Bit Reg316 (clk,x69, x69_0_1 );
 Register24Bit Reg317 (clk,x69_0_1, x69_0_2 );
 Register24Bit Reg318 (clk,x69_0_2, y6 );
 Register24Bit Reg319 (clk,x69, x69_1_1 );
 Register24Bit Reg320 (clk,x69_1_1, x69_1_2 );
 Register24Bit Reg321 (clk,x69_1_2, y144 );
 Register12Bit Reg322 (clk,x0, x74_36_1 );
 Register12Bit Reg323 (clk,x74_36_1, x74_36_2 );

 Adder24Bit Adder31(clk,  {x74_36_2[11],x74_36_2[11],x74_36_2[11],x74_36_2[11],x74_36_2[11],x74_36_2[11],x74_36_2[11],x74_36_2[11],x74_36_2[11],x74_36_2[11],x74_36_2[11],x74_36_2[11], x74_36_2[11: 0] },  { x8[18: 0], 5'b0 },x74); 

 Register25Bit Reg324 (clk,x74, x74_0_1 );
 Register25Bit Reg325 (clk,x74_0_1, y8 );
 Register12Bit Reg326 (clk,x0, x75_37_1 );
 Register12Bit Reg327 (clk,x75_37_1, x75_37_2 );

 Adder23Bit Adder32(clk,  {x75_37_2[11],x75_37_2[11],x75_37_2[11],x75_37_2[11],x75_37_2[11],x75_37_2[11],x75_37_2[11],x75_37_2[11],x75_37_2[11],x75_37_2[11],x75_37_2[11], x75_37_2[11: 0] },  { x6[17: 0], 5'b0 },x75); 

 Negator24Bit Neg18(clk, x75, x98 );
 Register24Bit Reg328 (clk,x98, y38 );
 Register12Bit Reg329 (clk,x0, x76_38_1 );
 Register12Bit Reg330 (clk,x76_38_1, x76_38_2 );

 Subtractor21Bit Sub42(clk, { x76_38_2[11: 0], 9'b0 }, {x8[18],x8[18], x8[18: 0] }, x76); 

 Register22Bit Reg331 (clk,x76, x76_0_1 );
 Register22Bit Reg332 (clk,x76_0_1, y46 );
 Register12Bit Reg333 (clk,x0, x77_39_1 );
 Register12Bit Reg334 (clk,x77_39_1, x77_39_2 );

 Subtractor19Bit Sub43(clk, { x77_39_2[11: 0], 7'b0 }, {x6[17], x6[17: 0] }, x77); 

 Register20Bit Reg335 (clk,x77, x77_0_1 );
 Register24Bit Reg336 (clk, {x77_0_1, 4'b0}, y66 );
 Register12Bit Reg337 (clk,x0, x78_40_1 );
 Register12Bit Reg338 (clk,x78_40_1, x78_40_2 );

 Subtractor21Bit Sub44(clk, { x11[17: 0], 3'b0 }, {x78_40_2[11],x78_40_2[11],x78_40_2[11],x78_40_2[11],x78_40_2[11],x78_40_2[11],x78_40_2[11],x78_40_2[11],x78_40_2[11], x78_40_2[11: 0] }, x78); 

 Register22Bit Reg339 (clk,x78, x78_0_1 );
 Register23Bit Reg340 (clk, {x78_0_1, 1'b0}, y67 );
 Register12Bit Reg341 (clk,x0, x79_41_1 );
 Register12Bit Reg342 (clk,x79_41_1, x79_41_2 );

 Adder22Bit Adder33(clk,  {x79_41_2[11],x79_41_2[11],x79_41_2[11],x79_41_2[11],x79_41_2[11],x79_41_2[11],x79_41_2[11],x79_41_2[11],x79_41_2[11],x79_41_2[11], x79_41_2[11: 0] },  { x11[17: 0], 4'b0 },x79); 

 Negator23Bit Neg19(clk, x79, x106 );
 Register23Bit Reg343 (clk,x106, y69 );
 Register12Bit Reg344 (clk,x0, x80_42_1 );
 Register12Bit Reg345 (clk,x80_42_1, x80_42_2 );

 Adder21Bit Adder34(clk,  {x80_42_2[11],x80_42_2[11],x80_42_2[11],x80_42_2[11],x80_42_2[11],x80_42_2[11],x80_42_2[11],x80_42_2[11],x80_42_2[11], x80_42_2[11: 0] },  { x11[17: 0], 3'b0 },x80); 

 Register22Bit Reg346 (clk,x80, x80_0_1 );
 Register23Bit Reg347 (clk, {x80_0_1, 1'b0}, y71 );
 Register12Bit Reg348 (clk,x0, x81_43_1 );
 Register12Bit Reg349 (clk,x81_43_1, x81_43_2 );

 Adder21Bit Adder35(clk,  {x81_43_2[11],x81_43_2[11],x81_43_2[11],x81_43_2[11],x81_43_2[11],x81_43_2[11],x81_43_2[11],x81_43_2[11],x81_43_2[11], x81_43_2[11: 0] },  { x11[17: 0], 3'b0 },x81); 

 Register22Bit Reg350 (clk,x81, x81_0_1 );
 Register23Bit Reg351 (clk, {x81_0_1, 1'b0}, y79 );
 Register12Bit Reg352 (clk,x0, x82_44_1 );
 Register12Bit Reg353 (clk,x82_44_1, x82_44_2 );

 Adder22Bit Adder36(clk,  {x82_44_2[11],x82_44_2[11],x82_44_2[11],x82_44_2[11],x82_44_2[11],x82_44_2[11],x82_44_2[11],x82_44_2[11],x82_44_2[11],x82_44_2[11], x82_44_2[11: 0] },  { x11[17: 0], 4'b0 },x82); 

 Negator23Bit Neg20(clk, x82, x108 );
 Register23Bit Reg354 (clk,x108, y81 );
 Register12Bit Reg355 (clk,x0, x83_45_1 );
 Register12Bit Reg356 (clk,x83_45_1, x83_45_2 );

 Subtractor21Bit Sub45(clk, { x11[17: 0], 3'b0 }, {x83_45_2[11],x83_45_2[11],x83_45_2[11],x83_45_2[11],x83_45_2[11],x83_45_2[11],x83_45_2[11],x83_45_2[11],x83_45_2[11], x83_45_2[11: 0] }, x83); 

 Register22Bit Reg357 (clk,x83, x83_0_1 );
 Register23Bit Reg358 (clk, {x83_0_1, 1'b0}, y83 );
 Register12Bit Reg359 (clk,x0, x84_46_1 );
 Register12Bit Reg360 (clk,x84_46_1, x84_46_2 );

 Subtractor19Bit Sub46(clk, { x84_46_2[11: 0], 7'b0 }, {x6[17], x6[17: 0] }, x84); 

 Register20Bit Reg361 (clk,x84, x84_0_1 );
 Register24Bit Reg362 (clk, {x84_0_1, 4'b0}, y84 );
 Register12Bit Reg363 (clk,x0, x85_47_1 );
 Register12Bit Reg364 (clk,x85_47_1, x85_47_2 );

 Subtractor21Bit Sub47(clk, { x85_47_2[11: 0], 9'b0 }, {x8[18],x8[18], x8[18: 0] }, x85); 

 Register22Bit Reg365 (clk,x85, x85_0_1 );
 Register22Bit Reg366 (clk,x85_0_1, y104 );
 Register12Bit Reg367 (clk,x0, x86_48_1 );
 Register12Bit Reg368 (clk,x86_48_1, x86_48_2 );

 Adder23Bit Adder37(clk,  {x86_48_2[11],x86_48_2[11],x86_48_2[11],x86_48_2[11],x86_48_2[11],x86_48_2[11],x86_48_2[11],x86_48_2[11],x86_48_2[11],x86_48_2[11],x86_48_2[11], x86_48_2[11: 0] },  { x6[17: 0], 5'b0 },x86); 

 Negator24Bit Neg21(clk, x86, x109 );
 Register24Bit Reg369 (clk,x109, y112 );
 Register12Bit Reg370 (clk,x0, x87_49_1 );
 Register12Bit Reg371 (clk,x87_49_1, x87_49_2 );

 Adder24Bit Adder38(clk,  {x87_49_2[11],x87_49_2[11],x87_49_2[11],x87_49_2[11],x87_49_2[11],x87_49_2[11],x87_49_2[11],x87_49_2[11],x87_49_2[11],x87_49_2[11],x87_49_2[11],x87_49_2[11], x87_49_2[11: 0] },  { x8[18: 0], 5'b0 },x87); 

 Register25Bit Reg372 (clk,x87, x87_0_1 );
 Register25Bit Reg373 (clk,x87_0_1, y142 );
 Register12Bit Reg374 (clk,x0, x0_50_1 );
 Register12Bit Reg375 (clk,x0_50_1, x0_50_2 );
 Register12Bit Reg376 (clk,x0_50_2, x0_50_3 );
 Register12Bit Reg377 (clk,x0_50_3, x0_50_4 );
 Register27Bit Reg378 (clk, {x0_50_4, 15'b0}, y75 );
 Register21Bit Reg379 (clk,y0, x110 );

 Adder25Bit Adder39(clk,  {x110[20],x110[20],x110[20],x110[20], x110[20: 0] },  { y1[24: 0]  }, x111); 

 Register26Bit Reg380 (clk,x111, x111_1 );

 Adder26Bit Adder40(clk,  { x111_1[25: 0] },  {y2[24], y2[24: 0]  }, x112); 

 Register27Bit Reg381 (clk,x112, x112_1 );

 Adder27Bit Adder41(clk,  { x112_1[26: 0] },  {y3[24],y3[24], y3[24: 0]  }, x113); 

 Register28Bit Reg382 (clk,x113, x113_1 );

 Adder28Bit Adder42(clk,  { x113_1[27: 0] },  {y4[24],y4[24],y4[24], y4[24: 0]  }, x114); 

 Register29Bit Reg383 (clk,x114, x114_1 );

 Adder29Bit Adder43(clk,  { x114_1[28: 0] },  {y5[22],y5[22],y5[22],y5[22],y5[22],y5[22], y5[22: 0]  }, x115); 

 Register29Bit Reg384 (clk,x115, x115_1 );

 Adder29Bit Adder44(clk,  { x115_1[28: 0] },  {y6[23],y6[23],y6[23],y6[23],y6[23], y6[23: 0]  }, x116); 

 Register29Bit Reg385 (clk,x116, x116_1 );

 Adder29Bit Adder45(clk,  { x116_1[28: 0] },  {y7[21],y7[21],y7[21],y7[21],y7[21],y7[21],y7[21], y7[21: 0]  }, x117); 

 Register29Bit Reg386 (clk,x117, x117_1 );

 Adder29Bit Adder46(clk,  { x117_1[28: 0] },  {y8[24],y8[24],y8[24],y8[24], y8[24: 0]  }, x118); 

 Register29Bit Reg387 (clk,x118, x118_1 );

 Adder29Bit Adder47(clk,  { x118_1[28: 0] },  {y9[22],y9[22],y9[22],y9[22],y9[22],y9[22], y9[22: 0]  }, x119); 

 Register29Bit Reg388 (clk,x119, x119_1 );

 Adder29Bit Adder48(clk,  { x119_1[28: 0] },  {y10[21],y10[21],y10[21],y10[21],y10[21],y10[21],y10[21], y10[21: 0]  }, x120); 

 Register29Bit Reg389 (clk,x120, x120_1 );

 Adder29Bit Adder49(clk,  { x120_1[28: 0] },  {y11[22],y11[22],y11[22],y11[22],y11[22],y11[22], y11[22: 0]  }, x121); 

 Register29Bit Reg390 (clk,x121, x121_1 );

 Adder29Bit Adder50(clk,  { x121_1[28: 0] },  {y12[22],y12[22],y12[22],y12[22],y12[22],y12[22], y12[22: 0]  }, x122); 

 Register29Bit Reg391 (clk,x122, x122_1 );

 Adder29Bit Adder51(clk,  { x122_1[28: 0] },  {y13[22],y13[22],y13[22],y13[22],y13[22],y13[22], y13[22: 0]  }, x123); 

 Register29Bit Reg392 (clk,x123, x123_1 );

 Adder29Bit Adder52(clk,  { x123_1[28: 0] },  {y14[21],y14[21],y14[21],y14[21],y14[21],y14[21],y14[21], y14[21: 0]  }, x124); 

 Register29Bit Reg393 (clk,x124, x124_1 );

 Adder29Bit Adder53(clk,  { x124_1[28: 0] },  {y15[22],y15[22],y15[22],y15[22],y15[22],y15[22], y15[22: 0]  }, x125); 

 Register29Bit Reg394 (clk,x125, x125_1 );

 Adder29Bit Adder54(clk,  { x125_1[28: 0] },  {y16[20],y16[20],y16[20],y16[20],y16[20],y16[20],y16[20],y16[20], y16[20: 0]  }, x126); 

 Register29Bit Reg395 (clk,x126, x126_1 );

 Adder29Bit Adder55(clk,  { x126_1[28: 0] },  {y17[22],y17[22],y17[22],y17[22],y17[22],y17[22], y17[22: 0]  }, x127); 

 Register29Bit Reg396 (clk,x127, x127_1 );

 Adder29Bit Adder56(clk,  { x127_1[28: 0] },  {y18[22],y18[22],y18[22],y18[22],y18[22],y18[22], y18[22: 0]  }, x128); 

 Register29Bit Reg397 (clk,x128, x128_1 );

 Adder29Bit Adder57(clk,  { x128_1[28: 0] },  {y19[23],y19[23],y19[23],y19[23],y19[23], y19[23: 0]  }, x129); 

 Register29Bit Reg398 (clk,x129, x129_1 );

 Adder29Bit Adder58(clk,  { x129_1[28: 0] },  {y20[21],y20[21],y20[21],y20[21],y20[21],y20[21],y20[21], y20[21: 0]  }, x130); 

 Register29Bit Reg399 (clk,x130, x130_1 );

 Adder29Bit Adder59(clk,  { x130_1[28: 0] },  {y21[21],y21[21],y21[21],y21[21],y21[21],y21[21],y21[21], y21[21: 0]  }, x131); 

 Register29Bit Reg400 (clk,x131, x131_1 );

 Adder29Bit Adder60(clk,  { x131_1[28: 0] },  {y22[21],y22[21],y22[21],y22[21],y22[21],y22[21],y22[21], y22[21: 0]  }, x132); 

 Register29Bit Reg401 (clk,x132, x132_1 );

 Adder29Bit Adder61(clk,  { x132_1[28: 0] },  {y23[21],y23[21],y23[21],y23[21],y23[21],y23[21],y23[21], y23[21: 0]  }, x133); 

 Register29Bit Reg402 (clk,x133, x133_1 );

 Adder29Bit Adder62(clk,  { x133_1[28: 0] },  {y24[21],y24[21],y24[21],y24[21],y24[21],y24[21],y24[21], y24[21: 0]  }, x134); 

 Register29Bit Reg403 (clk,x134, x134_1 );

 Adder29Bit Adder63(clk,  { x134_1[28: 0] },  {y25[21],y25[21],y25[21],y25[21],y25[21],y25[21],y25[21], y25[21: 0]  }, x135); 

 Register29Bit Reg404 (clk,x135, x135_1 );

 Adder29Bit Adder64(clk,  { x135_1[28: 0] },  {y26[21],y26[21],y26[21],y26[21],y26[21],y26[21],y26[21], y26[21: 0]  }, x136); 

 Register29Bit Reg405 (clk,x136, x136_1 );

 Adder29Bit Adder65(clk,  { x136_1[28: 0] },  {y27[21],y27[21],y27[21],y27[21],y27[21],y27[21],y27[21], y27[21: 0]  }, x137); 

 Register29Bit Reg406 (clk,x137, x137_1 );

 Adder29Bit Adder66(clk,  { x137_1[28: 0] },  {y28[21],y28[21],y28[21],y28[21],y28[21],y28[21],y28[21], y28[21: 0]  }, x138); 

 Register29Bit Reg407 (clk,x138, x138_1 );

 Adder29Bit Adder67(clk,  { x138_1[28: 0] },  {y29[21],y29[21],y29[21],y29[21],y29[21],y29[21],y29[21], y29[21: 0]  }, x139); 

 Register29Bit Reg408 (clk,x139, x139_1 );

 Adder29Bit Adder68(clk,  { x139_1[28: 0] },  {y30[20],y30[20],y30[20],y30[20],y30[20],y30[20],y30[20],y30[20], y30[20: 0]  }, x140); 

 Register29Bit Reg409 (clk,x140, x140_1 );

 Adder29Bit Adder69(clk,  { x140_1[28: 0] },  {y31[21],y31[21],y31[21],y31[21],y31[21],y31[21],y31[21], y31[21: 0]  }, x141); 

 Register29Bit Reg410 (clk,x141, x141_1 );

 Adder29Bit Adder70(clk,  { x141_1[28: 0] },  {y32[20],y32[20],y32[20],y32[20],y32[20],y32[20],y32[20],y32[20], y32[20: 0]  }, x142); 

 Register29Bit Reg411 (clk,x142, x142_1 );

 Adder29Bit Adder71(clk,  { x142_1[28: 0] },  {y33[21],y33[21],y33[21],y33[21],y33[21],y33[21],y33[21], y33[21: 0]  }, x143); 

 Register29Bit Reg412 (clk,x143, x143_1 );

 Adder29Bit Adder72(clk,  { x143_1[28: 0] },  {y34[21],y34[21],y34[21],y34[21],y34[21],y34[21],y34[21], y34[21: 0]  }, x144); 

 Register29Bit Reg413 (clk,x144, x144_1 );

 Adder29Bit Adder73(clk,  { x144_1[28: 0] },  {y35[21],y35[21],y35[21],y35[21],y35[21],y35[21],y35[21], y35[21: 0]  }, x145); 

 Register29Bit Reg414 (clk,x145, x145_1 );

 Adder29Bit Adder74(clk,  { x145_1[28: 0] },  {y36[20],y36[20],y36[20],y36[20],y36[20],y36[20],y36[20],y36[20], y36[20: 0]  }, x146); 

 Register29Bit Reg415 (clk,x146, x146_1 );

 Adder29Bit Adder75(clk,  { x146_1[28: 0] },  {y37[23],y37[23],y37[23],y37[23],y37[23], y37[23: 0]  }, x147); 

 Register29Bit Reg416 (clk,x147, x147_1 );

 Adder29Bit Adder76(clk,  { x147_1[28: 0] },  {y38[23],y38[23],y38[23],y38[23],y38[23], y38[23: 0]  }, x148); 

 Register29Bit Reg417 (clk,x148, x148_1 );

 Adder29Bit Adder77(clk,  { x148_1[28: 0] },  {y39[23],y39[23],y39[23],y39[23],y39[23], y39[23: 0]  }, x149); 

 Register29Bit Reg418 (clk,x149, x149_1 );

 Adder29Bit Adder78(clk,  { x149_1[28: 0] },  {y40[22],y40[22],y40[22],y40[22],y40[22],y40[22], y40[22: 0]  }, x150); 

 Register29Bit Reg419 (clk,x150, x150_1 );

 Adder29Bit Adder79(clk,  { x150_1[28: 0] },  {y41[23],y41[23],y41[23],y41[23],y41[23], y41[23: 0]  }, x151); 

 Register29Bit Reg420 (clk,x151, x151_1 );

 Adder29Bit Adder80(clk,  { x151_1[28: 0] },  {y42[21],y42[21],y42[21],y42[21],y42[21],y42[21],y42[21], y42[21: 0]  }, x152); 

 Register29Bit Reg421 (clk,x152, x152_1 );

 Adder29Bit Adder81(clk,  { x152_1[28: 0] },  {y43[22],y43[22],y43[22],y43[22],y43[22],y43[22], y43[22: 0]  }, x153); 

 Register29Bit Reg422 (clk,x153, x153_1 );

 Adder29Bit Adder82(clk,  { x153_1[28: 0] },  {y44[22],y44[22],y44[22],y44[22],y44[22],y44[22], y44[22: 0]  }, x154); 

 Register29Bit Reg423 (clk,x154, x154_1 );

 Adder29Bit Adder83(clk,  { x154_1[28: 0] },  {y45[22],y45[22],y45[22],y45[22],y45[22],y45[22], y45[22: 0]  }, x155); 

 Register29Bit Reg424 (clk,x155, x155_1 );

 Adder29Bit Adder84(clk,  { x155_1[28: 0] },  {y46[21],y46[21],y46[21],y46[21],y46[21],y46[21],y46[21], y46[21: 0]  }, x156); 

 Register29Bit Reg425 (clk,x156, x156_1 );

 Adder29Bit Adder85(clk,  { x156_1[28: 0] },  {y47[22],y47[22],y47[22],y47[22],y47[22],y47[22], y47[22: 0]  }, x157); 

 Register29Bit Reg426 (clk,x157, x157_1 );

 Adder29Bit Adder86(clk,  { x157_1[28: 0] },  {y48[22],y48[22],y48[22],y48[22],y48[22],y48[22], y48[22: 0]  }, x158); 

 Register29Bit Reg427 (clk,x158, x158_1 );

 Adder29Bit Adder87(clk,  { x158_1[28: 0] },  {y49[22],y49[22],y49[22],y49[22],y49[22],y49[22], y49[22: 0]  }, x159); 

 Register29Bit Reg428 (clk,x159, x159_1 );

 Adder29Bit Adder88(clk,  { x159_1[28: 0] },  {y50[22],y50[22],y50[22],y50[22],y50[22],y50[22], y50[22: 0]  }, x160); 

 Register29Bit Reg429 (clk,x160, x160_1 );

 Adder29Bit Adder89(clk,  { x160_1[28: 0] },  {y51[22],y51[22],y51[22],y51[22],y51[22],y51[22], y51[22: 0]  }, x161); 

 Register29Bit Reg430 (clk,x161, x161_1 );

 Adder29Bit Adder90(clk,  { x161_1[28: 0] },  {y52[23],y52[23],y52[23],y52[23],y52[23], y52[23: 0]  }, x162); 

 Register29Bit Reg431 (clk,x162, x162_1 );

 Adder29Bit Adder91(clk,  { x162_1[28: 0] },  {y53[22],y53[22],y53[22],y53[22],y53[22],y53[22], y53[22: 0]  }, x163); 

 Register29Bit Reg432 (clk,x163, x163_1 );

 Adder29Bit Adder92(clk,  { x163_1[28: 0] },  {y54[24],y54[24],y54[24],y54[24], y54[24: 0]  }, x164); 

 Register29Bit Reg433 (clk,x164, x164_1 );

 Adder29Bit Adder93(clk,  { x164_1[28: 0] },  {y55[22],y55[22],y55[22],y55[22],y55[22],y55[22], y55[22: 0]  }, x165); 

 Register29Bit Reg434 (clk,x165, x165_1 );

 Adder29Bit Adder94(clk,  { x165_1[28: 0] },  {y56[23],y56[23],y56[23],y56[23],y56[23], y56[23: 0]  }, x166); 

 Register29Bit Reg435 (clk,x166, x166_1 );

 Adder29Bit Adder95(clk,  { x166_1[28: 0] },  {y57[23],y57[23],y57[23],y57[23],y57[23], y57[23: 0]  }, x167); 

 Register29Bit Reg436 (clk,x167, x167_1 );

 Adder29Bit Adder96(clk,  { x167_1[28: 0] },  {y58[22],y58[22],y58[22],y58[22],y58[22],y58[22], y58[22: 0]  }, x168); 

 Register29Bit Reg437 (clk,x168, x168_1 );

 Adder29Bit Adder97(clk,  { x168_1[28: 0] },  {y59[23],y59[23],y59[23],y59[23],y59[23], y59[23: 0]  }, x169); 

 Register29Bit Reg438 (clk,x169, x169_1 );

 Adder29Bit Adder98(clk,  { x169_1[28: 0] },  {y60[23],y60[23],y60[23],y60[23],y60[23], y60[23: 0]  }, x170); 

 Register29Bit Reg439 (clk,x170, x170_1 );

 Adder29Bit Adder99(clk,  { x170_1[28: 0] },  {y61[22],y61[22],y61[22],y61[22],y61[22],y61[22], y61[22: 0]  }, x171); 

 Register29Bit Reg440 (clk,x171, x171_1 );

 Adder29Bit Adder100(clk,  { x171_1[28: 0] },  {y62[24],y62[24],y62[24],y62[24], y62[24: 0]  }, x172); 

 Register29Bit Reg441 (clk,x172, x172_1 );

 Adder29Bit Adder101(clk,  { x172_1[28: 0] },  {y63[23],y63[23],y63[23],y63[23],y63[23], y63[23: 0]  }, x173); 

 Register29Bit Reg442 (clk,x173, x173_1 );

 Adder29Bit Adder102(clk,  { x173_1[28: 0] },  {y64[24],y64[24],y64[24],y64[24], y64[24: 0]  }, x174); 

 Register29Bit Reg443 (clk,x174, x174_1 );

 Adder29Bit Adder103(clk,  { x174_1[28: 0] },  {y65[22],y65[22],y65[22],y65[22],y65[22],y65[22], y65[22: 0]  }, x175); 

 Register29Bit Reg444 (clk,x175, x175_1 );

 Adder29Bit Adder104(clk,  { x175_1[28: 0] },  {y66[23],y66[23],y66[23],y66[23],y66[23], y66[23: 0]  }, x176); 

 Register29Bit Reg445 (clk,x176, x176_1 );

 Adder29Bit Adder105(clk,  { x176_1[28: 0] },  {y67[22],y67[22],y67[22],y67[22],y67[22],y67[22], y67[22: 0]  }, x177); 

 Register29Bit Reg446 (clk,x177, x177_1 );

 Adder29Bit Adder106(clk,  { x177_1[28: 0] },  {y68[26],y68[26], y68[26: 0]  }, x178); 

 Register29Bit Reg447 (clk,x178, x178_1 );

 Adder29Bit Adder107(clk,  { x178_1[28: 0] },  {y69[22],y69[22],y69[22],y69[22],y69[22],y69[22], y69[22: 0]  }, x179); 

 Register29Bit Reg448 (clk,x179, x179_1 );

 Adder29Bit Adder108(clk,  { x179_1[28: 0] },  {y70[24],y70[24],y70[24],y70[24], y70[24: 0]  }, x180); 

 Register29Bit Reg449 (clk,x180, x180_1 );

 Adder29Bit Adder109(clk,  { x180_1[28: 0] },  {y71[22],y71[22],y71[22],y71[22],y71[22],y71[22], y71[22: 0]  }, x181); 

 Register29Bit Reg450 (clk,x181, x181_1 );

 Adder29Bit Adder110(clk,  { x181_1[28: 0] },  {y72[26],y72[26], y72[26: 0]  }, x182); 

 Register29Bit Reg451 (clk,x182, x182_1 );

 Adder29Bit Adder111(clk,  { x182_1[28: 0] },  {y73[22],y73[22],y73[22],y73[22],y73[22],y73[22], y73[22: 0]  }, x183); 

 Register29Bit Reg452 (clk,x183, x183_1 );

 Adder29Bit Adder112(clk,  { x183_1[28: 0] },  {y74[27], y74[27: 0]  }, x184); 

 Register29Bit Reg453 (clk,x184, x184_1 );

 Adder29Bit Adder113(clk,  { x184_1[28: 0] },  {y75[26],y75[26], y75[26: 0]  }, x185); 

 Register29Bit Reg454 (clk,x185, x185_1 );

 Adder29Bit Adder114(clk,  { x185_1[28: 0] },  {y76[27], y76[27: 0]  }, x186); 

 Register29Bit Reg455 (clk,x186, x186_1 );

 Adder29Bit Adder115(clk,  { x186_1[28: 0] },  {y77[22],y77[22],y77[22],y77[22],y77[22],y77[22], y77[22: 0]  }, x187); 

 Register29Bit Reg456 (clk,x187, x187_1 );

 Adder29Bit Adder116(clk,  { x187_1[28: 0] },  {y78[26],y78[26], y78[26: 0]  }, x188); 

 Register29Bit Reg457 (clk,x188, x188_1 );

 Adder29Bit Adder117(clk,  { x188_1[28: 0] },  {y79[22],y79[22],y79[22],y79[22],y79[22],y79[22], y79[22: 0]  }, x189); 

 Register29Bit Reg458 (clk,x189, x189_1 );

 Adder29Bit Adder118(clk,  { x189_1[28: 0] },  {y80[24],y80[24],y80[24],y80[24], y80[24: 0]  }, x190); 

 Register29Bit Reg459 (clk,x190, x190_1 );

 Adder29Bit Adder119(clk,  { x190_1[28: 0] },  {y81[22],y81[22],y81[22],y81[22],y81[22],y81[22], y81[22: 0]  }, x191); 

 Register29Bit Reg460 (clk,x191, x191_1 );

 Adder29Bit Adder120(clk,  { x191_1[28: 0] },  {y82[26],y82[26], y82[26: 0]  }, x192); 

 Register29Bit Reg461 (clk,x192, x192_1 );

 Adder29Bit Adder121(clk,  { x192_1[28: 0] },  {y83[22],y83[22],y83[22],y83[22],y83[22],y83[22], y83[22: 0]  }, x193); 

 Register29Bit Reg462 (clk,x193, x193_1 );

 Adder29Bit Adder122(clk,  { x193_1[28: 0] },  {y84[23],y84[23],y84[23],y84[23],y84[23], y84[23: 0]  }, x194); 

 Register29Bit Reg463 (clk,x194, x194_1 );

 Adder29Bit Adder123(clk,  { x194_1[28: 0] },  {y85[22],y85[22],y85[22],y85[22],y85[22],y85[22], y85[22: 0]  }, x195); 

 Register29Bit Reg464 (clk,x195, x195_1 );

 Adder29Bit Adder124(clk,  { x195_1[28: 0] },  {y86[24],y86[24],y86[24],y86[24], y86[24: 0]  }, x196); 

 Register29Bit Reg465 (clk,x196, x196_1 );

 Adder29Bit Adder125(clk,  { x196_1[28: 0] },  {y87[23],y87[23],y87[23],y87[23],y87[23], y87[23: 0]  }, x197); 

 Register29Bit Reg466 (clk,x197, x197_1 );

 Adder29Bit Adder126(clk,  { x197_1[28: 0] },  {y88[24],y88[24],y88[24],y88[24], y88[24: 0]  }, x198); 

 Register29Bit Reg467 (clk,x198, x198_1 );

 Adder29Bit Adder127(clk,  { x198_1[28: 0] },  {y89[22],y89[22],y89[22],y89[22],y89[22],y89[22], y89[22: 0]  }, x199); 

 Register29Bit Reg468 (clk,x199, x199_1 );

 Adder29Bit Adder128(clk,  { x199_1[28: 0] },  {y90[23],y90[23],y90[23],y90[23],y90[23], y90[23: 0]  }, x200); 

 Register29Bit Reg469 (clk,x200, x200_1 );

 Adder29Bit Adder129(clk,  { x200_1[28: 0] },  {y91[23],y91[23],y91[23],y91[23],y91[23], y91[23: 0]  }, x201); 

 Register29Bit Reg470 (clk,x201, x201_1 );

 Adder29Bit Adder130(clk,  { x201_1[28: 0] },  {y92[22],y92[22],y92[22],y92[22],y92[22],y92[22], y92[22: 0]  }, x202); 

 Register29Bit Reg471 (clk,x202, x202_1 );

 Adder29Bit Adder131(clk,  { x202_1[28: 0] },  {y93[23],y93[23],y93[23],y93[23],y93[23], y93[23: 0]  }, x203); 

 Register29Bit Reg472 (clk,x203, x203_1 );

 Adder29Bit Adder132(clk,  { x203_1[28: 0] },  {y94[23],y94[23],y94[23],y94[23],y94[23], y94[23: 0]  }, x204); 

 Register29Bit Reg473 (clk,x204, x204_1 );

 Adder29Bit Adder133(clk,  { x204_1[28: 0] },  {y95[22],y95[22],y95[22],y95[22],y95[22],y95[22], y95[22: 0]  }, x205); 

 Register29Bit Reg474 (clk,x205, x205_1 );

 Adder29Bit Adder134(clk,  { x205_1[28: 0] },  {y96[24],y96[24],y96[24],y96[24], y96[24: 0]  }, x206); 

 Register29Bit Reg475 (clk,x206, x206_1 );

 Adder29Bit Adder135(clk,  { x206_1[28: 0] },  {y97[22],y97[22],y97[22],y97[22],y97[22],y97[22], y97[22: 0]  }, x207); 

 Register29Bit Reg476 (clk,x207, x207_1 );

 Adder29Bit Adder136(clk,  { x207_1[28: 0] },  {y98[23],y98[23],y98[23],y98[23],y98[23], y98[23: 0]  }, x208); 

 Register29Bit Reg477 (clk,x208, x208_1 );

 Adder29Bit Adder137(clk,  { x208_1[28: 0] },  {y99[22],y99[22],y99[22],y99[22],y99[22],y99[22], y99[22: 0]  }, x209); 

 Register29Bit Reg478 (clk,x209, x209_1 );

 Adder29Bit Adder138(clk,  { x209_1[28: 0] },  {y100[22],y100[22],y100[22],y100[22],y100[22],y100[22], y100[22: 0]  }, x210); 

 Register29Bit Reg479 (clk,x210, x210_1 );

 Adder29Bit Adder139(clk,  { x210_1[28: 0] },  {y101[22],y101[22],y101[22],y101[22],y101[22],y101[22], y101[22: 0]  }, x211); 

 Register29Bit Reg480 (clk,x211, x211_1 );

 Adder29Bit Adder140(clk,  { x211_1[28: 0] },  {y102[22],y102[22],y102[22],y102[22],y102[22],y102[22], y102[22: 0]  }, x212); 

 Register29Bit Reg481 (clk,x212, x212_1 );

 Adder29Bit Adder141(clk,  { x212_1[28: 0] },  {y103[22],y103[22],y103[22],y103[22],y103[22],y103[22], y103[22: 0]  }, x213); 

 Register29Bit Reg482 (clk,x213, x213_1 );

 Adder29Bit Adder142(clk,  { x213_1[28: 0] },  {y104[21],y104[21],y104[21],y104[21],y104[21],y104[21],y104[21], y104[21: 0]  }, x214); 

 Register29Bit Reg483 (clk,x214, x214_1 );

 Adder29Bit Adder143(clk,  { x214_1[28: 0] },  {y105[22],y105[22],y105[22],y105[22],y105[22],y105[22], y105[22: 0]  }, x215); 

 Register29Bit Reg484 (clk,x215, x215_1 );

 Adder29Bit Adder144(clk,  { x215_1[28: 0] },  {y106[22],y106[22],y106[22],y106[22],y106[22],y106[22], y106[22: 0]  }, x216); 

 Register29Bit Reg485 (clk,x216, x216_1 );

 Adder29Bit Adder145(clk,  { x216_1[28: 0] },  {y107[22],y107[22],y107[22],y107[22],y107[22],y107[22], y107[22: 0]  }, x217); 

 Register29Bit Reg486 (clk,x217, x217_1 );

 Adder29Bit Adder146(clk,  { x217_1[28: 0] },  {y108[21],y108[21],y108[21],y108[21],y108[21],y108[21],y108[21], y108[21: 0]  }, x218); 

 Register29Bit Reg487 (clk,x218, x218_1 );

 Adder29Bit Adder147(clk,  { x218_1[28: 0] },  {y109[23],y109[23],y109[23],y109[23],y109[23], y109[23: 0]  }, x219); 

 Register29Bit Reg488 (clk,x219, x219_1 );

 Adder29Bit Adder148(clk,  { x219_1[28: 0] },  {y110[22],y110[22],y110[22],y110[22],y110[22],y110[22], y110[22: 0]  }, x220); 

 Register29Bit Reg489 (clk,x220, x220_1 );

 Adder29Bit Adder149(clk,  { x220_1[28: 0] },  {y111[23],y111[23],y111[23],y111[23],y111[23], y111[23: 0]  }, x221); 

 Register29Bit Reg490 (clk,x221, x221_1 );

 Adder29Bit Adder150(clk,  { x221_1[28: 0] },  {y112[23],y112[23],y112[23],y112[23],y112[23], y112[23: 0]  }, x222); 

 Register29Bit Reg491 (clk,x222, x222_1 );

 Adder29Bit Adder151(clk,  { x222_1[28: 0] },  {y113[23],y113[23],y113[23],y113[23],y113[23], y113[23: 0]  }, x223); 

 Register29Bit Reg492 (clk,x223, x223_1 );

 Adder29Bit Adder152(clk,  { x223_1[28: 0] },  {y114[20],y114[20],y114[20],y114[20],y114[20],y114[20],y114[20],y114[20], y114[20: 0]  }, x224); 

 Register29Bit Reg493 (clk,x224, x224_1 );

 Adder29Bit Adder153(clk,  { x224_1[28: 0] },  {y115[21],y115[21],y115[21],y115[21],y115[21],y115[21],y115[21], y115[21: 0]  }, x225); 

 Register29Bit Reg494 (clk,x225, x225_1 );

 Adder29Bit Adder154(clk,  { x225_1[28: 0] },  {y116[21],y116[21],y116[21],y116[21],y116[21],y116[21],y116[21], y116[21: 0]  }, x226); 

 Register29Bit Reg495 (clk,x226, x226_1 );

 Adder29Bit Adder155(clk,  { x226_1[28: 0] },  {y117[21],y117[21],y117[21],y117[21],y117[21],y117[21],y117[21], y117[21: 0]  }, x227); 

 Register29Bit Reg496 (clk,x227, x227_1 );

 Adder29Bit Adder156(clk,  { x227_1[28: 0] },  {y118[20],y118[20],y118[20],y118[20],y118[20],y118[20],y118[20],y118[20], y118[20: 0]  }, x228); 

 Register29Bit Reg497 (clk,x228, x228_1 );

 Adder29Bit Adder157(clk,  { x228_1[28: 0] },  {y119[21],y119[21],y119[21],y119[21],y119[21],y119[21],y119[21], y119[21: 0]  }, x229); 

 Register29Bit Reg498 (clk,x229, x229_1 );

 Adder29Bit Adder158(clk,  { x229_1[28: 0] },  {y120[20],y120[20],y120[20],y120[20],y120[20],y120[20],y120[20],y120[20], y120[20: 0]  }, x230); 

 Register29Bit Reg499 (clk,x230, x230_1 );

 Adder29Bit Adder159(clk,  { x230_1[28: 0] },  {y121[21],y121[21],y121[21],y121[21],y121[21],y121[21],y121[21], y121[21: 0]  }, x231); 

 Register29Bit Reg500 (clk,x231, x231_1 );

 Adder29Bit Adder160(clk,  { x231_1[28: 0] },  {y122[21],y122[21],y122[21],y122[21],y122[21],y122[21],y122[21], y122[21: 0]  }, x232); 

 Register29Bit Reg501 (clk,x232, x232_1 );

 Adder29Bit Adder161(clk,  { x232_1[28: 0] },  {y123[21],y123[21],y123[21],y123[21],y123[21],y123[21],y123[21], y123[21: 0]  }, x233); 

 Register29Bit Reg502 (clk,x233, x233_1 );

 Adder29Bit Adder162(clk,  { x233_1[28: 0] },  {y124[21],y124[21],y124[21],y124[21],y124[21],y124[21],y124[21], y124[21: 0]  }, x234); 

 Register29Bit Reg503 (clk,x234, x234_1 );

 Adder29Bit Adder163(clk,  { x234_1[28: 0] },  {y125[21],y125[21],y125[21],y125[21],y125[21],y125[21],y125[21], y125[21: 0]  }, x235); 

 Register29Bit Reg504 (clk,x235, x235_1 );

 Adder29Bit Adder164(clk,  { x235_1[28: 0] },  {y126[21],y126[21],y126[21],y126[21],y126[21],y126[21],y126[21], y126[21: 0]  }, x236); 

 Register29Bit Reg505 (clk,x236, x236_1 );

 Adder29Bit Adder165(clk,  { x236_1[28: 0] },  {y127[21],y127[21],y127[21],y127[21],y127[21],y127[21],y127[21], y127[21: 0]  }, x237); 

 Register29Bit Reg506 (clk,x237, x237_1 );

 Adder29Bit Adder166(clk,  { x237_1[28: 0] },  {y128[21],y128[21],y128[21],y128[21],y128[21],y128[21],y128[21], y128[21: 0]  }, x238); 

 Register29Bit Reg507 (clk,x238, x238_1 );

 Adder29Bit Adder167(clk,  { x238_1[28: 0] },  {y129[21],y129[21],y129[21],y129[21],y129[21],y129[21],y129[21], y129[21: 0]  }, x239); 

 Register29Bit Reg508 (clk,x239, x239_1 );

 Adder29Bit Adder168(clk,  { x239_1[28: 0] },  {y130[21],y130[21],y130[21],y130[21],y130[21],y130[21],y130[21], y130[21: 0]  }, x240); 

 Register29Bit Reg509 (clk,x240, x240_1 );

 Adder29Bit Adder169(clk,  { x240_1[28: 0] },  {y131[23],y131[23],y131[23],y131[23],y131[23], y131[23: 0]  }, x241); 

 Register29Bit Reg510 (clk,x241, x241_1 );

 Adder29Bit Adder170(clk,  { x241_1[28: 0] },  {y132[22],y132[22],y132[22],y132[22],y132[22],y132[22], y132[22: 0]  }, x242); 

 Register29Bit Reg511 (clk,x242, x242_1 );

 Adder29Bit Adder171(clk,  { x242_1[28: 0] },  {y133[22],y133[22],y133[22],y133[22],y133[22],y133[22], y133[22: 0]  }, x243); 

 Register29Bit Reg512 (clk,x243, x243_1 );

 Adder29Bit Adder172(clk,  { x243_1[28: 0] },  {y134[20],y134[20],y134[20],y134[20],y134[20],y134[20],y134[20],y134[20], y134[20: 0]  }, x244); 

 Register29Bit Reg513 (clk,x244, x244_1 );

 Adder29Bit Adder173(clk,  { x244_1[28: 0] },  {y135[22],y135[22],y135[22],y135[22],y135[22],y135[22], y135[22: 0]  }, x245); 

 Register29Bit Reg514 (clk,x245, x245_1 );

 Adder29Bit Adder174(clk,  { x245_1[28: 0] },  {y136[21],y136[21],y136[21],y136[21],y136[21],y136[21],y136[21], y136[21: 0]  }, x246); 

 Register29Bit Reg515 (clk,x246, x246_1 );

 Adder29Bit Adder175(clk,  { x246_1[28: 0] },  {y137[22],y137[22],y137[22],y137[22],y137[22],y137[22], y137[22: 0]  }, x247); 

 Register29Bit Reg516 (clk,x247, x247_1 );

 Adder29Bit Adder176(clk,  { x247_1[28: 0] },  {y138[22],y138[22],y138[22],y138[22],y138[22],y138[22], y138[22: 0]  }, x248); 

 Register29Bit Reg517 (clk,x248, x248_1 );

 Adder29Bit Adder177(clk,  { x248_1[28: 0] },  {y139[22],y139[22],y139[22],y139[22],y139[22],y139[22], y139[22: 0]  }, x249); 

 Register29Bit Reg518 (clk,x249, x249_1 );

 Adder29Bit Adder178(clk,  { x249_1[28: 0] },  {y140[21],y140[21],y140[21],y140[21],y140[21],y140[21],y140[21], y140[21: 0]  }, x250); 

 Register29Bit Reg519 (clk,x250, x250_1 );

 Adder29Bit Adder179(clk,  { x250_1[28: 0] },  {y141[22],y141[22],y141[22],y141[22],y141[22],y141[22], y141[22: 0]  }, x251); 

 Register29Bit Reg520 (clk,x251, x251_1 );

 Adder29Bit Adder180(clk,  { x251_1[28: 0] },  {y142[24],y142[24],y142[24],y142[24], y142[24: 0]  }, x252); 

 Register29Bit Reg521 (clk,x252, x252_1 );

 Adder29Bit Adder181(clk,  { x252_1[28: 0] },  {y143[21],y143[21],y143[21],y143[21],y143[21],y143[21],y143[21], y143[21: 0]  }, x253); 

 Register29Bit Reg522 (clk,x253, x253_1 );

 Adder29Bit Adder182(clk,  { x253_1[28: 0] },  {y144[23],y144[23],y144[23],y144[23],y144[23], y144[23: 0]  }, x254); 

 Register29Bit Reg523 (clk,x254, x254_1 );

 Adder29Bit Adder183(clk,  { x254_1[28: 0] },  {y145[22],y145[22],y145[22],y145[22],y145[22],y145[22], y145[22: 0]  }, x255); 

 Register29Bit Reg524 (clk,x255, x255_1 );

 Adder29Bit Adder184(clk,  { x255_1[28: 0] },  {y146[24],y146[24],y146[24],y146[24], y146[24: 0]  }, x256); 

 Register29Bit Reg525 (clk,x256, x256_1 );

 Adder29Bit Adder185(clk,  { x256_1[28: 0] },  {y147[24],y147[24],y147[24],y147[24], y147[24: 0]  }, x257); 

 Register29Bit Reg526 (clk,x257, x257_1 );

 Adder29Bit Adder186(clk,  { x257_1[28: 0] },  {y148[24],y148[24],y148[24],y148[24], y148[24: 0]  }, x258); 

 Register29Bit Reg527 (clk,x258, x258_1 );

 Adder29Bit Adder187(clk,  { x258_1[28: 0] },  {y149[24],y149[24],y149[24],y149[24], y149[24: 0]  }, x259); 

 Register29Bit Reg528 (clk,x259, x259_1 );

 Adder29Bit Adder188(clk,  { x259_1[28: 0] },  {y150[20],y150[20],y150[20],y150[20],y150[20],y150[20],y150[20],y150[20], y150[20: 0]  }, Out_Y_wire); 

 endmodule 



module Adder21Bit (clk, In1, In2, AddOut);
 input clk;
 input [20:0] In1, In2; 

 output [21:0] AddOut;

 reg [21 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder22Bit (clk, In1, In2, AddOut);
 input clk;
 input [21:0] In1, In2; 

 output [22:0] AddOut;

 reg [22 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder23Bit (clk, In1, In2, AddOut);
 input clk;
 input [22:0] In1, In2; 

 output [23:0] AddOut;

 reg [23 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder17Bit (clk, In1, In2, AddOut);
 input clk;
 input [16:0] In1, In2; 

 output [17:0] AddOut;

 reg [17 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder18Bit (clk, In1, In2, AddOut);
 input clk;
 input [17:0] In1, In2; 

 output [18:0] AddOut;

 reg [18 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder24Bit (clk, In1, In2, AddOut);
 input clk;
 input [23:0] In1, In2; 

 output [24:0] AddOut;

 reg [24 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder19Bit (clk, In1, In2, AddOut);
 input clk;
 input [18:0] In1, In2; 

 output [19:0] AddOut;

 reg [19 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder20Bit (clk, In1, In2, AddOut);
 input clk;
 input [19:0] In1, In2; 

 output [20:0] AddOut;

 reg [20 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder14Bit (clk, In1, In2, AddOut);
 input clk;
 input [13:0] In1, In2; 

 output [14:0] AddOut;

 reg [14 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder15Bit (clk, In1, In2, AddOut);
 input clk;
 input [14:0] In1, In2; 

 output [15:0] AddOut;

 reg [15 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder25Bit (clk, In1, In2, AddOut);
 input clk;
 input [24:0] In1, In2; 

 output [25:0] AddOut;

 reg [25 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder26Bit (clk, In1, In2, AddOut);
 input clk;
 input [25:0] In1, In2; 

 output [26:0] AddOut;

 reg [26 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder27Bit (clk, In1, In2, AddOut);
 input clk;
 input [26:0] In1, In2; 

 output [27:0] AddOut;

 reg [27 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder28Bit (clk, In1, In2, AddOut);
 input clk;
 input [27:0] In1, In2; 

 output [28:0] AddOut;

 reg [28 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder29Bit (clk, In1, In2, AddOut);
 input clk;
 input [28:0] In1, In2; 

 output [28:0] AddOut;

 reg [28 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule



module Subtractor14Bit (clk, In1, In2, SubOut);
 input clk;
 input [13:0] In1, In2;
 output [14 :0] SubOut;

 reg [14 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule

module Subtractor17Bit (clk, In1, In2, SubOut);
 input clk;
 input [16:0] In1, In2;
 output [17 :0] SubOut;

 reg [17 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule

module Subtractor22Bit (clk, In1, In2, SubOut);
 input clk;
 input [21:0] In1, In2;
 output [22 :0] SubOut;

 reg [22 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule

module Subtractor24Bit (clk, In1, In2, SubOut);
 input clk;
 input [23:0] In1, In2;
 output [24 :0] SubOut;

 reg [24 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule

module Subtractor21Bit (clk, In1, In2, SubOut);
 input clk;
 input [20:0] In1, In2;
 output [21 :0] SubOut;

 reg [21 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule

module Subtractor19Bit (clk, In1, In2, SubOut);
 input clk;
 input [18:0] In1, In2;
 output [19 :0] SubOut;

 reg [19 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule

module Subtractor23Bit (clk, In1, In2, SubOut);
 input clk;
 input [22:0] In1, In2;
 output [23 :0] SubOut;

 reg [23 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule

module Subtractor18Bit (clk, In1, In2, SubOut);
 input clk;
 input [17:0] In1, In2;
 output [18 :0] SubOut;

 reg [18 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule

module Subtractor20Bit (clk, In1, In2, SubOut);
 input clk;
 input [19:0] In1, In2;
 output [20 :0] SubOut;

 reg [20 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule

module Subtractor15Bit (clk, In1, In2, SubOut);
 input clk;
 input [14:0] In1, In2;
 output [15 :0] SubOut;

 reg [15 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule

module Subtractor16Bit (clk, In1, In2, SubOut);
 input clk;
 input [15:0] In1, In2;
 output [16 :0] SubOut;

 reg [16 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule



module Register23Bit (clk, In1, RegOut);
 input clk;
 input [22:0] In1;
 output [22 :0] RegOut;

 reg [22 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register22Bit (clk, In1, RegOut);
 input clk;
 input [21:0] In1;
 output [21 :0] RegOut;

 reg [21 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register24Bit (clk, In1, RegOut);
 input clk;
 input [23:0] In1;
 output [23 :0] RegOut;

 reg [23 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register25Bit (clk, In1, RegOut);
 input clk;
 input [24:0] In1;
 output [24 :0] RegOut;

 reg [24 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register20Bit (clk, In1, RegOut);
 input clk;
 input [19:0] In1;
 output [19 :0] RegOut;

 reg [19 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register19Bit (clk, In1, RegOut);
 input clk;
 input [18:0] In1;
 output [18 :0] RegOut;

 reg [18 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register21Bit (clk, In1, RegOut);
 input clk;
 input [20:0] In1;
 output [20 :0] RegOut;

 reg [20 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register27Bit (clk, In1, RegOut);
 input clk;
 input [26:0] In1;
 output [26 :0] RegOut;

 reg [26 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register28Bit (clk, In1, RegOut);
 input clk;
 input [27:0] In1;
 output [27 :0] RegOut;

 reg [27 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register18Bit (clk, In1, RegOut);
 input clk;
 input [17:0] In1;
 output [17 :0] RegOut;

 reg [17 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register15Bit (clk, In1, RegOut);
 input clk;
 input [14:0] In1;
 output [14 :0] RegOut;

 reg [14 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register12Bit (clk, In1, RegOut);
 input clk;
 input [11:0] In1;
 output [11 :0] RegOut;

 reg [11 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register26Bit (clk, In1, RegOut);
 input clk;
 input [25:0] In1;
 output [25 :0] RegOut;

 reg [25 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register29Bit (clk, In1, RegOut);
 input clk;
 input [28:0] In1;
 output [28 :0] RegOut;

 reg [28 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule



module Negator23Bit (clk, In1, NegOut);
 input clk;
 input [22:0] In1;
 output [22 :0] NegOut;

 reg [22 :0] NegOut; 

always @(posedge clk)
begin
NegOut <= -(In1);
end
endmodule

module Negator24Bit (clk, In1, NegOut);
 input clk;
 input [23:0] In1;
 output [23 :0] NegOut;

 reg [23 :0] NegOut; 

always @(posedge clk)
begin
NegOut <= -(In1);
end
endmodule

module Negator21Bit (clk, In1, NegOut);
 input clk;
 input [20:0] In1;
 output [20 :0] NegOut;

 reg [20 :0] NegOut; 

always @(posedge clk)
begin
NegOut <= -(In1);
end
endmodule

module Negator20Bit (clk, In1, NegOut);
 input clk;
 input [19:0] In1;
 output [19 :0] NegOut;

 reg [19 :0] NegOut; 

always @(posedge clk)
begin
NegOut <= -(In1);
end
endmodule

module Negator22Bit (clk, In1, NegOut);
 input clk;
 input [21:0] In1;
 output [21 :0] NegOut;

 reg [21 :0] NegOut; 

always @(posedge clk)
begin
NegOut <= -(In1);
end
endmodule

module Negator25Bit (clk, In1, NegOut);
 input clk;
 input [24:0] In1;
 output [24 :0] NegOut;

 reg [24 :0] NegOut; 

always @(posedge clk)
begin
NegOut <= -(In1);
end
endmodule

module Negator15Bit (clk, In1, NegOut);
 input clk;
 input [14:0] In1;
 output [14 :0] NegOut;

 reg [14 :0] NegOut; 

always @(posedge clk)
begin
NegOut <= -(In1);
end
endmodule
