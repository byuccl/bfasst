
module chip (input \dd_pad_i[11] , input io_0_3_0, input io_0_3_1, input io_0_4_0, input io_0_4_1, input \wb_sel_i[0] , input wb_stb_i, input io_0_6_0, output io_0_6_1, input arst_i, input io_0_7_1, input \wb_sel_i[3] , output diown_pad_o, output dmarq_pad_i, input \wb_sel_i[1] , input iordy_pad_i, input wb_cyc_i, input DMA_req, input wb_inta_o, input \dd_pad_i[9] , input \dd_pad_i[1] , input \dd_pad_i[14] , input \dd_pad_i[6] , input \dd_pad_i[8] , input \dd_pad_i[13] , input \dd_pad_i[0] , input \dd_pad_i[10] , input \dd_pad_i[15] , input io_33_7_0, input io_31_0_1, output dmackn_pad_o, input io_33_13_0, input \dd_pad_i[3] , input \dd_pad_i[5] , input wb_we_i, input \dd_pad_i[7] , input \wb_dat_i[16] , input \dd_pad_i[2] , input \wb_dat_i[4] , input \wb_dat_i[27] , input wb_clk_i, input \wb_dat_i[30] , input \dd_pad_i[12] , input \wb_dat_i[14] , input \wb_dat_i[18] , input \wb_dat_i[24] , input \wb_dat_i[23] , input \wb_dat_i[17] , input \wb_dat_i[25] , input \wb_dat_i[11] , input \wb_dat_i[20] , input io_33_1_1, output \wb_dat_o[7] , input \wb_dat_i[0] , input \wb_dat_i[21] , input \wb_dat_i[5] , input io_33_5_0, output cs0n_pad_o, input \wb_dat_o[5] , input \wb_dat_i[22] , input \wb_dat_i[19] , input \wb_adr_i[4] , output io_14_33_0, output \dd_pad_o[9] , output \dd_pad_o[11] , output \dd_pad_o[14] , input io_33_9_0, input \wb_dat_i[8] , input io_33_16_1, input io_33_14_0, output \da_pad_o[1] , output \dd_pad_o[2] , output \dd_pad_o[8] , output \wb_dat_i[12] , output \dd_pad_o[5] , input io_33_17_0, output \da_pad_o[2] , input io_33_8_0, output io_33_23_0, input io_33_15_1, input io_33_19_0, output \dd_pad_o[3] , output \dd_pad_o[13] , output \dd_pad_o[12] , output io_27_33_1, input \wb_adr_i[5] , output io_18_33_0, output wb_rty_o, output \wb_dat_o[30] , output \wb_dat_i[1] , output dd_padoe_o, output \dd_pad_o[6] , output \wb_dat_i[29] , output resetn_pad_o, output io_33_21_0, output \wb_dat_o[21] , output \wb_dat_o[19] , input \wb_adr_i[3] , output \wb_dat_o[8] , output \wb_dat_o[18] , output \wb_dat_o[28] , output \dd_pad_o[15] , input \wb_dat_i[2] , output \wb_dat_o[24] , output \wb_dat_o[6] , output io_21_33_0, output \wb_dat_o[15] , output \wb_dat_o[0] , output \wb_dat_o[3] , output io_33_28_0, output diorn_pad_o, output io_33_30_0, output \wb_dat_o[16] , output \dd_pad_o[0] , output cs1n_pad_o, output \wb_dat_o[29] , output \wb_dat_o[23] , output io_33_24_0, output \wb_dat_i[3] , output \wb_dat_o[9] , output \wb_dat_o[25] , output \wb_dat_o[27] , output \wb_dat_o[1] , output \wb_dat_i[28] , output \wb_dat_o[31] , output \wb_dat_o[11] , output \wb_dat_o[4] , output io_33_27_0, output \wb_dat_o[26] , output wb_err_o, input \dd_pad_i[4] , input \wb_dat_o[20] , input wb_ack_o, input \da_pad_o[0] , input \wb_dat_i[31] , input DMA_Ack, input \dd_pad_o[4] , input wb_rst_i, input \wb_dat_i[13] , input \wb_dat_i[10] , input \wb_dat_o[10] , input \wb_dat_i[7] , input \dd_pad_o[7] , input \wb_dat_i[9] , input intrq_pad_i, input \wb_dat_o[13] , input \wb_adr_i[6] , input \wb_adr_i[2] , input \wb_sel_i[2] , input \wb_dat_o[22] , input \wb_dat_i[26] , input \dd_pad_o[1] , input \wb_dat_i[6] , input \wb_dat_o[2] , input \wb_dat_o[17] , input \wb_dat_o[14] , input \wb_dat_i[15] , input \dd_pad_o[10] , input \wb_dat_o[12] );

wire n1, n2, \dd_pad_i[11] , n4, n5, n6, io_0_3_0, io_0_3_1, io_0_4_0, io_0_4_1;
wire \wb_sel_i[0] , wb_stb_i, io_0_6_0, arst_i, io_0_7_1, n17, \wb_sel_i[3] , \wb_sel_i[1] , iordy_pad_i, wb_cyc_i;
wire DMA_req, wb_inta_o, \dd_pad_i[9] , \dd_pad_i[1] , \dd_pad_i[14] , \dd_pad_i[6] , \dd_pad_i[8] , n33, n34, n35;
wire n36, n37, n38, n39, n44, \dd_pad_i[13] , \dd_pad_i[0] , n53, n54, n62;
wire \dd_pad_i[10] , \dd_pad_i[15] , n65, n67, n68, n70, n71, io_33_7_0, n73, io_31_0_1;
wire n77, n79, io_33_13_0, \dd_pad_i[3] , \dd_pad_i[5] , n83, wb_we_i, \dd_pad_i[7] , n96, \wb_dat_i[16] ;
wire \dd_pad_i[2] , n104, \wb_dat_i[4] , n112, n113, \wb_dat_i[27] , wb_clk_i, n118, \wb_dat_i[30] , \dd_pad_i[12] ;
wire \wb_dat_i[14] , \wb_dat_i[18] , n130, \wb_dat_i[24] , \wb_dat_i[23] , n134, n136, \wb_dat_i[17] , \wb_dat_i[25] , \wb_dat_i[11] ;
wire \wb_dat_i[20] , io_33_1_1, \wb_dat_o[7] , n144, n145, n146, n147, n148, n149, n150;
wire n153, n156, n157, n158, n159, n160, n161, n162, n163, n165;
wire \wb_dat_i[0] , n170, n171, n172, n175, \wb_dat_i[21] , \wb_dat_i[5] , n183, n186, n187;
wire n188, n189, n190, n191, n192, n194, io_33_5_0, n205, n211, n212;
wire n213, n214, n215, n216, n217, n219, \wb_dat_o[5] , n227, \wb_dat_i[22] , \wb_dat_i[19] ;
wire n237, n247, n248, n249, n250, n251, n252, n253, n254, n255;
wire n256, n257, n259, n260, n265, n275, n276, n277, n278, n279;
wire n281, n282, n283, n284, n286, n289, n290, n291, n292, n293;
wire n294, n295, n296, n297, n298, n299, n300, \wb_adr_i[4] , n307, n312;
wire n318, n321, n322, n323, n324, n325, n326, n327, n329, n331;
wire n345, n346, n349, n350, n351, io_33_9_0, n356, n358, n359, n361;
wire n362, n367, n368, n369, n370, n371, n372, n373, n374, \wb_dat_i[8] ;
wire n379, n389, n390, n393, n394, n395, n396, n397, n403, n404;
wire n405, n406, n409, n410, n411, n412, n413, n424, io_33_16_1, n429;
wire io_33_14_0, n437, n438, n441, n448, n450, n451, n458, n459, n460;
wire n461, io_33_17_0, n465, n466, n467, n468, n470, n471, n477, n478;
wire n479, n480, n481, n482, n484, n485, n486, n487, n488, n489;
wire n490, n491, n492, n493, n494, n495, n496, n497, n499, n500;
wire n501, n502, io_33_8_0, n506, n512, n513, n516, n517, io_33_23_0, io_33_15_1;
wire io_33_19_0, n549, n550, n552, n555, n556, n557, n558, n561, n562;
wire n563, n564, n565, n566, n577, n578, n586, n588, n589, n590;
wire n591, n592, n594, n595, n596, n597, n598, \wb_adr_i[5] , n604, n605;
wire n606, io_18_33_0, wb_rty_o, n609, n613, \wb_dat_i[1] , n616, n628, n629, n630;
wire n631, n632, n638, n644, n649, n652, n653, n654, n655, n656;
wire n660, n663, n667, n668, n669, n670, n671, n672, n673, n674;
wire n680, n682, n684, n694, n695, n696, n701, n704, n705, n708;
wire n711, n712, n714, n716, n717, n718, n721, n722, n723, n724;
wire n727, n730, n732, n733, n738, n739, n740, n741, n742, n743;
wire n744, n745, n746, n748, n751, n752, n753, n754, n756, n758;
wire n759, n760, io_33_21_0, n762, n763, n765, n766, n767, n768, n770;
wire \wb_dat_o[21] , \wb_dat_o[19] , n777, n778, n785, n786, n787, n792, n794, n798;
wire \wb_adr_i[3] , n807, n808, n809, \wb_dat_o[8] , n811, n812, n816, n817, n818;
wire n820, n821, \wb_dat_o[18] , n824, n825, n832, n834, n836, n837, n840;
wire n841, n864, n867, n870, \dd_pad_o[15] , n876, \wb_dat_i[2] , n882, n884, n888;
wire n892, n893, n894, n895, n896, n898, n899, n909, n911, n913;
wire n917, n922, n923, n924, n927, n929, \wb_dat_o[15] , n932, n934, n935;
wire n936, n939, n956, n957, n958, n980, n983, n985, n988, n989;
wire n999, n1000, n1002, n1003, n1008, n1009, n1010, n1014, n1015, n1016;
wire n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1030, n1031, n1032;
wire n1033, n1034, n1035, n1036, n1047, n1048, n1049, n1050, n1051, n1052;
wire n1054, n1055, n1057, n1058, n1059, n1062, n1065, n1074, n1086, n1087;
wire n1104, n1106, n1107, n1116, n1117, n1118, n1122, n1123, n1124, n1131;
wire n1132, n1133, n1140, n1141, \wb_dat_o[0] , n1144, n1145, n1146, n1147, n1149;
wire n1150, n1151, n1152, n1154, n1155, n1156, n1157, n1158, n1159, n1160;
wire n1161, n1162, n1163, n1165, n1166, n1172, n1173, n1174, n1175, n1176;
wire n1178, n1192, n1193, n1195, n1199, n1203, n1204, n1207, n1211, n1212;
wire n1213, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224;
wire n1225, n1226, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1238;
wire n1239, n1240, n1241, n1243, n1244, n1250, n1251, n1261, n1262, n1263;
wire n1266, n1267, n1268, n1270, n1271, n1272, n1273, n1276, n1277, n1278;
wire n1279, n1281, n1282, n1283, n1284, n1285, n1286, \wb_dat_o[3] , n1289, n1291;
wire n1292, n1293, n1296, n1301, n1302, n1303, n1306, n1309, io_33_28_0, n1312;
wire n1313, n1316, n1317, n1318, n1319, n1320, n1322, n1324, n1325, n1326;
wire n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336;
wire n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, diorn_pad_o;
wire n1348, n1349, io_33_30_0, n1352, n1353, n1354, n1356, n1357, \wb_dat_o[16] , n1360;
wire n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1373, n1374;
wire n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1384, n1387;
wire \dd_pad_o[0] , n1390, n1391, n1392, n1393, cs1n_pad_o, n1397, n1398, n1399, n1401;
wire n1402, n1403, n1405, n1406, n1407, n1408, n1409, \wb_dat_o[29] , n1411, n1412;
wire n1413, n1415, n1417, n1418, n1419, n1420, n1426, \wb_dat_o[23] , n1429, n1430;
wire n1431, n1432, n1433, n1434, n1435, io_33_24_0, n1438, n1439, \wb_dat_i[3] , n1441;
wire n1442, n1443, n1444, n1446, n1447, n1448, n1449, n1450, \wb_dat_o[9] , n1452;
wire n1453, \wb_dat_o[25] , n1456, \wb_dat_o[27] , n1458, \wb_dat_o[1] , n1460, n1462, n1463, \wb_dat_i[28] ;
wire n1466, n1468, n1470, n1471, n1473, n1474, n1475, n1476, n1477, n1479;
wire n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489;
wire n1490, n1491, n1492, n1493, n1494, n1495, \wb_dat_o[31] , n1498, n1499, \wb_dat_o[11] ;
wire \wb_dat_o[4] , n1502, n1503, n1504, n1505, io_33_27_0, n1507, n1508, n1509, n1511;
wire n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521;
wire n1522, n1523, \wb_dat_o[26] , wb_err_o, n1526, n1527, n1528, n1529, n1530, n1531;
wire n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541;
wire n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551;
wire n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561;
wire n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571;
wire n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581;
wire n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591;
wire n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601;
wire n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611;
wire n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621;
wire n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631;
wire n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641;
wire n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651;
wire n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661;
wire n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671;
wire n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681;
wire n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691;
wire n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701;
wire n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711;
wire n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721;
wire n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731;
wire n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741;
wire n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751;
wire n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761;
wire n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771;
wire n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781;
wire n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791;
wire n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801;
wire n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811;
wire n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821;
wire n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831;
wire n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841;
wire n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851;
wire n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861;
wire n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871;
wire n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881;
wire n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891;
wire n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901;
wire n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911;
wire n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921;
wire n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931;
wire n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941;
wire n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951;
wire n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961;
wire n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971;
wire n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981;
wire n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991;
wire n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001;
wire n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011;
wire n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021;
wire n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031;
wire n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041;
wire n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051;
wire n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061;
wire n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071;
wire n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081;
wire n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091;
wire n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101;
wire n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111;
wire n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121;
wire n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131;
wire n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141;
wire n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151;
wire n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161;
wire n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171;
wire n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181;
wire n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191;
wire n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201;
wire n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211;
wire n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221;
wire n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231;
wire n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241;
wire n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251;
wire n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261;
wire n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271;
wire n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281;
wire n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291;
wire n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301;
wire n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311;
wire n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321;
wire n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331;
wire n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341;
wire n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351;
wire n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361;
wire n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371;
wire n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381;
wire n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391;
wire n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401;
wire n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411;
wire n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421;
wire n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431;
wire n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441;
wire n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451;
wire n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461;
wire n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471;
wire n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481;
wire n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491;
wire n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501;
wire n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511;
wire n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521;
wire n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531;
wire n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541;
wire n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551;
wire n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561;
wire n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571;
wire n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581;
wire n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591;
wire n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601;
wire n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611;
wire n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621;
wire n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631;
wire n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641;
wire n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651;
wire n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661;
wire n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671;
wire n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681;
wire n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691;
wire n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701;
wire n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711;
wire n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721;
wire n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731;
wire n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741;
wire n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751;
wire n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761;
wire n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771;
wire n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781;
wire n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791;
wire n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801;
wire n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811;
wire n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821;
wire n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831;
wire n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841;
wire n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851;
wire n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861;
wire n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871;
wire n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881;
wire n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891;
wire n2892, n2893, n2894, n2895;
reg io_0_6_1 = 0, diown_pad_o = 0, dmarq_pad_i = 0, n24 = 0, n31 = 0, n40 = 0, n41 = 0, n42 = 0, n43 = 0, n45 = 0;
reg n48 = 0, n49 = 0, n50 = 0, n51 = 0, n52 = 0, n55 = 0, n56 = 0, n57 = 0, n58 = 0, n59 = 0;
reg n60 = 0, n61 = 0, n66 = 0, n69 = 0, n75 = 0, dmackn_pad_o = 0, n78 = 0, n84 = 0, n85 = 0, n86 = 0;
reg n89 = 0, n90 = 0, n91 = 0, n92 = 0, n93 = 0, n94 = 0, n95 = 0, n97 = 0, n100 = 0, n101 = 0;
reg n102 = 0, n103 = 0, n105 = 0, n106 = 0, n107 = 0, n109 = 0, n110 = 0, n111 = 0, n114 = 0, n115 = 0;
reg n119 = 0, n122 = 0, n123 = 0, n124 = 0, n125 = 0, n126 = 0, n129 = 0, n131 = 0, n135 = 0, n141 = 0;
reg n151 = 0, n152 = 0, n154 = 0, n155 = 0, n164 = 0, n166 = 0, n168 = 0, n169 = 0, n173 = 0, n174 = 0;
reg n176 = 0, n177 = 0, n180 = 0, n181 = 0, n182 = 0, n184 = 0, n185 = 0, n193 = 0, n195 = 0, n196 = 0;
reg n197 = 0, n198 = 0, n199 = 0, n200 = 0, n202 = 0, n203 = 0, n204 = 0, n206 = 0, n207 = 0, n208 = 0;
reg n209 = 0, n210 = 0, cs0n_pad_o = 0, n220 = 0, n221 = 0, n222 = 0, n223 = 0, n224 = 0, n225 = 0, n228 = 0;
reg n229 = 0, n230 = 0, n231 = 0, n232 = 0, n233 = 0, n234 = 0, n238 = 0, n239 = 0, n240 = 0, n241 = 0;
reg n242 = 0, n243 = 0, n244 = 0, n245 = 0, n246 = 0, n258 = 0, n261 = 0, n262 = 0, n263 = 0, n264 = 0;
reg n266 = 0, n267 = 0, n268 = 0, n269 = 0, n270 = 0, n271 = 0, n272 = 0, n273 = 0, n274 = 0, n280 = 0;
reg n285 = 0, n287 = 0, n288 = 0, n301 = 0, n302 = 0, n303 = 0, n305 = 0, io_14_33_0 = 0, n308 = 0, n309 = 0;
reg n310 = 0, n311 = 0, n313 = 0, n314 = 0, n315 = 0, n316 = 0, n317 = 0, n319 = 0, n320 = 0, n328 = 0;
reg n330 = 0, n332 = 0, n333 = 0, n334 = 0, n335 = 0, \dd_pad_o[9]  = 0, n337 = 0, n338 = 0, \dd_pad_o[11]  = 0, \dd_pad_o[14]  = 0;
reg n341 = 0, n342 = 0, n343 = 0, n344 = 0, n347 = 0, n348 = 0, n352 = 0, n353 = 0, n355 = 0, n357 = 0;
reg n360 = 0, n363 = 0, n364 = 0, n365 = 0, n366 = 0, n376 = 0, n377 = 0, n378 = 0, n380 = 0, n381 = 0;
reg n382 = 0, n383 = 0, n384 = 0, n385 = 0, n386 = 0, n387 = 0, n388 = 0, n391 = 0, n392 = 0, n398 = 0;
reg n399 = 0, n400 = 0, n401 = 0, n402 = 0, n407 = 0, n408 = 0, n414 = 0, n415 = 0, n416 = 0, n417 = 0;
reg n418 = 0, n419 = 0, n420 = 0, n421 = 0, n422 = 0, n423 = 0, n425 = 0, n427 = 0, n428 = 0, n430 = 0;
reg n431 = 0, n432 = 0, n433 = 0, n434 = 0, \da_pad_o[1]  = 0, \dd_pad_o[2]  = 0, n440 = 0, n442 = 0, \dd_pad_o[8]  = 0, \wb_dat_i[12]  = 0;
reg \dd_pad_o[5]  = 0, n446 = 0, n447 = 0, n449 = 0, n452 = 0, n453 = 0, n454 = 0, n455 = 0, n456 = 0, n457 = 0;
reg n462 = 0, n464 = 0, \da_pad_o[2]  = 0, n472 = 0, n473 = 0, n474 = 0, n475 = 0, n476 = 0, n483 = 0, n498 = 0;
reg n504 = 0, n505 = 0, n507 = 0, n508 = 0, n509 = 0, n510 = 0, n511 = 0, n514 = 0, n515 = 0, n518 = 0;
reg n519 = 0, n520 = 0, n521 = 0, n522 = 0, n523 = 0, n525 = 0, n526 = 0, n529 = 0, n530 = 0, n531 = 0;
reg n532 = 0, n533 = 0, n534 = 0, n535 = 0, n536 = 0, n537 = 0, n538 = 0, n539 = 0, n540 = 0, n541 = 0;
reg n542 = 0, n543 = 0, n544 = 0, n545 = 0, n546 = 0, n547 = 0, n548 = 0, \dd_pad_o[3]  = 0, n553 = 0, \dd_pad_o[13]  = 0;
reg \dd_pad_o[12]  = 0, n560 = 0, n567 = 0, n568 = 0, n569 = 0, n570 = 0, n571 = 0, n572 = 0, n573 = 0, n574 = 0;
reg n575 = 0, n576 = 0, n579 = 0, n580 = 0, n581 = 0, n582 = 0, n583 = 0, n584 = 0, n585 = 0, n587 = 0;
reg io_27_33_1 = 0, n599 = 0, n600 = 0, n601 = 0, n603 = 0, n610 = 0, n611 = 0, n612 = 0, \wb_dat_o[30]  = 0, dd_padoe_o = 0;
reg n618 = 0, n619 = 0, n620 = 0, n621 = 0, n622 = 0, n623 = 0, n624 = 0, n625 = 0, n626 = 0, n627 = 0;
reg n633 = 0, n634 = 0, n635 = 0, n636 = 0, n637 = 0, n639 = 0, n640 = 0, n641 = 0, n642 = 0, n643 = 0;
reg n645 = 0, n646 = 0, n647 = 0, n648 = 0, n650 = 0, n651 = 0, n657 = 0, n658 = 0, n659 = 0, \dd_pad_o[6]  = 0;
reg n662 = 0, n664 = 0, n665 = 0, n666 = 0, n675 = 0, n676 = 0, n677 = 0, n678 = 0, n679 = 0, n681 = 0;
reg n683 = 0, n685 = 0, n686 = 0, n687 = 0, n688 = 0, n689 = 0, \wb_dat_i[29]  = 0, n691 = 0, n692 = 0, n693 = 0;
reg n697 = 0, n698 = 0, n699 = 0, n700 = 0, resetn_pad_o = 0, n703 = 0, n706 = 0, n707 = 0, n709 = 0, n710 = 0;
reg n713 = 0, n715 = 0, n719 = 0, n720 = 0, n725 = 0, n726 = 0, n728 = 0, n729 = 0, n731 = 0, n734 = 0;
reg n735 = 0, n736 = 0, n737 = 0, n747 = 0, n749 = 0, n750 = 0, n755 = 0, n757 = 0, n764 = 0, n769 = 0;
reg n772 = 0, n773 = 0, n774 = 0, n775 = 0, n779 = 0, n780 = 0, n781 = 0, n782 = 0, n783 = 0, n784 = 0;
reg n788 = 0, n789 = 0, n790 = 0, n791 = 0, n793 = 0, n795 = 0, n796 = 0, n797 = 0, n799 = 0, n800 = 0;
reg n801 = 0, n802 = 0, n803 = 0, n804 = 0, n805 = 0, n813 = 0, n814 = 0, n815 = 0, n819 = 0, \wb_dat_o[28]  = 0;
reg n826 = 0, n827 = 0, n828 = 0, n829 = 0, n830 = 0, n831 = 0, n833 = 0, n835 = 0, n838 = 0, n839 = 0;
reg n842 = 0, n843 = 0, n844 = 0, n845 = 0, n846 = 0, n847 = 0, n848 = 0, n849 = 0, n850 = 0, n851 = 0;
reg n852 = 0, n853 = 0, n854 = 0, n855 = 0, n856 = 0, n857 = 0, n858 = 0, n859 = 0, n860 = 0, n861 = 0;
reg n862 = 0, n863 = 0, n865 = 0, n866 = 0, n868 = 0, n869 = 0, n871 = 0, n872 = 0, n873 = 0, n874 = 0;
reg n877 = 0, n879 = 0, n880 = 0, n881 = 0, n883 = 0, n885 = 0, n886 = 0, n887 = 0, n889 = 0, n890 = 0;
reg n891 = 0, n897 = 0, n900 = 0, n901 = 0, n902 = 0, n903 = 0, n904 = 0, n905 = 0, n906 = 0, n907 = 0;
reg n908 = 0, \wb_dat_o[24]  = 0, \wb_dat_o[6]  = 0, io_21_33_0 = 0, n915 = 0, n916 = 0, n918 = 0, n919 = 0, n920 = 0, n921 = 0;
reg n925 = 0, n926 = 0, n928 = 0, n931 = 0, n933 = 0, n937 = 0, n938 = 0, n940 = 0, n941 = 0, n942 = 0;
reg n943 = 0, n944 = 0, n945 = 0, n946 = 0, n947 = 0, n948 = 0, n949 = 0, n950 = 0, n951 = 0, n952 = 0;
reg n953 = 0, n954 = 0, n955 = 0, n959 = 0, n960 = 0, n961 = 0, n962 = 0, n963 = 0, n964 = 0, n965 = 0;
reg n966 = 0, n967 = 0, n968 = 0, n969 = 0, n970 = 0, n971 = 0, n972 = 0, n973 = 0, n974 = 0, n975 = 0;
reg n976 = 0, n977 = 0, n978 = 0, n979 = 0, n981 = 0, n982 = 0, n984 = 0, n986 = 0, n987 = 0, n990 = 0;
reg n991 = 0, n992 = 0, n993 = 0, n994 = 0, n995 = 0, n996 = 0, n997 = 0, n998 = 0, n1001 = 0, n1004 = 0;
reg n1005 = 0, n1006 = 0, n1007 = 0, n1011 = 0, n1012 = 0, n1013 = 0, n1017 = 0, n1018 = 0, n1026 = 0, n1027 = 0;
reg n1028 = 0, n1029 = 0, n1037 = 0, n1038 = 0, n1039 = 0, n1040 = 0, n1041 = 0, n1042 = 0, n1043 = 0, n1044 = 0;
reg n1045 = 0, n1046 = 0, n1053 = 0, n1056 = 0, n1060 = 0, n1061 = 0, n1063 = 0, n1064 = 0, n1066 = 0, n1067 = 0;
reg n1068 = 0, n1069 = 0, n1070 = 0, n1071 = 0, n1072 = 0, n1073 = 0, n1075 = 0, n1076 = 0, n1077 = 0, n1078 = 0;
reg n1079 = 0, n1080 = 0, n1081 = 0, n1082 = 0, n1083 = 0, n1084 = 0, n1085 = 0, n1088 = 0, n1089 = 0, n1090 = 0;
reg n1091 = 0, n1092 = 0, n1093 = 0, n1094 = 0, n1095 = 0, n1096 = 0, n1097 = 0, n1098 = 0, n1099 = 0, n1100 = 0;
reg n1101 = 0, n1102 = 0, n1103 = 0, n1105 = 0, n1108 = 0, n1109 = 0, n1110 = 0, n1111 = 0, n1112 = 0, n1113 = 0;
reg n1114 = 0, n1115 = 0, n1119 = 0, n1120 = 0, n1121 = 0, n1125 = 0, n1126 = 0, n1127 = 0, n1128 = 0, n1129 = 0;
reg n1130 = 0, n1134 = 0, n1135 = 0, n1136 = 0, n1137 = 0, n1138 = 0, n1139 = 0, n1143 = 0, n1148 = 0, n1153 = 0;
reg n1164 = 0, n1167 = 0, n1168 = 0, n1169 = 0, n1170 = 0, n1171 = 0, n1177 = 0, n1179 = 0, n1180 = 0, n1181 = 0;
reg n1182 = 0, n1183 = 0, n1184 = 0, n1185 = 0, n1186 = 0, n1187 = 0, n1188 = 0, n1189 = 0, n1190 = 0, n1191 = 0;
reg n1194 = 0, n1196 = 0, n1197 = 0, n1198 = 0, n1200 = 0, n1201 = 0, n1202 = 0, n1205 = 0, n1206 = 0, n1208 = 0;
reg n1209 = 0, n1210 = 0, n1214 = 0, n1215 = 0, n1227 = 0, n1228 = 0, n1236 = 0, n1237 = 0, n1242 = 0, n1245 = 0;
reg n1246 = 0, n1247 = 0, n1248 = 0, n1249 = 0, n1252 = 0, n1253 = 0, n1254 = 0, n1255 = 0, n1256 = 0, n1257 = 0;
reg n1258 = 0, n1259 = 0, n1260 = 0, n1264 = 0, n1265 = 0, n1269 = 0, n1274 = 0, n1275 = 0, n1280 = 0, n1288 = 0;
reg n1290 = 0, n1294 = 0, n1295 = 0, n1297 = 0, n1298 = 0, n1299 = 0, n1300 = 0, n1304 = 0, n1305 = 0, n1307 = 0;
reg n1308 = 0, n1310 = 0, n1314 = 0, n1315 = 0, n1321 = 0, n1323 = 0, n1347 = 0, n1351 = 0, n1355 = 0, n1359 = 0;
reg n1369 = 0, n1370 = 0, n1371 = 0, n1372 = 0, n1383 = 0, n1385 = 0, n1386 = 0, n1388 = 0, n1394 = 0, n1395 = 0;
reg n1400 = 0, n1404 = 0, n1414 = 0, n1416 = 0, n1421 = 0, n1422 = 0, n1423 = 0, n1424 = 0, n1425 = 0, n1428 = 0;
reg n1437 = 0, n1445 = 0, n1455 = 0, n1461 = 0, n1465 = 0, n1467 = 0, n1469 = 0, n1472 = 0, n1478 = 0, n1497 = 0;
reg n1510 = 0;
assign n1547 = 1;
assign n1556 = 1;
assign n2277 = 1;
assign n2319 = 1;
assign n2542 = 1;
assign n2713 = 1;
assign n2823 = 1;

assign n1546 = /* LUT    2 24  0 */ 1'b0;
assign n1555 = /* LUT    7 17  0 */ 1'b0;
assign n186  = /* LUT    1 20  3 */ 1'b1;
assign n2276 = /* LUT    4 20  0 */ 1'b0;
assign n2318 = /* LUT    1 18  0 */ 1'b0;
assign n2541 = /* LUT   12 18  0 */ 1'b0;
assign n2712 = /* LUT    2 21  0 */ 1'b0;
assign n2822 = /* LUT    2 17  0 */ 1'b0;
assign n1527 = /* LUT    4 25  6 */ io_33_14_0;
assign n1528 = /* LUT    4 22  7 */ (n502 ? (n514 ? n84 : 1'b0) : 1'b1);
assign n1529 = /* LUT    9 25  2 */ (n827 ? (n828 ? 1'b1 : n130) : (n828 ? !n130 : 1'b0));
assign n1530 = /* LUT   13 27  1 */ (n130 ? n769 : n968);
assign n1160 = /* LUT   11 23  0 */ (n677 ? n1075 : n1159);
assign n1443 = /* LUT   16 19  4 */ (n708 ? n689 : 1'b0);
assign n1533 = /* LUT   10 21  3 */ (n815 ? !n1048 : (n1048 ? 1'b0 : !n798));
assign n1534 = /* LUT    2 20  7 */ (n173 ? !io_33_1_1 : 1'b0);
assign n1535 = /* LUT   20 23  7 */ (n107 ? (n1462 ? 1'b1 : (n701 ? 1'b1 : n1392)) : (n1462 ? 1'b1 : n1392));
assign n1536 = /* LUT   12 27  5 */ (n130 ? n779 : n964);
assign n1537 = /* LUT   15 28  5 */ (n1275 ? (n862 ? 1'b1 : !n666) : (n862 ? n666 : 1'b0));
assign n1538 = /* LUT   13 31  6 */ (n666 ? n1257 : n1246);
assign n1539 = /* LUT   12 22  5 */ (n100 ? (n1239 ? (n286 ? 1'b1 : \wb_adr_i[5] ) : \wb_adr_i[5] ) : (n1239 ? n286 : 1'b0));
assign n1540 = /* LUT    1 22  3 */ (\dd_pad_i[12]  ? !io_33_1_1 : 1'b0);
assign n1541 = /* LUT    4 24  1 */ (n118 ? 1'b0 : io_33_17_0);
assign n1542 = /* LUT    4 21  6 */ (n384 ? 1'b1 : (n385 ? 1'b1 : n391));
assign n957  = /* LUT    9 26  3 */ (n130 ? (n541 ? 1'b0 : !n376) : (n541 ? (n376 ? !n432 : 1'b0) : (n376 ? !n432 : 1'b1)));
assign n1544 = /* LUT   13 28  0 */ (n1102 ? (n851 ? 1'b1 : !n666) : (n851 ? n666 : 1'b0));
assign n1548 = /* LUT   11 20  1 */ (n1139 ? (n1037 ? 1'b0 : n893) : (n892 ? 1'b1 : (n1037 ? 1'b0 : n893)));
assign n1549 = /* LUT   16 18  7 */ (io_33_16_1 ? 1'b1 : io_33_1_1);
assign n1030 = /* LUT   10 20  0 */ (n893 ? (n892 ? (n906 ? !n907 : 1'b1) : !n907) : (n892 ? !n906 : 1'b0));
assign n393  = /* LUT    3 21  4 */ (n379 ? 1'b1 : (n202 ? (n79 ? 1'b1 : n182) : 1'b1));
assign n1551 = /* LUT    2 23  6 */ (n215 ? (io_33_1_1 ? !n205 : (n205 ? n110 : 1'b1)) : (io_33_1_1 ? 1'b0 : (n205 ? n110 : 1'b0)));
assign n1552 = /* LUT   12 26  6 */ (n1181 ? (n856 ? 1'b1 : !n666) : (n856 ? n666 : 1'b0));
assign n1553 = /* LUT   17 21  5 */ (n1480 ? 1'b1 : (n1491 ? 1'b1 : (n1449 ? 1'b1 : n1262)));
assign n1557 = /* LUT    9 22  6 */ wb_inta_o;
assign n1558 = /* LUT    7 28  7 */ (n729 ? (n774 ? 1'b1 : !n666) : (n774 ? n666 : 1'b0));
assign n1559 = /* LUT   14 26  2 */ (n130 ? \wb_sel_i[1]  : wb_cyc_i);
assign n1560 = /* LUT   12 21  4 */ (io_33_1_1 ? 1'b0 : \wb_dat_i[24] );
assign n1326 = /* LUT   13 29  3 */ (n666 ? n232 : n1198);
assign n1562 = /* LUT    3 17  1 */ (n144 ? (io_33_1_1 ? 1'b1 : (n43 ? 1'b1 : !n254)) : (io_33_1_1 ? n254 : (n43 ? n254 : 1'b0)));
assign n1563 = /* LUT   14 25  4 */ (n677 ? n980 : n1062);
assign n1564 = /* LUT    6 21  2 */ (n483 ? 1'b1 : n319);
assign n1565 = /* LUT   11 21  6 */ (n897 ? (n692 ? (n104 ? 1'b1 : n96) : n104) : (n692 ? n96 : 1'b0));
assign n1566 = /* LUT    5 19  3 */ (n471 ? (n589 ? (n180 ? !io_33_1_1 : 1'b0) : !io_33_1_1) : (n589 ? 1'b0 : !io_33_1_1));
assign n1567 = /* LUT   10 23  1 */ (n720 ? (n764 ? 1'b1 : !n130) : (n764 ? n130 : 1'b0));
assign n1568 = /* LUT   15 26  6 */ (n1342 ? 1'b0 : (n1420 ? 1'b0 : (n817 ? 1'b0 : !n1418)));
assign n1569 = /* LUT   15 17  7 */ (io_33_1_1 ? 1'b0 : io_33_13_0);
assign n1570 = /* LUT    7 21  5 */ (io_33_1_1 ? 1'b0 : io_33_16_1);
assign n1571 = /* LUT    3 18  5 */ (n357 ? 1'b1 : (n261 ? 1'b1 : n52));
assign n1572 = /* LUT   12 25  7 */ (n826 ? (n122 ? 1'b1 : n666) : (n122 ? !n666 : 1'b0));
assign n1573 = /* LUT    1 19  1 */ wb_we_i;
assign n1574 = /* LUT   10 25  0 */ (n845 ? (n944 ? 1'b1 : n666) : (n944 ? !n666 : 1'b0));
assign n1575 = /* LUT    4 19  7 */ (n466 ? (n482 ? (n288 ? !io_33_1_1 : 1'b0) : !io_33_1_1) : (n482 ? 1'b0 : !io_33_1_1));
assign n1576 = /* LUT    7 22  1 */ (io_33_1_1 ? 1'b0 : !n706);
assign n1577 = /* LUT    9 23  1 */ (n675 ? (n821 ? 1'b0 : \wb_adr_i[3] ) : (n934 ? 1'b0 : \wb_adr_i[3] ));
assign n1578 = /* LUT   12 15  2 */ (io_33_7_0 ? !\wb_dat_i[2]  : 1'b0);
assign n1579 = /* LUT   14 21  3 */ (\wb_dat_i[18]  ? !io_33_1_1 : 1'b0);
assign n1580 = /* LUT    6 26  0 */ (n130 ? (n419 ? !n628 : (n628 ? 1'b0 : !n376)) : !n628);
assign n1581 = /* LUT   11 17  3 */ (n1003 ? 1'b0 : (n798 ? n993 : 1'b1));
assign n1582 = /* LUT   15 21  4 */ (n916 ? (n919 ? 1'b0 : n1338) : (n919 ? n1285 : (n1285 ? 1'b1 : n1338)));
assign n1583 = /* LUT   13 30  2 */ (n677 ? n1327 : n1272);
assign n1584 = /* LUT    2 17  7 */ (n253 ? n245 : !n245);
assign n695  = /* LUT    6 20  1 */ (n258 ? 1'b0 : n694);
assign n1585 = /* LUT   11 18  7 */ (n685 ? !n1124 : (n1124 ? 1'b0 : !n798));
assign n1586 = /* LUT    5 20  2 */ (n595 ? !n597 : (n597 ? 1'b0 : (n319 ? 1'b1 : n483)));
assign n1587 = /* LUT   15 27  5 */ (n338 ? (n781 ? 1'b1 : n130) : (n781 ? !n130 : 1'b0));
assign n1588 = /* LUT   11 32  5 */ (n130 ? n526 : n633);
assign n1589 = /* LUT   15 22  6 */ (io_33_1_1 ? 1'b0 : \wb_dat_i[4] );
assign n1590 = /* LUT    9 19  6 */ (n75 ? (n800 ? 1'b1 : n802) : 1'b1);
assign n1591 = /* LUT    3 19  6 */ (n37 ? (io_33_1_1 ? !n254 : (n365 ? 1'b1 : !n254)) : (io_33_1_1 ? 1'b0 : (n365 ? n254 : 1'b0)));
assign n1592 = /* LUT   12 24  0 */ (n666 ? n1069 : n1164);
assign n1593 = /* LUT   17 23  3 */ (n1309 ? (n1086 ? 1'b1 : !n677) : (n1086 ? n677 : 1'b0));
assign n1594 = /* LUT   10 24  3 */ (n666 ? n952 : n940);
assign n468  = /* LUT    4 18  4 */ (n356 ? (io_33_1_1 ? 1'b1 : n352) : (io_33_1_1 ? 1'b1 : (n352 ? 1'b1 : n263)));
assign n1596 = /* LUT    7 23  2 */ (\wb_dat_i[5]  ? !io_33_1_1 : 1'b0);
assign n1597 = /* LUT   14 20  0 */ (n815 ? (n1338 ? !n918 : 1'b0) : (n1285 ? 1'b1 : (n1338 ? !n918 : 1'b0)));
assign n1598 = /* LUT   11 30  2 */ (n526 ? (n633 ? 1'b1 : n130) : (n633 ? !n130 : 1'b0));
assign n1599 = /* LUT   16 28  6 */ (n1375 ? (n1422 ? 1'b1 : !n677) : (n1422 ? n677 : 1'b0));
assign n1600 = /* LUT   14 27  6 */ (n666 ? n1259 : n1310);
assign n1268 = /* LUT   12 28  5 */ (n1196 ? (n1267 ? 1'b1 : n677) : (n1267 ? !n677 : 1'b0));
assign n1133 = /* LUT   11 19  4 */ (n798 ? (n892 ? (n1130 ? !n1127 : 1'b1) : !n1127) : (n892 ? !n1130 : 1'b0));
assign n605  = /* LUT    5 21  1 */ (n75 ? (n604 ? n499 : 1'b0) : (n604 ? 1'b0 : (n499 ? !n473 : 1'b0)));
assign n1604 = /* LUT   15 24  4 */ (n441 ? (n1412 ? 1'b1 : n677) : (n1412 ? !n677 : 1'b0));
assign n1605 = /* LUT   15 23  5 */ (n286 ? (n708 ? (n1313 ? 1'b1 : n1042) : n1313) : (n708 ? n1042 : 1'b0));
assign n1606 = /* LUT    7 27  7 */ (n710 ? 1'b0 : (n709 ? 1'b0 : (n408 ? n686 : 1'b0)));
assign n1607 = /* LUT   12 31  1 */ (n677 ? n1213 : n1281);
assign n1608 = /* LUT   17 16  2 */ (n104 ? (n517 ? 1'b1 : io_33_1_1) : io_33_1_1);
assign n1609 = /* LUT   22 20  6 */ (\wb_adr_i[3]  ? 1'b0 : \wb_dat_i[2] );
assign n1610 = /* LUT    7 20  3 */ (\wb_dat_i[22]  ? !io_33_1_1 : 1'b0);
assign n1611 = /* LUT    9 17  3 */ (n78 ? (n258 ? 1'b0 : !io_33_1_1) : 1'b0);
assign n1612 = /* LUT   14 23  1 */ (io_33_19_0 ? !io_33_1_1 : 1'b0);
assign n1613 = /* LUT    1 18  7 */ (n162 ? n154 : !n154);
assign n1216 = /* LUT   11 31  1 */ (n666 ? n772 : n945);
assign n1615 = /* LUT   16 22  4 */ (io_33_1_1 ? 1'b0 : \dd_pad_i[2] );
assign n1616 = /* LUT   16 27  7 */ (n677 ? n1425 : n1324);
assign n1617 = /* LUT    6 22  7 */ (wb_stb_i ? (n17 ? 1'b0 : (io_0_6_0 ? wb_we_i : 1'b0)) : 1'b0);
assign n613  = /* LUT    5 22  0 */ (n320 ? io_33_1_1 : 1'b1);
assign n1618 = /* LUT   15 25  3 */ (n96 ? (n388 ? 1'b1 : (n1359 ? \wb_adr_i[5]  : 1'b0)) : (n1359 ? \wb_adr_i[5]  : 1'b0));
assign n1619 = /* LUT   13 18  3 */ (n377 ? (n1005 ? (n465 ? 1'b1 : n104) : n465) : (n1005 ? n104 : 1'b0));
assign n1620 = /* LUT   15 20  4 */ (io_33_1_1 ? 1'b0 : io_33_19_0);
assign n1621 = /* LUT    3 26  1 */ (io_33_1_1 ? 1'b0 : \wb_dat_i[25] );
assign n1622 = /* LUT   12 30  2 */ (n964 ? (n779 ? 1'b1 : !n130) : (n779 ? n130 : 1'b0));
assign n1623 = /* LUT    5 24  3 */ (\wb_dat_i[23]  ? !n118 : 1'b0);
assign n1624 = /* LUT   10 26  5 */ (n633 ? (n526 ? 1'b1 : n130) : (n526 ? !n130 : 1'b0));
assign n1625 = /* LUT    9 18  2 */ (n166 ? n67 : n894);
assign n1626 = /* LUT   14 29  7 */ (n666 ? n662 : n1383);
assign n1627 = /* LUT   14 22  6 */ (n677 ? n1066 : n1173);
assign n1628 = /* LUT   11 28  0 */ (n968 ? (n769 ? 1'b1 : n130) : (n769 ? !n130 : 1'b0));
assign n1629 = /* LUT   16 21  5 */ (n998 ? (n1453 ? 1'b1 : (n1397 ? 1'b1 : n758)) : (n1453 ? 1'b1 : n1397));
assign n1471 = /* LUT   16 26  4 */ (n677 ? n864 : n1368);
assign n1631 = /* LUT    9 28  1 */ (n636 ? (n634 ? 1'b1 : !n130) : (n634 ? n130 : 1'b0));
assign n405  = /* LUT    3 22  4 */ (n209 ? 1'b0 : (n210 ? 1'b0 : !n220));
assign n1632 = /* LUT   18 24  2 */ (n1519 ? 1'b0 : (n1520 ? 1'b0 : (n1470 ? 1'b0 : !n1432)));
assign n1633 = /* LUT    6 17  6 */ (n673 ? (io_33_1_1 ? !n450 : (n450 ? n575 : 1'b1)) : (io_33_1_1 ? 1'b0 : (n450 ? n575 : 1'b0)));
assign n1634 = /* LUT   10 30  2 */ (n130 ? n978 : n1105);
assign n1635 = /* LUT    4 20  7 */ (n497 ? n383 : !n383);
assign n1636 = /* LUT   13 19  4 */ (\wb_dat_i[19]  ? !io_33_1_1 : 1'b0);
assign n1435 = /* LUT   15 30  2 */ (n677 ? n1424 : n1322);
assign n1638 = /* LUT   14 18  3 */ (io_33_1_1 ? 1'b1 : \wb_dat_i[19] );
assign n1639 = /* LUT   12 29  3 */ (n666 ? n863 : n1200);
assign n1640 = /* LUT    1 20  4 */ (n182 ? !n186 : n186);
assign n1641 = /* LUT   19 25  6 */ (n1507 ? 1'b0 : (n1526 ? 1'b0 : (n817 ? 1'b0 : !n1426)));
assign n1479 = /* LUT   17 18  0 */ (n599 ? (n708 ? 1'b1 : (n512 ? n750 : 1'b0)) : (n512 ? n750 : 1'b0));
assign n1643 = /* LUT    5 25  0 */ (n636 ? (n634 ? 1'b1 : !n130) : (n634 ? n130 : 1'b0));
assign n1644 = /* LUT   10 29  4 */ (n130 ? n769 : n968);
assign n1645 = /* LUT    4 23  3 */ (n297 ? (io_33_1_1 ? 1'b0 : n176) : (io_33_1_1 ? 1'b0 : (n176 ? 1'b1 : n402)));
assign n1646 = /* LUT   14 28  4 */ (n547 ? (n962 ? 1'b1 : !n130) : (n962 ? n130 : 1'b0));
assign n1647 = /* LUT    6 29  5 */ (n287 ? (io_33_1_1 ? 1'b0 : n653) : (io_33_1_1 ? 1'b0 : n642));
assign n1151 = /* LUT   11 22  6 */ (n1078 ? (n767 ? 1'b1 : n677) : (n767 ? !n677 : 1'b0));
assign n1649 = /* LUT   11 29  7 */ (n130 ? n874 : n872);
assign n1650 = /* LUT    9 29  2 */ (n130 ? n538 : n635);
assign n1651 = /* LUT   13 23  1 */ (n169 ? n1169 : n1294);
assign n1652 = /* LUT    3 23  7 */ (n307 ? 1'b0 : (n258 ? !n78 : (n78 ? 1'b0 : !n390)));
assign n1653 = /* LUT    2 21  3 */ (n291 ? (n67 ? n193 : !n193) : (n67 ? !n193 : n193));
assign n1654 = /* LUT    7 29  6 */ (n635 ? (n538 ? 1'b1 : !n130) : (n538 ? n130 : 1'b0));
assign n1655 = /* LUT   18 27  3 */ (n675 ? (n1522 ? 1'b0 : \wb_adr_i[3] ) : (n1505 ? 1'b0 : \wb_adr_i[3] ));
assign n1656 = /* LUT   10 17  3 */ (n899 ? 1'b0 : (n998 ? 1'b1 : !n798));
assign n1657 = /* LUT   13 20  5 */ (io_33_1_1 ? 1'b0 : \wb_dat_i[16] );
assign n1658 = /* LUT    3 24  3 */ (\wb_dat_i[4]  ? !n118 : 1'b0);
assign n1659 = /* LUT    5 15  6 */ \dd_pad_i[10] ;
assign n1660 = /* LUT    5 26  1 */ io_33_15_1;
assign n1661 = /* LUT   11 25  4 */ (n764 ? (n720 ? 1'b1 : !n130) : (n720 ? n130 : 1'b0));
assign n1662 = /* LUT   16 16  7 */ (\wb_dat_i[0]  ? !io_33_1_1 : 1'b0);
assign n1663 = /* LUT   10 28  7 */ (n719 ? (n643 ? 1'b1 : !n130) : (n643 ? n130 : 1'b0));
assign n1664 = /* LUT    4 22  0 */ (n300 ? (io_33_1_1 ? 1'b1 : n515) : n68);
assign n1665 = /* LUT   11 26  6 */ (n130 ? n849 : n850);
assign n1666 = /* LUT   16 19  3 */ (io_33_1_1 ? 1'b0 : \wb_dat_i[22] );
assign n1667 = /* LUT    9 30  3 */ (n666 ? n736 : n868);
assign n1668 = /* LUT   13 24  0 */ (n130 ? n874 : n872);
assign n1669 = /* LUT   15 14  1 */ (io_33_14_0 ? !io_33_1_1 : 1'b0);
assign n1670 = /* LUT    3 20  6 */ (n163 ? (io_33_1_1 ? 1'b0 : n199) : n190);
assign n277  = /* LUT    2 20  0 */ (n151 ? 1'b1 : (n269 ? 1'b1 : (n267 ? 1'b1 : n268)));
assign n1672 = /* LUT    6 19  4 */ \wb_dat_i[19] ;
assign n1673 = /* LUT    4 10  6 */ \wb_sel_i[3] ;
assign n1674 = /* LUT   10 16  0 */ (n881 ? (n880 ? (n758 ? 1'b1 : n512) : n512) : (n880 ? n758 : 1'b0));
assign n1675 = /* LUT   15 28  0 */ (n677 ? n1252 : n1373);
assign n1676 = /* LUT   13 21  6 */ (n169 ? n1026 : n86);
assign n1677 = /* LUT    1 22  6 */ (io_33_1_1 ? 1'b0 : \wb_dat_i[27] );
assign n1678 = /* LUT    5 27  6 */ (n130 ? n430 : n428);
assign n1679 = /* LUT   22 16  2 */ (n758 ? (n517 ? 1'b1 : io_33_1_1) : io_33_1_1);
assign n1680 = /* LUT   16 31  6 */ (n1107 ? (n663 ? 1'b1 : !n675) : (n663 ? n675 : 1'b0));
assign n1681 = /* LUT    4 21  1 */ (n300 ? (io_33_1_1 ? 1'b1 : n302) : n369);
assign n1682 = /* LUT    2 24  5 */ (n325 ? (n67 ? n209 : !n209) : (n67 ? !n209 : n209));
assign n1683 = /* LUT   14 19  5 */ (\wb_dat_i[5]  ? !io_33_1_1 : 1'b0);
assign n1141 = /* LUT   11 20  4 */ (n892 ? (n1119 ? !n386 : (n893 ? 1'b1 : !n386)) : (n1119 ? 1'b0 : n893));
assign n1685 = /* LUT   11 27  5 */ (n526 ? (n633 ? 1'b1 : n130) : (n633 ? !n130 : 1'b0));
assign n1686 = /* LUT   13 25  3 */ n635;
assign n1687 = /* LUT    3 21  1 */ (n317 ? 1'b0 : n280);
assign n312  = /* LUT    2 23  1 */ (n176 ? 1'b1 : io_33_1_1);
assign n1688 = /* LUT   10 19  1 */ (n471 ? (n506 ? 1'b0 : n75) : (n506 ? 1'b0 : (n362 ? !n75 : n75)));
assign n1689 = /* LUT    7 28  2 */ (n130 ? n720 : n764);
assign n1690 = /* LUT   14 26  7 */ n874;
assign n1691 = /* LUT   14 15  0 */ (io_33_13_0 ? !io_33_1_1 : 1'b0);
assign n1692 = /* LUT    1 23  1 */ \dd_pad_i[0] ;
assign n1693 = /* LUT    7 18  1 */ (n118 ? 1'b0 : (n684 ? n666 : n677));
assign n1694 = /* LUT    9 27  1 */ (n337 ? (n131 ? 1'b1 : n130) : (n131 ? !n130 : 1'b0));
assign n1695 = /* LUT    3 17  6 */ (n149 ? (io_33_1_1 ? !n254 : (n254 ? n41 : 1'b1)) : (io_33_1_1 ? 1'b0 : (n254 ? n41 : 1'b0)));
assign n1696 = /* LUT   14 25  3 */ (n130 ? n781 : n338);
assign n1697 = /* LUT    6 30  0 */ (n557 ? (io_33_1_1 ? 1'b0 : (n287 ? 1'b1 : n646)) : (io_33_1_1 ? 1'b0 : (n287 ? 1'b0 : n646)));
assign n1698 = /* LUT   11 21  3 */ (n959 ? (n782 ? (n96 ? 1'b1 : n104) : n96) : (n782 ? n104 : 1'b0));
assign n1699 = /* LUT   11 24  4 */ (n666 ? n951 : n1063);
assign n1700 = /* LUT    4 26  3 */ (\wb_dat_i[17]  ? !n118 : 1'b0);
assign n1701 = /* LUT    9 24  5 */ n634;
assign n358  = /* LUT    3 18  0 */ (n255 ? 1'b1 : (n166 ? 1'b1 : (n165 ? 1'b1 : !n51)));
assign n1523 = /* LUT   18 28  6 */ (n688 ? n708 : 1'b0);
assign n1703 = /* LUT   16 15  0 */ (io_33_14_0 ? !io_33_1_1 : 1'b0);
assign n1704 = /* LUT    5 16  2 */ (n152 ? !n448 : (n565 ? !n448 : (n448 ? 1'b0 : !n352)));
assign n1705 = /* LUT   10 25  7 */ (n130 ? n874 : n872);
assign n1706 = /* LUT   10 18  6 */ (n892 ? (n1014 ? (n897 ? !n1011 : 1'b1) : !n897) : (n1014 ? !n1011 : 1'b0));
assign n1707 = /* LUT   20 27  3 */ (io_33_1_1 ? 1'b0 : io_33_9_0);
assign n1708 = /* LUT   14 21  6 */ (io_33_1_1 ? 1'b0 : io_33_19_0);
assign n1709 = /* LUT   12 20  0 */ (\dd_pad_i[2]  ? 1'b1 : io_33_1_1);
assign n1710 = /* LUT    6 26  5 */ (n631 ? 1'b0 : (n328 ? 1'b1 : (n376 ? !n130 : 1'b1)));
assign n753  = /* LUT    7 19  2 */ (n686 ? (n752 ? 1'b1 : !n666) : (n752 ? 1'b1 : n666));
assign n1711 = /* LUT    9 20  0 */ \wb_dat_i[2] ;
assign n1712 = /* LUT   14 24  0 */ (n1297 ? (n814 ? 1'b0 : n762) : (n814 ? n746 : (n746 ? 1'b1 : n762)));
assign n1713 = /* LUT    2  7  4 */ (io_0_3_1 ? (io_0_4_1 ? (io_0_3_0 ? !io_0_4_0 : 1'b1) : 1'b1) : 1'b1);
assign n1714 = /* LUT    6 25  1 */ (n130 ? (n376 ? 1'b0 : !n539) : (n376 ? !n520 : !n539));
assign n1123 = /* LUT   11 18  2 */ (n749 ? (n750 ? 1'b0 : n893) : (n892 ? 1'b1 : (n750 ? 1'b0 : n893)));
assign n1716 = /* LUT    4 25  2 */ io_33_17_0;
assign n1717 = /* LUT   10 22  3 */ (n75 ? n803 : n579);
assign n1718 = /* LUT    9 25  6 */ (n666 ? n843 : n835);
assign n1719 = /* LUT   13 27  5 */ (n130 ? n966 : n847);
assign n1720 = /* LUT    3 19  3 */ (n254 ? (io_33_1_1 ? 1'b0 : n274) : n34);
assign n1721 = /* LUT    5 17  1 */ io_33_14_0;
assign n1722 = /* LUT   10 24  4 */ (n719 ? (n643 ? 1'b1 : n130) : (n643 ? !n130 : 1'b0));
assign n1723 = /* LUT   10 21  7 */ (n757 ? !n1050 : (n1050 ? 1'b0 : !n893));
assign n1724 = /* LUT   12 27  1 */ (n130 ? n131 : n337);
assign n1725 = /* LUT   17 20  2 */ (wb_clk_i ? !io_33_1_1 : 1'b0);
assign n1477 = /* LUT   16 28  3 */ (n985 ? (n677 ? 1'b1 : n1306) : (n677 ? 1'b0 : n1306));
assign n1727 = /* LUT    7 16  3 */ (io_33_1_1 ? 1'b1 : \wb_dat_o[5] );
assign n1728 = /* LUT    9 21  3 */ (n708 ? (n601 ? 1'b1 : (n908 ? n512 : 1'b0)) : (n908 ? n512 : 1'b0));
assign n1729 = /* LUT   13 31  2 */ (n1278 ? (n1331 ? 1'b1 : !n675) : (n1331 ? n675 : 1'b0));
assign n1730 = /* LUT   18 22  5 */ (n272 ? (n1337 ? !io_33_7_0 : 1'b0) : 1'b0);
assign n1731 = /* LUT   14 27  1 */ (n968 ? (n769 ? 1'b1 : n130) : (n769 ? !n130 : 1'b0));
assign n1732 = /* LUT    6 24  2 */ (n130 ? n521 : n328);
assign n1733 = /* LUT   11 19  1 */ (n1126 ? !n1131 : (n1131 ? 1'b0 : !n798));
assign n1734 = /* LUT    4 24  5 */ (n118 ? 1'b0 : \wb_dat_i[25] );
assign n1735 = /* LUT    9 26  7 */ (n130 ? (n958 ? 1'b0 : (n376 ? n417 : 1'b1)) : !n958);
assign n1320 = /* LUT   13 28  4 */ (n1185 ? (n1237 ? 1'b1 : n666) : (n1237 ? !n666 : 1'b0));
assign n1737 = /* LUT   18 21  1 */ (\wb_dat_i[2]  ? (io_33_8_0 ? (n1486 ? !io_33_7_0 : 1'b0) : 1'b0) : 1'b0);
assign n1738 = /* LUT   17 27  0 */ (n762 ? (n1053 ? (n1472 ? 1'b0 : n746) : 1'b1) : (n1472 ? 1'b0 : n746));
assign n577  = /* LUT    5 18  0 */ (n568 ? 1'b1 : (n476 ? 1'b1 : (n571 ? 1'b1 : n572)));
assign n1739 = /* LUT   10 27  5 */ (io_33_1_1 ? 1'b0 : io_33_17_0);
assign n1740 = /* LUT   10 20  4 */ (n1017 ? !n1031 : (n1031 ? 1'b0 : !n798));
assign n1741 = /* LUT   12 26  2 */ (n130 ? n779 : n964);
assign n1742 = /* LUT   17 21  1 */ (\wb_dat_i[2]  ? 1'b0 : (io_33_8_0 ? 1'b0 : (io_33_7_0 ? n1486 : 1'b0)));
assign n1743 = /* LUT    1 18  2 */ (n157 ? (n67 ? n59 : !n59) : (n67 ? !n59 : n59));
assign n1744 = /* LUT   16 27  2 */ (n872 ? (n874 ? 1'b1 : n130) : (n874 ? !n130 : 1'b0));
assign n1745 = /* LUT    7 17  4 */ (n742 ? (n67 ? n570 : !n570) : (n67 ? !n570 : n570));
assign n1746 = /* LUT    9 22  2 */ (n816 ? 1'b1 : (n923 ? 1'b1 : (n824 ? 1'b1 : n592)));
assign n723  = /* LUT    6 27  3 */ (n427 ? (n376 ? 1'b0 : !n624) : (n376 ? !n130 : !n624));
assign n1748 = /* LUT   13 18  6 */ (n701 ? (n611 ? 1'b1 : (n512 ? n902 : 1'b0)) : (n512 ? n902 : 1'b0));
assign n1749 = /* LUT    5 24  6 */ (n118 ? 1'b0 : io_33_13_0);
assign n1750 = /* LUT    5 19  7 */ (n471 ? (n485 ? 1'b1 : n489) : (n485 ? !n75 : (n489 ? !n75 : 1'b0)));
assign n1751 = /* LUT   10 26  2 */ (n130 ? n337 : n131);
assign n1752 = /* LUT   10 23  5 */ (n780 ? (n234 ? 1'b1 : n130) : (n234 ? !n130 : 1'b0));
assign n1753 = /* LUT    7 21  1 */ (io_33_1_1 ? 1'b0 : \wb_dat_o[5] );
assign n1345 = /* LUT   14 22  3 */ (n994 ? (n708 ? (n1294 ? 1'b1 : n512) : n512) : (n708 ? n1294 : 1'b0));
assign n1755 = /* LUT   12 25  3 */ (n1084 ? (n1088 ? 1'b1 : !n666) : (n1088 ? n666 : 1'b0));
assign n1493 = /* LUT   17 22  0 */ (n97 ? n701 : 1'b0);
assign n1757 = /* LUT    4 19  3 */ (n362 ? 1'b1 : (n452 ? (n458 ? 1'b1 : n273) : 1'b1));
assign n1758 = /* LUT    9 28  4 */ (n130 ? n849 : n850);
assign n935  = /* LUT    9 23  5 */ (n931 ? (n746 ? !n819 : 1'b0) : (n762 ? 1'b1 : (n746 ? !n819 : 1'b0)));
assign n1760 = /* LUT   10 30  7 */ (n720 ? (n764 ? 1'b1 : !n130) : (n764 ? n130 : 1'b0));
assign n1761 = /* LUT   13 19  1 */ (io_33_9_0 ? !io_33_1_1 : 1'b0);
assign n1762 = /* LUT   15 21  0 */ (n901 ? (n1127 ? 1'b0 : n1285) : (n1127 ? n1338 : (n1285 ? 1'b1 : n1338)));
assign n1763 = /* LUT   13 30  6 */ (n130 ? n847 : n966);
assign n1764 = /* LUT    2 17  3 */ (n249 ? (n67 ? n241 : !n241) : (n67 ? !n241 : n241));
assign n1765 = /* LUT   10 32  5 */ (n130 ? n781 : n338);
assign n1766 = /* LUT    5 20  6 */ (n345 ? (wb_we_i ? 1'b1 : !n286) : 1'b1);
assign n1767 = /* LUT   15 27  1 */ (n964 ? (n779 ? 1'b1 : n130) : (n779 ? !n130 : 1'b0));
assign n1768 = /* LUT    7 26  0 */ (n523 ? (n376 ? 1'b0 : !n544) : (n376 ? !n130 : !n544));
assign n1769 = /* LUT    9 19  2 */ (n75 ? n801 : n791);
assign n1770 = /* LUT   12 19  5 */ (n798 ? (n1230 ? 1'b0 : n805) : !n1230);
assign n1771 = /* LUT   12 24  4 */ (n130 ? n828 : n827);
assign n1772 = /* LUT   16 25  0 */ (n1414 ? (n762 ? !n1130 : 1'b0) : (n762 ? (n746 ? 1'b1 : !n1130) : n746));
assign n1773 = /* LUT    4 18  0 */ (n180 ? 1'b1 : (io_33_1_1 ? 1'b1 : (n356 ? 1'b0 : n263)));
assign n1774 = /* LUT   13 23  6 */ (n1247 ? (n666 ? n953 : 1'b1) : (n666 ? n953 : 1'b0));
assign n1775 = /* LUT    7 23  6 */ (io_33_14_0 ? !io_33_1_1 : 1'b0);
assign n1776 = /* LUT   16 23  3 */ (n1404 ? \wb_adr_i[5]  : 1'b0);
assign n1777 = /* LUT   10 17  6 */ (n798 ? (n1000 ? 1'b0 : n679) : !n1000);
assign n1778 = /* LUT   12 28  1 */ (n1241 ? (n1266 ? 1'b1 : !n677) : (n1266 ? n677 : 1'b0));
assign n1779 = /* LUT   17 19  4 */ (n1441 ? 1'b1 : (n1482 ? 1'b1 : (n1444 ? 1'b1 : n1446)));
assign n1780 = /* LUT    5 26  4 */ \wb_dat_o[5] ;
assign n1781 = /* LUT    5 21  5 */ (n510 ? 1'b0 : (wb_we_i ? (n509 ? 1'b0 : n473) : 1'b0));
assign n1782 = /* LUT   10 28  0 */ (n130 ? n547 : n962);
assign n1411 = /* LUT   15 24  0 */ (n675 ? (n1353 ? 1'b0 : \wb_adr_i[3] ) : (\wb_adr_i[3]  ? !n1352 : 1'b0));
assign n1784 = /* LUT    7 27  3 */ (n710 ? (n709 ? 1'b0 : (n408 ? !n686 : 1'b0)) : 1'b0);
assign n1785 = /* LUT   12 18  6 */ (n1225 ? (n67 ? n886 : !n886) : (n67 ? !n886 : n886));
assign n1786 = /* LUT   12 31  5 */ (n975 ? (n1101 ? 1'b1 : n666) : (n1101 ? !n666 : 1'b0));
assign n1284 = /* LUT   12 32  0 */ (n866 ? (n1096 ? 1'b1 : !n666) : (n1096 ? n666 : 1'b0));
assign n1788 = /* LUT    9 30  6 */ (n869 ? (n873 ? 1'b1 : !n666) : (n873 ? n666 : 1'b0));
assign n1789 = /* LUT   13 24  7 */ (n538 ? (n635 ? 1'b1 : !n130) : (n635 ? n130 : 1'b0));
assign n1790 = /* LUT    7 20  7 */ (wb_clk_i ? !io_33_1_1 : 1'b0);
assign n1458 = /* LUT   16 22  0 */ (n1134 ? (n96 ? (n104 ? 1'b1 : n1400) : n104) : (n96 ? n1400 : 1'b0));
assign n1792 = /* LUT   10 16  5 */ (io_33_1_1 ? 1'b1 : (n517 ? (n465 ? !io_33_5_0 : 1'b0) : 1'b0));
assign n1793 = /* LUT   13 21  3 */ (n679 ? (n1169 ? (n701 ? 1'b1 : n758) : n758) : (n1169 ? n701 : 1'b0));
assign n1794 = /* LUT    3 25  1 */ (n130 ? n131 : n337);
assign n1795 = /* LUT    5 27  3 */ (n432 ? (n126 ? 1'b1 : n130) : (n126 ? !n130 : 1'b0));
assign n1796 = /* LUT    5 22  4 */ (io_33_1_1 ? 1'b0 : n473);
assign n1797 = /* LUT   10 31  1 */ (n130 ? n781 : n338);
assign n763  = /* LUT    7 24  2 */ (n709 ? !n710 : n710);
assign n1799 = /* LUT   12 17  7 */ (io_33_1_1 ? 1'b1 : \wb_dat_i[20] );
assign n1800 = /* LUT   14 19  0 */ (io_33_1_1 ? 1'b1 : \dd_pad_i[2] );
assign n1801 = /* LUT   12 30  6 */ (n677 ? n1207 : n1276);
assign n1802 = /* LUT    4 27  7 */ (n75 ? n535 : n423);
assign n1803 = /* LUT   13 25  4 */ (n130 ? \dd_pad_i[1]  : wb_inta_o);
assign n1804 = /* LUT    9 18  6 */ (n892 ? (n799 ? !n879 : (n879 ? n893 : 1'b1)) : (n799 ? 1'b0 : n893));
assign n1805 = /* LUT   14 29  3 */ (n666 ? n1090 : n1321);
assign n1452 = /* LUT   16 21  1 */ (n91 ? (n286 ? (n708 ? 1'b1 : n929) : n708) : (n286 ? n929 : 1'b0));
assign n1020 = /* LUT   10 19  4 */ (n895 ? (n1019 ? 1'b1 : n791) : (n1019 ? !n791 : 1'b0));
assign n1807 = /* LUT   15 29  4 */ (n1269 ? (n1434 ? 1'b1 : n677) : (n1434 ? !n677 : 1'b0));
assign n1292 = /* LUT   13 22  2 */ (n675 ? n1234 : n1291);
assign n1809 = /* LUT    3 22  0 */ (n301 ? (io_33_1_1 ? 1'b1 : (n287 ? !n288 : 1'b0)) : (io_33_1_1 ? 1'b1 : (n287 ? !n288 : 1'b1)));
assign n1810 = /* LUT    4 20  3 */ (n493 ? (n67 ? n385 : !n385) : (n67 ? !n385 : n385));
assign n1811 = /* LUT    7 18  4 */ (n377 ? (n376 ? (n714 ? !n118 : 1'b0) : !n118) : (n714 ? !n118 : 1'b0));
assign n1812 = /* LUT    9 27  6 */ (n130 ? n720 : n764);
assign n766  = /* LUT    7 25  5 */ (n377 ? 1'b0 : (n286 ? n517 : 1'b0));
assign n1813 = /* LUT   12 16  0 */ (\wb_dat_i[8]  ? !io_33_1_1 : 1'b0);
assign n1814 = /* LUT   12 29  7 */ (n827 ? (n828 ? 1'b1 : !n130) : (n828 ? n130 : 1'b0));
assign n1815 = /* LUT    4 26  4 */ (n118 ? 1'b0 : \wb_dat_i[21] );
assign n1816 = /* LUT    4 23  7 */ (n396 ? 1'b1 : (n397 ? (diown_pad_o ? 1'b1 : n389) : 1'b0));
assign n1817 = /* LUT    9 24  0 */ (n130 ? \dd_pad_i[6]  : \dd_pad_i[0] );
assign n1818 = /* LUT   13 26  5 */ n962;
assign n1819 = /* LUT   14 28  0 */ (n1253 ? (n1314 ? 1'b1 : n666) : (n1314 ? !n666 : 1'b0));
assign n1820 = /* LUT    2 22  3 */ (n221 ? (n102 ? 1'b1 : !n169) : (n102 ? n169 : 1'b0));
assign n1821 = /* LUT   10 18  3 */ (n751 ? (n997 ? (io_33_1_1 ? !n460 : 1'b1) : !n460) : (n997 ? (io_33_1_1 ? 1'b0 : n460) : 1'b0));
assign n1822 = /* LUT   15 18  5 */ (io_33_1_1 ? 1'b1 : \wb_dat_i[21] );
assign n412  = /* LUT    3 23  3 */ (n259 ? io_33_1_1 : (n154 ? io_33_1_1 : 1'b1));
assign n1823 = /* LUT    2 21  7 */ (n295 ? n66 : !n66);
assign n777  = /* LUT    7 29  2 */ (n677 ? n734 : n717);
assign n1825 = /* LUT   12 20  5 */ (io_33_1_1 ? 1'b0 : \wb_dat_i[5] );
assign n660  = /* LUT    5 29  1 */ (n75 ? n536 : n225);
assign n1827 = /* LUT    7 19  7 */ (n377 ? (n686 ? (n317 ? 1'b1 : !n677) : (n317 ? 1'b1 : n677)) : (n686 ? (n317 ? 1'b0 : !n677) : (n317 ? 1'b0 : n677)));
assign n1828 = /* LUT    9 20  7 */ \wb_dat_i[19] ;
assign n1829 = /* LUT    3 24  7 */ (\dd_pad_i[2]  ? !n118 : 1'b0);
assign n1830 = /* LUT   12 23  1 */ (n1035 ? 1'b1 : (n1243 ? 1'b1 : (n711 ? 1'b1 : n1065)));
assign n1831 = /* LUT   11 25  0 */ (n849 ? (n850 ? 1'b1 : !n130) : (n850 ? n130 : 1'b0));
assign n1832 = /* LUT    4 25  5 */ \wb_dat_i[0] ;
assign n516  = /* LUT    4 22  4 */ (n84 ? (n514 ? (io_33_1_1 ? 1'b0 : n317) : 1'b0) : 1'b0);
assign n1834 = /* LUT    9 25  3 */ (n833 ? (n666 ? n846 : 1'b1) : (n666 ? n846 : 1'b0));
assign n1835 = /* LUT   13 27  2 */ (n978 ? (n1105 ? 1'b1 : n130) : (n1105 ? !n130 : 1'b0));
assign n1836 = /* LUT    6 28  2 */ (n287 ? (n732 ? !io_33_1_1 : 1'b0) : (n640 ? !io_33_1_1 : 1'b0));
assign n1161 = /* LUT   11 23  1 */ (n1160 ? (n1057 ? 1'b1 : n675) : (n1057 ? !n675 : 1'b0));
assign n1048 = /* LUT   10 21  2 */ (n892 ? (n918 ? !n931 : (n893 ? 1'b1 : !n931)) : (n918 ? 1'b0 : n893));
assign n1839 = /* LUT   15 19  6 */ (dmarq_pad_i ? (n1391 ? 1'b1 : (n465 ? 1'b1 : n513)) : (n1391 ? 1'b1 : n513));
assign n1840 = /* LUT    3 20  2 */ (n163 ? (io_33_1_1 ? 1'b0 : n195) : n187);
assign n1841 = /* LUT    2 20  4 */ (n69 ? 1'b1 : (n174 ? (n266 ? 1'b1 : n193) : 1'b1));
assign n1842 = /* LUT   12 27  4 */ (n964 ? (n779 ? 1'b1 : n130) : (n779 ? !n130 : 1'b0));
assign n1843 = /* LUT    5 30  0 */ (n654 ? (io_33_1_1 ? 1'b0 : (n287 ? 1'b1 : n553)) : (io_33_1_1 ? 1'b0 : (n287 ? 1'b0 : n553)));
assign n909  = /* LUT    9 21  4 */ (n792 ? 1'b0 : (n470 ? (n362 ? n616 : 1'b0) : 1'b0));
assign n1845 = /* LUT   13 31  7 */ \dd_pad_i[13] ;
assign n1846 = /* LUT   12 22  2 */ (io_33_1_1 ? 1'b0 : \wb_dat_i[21] );
assign n1847 = /* LUT    1 22  2 */ (io_33_1_1 ? 1'b0 : \wb_dat_i[5] );
assign n1848 = /* LUT    4 24  2 */ (\wb_dat_i[16]  ? !n118 : 1'b0);
assign n1849 = /* LUT    4 21  5 */ (n300 ? (io_33_1_1 ? 1'b0 : n85) : n368);
assign n1850 = /* LUT    9 26  2 */ (n376 ? (n956 ? 1'b0 : (n431 ? 1'b1 : !n130)) : !n956);
assign n1851 = /* LUT   13 28  3 */ (n675 ? (n1319 ? n286 : 1'b0) : (n286 ? n1263 : 1'b0));
assign n1852 = /* LUT    2 24  1 */ (n321 ? (n67 ? n204 : !n204) : (n67 ? !n204 : n204));
assign n1853 = /* LUT   11 20  0 */ (n892 ? (n1038 ? !n1138 : (n893 ? 1'b1 : !n1138)) : (n1038 ? 1'b0 : n893));
assign n1854 = /* LUT   10 20  1 */ (n798 ? (n1030 ? 1'b0 : n959) : !n1030);
assign n1855 = /* LUT   15 15  6 */ (n1386 ? (n1007 ? (n512 ? 1'b1 : n701) : n701) : (n1007 ? n512 : 1'b0));
assign n1856 = /* LUT    3 21  5 */ (io_33_1_1 ? 1'b0 : (n393 ? n392 : 1'b0));
assign n1857 = /* LUT    2 23  5 */ (n214 ? (io_33_1_1 ? !n205 : (n109 ? 1'b1 : !n205)) : (io_33_1_1 ? 1'b0 : (n109 ? n205 : 1'b0)));
assign n1858 = /* LUT   20 22  5 */ (n701 ? (n106 ? 1'b1 : (n1155 ? 1'b1 : n1401)) : (n1155 ? 1'b1 : n1401));
assign n1859 = /* LUT   12 26  7 */ (n666 ? n442 : n1171);
assign n1860 = /* LUT   17 24  1 */ (n1466 ? 1'b1 : (n1502 ? 1'b1 : (n461 ? 1'b1 : n562)));
assign n1861 = /* LUT    7 17  1 */ (n739 ? (n67 ? n567 : !n567) : (n67 ? !n567 : n567));
assign n1862 = /* LUT    9 22  5 */ (n677 ? n825 : n760);
assign n1863 = /* LUT    7 28  6 */ (n130 ? n643 : n719);
assign n1864 = /* LUT   14 26  3 */ n781;
assign n1865 = /* LUT   12 21  3 */ (\wb_dat_i[18]  ? !io_33_1_1 : 1'b0);
assign n1866 = /* LUT   13 29  0 */ (n968 ? (n769 ? 1'b1 : n130) : (n769 ? !n130 : 1'b0));
assign n1867 = /* LUT   14 25  7 */ (n675 ? n1366 : n1301);
assign n1868 = /* LUT    3 17  2 */ (n145 ? (io_33_1_1 ? 1'b1 : (n254 ? n42 : 1'b1)) : (io_33_1_1 ? n254 : (n254 ? n42 : 1'b0)));
assign n1869 = /* LUT    6 21  5 */ (n599 ? (n699 ? 1'b1 : !n169) : (n699 ? n169 : 1'b0));
assign n1870 = /* LUT   11 21  7 */ (n96 ? (n906 ? 1'b1 : (n783 ? n104 : 1'b0)) : (n783 ? n104 : 1'b0));
assign n1871 = /* LUT   16 17  5 */ (io_33_1_1 ? 1'b0 : \wb_adr_i[4] );
assign n1872 = /* LUT   10 23  0 */ (n130 ? n720 : n764);
assign n1873 = /* LUT   13 15  1 */ (io_33_1_1 ? 1'b0 : \wb_dat_o[5] );
assign n1874 = /* LUT   15 17  0 */ (\wb_dat_i[30]  ? !io_33_1_1 : 1'b0);
assign n1875 = /* LUT    7 21  6 */ (io_33_5_0 ? !io_33_1_1 : 1'b0);
assign n1876 = /* LUT   18 19  3 */ (n462 ? (n758 ? 1'b1 : (n1016 ? 1'b1 : n1219)) : (n1016 ? 1'b1 : n1219));
assign n1877 = /* LUT    3 18  4 */ (n254 ? (io_33_1_1 ? 1'b0 : n355) : n39);
assign n1878 = /* LUT   12 25  6 */ (n666 ? n440 : n433);
assign n1879 = /* LUT   17 25  2 */ DMA_req;
assign n1880 = /* LUT   10 25  3 */ (n666 ? n857 : n946);
assign n482  = /* LUT    4 19  6 */ (n275 ? n67 : n481);
assign n1882 = /* LUT    7 22  0 */ (n616 ? !io_33_1_1 : 1'b0);
assign n1883 = /* LUT    9 23  2 */ (io_33_1_1 ? 1'b0 : \wb_dat_i[17] );
assign n1884 = /* LUT   14 21  2 */ (io_33_1_1 ? 1'b0 : \wb_dat_i[16] );
assign n1885 = /* LUT    6 26  1 */ (n317 ? (n280 ? 1'b1 : n376) : n376);
assign n1117 = /* LUT   11 17  4 */ (n892 ? (n890 ? !n1006 : (n1006 ? n798 : 1'b1)) : (n890 ? 1'b0 : n798));
assign n1887 = /* LUT   15 21  5 */ (n1044 ? (n757 ? 1'b0 : n1338) : (n757 ? n1285 : (n1338 ? 1'b1 : n1285)));
assign n1327 = /* LUT   13 30  1 */ (n666 ? n1095 : n1098);
assign n1889 = /* LUT    2 17  6 */ (n252 ? (n67 ? n244 : !n244) : (n67 ? !n244 : n244));
assign n1357 = /* LUT   14 24  4 */ (n666 ? n1186 : n938);
assign n696  = /* LUT    6 20  6 */ (n319 ? !io_33_1_1 : 1'b0);
assign n1891 = /* LUT    6 25  5 */ (n130 ? (n543 ? 1'b0 : !n376) : (n543 ? (n376 ? !n521 : 1'b0) : (n376 ? !n521 : 1'b1)));
assign n1124 = /* LUT   11 18  6 */ (n363 ? (n908 ? 1'b0 : n893) : (n892 ? 1'b1 : (n908 ? 1'b0 : n893)));
assign n1893 = /* LUT   13 16  0 */ (io_33_1_1 ? 1'b0 : io_33_5_0);
assign n1894 = /* LUT   15 22  1 */ (io_33_1_1 ? 1'b0 : io_33_19_0);
assign n1895 = /* LUT    9 19  7 */ \wb_dat_i[2] ;
assign n1896 = /* LUT   12 24  1 */ (n827 ? (n828 ? 1'b1 : n130) : (n828 ? !n130 : 1'b0));
assign n1897 = /* LUT   17 26  3 */ (n666 ? n1260 : n1245);
assign n1898 = /* LUT   10 24  0 */ (n942 ? (n937 ? 1'b1 : n666) : (n937 ? !n666 : 1'b0));
assign n1899 = /* LUT    4 18  5 */ (n468 ? 1'b1 : (n53 ? 1'b0 : !n356));
assign n1900 = /* LUT    7 23  3 */ (io_33_1_1 ? 1'b0 : \wb_dat_i[8] );
assign n1901 = /* LUT   11 30  5 */ (n130 ? n634 : n636);
assign n1902 = /* LUT   16 23  6 */ (n789 ? (n758 ? 1'b1 : (n104 ? n1110 : 1'b0)) : (n104 ? n1110 : 1'b0));
assign n1903 = /* LUT   14 27  5 */ (n1105 ? (n978 ? 1'b1 : !n130) : (n978 ? n130 : 1'b0));
assign n1904 = /* LUT   12 28  6 */ (n1203 ? (n1268 ? 1'b1 : !n675) : (n1268 ? n675 : 1'b0));
assign n1905 = /* LUT    6 24  6 */ (n130 ? n520 : n419);
assign n1906 = /* LUT   11 19  5 */ (n893 ? (n1133 ? 1'b0 : n901) : !n1133);
assign n1907 = /* LUT   13 17  3 */ (\wb_dat_i[4]  ? !io_33_1_1 : 1'b0);
assign n1908 = /* LUT   15 23  2 */ (n1028 ? (n1408 ? 1'b1 : (n1349 ? 1'b1 : n701)) : (n1408 ? 1'b1 : n1349));
assign n1909 = /* LUT    7 27  4 */ (n686 ? (n408 ? (n709 ? !n710 : 1'b0) : 1'b0) : 1'b0);
assign n1910 = /* LUT   18 21  5 */ (\wb_dat_i[2]  ? (io_33_8_0 ? (\wb_adr_i[3]  ? 1'b0 : io_33_7_0) : \wb_adr_i[3] ) : (io_33_8_0 ? (\wb_adr_i[3]  ? 1'b1 : io_33_7_0) : \wb_adr_i[3] ));
assign n1281 = /* LUT   12 31  0 */ (n848 ? (n666 ? 1'b1 : n838) : (n666 ? 1'b0 : n838));
assign n1912 = /* LUT    4 17  4 */ (n257 ? 1'b1 : (n256 ? (n171 ? 1'b1 : n173) : 1'b0));
assign n1913 = /* LUT    7 20  2 */ (io_33_1_1 ? 1'b0 : io_33_13_0);
assign n1914 = /* LUT    9 17  0 */ (n884 ? 1'b0 : (n798 ? n664 : 1'b1));
assign n1915 = /* LUT   14 23  0 */ (io_33_1_1 ? 1'b0 : io_33_16_1);
assign n1916 = /* LUT    1 18  6 */ (n161 ? (n67 ? n61 : !n61) : (n67 ? !n61 : n61));
assign n1917 = /* LUT   11 31  6 */ (n849 ? (n850 ? 1'b1 : !n130) : (n850 ? n130 : 1'b0));
assign n1918 = /* LUT   16 22  5 */ (n708 ? (n93 ? 1'b1 : (n558 ? n286 : 1'b0)) : (n558 ? n286 : 1'b0));
assign n1919 = /* LUT    2 19  4 */ (n169 ? n103 : n91);
assign n1920 = /* LUT    6 22  0 */ (n17 ? 1'b1 : !\wb_adr_i[5] );
assign n1921 = /* LUT    6 27  7 */ (n644 ? 1'b0 : (n376 ? (n125 ? 1'b1 : !n130) : 1'b1));
assign n1922 = /* LUT   13 18  2 */ (n890 ? (n1006 ? (n104 ? 1'b1 : n758) : n758) : (n1006 ? n104 : 1'b0));
assign n1923 = /* LUT    7 24  5 */ (n706 ? 1'b1 : io_33_1_1);
assign n1924 = /* LUT   18 20  6 */ (n1212 ? 1'b1 : (n1513 ? 1'b1 : (n1483 ? 1'b1 : n1484)));
assign n1925 = /* LUT   12 30  3 */ (n666 ? n1097 : n1099);
assign n1926 = /* LUT    5 24  2 */ (n118 ? 1'b0 : \wb_dat_i[11] );
assign n1927 = /* LUT   10 26  6 */ (n130 ? n719 : n643);
assign n894  = /* LUT    9 18  1 */ (n357 ? 1'b1 : (n51 ? (n52 ? 1'b1 : n261) : 1'b1));
assign n1929 = /* LUT   11 28  7 */ (n130 ? n634 : n636);
assign n1453 = /* LUT   16 21  4 */ (n1018 ? (n104 ? 1'b1 : (n96 ? n1395 : 1'b0)) : (n96 ? n1395 : 1'b0));
assign n1931 = /* LUT   16 26  5 */ (n675 ? (n1367 ? 1'b0 : \wb_adr_i[3] ) : (n1471 ? 1'b0 : \wb_adr_i[3] ));
assign n1932 = /* LUT    9 28  0 */ (n130 ? n719 : n643);
assign n1933 = /* LUT    3 22  7 */ (n284 ? (n281 ? 1'b1 : !n297) : (n281 ? n297 : 1'b0));
assign n1934 = /* LUT   10 30  3 */ (n538 ? (n635 ? 1'b1 : !n130) : (n635 ? n130 : 1'b0));
assign n1935 = /* LUT   13 19  5 */ (\wb_dat_i[21]  ? !io_33_1_1 : 1'b0);
assign n1936 = /* LUT    7 25  2 */ (n130 ? n337 : n131);
assign n1937 = /* LUT   14 18  4 */ (io_33_1_1 ? 1'b1 : \wb_dat_i[11] );
assign n1938 = /* LUT   12 29  2 */ (n130 ? n769 : n968);
assign n1939 = /* LUT    1 20  7 */ (n152 ? !n67 : n67);
assign n1940 = /* LUT    5 25  1 */ (n130 ? n538 : n635);
assign n1941 = /* LUT   10 29  7 */ (n719 ? (n643 ? 1'b1 : !n130) : (n643 ? n130 : 1'b0));
assign n1942 = /* LUT    4 23  2 */ (n282 ? (n283 ? 1'b1 : !n297) : (n283 ? n297 : 1'b0));
assign n1943 = /* LUT   14 28  5 */ (n130 ? n547 : n962);
assign n1229 = /* LUT   12 19  1 */ (n892 ? (n1004 ? !n1136 : (n798 ? 1'b1 : !n1136)) : (n1004 ? 1'b0 : n798));
assign n1945 = /* LUT   11 29  0 */ (n968 ? (n769 ? 1'b1 : n130) : (n769 ? !n130 : 1'b0));
assign n1946 = /* LUT   16 20  3 */ (n1139 ? (n104 ? 1'b1 : (n96 ? n1394 : 1'b0)) : (n96 ? n1394 : 1'b0));
assign n1947 = /* LUT   21 19  4 */ (\wb_adr_i[3]  ? 1'b0 : io_33_8_0);
assign n1948 = /* LUT    9 29  3 */ (n538 ? (n635 ? 1'b1 : !n130) : (n635 ? n130 : 1'b0));
assign n1949 = /* LUT   13 23  2 */ (n1242 ? (n1249 ? 1'b1 : !n169) : (n1249 ? n169 : 1'b0));
assign n1950 = /* LUT    3 23  4 */ (n362 ? (n412 ? 1'b0 : (n219 ? n308 : 1'b1)) : (n412 ? 1'b0 : n308));
assign n1951 = /* LUT    2 21  2 */ (n290 ? (n67 ? n151 : !n151) : (n67 ? !n151 : n151));
assign n1952 = /* LUT    7 29  7 */ (n130 ? n635 : n538);
assign n1522 = /* LUT   18 27  2 */ (n1423 ? (n768 ? 1'b1 : n677) : (n768 ? !n677 : 1'b0));
assign n1954 = /* LUT    6 16  2 */ (n450 ? (io_33_1_1 ? 1'b0 : n457) : n668);
assign n1955 = /* LUT   10 17  2 */ (n888 ? 1'b0 : (n790 ? 1'b1 : !n893));
assign n1956 = /* LUT   13 20  4 */ (\dd_pad_i[7]  ? !io_33_1_1 : 1'b0);
assign n1957 = /* LUT    3 24  2 */ (n118 ? 1'b0 : \dd_pad_i[12] );
assign n1958 = /* LUT    1 21  4 */ (n69 ? !n67 : n67);
assign n1959 = /* LUT    5 26  0 */ \wb_dat_i[21] ;
assign n1960 = /* LUT   11 25  5 */ (n130 ? n234 : n780);
assign n1961 = /* LUT   10 28  4 */ (n130 ? n526 : n633);
assign n1962 = /* LUT    4 22  1 */ (n371 ? (io_33_1_1 ? 1'b1 : (n309 ? 1'b1 : !n300)) : (io_33_1_1 ? n300 : (n309 ? n300 : 1'b0)));
assign n1963 = /* LUT   12 18  2 */ (n1221 ? (n67 ? n475 : !n475) : (n67 ? !n475 : n475));
assign n1964 = /* LUT    6 28  7 */ (n75 ? n530 : n584);
assign n1965 = /* LUT   11 26  1 */ (n337 ? (n131 ? 1'b1 : !n130) : (n131 ? n130 : 1'b0));
assign n1966 = /* LUT    9 30  2 */ (n130 ? n538 : n635);
assign n1967 = /* LUT   13 24  3 */ (n634 ? (n636 ? 1'b1 : n130) : (n636 ? !n130 : 1'b0));
assign n1968 = /* LUT    3 20  5 */ (n189 ? (io_33_1_1 ? 1'b1 : (n198 ? 1'b1 : !n163)) : (io_33_1_1 ? n163 : (n198 ? n163 : 1'b0)));
assign n278  = /* LUT    2 20  1 */ (n175 ? 1'b1 : (n277 ? 1'b1 : n66));
assign n1969 = /* LUT   18 26  5 */ (n675 ? (n1509 ? 1'b0 : \wb_adr_i[3] ) : (n1419 ? 1'b0 : \wb_adr_i[3] ));
assign n1970 = /* LUT    6 19  3 */ \wb_dat_i[22] ;
assign n1971 = /* LUT    1 22  5 */ (\dd_pad_i[2]  ? !io_33_1_1 : 1'b0);
assign n1972 = /* LUT    5 27  7 */ (n229 ? (n427 ? 1'b1 : !n130) : (n427 ? n130 : 1'b0));
assign n1973 = /* LUT   10 31  5 */ (n130 ? n978 : n1105);
assign n1974 = /* LUT    4 21  0 */ (n380 ? 1'b1 : (n383 ? 1'b1 : (n381 ? 1'b1 : n382)));
assign n1975 = /* LUT   12 17  3 */ (io_33_1_1 ? 1'b1 : \wb_dat_i[22] );
assign n1976 = /* LUT   14 19  4 */ (io_33_1_1 ? 1'b0 : wb_clk_i);
assign n1977 = /* LUT   11 27  2 */ (n130 ? n847 : n966);
assign n550  = /* LUT    4 27  3 */ (n75 ? n534 : n422);
assign n1979 = /* LUT   13 25  0 */ (n130 ? \dd_pad_i[9]  : \dd_pad_i[14] );
assign n1980 = /* LUT    3 21  2 */ (n379 ? 1'b0 : (n202 ? (n79 ? 1'b0 : !n182) : 1'b0));
assign n1981 = /* LUT    2 23  0 */ (n205 ? (io_33_1_1 ? 1'b0 : n203) : n211);
assign n1982 = /* LUT   10 19  0 */ (n75 ? (io_33_1_1 ? 1'b0 : n800) : (io_33_1_1 ? 1'b0 : n795));
assign n1983 = /* LUT   15 29  0 */ (n1381 ? (n1192 ? 1'b1 : !n677) : (n1192 ? n677 : 1'b0));
assign n1984 = /* LUT   13 22  6 */ \dd_pad_i[8] ;
assign n1985 = /* LUT    7 28  1 */ (n720 ? (n764 ? 1'b1 : !n130) : (n764 ? n130 : 1'b0));
assign n1986 = /* LUT    1 23  2 */ \dd_pad_i[14] ;
assign n1987 = /* LUT    7 18  0 */ (n684 ? (n748 ? 1'b0 : !n118) : (n666 ? !n118 : 1'b0));
assign n1988 = /* LUT    9 27  2 */ (n130 ? n827 : n828);
assign n1989 = /* LUT   14 25  2 */ (n338 ? (n781 ? 1'b1 : n130) : (n781 ? !n130 : 1'b0));
assign n1990 = /* LUT    3 17  7 */ (n150 ? (io_33_1_1 ? !n254 : (n347 ? 1'b1 : !n254)) : (io_33_1_1 ? 1'b0 : (n347 ? n254 : 1'b0)));
assign n1991 = /* LUT   11 24  3 */ (n949 ? (n1061 ? 1'b1 : n666) : (n1061 ? !n666 : 1'b0));
assign n1992 = /* LUT    4 26  0 */ (n118 ? 1'b0 : \wb_dat_i[18] );
assign n1993 = /* LUT    9 24  4 */ (n130 ? \dd_pad_i[8]  : \dd_pad_i[13] );
assign n1994 = /* LUT   13 26  1 */ n966;
assign n1995 = /* LUT    3 18  3 */ (n38 ? (io_33_1_1 ? !n254 : (n55 ? 1'b1 : !n254)) : (io_33_1_1 ? 1'b0 : (n55 ? n254 : 1'b0)));
assign n1996 = /* LUT   18 28  7 */ (n1475 ? 1'b1 : (n1523 ? 1'b1 : (n1481 ? 1'b1 : n1473)));
assign n566  = /* LUT    5 16  5 */ (n447 ? 1'b1 : (n449 ? 1'b0 : !n472));
assign n1997 = /* LUT   10 25  6 */ (n954 ? (n947 ? 1'b1 : n666) : (n947 ? !n666 : 1'b0));
assign n1998 = /* LUT   10 18  7 */ (n995 ? (n1010 ? 1'b1 : n460) : (n1010 ? (io_33_1_1 ? 1'b1 : !n460) : (io_33_1_1 ? n460 : 1'b0)));
assign n1999 = /* LUT   12 20  1 */ (io_33_1_1 ? 1'b1 : \wb_dat_i[27] );
assign n2000 = /* LUT    6 26  6 */ (n716 ? 1'b0 : (n314 ? 1'b1 : (n130 ? !n376 : 1'b1)));
assign n2001 = /* LUT    5 29  5 */ (n75 ? n455 : n334);
assign n2002 = /* LUT    7 19  3 */ (n465 ? (n753 ? (n683 ? \wb_adr_i[5]  : 1'b0) : 1'b1) : (n683 ? \wb_adr_i[5]  : 1'b0));
assign n2003 = /* LUT    9 20  3 */ \wb_adr_i[3] ;
assign n2004 = /* LUT   12 23  5 */ \dd_pad_i[6] ;
assign n2005 = /* LUT    6 25  0 */ (n217 ? (io_33_1_1 ? !n205 : (n205 ? n665 : 1'b1)) : (io_33_1_1 ? 1'b0 : (n205 ? n665 : 1'b0)));
assign n1055 = /* LUT   10 22  4 */ (n580 ? (n804 ? 1'b1 : !n75) : (n804 ? n75 : 1'b0));
assign n2007 = /* LUT    9 25  7 */ (n130 ? n635 : n538);
assign n2008 = /* LUT   13 27  6 */ (n872 ? (n874 ? 1'b1 : n130) : (n874 ? !n130 : 1'b0));
assign n367  = /* LUT    3 19  0 */ (n58 ? 1'b1 : (n180 ? (n56 ? 1'b1 : n155) : 1'b1));
assign n2010 = /* LUT   16 14  0 */ (io_33_14_0 ? !io_33_1_1 : 1'b0);
assign n2011 = /* LUT   10 24  5 */ (n130 ? n643 : n719);
assign n1050 = /* LUT   10 21  6 */ (n892 ? (n1044 ? !n915 : (n798 ? 1'b1 : !n915)) : (n1044 ? 1'b0 : n798));
assign n1390 = /* LUT   15 19  2 */ (n287 ? (n992 ? (n465 ? 1'b1 : n104) : n465) : (n992 ? n104 : 1'b0));
assign n2014 = /* LUT   12 27  0 */ (n636 ? (n634 ? 1'b1 : !n130) : (n634 ? n130 : 1'b0));
assign n2015 = /* LUT   17 20  5 */ (n675 ? n1166 : n1193);
assign n2016 = /* LUT    2 11  6 */ io_0_7_1;
assign n2017 = /* LUT    9 21  0 */ (n262 ? (n758 ? 1'b1 : (n699 ? n701 : 1'b0)) : (n699 ? n701 : 1'b0));
assign n1332 = /* LUT   13 31  3 */ (n986 ? (n976 ? 1'b1 : !n666) : (n976 ? n666 : 1'b0));
assign n1517 = /* LUT   18 22  6 */ (io_33_7_0 ? (\wb_adr_i[3]  ? (\wb_adr_i[5]  ? 1'b0 : !n1489) : 1'b0) : 1'b0);
assign n2019 = /* LUT   14 27  0 */ (n666 ? n950 : n1304);
assign n2020 = /* LUT    6 24  3 */ (n523 ? (n314 ? 1'b1 : n130) : (n314 ? !n130 : 1'b0));
assign n2021 = /* LUT    4 24  6 */ (\wb_dat_i[8]  ? !n118 : 1'b0);
assign n958  = /* LUT    9 26  6 */ (n119 ? (n376 ? 1'b0 : !n546) : (n376 ? !n130 : !n546));
assign n2023 = /* LUT   13 28  7 */ (n130 ? n636 : n634);
assign n2024 = /* LUT   18 21  0 */ (n386 ? n104 : 1'b0);
assign n2025 = /* LUT   10 27  4 */ (\wb_dat_o[5]  ? !io_33_1_1 : 1'b0);
assign n2026 = /* LUT   10 20  5 */ (n169 ? n904 : n688);
assign n2027 = /* LUT    3 30  0 */ n131;
assign n2028 = /* LUT   12 26  3 */ (n666 ? n977 : n1180);
assign n2029 = /* LUT   17 21  6 */ (io_33_8_0 ? (io_33_7_0 ? 1'b0 : (n1486 ? !\wb_dat_i[2]  : 1'b0)) : 1'b0);
assign n2030 = /* LUT    1 18  1 */ (n156 ? (n67 ? n56 : !n56) : (n67 ? !n56 : n56));
assign n2031 = /* LUT    7 17  5 */ (n743 ? (n67 ? n571 : !n571) : (n67 ? !n571 : n571));
assign n923  = /* LUT    9 22  1 */ (n90 ? (n922 ? 1'b1 : (n708 ? 1'b1 : n811)) : (n922 ? 1'b1 : n811));
assign n2033 = /* LUT    6 27  2 */ (n130 ? (n722 ? 1'b0 : (n376 ? n428 : 1'b1)) : !n722);
assign n2034 = /* LUT   13 18  5 */ (n1112 ? (n701 ? (n904 ? 1'b1 : n512) : n512) : (n701 ? n904 : 1'b0));
assign n2035 = /* LUT   13 29  4 */ (n1326 ? (n1270 ? 1'b1 : n677) : (n1270 ? !n677 : 1'b0));
assign n2036 = /* LUT    6 21  1 */ (n89 ? (n697 ? 1'b1 : !n169) : (n697 ? n169 : 1'b0));
assign n2037 = /* LUT    5 19  0 */ (n270 ? (io_33_1_1 ? 1'b0 : (n75 ? n587 : 1'b1)) : (io_33_1_1 ? 1'b0 : (n75 ? n587 : 1'b0)));
assign n2038 = /* LUT   10 26  3 */ (n338 ? (n781 ? 1'b1 : !n130) : (n781 ? n130 : 1'b0));
assign n2039 = /* LUT   10 23  4 */ (n677 ? n928 : n1058);
assign n1420 = /* LUT   15 26  5 */ (n1138 ? (n1369 ? 1'b0 : n746) : (n762 ? 1'b1 : (n1369 ? 1'b0 : n746)));
assign n2041 = /* LUT    7 21  2 */ (\wb_dat_i[20]  ? !io_33_1_1 : 1'b0);
assign n2042 = /* LUT   12 25  2 */ (n130 ? n131 : n337);
assign n2043 = /* LUT    4 19  2 */ (n287 ? (n360 ? io_33_1_1 : 1'b1) : (io_33_1_1 ? 1'b1 : !n392));
assign n2044 = /* LUT    9 23  6 */ (n818 ? 1'b0 : (n935 ? 1'b0 : (n932 ? 1'b0 : !n817)));
assign n1521 = /* LUT   18 24  4 */ (n1176 ? (n675 ? 1'b1 : n1460) : (n675 ? 1'b0 : n1460));
assign n1116 = /* LUT   11 17  0 */ (n892 ? (n1111 ? !n1110 : (n893 ? 1'b1 : !n1110)) : (n1111 ? 1'b0 : n893));
assign n2047 = /* LUT    5 23  5 */ (io_33_1_1 ? 1'b0 : \wb_dat_i[23] );
assign n2048 = /* LUT   13 19  2 */ (io_33_1_1 ? 1'b0 : io_33_13_0);
assign n2049 = /* LUT   13 30  5 */ (n286 ? (n1329 ? (n675 ? 1'b1 : n1273) : (n675 ? 1'b0 : n1273)) : 1'b0);
assign n2050 = /* LUT    2 17  2 */ (n248 ? (n67 ? n240 : !n240) : (n67 ? !n240 : n240));
assign n2051 = /* LUT   18 23  2 */ (n105 ? (n1518 ? 1'b1 : (n701 ? 1'b1 : n1492)) : (n1518 ? 1'b1 : n1492));
assign n2052 = /* LUT    6 20  2 */ (n409 ? n695 : (n695 ? (n410 ? !n317 : 1'b0) : 1'b0));
assign n597  = /* LUT    5 20  1 */ (n474 ? !n473 : (n473 ? n320 : 1'b1));
assign n2054 = /* LUT   10 29  2 */ (n130 ? n874 : n872);
assign n2055 = /* LUT   15 27  6 */ (n130 ? n781 : n338);
assign n2056 = /* LUT   15 22  5 */ (io_33_1_1 ? 1'b0 : \wb_dat_i[8] );
assign n2057 = /* LUT    7 26  3 */ (n130 ? (n376 ? 1'b0 : !n620) : (n376 ? !n414 : !n620));
assign n898  = /* LUT    9 19  3 */ (n802 ? (n795 ? 1'b1 : n75) : (n800 ? (n795 ? 1'b1 : n75) : (n795 ? !n75 : 1'b0)));
assign n1230 = /* LUT   12 19  4 */ (n893 ? (n892 ? (n990 ? !n1228 : 1'b1) : !n1228) : (n892 ? !n990 : 1'b0));
assign n1251 = /* LUT   12 24  5 */ (n1100 ? (n955 ? 1'b1 : !n666) : (n955 ? n666 : 1'b0));
assign n1499 = /* LUT   17 23  0 */ (n1029 ? (n877 ? (n512 ? 1'b1 : n708) : n512) : (n877 ? n708 : 1'b0));
assign n2062 = /* LUT    4 18  1 */ (n263 ? (io_33_1_1 ? 1'b0 : n356) : (n53 ? 1'b0 : (io_33_1_1 ? 1'b0 : n356)));
assign n2063 = /* LUT    9 29  4 */ (n130 ? n964 : n779);
assign n2064 = /* LUT   13 23  7 */ (n666 ? n1068 : n948);
assign n2065 = /* LUT    7 23  7 */ (io_33_13_0 ? !io_33_1_1 : 1'b0);
assign n2066 = /* LUT   11 30  1 */ (n130 ? n966 : n847);
assign n2067 = /* LUT   13 20  3 */ (io_33_1_1 ? 1'b0 : \wb_dat_i[5] );
assign n2068 = /* LUT   12 28  2 */ (n849 ? (n850 ? 1'b1 : n130) : (n850 ? !n130 : 1'b0));
assign n2069 = /* LUT   17 19  5 */ (n101 ? (n286 ? (n1447 ? 1'b1 : \wb_adr_i[5] ) : \wb_adr_i[5] ) : (n286 ? n1447 : 1'b0));
assign n2070 = /* LUT    5 21  2 */ (n500 ? (n605 ? 1'b1 : !n499) : (n605 ? 1'b1 : (n501 ? !n499 : 1'b0)));
assign n2071 = /* LUT   10 28  1 */ (n962 ? (n547 ? 1'b1 : n130) : (n547 ? !n130 : 1'b0));
assign n770  = /* LUT    7 27  0 */ (n376 ? (n316 ? 1'b0 : !n130) : !n626);
assign n2073 = /* LUT   12 18  7 */ (n1226 ? n887 : !n887);
assign n2074 = /* LUT   12 31  4 */ (n1211 ? (n1283 ? n286 : (n286 ? !n675 : 1'b0)) : (n1283 ? (n286 ? n675 : 1'b0) : 1'b0));
assign n2075 = /* LUT   12 32  1 */ (n1218 ? (n1284 ? 1'b1 : !n677) : (n1284 ? n677 : 1'b0));
assign n2076 = /* LUT   16 24  0 */ (n1299 ? (n1317 ? 1'b1 : n677) : (n1317 ? !n677 : 1'b0));
assign n2077 = /* LUT    9 30  5 */ (n234 ? (n780 ? 1'b1 : n130) : (n780 ? !n130 : 1'b0));
assign n2078 = /* LUT   13 24  6 */ (n130 ? n538 : n635);
assign n2079 = /* LUT    7 20  6 */ (io_33_15_1 ? !io_33_1_1 : 1'b0);
assign n2080 = /* LUT   11 31  2 */ (n1079 ? (n1216 ? 1'b1 : n677) : (n1216 ? !n677 : 1'b0));
assign n2081 = /* LUT   16 22  1 */ (n1115 ? (n1458 ? 1'b1 : (n758 ? 1'b1 : n1399)) : (n1458 ? 1'b1 : n1399));
assign n2082 = /* LUT    6 22  4 */ (\wb_adr_i[5]  ? (n17 ? 1'b0 : n596) : 1'b0);
assign n2083 = /* LUT   17 28  4 */ (n675 ? (n286 ? n1374 : 1'b0) : (n1508 ? n286 : 1'b0));
assign n2084 = /* LUT    5 22  3 */ (n473 ? !io_33_1_1 : 1'b0);
assign n2085 = /* LUT   10 31  0 */ (n987 ? (n981 ? 1'b1 : n666) : (n981 ? !n666 : 1'b0));
assign n1417 = /* LUT   15 25  0 */ (n1361 ? (n675 ? (n1363 ? n286 : 1'b0) : n286) : (n675 ? (n1363 ? n286 : 1'b0) : 1'b0));
assign n2087 = /* LUT    3  7  7 */ (io_0_4_1 ? io_0_3_0 : 1'b0);
assign n2088 = /* LUT   15 20  7 */ (\dd_pad_i[12]  ? !io_33_1_1 : 1'b0);
assign n2089 = /* LUT    7 24  1 */ (n118 ? 1'b0 : (n709 ? (n408 ? n686 : 1'b1) : (n408 ? n686 : 1'b0)));
assign n2090 = /* LUT   12 17  6 */ (\wb_dat_i[11]  ? 1'b1 : io_33_1_1);
assign n2091 = /* LUT   12 30  7 */ (n130 ? n847 : n966);
assign n2092 = /* LUT   13 25  5 */ n780;
assign n2093 = /* LUT   14 29  2 */ (n978 ? (n1105 ? 1'b1 : n130) : (n1105 ? !n130 : 1'b0));
assign n2094 = /* LUT   11 28  3 */ (n130 ? n1105 : n978);
assign n2095 = /* LUT   16 21  0 */ (io_33_1_1 ? 1'b0 : \dd_pad_i[12] );
assign n1291 = /* LUT   13 22  1 */ (n677 ? n134 : n1240);
assign n2097 = /* LUT    3 22  3 */ (n202 ? 1'b1 : (n404 ? 1'b1 : io_33_1_1));
assign n2098 = /* LUT    6 17  5 */ (n672 ? (io_33_1_1 ? !n450 : (n353 ? 1'b1 : !n450)) : (io_33_1_1 ? 1'b0 : (n353 ? n450 : 1'b0)));
assign n2099 = /* LUT    4 20  4 */ (n494 ? (n391 ? n67 : !n67) : (n391 ? !n67 : n67));
assign n2100 = /* LUT    7 18  7 */ (n484 ? (n488 ? (n388 ? 1'b1 : n505) : n505) : 1'b0);
assign n2101 = /* LUT    9 27  7 */ (n720 ? (n764 ? 1'b1 : !n130) : (n764 ? n130 : 1'b0));
assign n2102 = /* LUT    7 25  6 */ (n706 ? 1'b1 : (n766 ? 1'b1 : io_33_1_1));
assign n2103 = /* LUT   12 16  1 */ (io_33_1_1 ? 1'b0 : \wb_dat_i[4] );
assign n2104 = /* LUT   14 18  0 */ (io_33_1_1 ? 1'b1 : \wb_adr_i[4] );
assign n2105 = /* LUT   12 29  6 */ (n1202 ? (n853 ? 1'b1 : !n666) : (n853 ? n666 : 1'b0));
assign n2106 = /* LUT    4 26  5 */ (io_33_15_1 ? !n118 : 1'b0);
assign n2107 = /* LUT    4 23  6 */ (n1 ? (n173 ? 1'b0 : !io_33_1_1) : 1'b0);
assign n2108 = /* LUT    9 24  3 */ n828;
assign n2109 = /* LUT   13 26  4 */ (n130 ? \dd_pad_i[3]  : \dd_pad_i[10] );
assign n1377 = /* LUT   14 28  1 */ (n666 ? n659 : n1201);
assign n2111 = /* LUT    2 22  4 */ (n169 ? n303 : n272);
assign n2112 = /* LUT   11 22  5 */ (n675 ? !n677 : n677);
assign n2113 = /* LUT   11 29  4 */ (n636 ? (n634 ? 1'b1 : n130) : (n634 ? !n130 : 1'b0));
assign n2114 = /* LUT   15 18  4 */ (\wb_dat_i[19]  ? 1'b1 : io_33_1_1);
assign n2115 = /* LUT    3 23  0 */ (n390 ? (n287 ? !n307 : 1'b0) : (n287 ? !n307 : (n77 ? 1'b0 : !n307)));
assign n2116 = /* LUT    2 21  6 */ (n294 ? (n67 ? n269 : !n269) : (n67 ? !n269 : n269));
assign n2117 = /* LUT    7 29  3 */ (n675 ? (n777 ? n286 : 1'b0) : (n136 ? n286 : 1'b0));
assign n2118 = /* LUT   12 20  6 */ (\dd_pad_i[7]  ? !io_33_1_1 : 1'b0);
assign n754  = /* LUT    7 19  4 */ (n675 ? (n698 ? (n677 ? !n693 : n693) : 1'b1) : (n698 ? 1'b1 : (n677 ? !n693 : n693)));
assign n2120 = /* LUT    9 20  6 */ \wb_dat_i[22] ;
assign n2121 = /* LUT    3 24  6 */ (n118 ? 1'b0 : \wb_adr_i[4] );
assign n1243 = /* LUT   12 23  0 */ (n1153 ? (n286 ? (n1152 ? 1'b1 : \wb_adr_i[5] ) : \wb_adr_i[5] ) : (n286 ? n1152 : 1'b0));
assign n2123 = /* LUT   11 25  1 */ (n130 ? n849 : n850);
assign n2124 = /* LUT    4 25  4 */ \wb_dat_i[4] ;
assign n2125 = /* LUT    4 22  5 */ (n377 ? 1'b0 : (n516 ? (io_31_0_1 ? 1'b0 : !n511) : 1'b0));
assign n2126 = /* LUT    9 25  0 */ (n666 ? n842 : n831);
assign n2127 = /* LUT   13 27  3 */ (n130 ? n1105 : n978);
assign n2128 = /* LUT    6 28  3 */ (n75 ? n529 : n583);
assign n2129 = /* LUT   11 23  6 */ (n677 ? n1157 : n936);
assign n2130 = /* LUT   11 26  5 */ (n827 ? (n828 ? 1'b1 : !n130) : (n828 ? n130 : 1'b0));
assign n2131 = /* LUT    2 20  5 */ (n276 ? (n174 ? 1'b1 : io_33_1_1) : 1'b1);
assign n2132 = /* LUT   12 27  7 */ (n130 ? n847 : n966);
assign n2133 = /* LUT    6 19  7 */ wb_clk_i;
assign n2134 = /* LUT   15 28  3 */ (n1210 ? (n1433 ? 1'b1 : n677) : (n1433 ? !n677 : 1'b0));
assign n2135 = /* LUT    9 21  5 */ (n471 ? n169 : (n909 ? n438 : n169));
assign n2136 = /* LUT    7 31  4 */ (n130 ? n131 : n337);
assign n2137 = /* LUT   12 22  3 */ (n610 ? (n600 ? (n701 ? 1'b1 : n708) : n701) : (n600 ? n708 : 1'b0));
assign n2138 = /* LUT    4 24  3 */ (n118 ? 1'b0 : io_33_5_0);
assign n2139 = /* LUT    4 21  4 */ (n374 ? (io_33_1_1 ? !n300 : (n400 ? 1'b1 : !n300)) : (io_33_1_1 ? 1'b0 : (n400 ? n300 : 1'b0)));
assign n956  = /* LUT    9 26  1 */ (n130 ? (n619 ? 1'b0 : !n376) : (n619 ? (n376 ? !n416 : 1'b0) : (n376 ? !n416 : 1'b1)));
assign n1319 = /* LUT   13 28  2 */ (n677 ? n1264 : n1318);
assign n2142 = /* LUT    2 24  6 */ (n326 ? (n210 ? n67 : !n67) : (n210 ? !n67 : n67));
assign n2143 = /* LUT   11 20  7 */ (n1135 ? (n905 ? 1'b0 : n893) : (n892 ? 1'b1 : (n905 ? 1'b0 : n893)));
assign n2144 = /* LUT   17 27  6 */ (n675 ? (\wb_adr_i[3]  ? !n1325 : 1'b0) : (n1380 ? 1'b0 : \wb_adr_i[3] ));
assign n2145 = /* LUT   11 27  6 */ (n130 ? n633 : n526);
assign n2146 = /* LUT    3 21  6 */ (n317 ? (io_33_1_1 ? 1'b0 : (n392 ? n276 : 1'b0)) : !io_33_1_1);
assign n2147 = /* LUT    2 23  4 */ (n213 ? (io_33_1_1 ? !n205 : (n205 ? n114 : 1'b1)) : (io_33_1_1 ? 1'b0 : (n205 ? n114 : 1'b0)));
assign n2148 = /* LUT   12 26  4 */ (n130 ? n874 : n872);
assign n1502 = /* LUT   17 24  0 */ (n228 ? (\wb_adr_i[5]  ? (n96 ? 1'b1 : n1465) : n96) : (\wb_adr_i[5]  ? n1465 : 1'b0));
assign n2150 = /* LUT    7 17  2 */ (n740 ? (n67 ? n568 : !n568) : (n67 ? !n568 : n568));
assign n2151 = /* LUT    9 22  4 */ (n675 ? (n924 ? n286 : 1'b0) : (n286 ? n812 : 1'b0));
assign n2152 = /* LUT    7 28  5 */ (n643 ? (n719 ? 1'b1 : !n130) : (n719 ? n130 : 1'b0));
assign n2153 = /* LUT   14 26  4 */ (n130 ? DMA_req : iordy_pad_i);
assign n2154 = /* LUT   12 21  2 */ (io_33_1_1 ? 1'b0 : \wb_dat_i[14] );
assign n2155 = /* LUT   19 20  0 */ (io_33_1_1 ? 1'b0 : io_33_19_0);
assign n2156 = /* LUT   13 29  1 */ (n130 ? n769 : n968);
assign n2157 = /* LUT   12 11  1 */ (io_33_1_1 ? 1'b0 : \wb_dat_i[0] );
assign n1366 = /* LUT   14 25  6 */ (n1300 ? (n1365 ? 1'b1 : n677) : (n1365 ? !n677 : 1'b0));
assign n2159 = /* LUT    3 17  3 */ (n146 ? (io_33_1_1 ? !n254 : (n246 ? 1'b1 : !n254)) : (io_33_1_1 ? 1'b0 : (n246 ? n254 : 1'b0)));
assign n2160 = /* LUT    6 21  4 */ (n169 ? n691 : n689);
assign n2161 = /* LUT   11 24  7 */ (n1072 ? (n1064 ? 1'b1 : n666) : (n1064 ? !n666 : 1'b0));
assign n2162 = /* LUT   15 17  1 */ (\dd_pad_i[12]  ? !io_33_1_1 : 1'b0);
assign n2163 = /* LUT    7 21  7 */ (io_33_1_1 ? 1'b0 : \wb_dat_i[5] );
assign n2164 = /* LUT    3 18  7 */ (n349 ? 1'b1 : (n356 ? 1'b0 : !n53));
assign n2165 = /* LUT   12 25  5 */ (n135 ? (n715 ? 1'b1 : n666) : (n715 ? !n666 : 1'b0));
assign n565  = /* LUT    5 16  1 */ (n239 ? 1'b1 : (n564 ? 1'b1 : (n241 ? 1'b1 : n242)));
assign n2167 = /* LUT   10 25  2 */ (n850 ? (n849 ? 1'b1 : n130) : (n849 ? !n130 : 1'b0));
assign n2168 = /* LUT    9 23  3 */ (n933 ? (n830 ? 1'b1 : !n666) : (n830 ? n666 : 1'b0));
assign n2169 = /* LUT   14 21  5 */ (io_33_1_1 ? 1'b0 : \wb_dat_i[23] );
assign n2170 = /* LUT    6 26  2 */ (n522 ? !n629 : (n130 ? (n629 ? 1'b0 : !n376) : !n629));
assign n2171 = /* LUT   11 17  5 */ (n891 ? !n1117 : (n1117 ? 1'b0 : !n893));
assign n2172 = /* LUT   15 21  6 */ (n1285 ? (n1227 ? (n1038 ? 1'b0 : n1338) : 1'b1) : (n1038 ? 1'b0 : n1338));
assign n2173 = /* LUT   13 30  0 */ (n1209 ? (n1191 ? 1'b1 : !n666) : (n1191 ? n666 : 1'b0));
assign n2174 = /* LUT   14 24  5 */ (n677 ? n1087 : n1357);
assign n2175 = /* LUT    6 20  7 */ (n257 ? 1'b1 : (n696 ? (n171 ? 1'b1 : !n395) : 1'b0));
assign n2176 = /* LUT    6 25  4 */ (n376 ? (n519 ? 1'b0 : !n130) : !n542);
assign n2177 = /* LUT   11 18  1 */ (n893 ? (n1122 ? 1'b0 : n1120) : !n1122);
assign n2178 = /* LUT   10 22  0 */ (n913 ? (io_33_1_1 ? 1'b0 : (n287 ? 1'b1 : n637)) : (io_33_1_1 ? 1'b0 : (n287 ? 1'b0 : n637)));
assign n2179 = /* LUT   15 22  0 */ (io_33_1_1 ? 1'b0 : \wb_dat_i[23] );
assign n2180 = /* LUT    3 19  4 */ (n366 ? (n36 ? (io_33_1_1 ? !n254 : 1'b1) : (io_33_1_1 ? 1'b0 : n254)) : (n36 ? !n254 : 1'b0));
assign n1250 = /* LUT   12 24  2 */ (n666 ? n1109 : n1085);
assign n2182 = /* LUT    5 17  2 */ io_33_9_0;
assign n2183 = /* LUT   10 24  1 */ (n130 ? n337 : n131);
assign n2184 = /* LUT    7 23  0 */ (io_33_5_0 ? 1'b1 : io_33_1_1);
assign n2185 = /* LUT   11 30  4 */ (n636 ? (n634 ? 1'b1 : n130) : (n634 ? !n130 : 1'b0));
assign n1476 = /* LUT   16 28  0 */ (n89 ? n708 : 1'b0);
assign n1516 = /* LUT   18 22  2 */ (n747 ? n512 : 1'b0);
assign n2188 = /* LUT   14 27  4 */ (n130 ? n1105 : n978);
assign n2189 = /* LUT   12 28  7 */ (n960 ? (n974 ? 1'b1 : !n666) : (n974 ? n666 : 1'b0));
assign n2190 = /* LUT    6 24  7 */ (n518 ? (n522 ? 1'b1 : n130) : (n522 ? !n130 : 1'b0));
assign n1132 = /* LUT   11 19  2 */ (n387 ? (n902 ? 1'b0 : n893) : (n892 ? 1'b1 : (n902 ? 1'b0 : n893)));
assign n2192 = /* LUT   13 17  0 */ (io_33_1_1 ? 1'b0 : \wb_dat_i[30] );
assign n2193 = /* LUT   15 23  3 */ (\wb_dat_i[23]  ? !io_33_1_1 : 1'b0);
assign n2194 = /* LUT    7 27  5 */ (n710 ? (n709 ? (n408 ? !n686 : 1'b0) : 1'b0) : 1'b0);
assign n2195 = /* LUT   18 21  4 */ (n1455 ? (n1515 ? 1'b1 : (n104 ? n1135 : 1'b0)) : (n104 ? n1135 : 1'b0));
assign n1283 = /* LUT   12 31  3 */ (n677 ? n1214 : n1282);
assign n2197 = /* LUT    5 18  3 */ (n458 ? io_33_1_1 : n578);
assign n2198 = /* LUT   10 27  0 */ (n96 ? (n517 ? 1'b1 : io_33_1_1) : io_33_1_1);
assign n2199 = /* LUT    7 20  1 */ (io_33_1_1 ? 1'b0 : io_33_9_0);
assign n2200 = /* LUT    9 17  1 */ (n787 ? 1'b0 : (n788 ? 1'b1 : !n798));
assign n2201 = /* LUT   14 23  7 */ (io_33_1_1 ? 1'b0 : \wb_dat_i[0] );
assign n2202 = /* LUT   17 21  2 */ (n1337 ? (n285 ? (n1485 ? 1'b1 : !io_33_7_0) : n1485) : n1485);
assign n2203 = /* LUT    1 18  5 */ (n160 ? (n67 ? n57 : !n57) : (n67 ? !n57 : n57));
assign n2204 = /* LUT   11 31  7 */ (n130 ? n849 : n850);
assign n2205 = /* LUT   16 27  1 */ (n130 ? n1105 : n978);
assign n704  = /* LUT    6 22  1 */ (wb_stb_i ? (io_0_6_0 ? 1'b1 : \wb_adr_i[5] ) : \wb_adr_i[5] );
assign n2206 = /* LUT    6 27  6 */ (n130 ? (n724 ? 1'b0 : (n376 ? n129 : 1'b1)) : !n724);
assign n2207 = /* LUT   11 16  3 */ (io_33_17_0 ? !io_33_1_1 : 1'b0);
assign n2208 = /* LUT    9 13  7 */ (n169 ? n398 : n877);
assign n2209 = /* LUT   15 20  2 */ (io_33_1_1 ? 1'b0 : \wb_dat_i[24] );
assign n2210 = /* LUT    7 24  4 */ (n709 ? (n408 ? !n118 : (n710 ? !n118 : 1'b0)) : (n408 ? 1'b0 : (n710 ? !n118 : 1'b0)));
assign n2211 = /* LUT   18 20  7 */ (io_33_8_0 ? 1'b0 : (n1337 ? io_33_7_0 : 1'b0));
assign n2212 = /* LUT   12 30  0 */ (n1189 ? (n1205 ? 1'b1 : n666) : (n1205 ? !n666 : 1'b0));
assign n2213 = /* LUT    5 24  5 */ (io_33_16_1 ? !n118 : 1'b0);
assign n590  = /* LUT    5 19  4 */ (n259 ? 1'b1 : n154);
assign n2214 = /* LUT   10 26  7 */ (n719 ? (n643 ? 1'b1 : !n130) : (n643 ? n130 : 1'b0));
assign n2215 = /* LUT   15 26  1 */ (n1188 ? (n666 ? 1'b1 : n1248) : (n666 ? 1'b0 : n1248));
assign n2216 = /* LUT    9 18  0 */ (n667 ? (io_33_1_1 ? !n450 : (n450 ? n797 : 1'b1)) : (io_33_1_1 ? 1'b0 : (n450 ? n797 : 1'b0)));
assign n1343 = /* LUT   14 22  0 */ (n677 ? n727 : n939);
assign n2218 = /* LUT    6 18  6 */ (n460 ? (io_33_1_1 ? 1'b1 : n681) : n680);
assign n2219 = /* LUT   17 22  3 */ (\wb_dat_i[27]  ? !io_33_1_1 : 1'b0);
assign n2220 = /* LUT   11 28  6 */ (n872 ? (n874 ? 1'b1 : n130) : (n874 ? !n130 : 1'b0));
assign n2221 = /* LUT    9 28  3 */ (n827 ? (n828 ? 1'b1 : !n130) : (n828 ? n130 : 1'b0));
assign n2222 = /* LUT    3 22  6 */ (n296 ? n406 : io_33_1_1);
assign n2223 = /* LUT   10 30  4 */ (n130 ? n964 : n779);
assign n2224 = /* LUT   13 19  6 */ (io_33_1_1 ? 1'b0 : io_33_15_1);
assign n2225 = /* LUT    7 25  3 */ (n666 ? n537 : n713);
assign n2226 = /* LUT   14 18  5 */ (io_33_1_1 ? 1'b1 : \wb_dat_i[20] );
assign n2227 = /* LUT   12 29  1 */ (n769 ? (n968 ? 1'b1 : !n130) : (n968 ? n130 : 1'b0));
assign n2228 = /* LUT    1 20  6 */ (n58 ? !n67 : n67);
assign n2229 = /* LUT    5 20  5 */ (n484 ? (n505 ? 1'b0 : (n509 ? 1'b0 : n388)) : 1'b0);
assign n2230 = /* LUT   10 29  6 */ (n130 ? n719 : n643);
assign n2231 = /* LUT   15 27  2 */ (n130 ? n779 : n964);
assign n2232 = /* LUT   12 19  0 */ (n1024 ? 1'b0 : (n1115 ? 1'b1 : !n798));
assign n2233 = /* LUT   14 17  1 */ (io_33_9_0 ? !io_33_1_1 : 1'b0);
assign n2234 = /* LUT    6 29  7 */ (n556 ? (io_33_1_1 ? 1'b0 : (n287 ? 1'b1 : n647)) : (io_33_1_1 ? 1'b0 : (n287 ? 1'b0 : n647)));
assign n2235 = /* LUT   11 29  1 */ (n130 ? n847 : n966);
assign n2236 = /* LUT   16 25  3 */ (n666 ? n1255 : n1308);
assign n2237 = /* LUT    9 29  0 */ (n130 ? n234 : n780);
assign n2238 = /* LUT   13 23  3 */ (n169 ? n1167 : n1290);
assign n413  = /* LUT    3 23  5 */ (n75 ? n364 : n48);
assign n2240 = /* LUT    1 27  4 */ \wb_dat_o[5] ;
assign n1000 = /* LUT   10 17  5 */ (n892 ? (n994 ? !n991 : (n893 ? 1'b1 : !n991)) : (n994 ? 1'b0 : n893));
assign n2242 = /* LUT   13 20  7 */ (io_33_1_1 ? 1'b0 : \wb_dat_i[25] );
assign n2243 = /* LUT    3 24  1 */ (\wb_dat_i[14]  ? !n118 : 1'b0);
assign n2244 = /* LUT    1 21  5 */ n24;
assign n2245 = /* LUT   17 19  1 */ (n1120 ? (n691 ? (n701 ? 1'b1 : n512) : n512) : (n691 ? n701 : 1'b0));
assign n2246 = /* LUT    5 26  7 */ \wb_dat_i[4] ;
assign n2247 = /* LUT   11 25  6 */ (n338 ? (n781 ? 1'b1 : n130) : (n781 ? !n130 : 1'b0));
assign n2248 = /* LUT    5 21  6 */ (n473 ? (n509 ? !n474 : 1'b0) : (n509 ? !n474 : 1'b1));
assign n2249 = /* LUT   10 28  5 */ (n968 ? (n769 ? 1'b1 : !n130) : (n769 ? n130 : 1'b0));
assign n1412 = /* LUT   15 24  3 */ (n666 ? n1073 : n1177);
assign n2251 = /* LUT   12 18  3 */ (n1222 ? (n67 ? n261 : !n261) : (n67 ? !n261 : n261));
assign n2252 = /* LUT   11 26  0 */ (n130 ? n337 : n131);
assign n2253 = /* LUT    9 30  1 */ (n538 ? (n635 ? 1'b1 : !n130) : (n635 ? n130 : 1'b0));
assign n2254 = /* LUT   13 24  2 */ (n130 ? n636 : n634);
assign n2255 = /* LUT    3 20  4 */ (n163 ? (io_33_1_1 ? 1'b0 : n378) : n188);
assign n2256 = /* LUT   12 13  7 */ (io_33_1_1 ? 1'b0 : \wb_adr_i[4] );
assign n2257 = /* LUT   18 26  6 */ (n1468 ? (n649 ? 1'b1 : !n677) : (n649 ? n677 : 1'b0));
assign n2258 = /* LUT    6 19  2 */ \wb_adr_i[4] ;
assign n2259 = /* LUT   10 16  6 */ (io_33_5_0 ? !io_33_1_1 : 1'b0);
assign n2260 = /* LUT    1 22  4 */ (io_33_1_1 ? 1'b0 : \wb_dat_i[20] );
assign n2261 = /* LUT   17 28  0 */ (\wb_adr_i[5]  ? (n96 ? (n1467 ? 1'b1 : n707) : n1467) : (n96 ? n707 : 1'b0));
assign n2262 = /* LUT    5 27  0 */ (n130 ? n425 : n129);
assign n2263 = /* LUT    5 22  7 */ (n394 ? 1'b0 : (n181 ? 1'b1 : (n511 ? n317 : 1'b0)));
assign n2264 = /* LUT   10 31  4 */ (n984 ? (n972 ? 1'b1 : !n666) : (n972 ? n666 : 1'b0));
assign n2265 = /* LUT   15 25  4 */ (n1204 ? (n1178 ? 1'b1 : !n677) : (n1178 ? n677 : 1'b0));
assign n2266 = /* LUT   12 17  2 */ (io_33_17_0 ? !io_33_1_1 : 1'b0);
assign n2267 = /* LUT   14 19  3 */ (io_33_15_1 ? !io_33_1_1 : 1'b0);
assign n2268 = /* LUT   11 27  3 */ (n966 ? (n847 ? 1'b1 : n130) : (n847 ? !n130 : 1'b0));
assign n2269 = /* LUT    4 27  2 */ (n287 ? (n549 ? !io_33_1_1 : 1'b0) : (n230 ? !io_33_1_1 : 1'b0));
assign n2270 = /* LUT    9 31  6 */ (n130 ? n633 : n526);
assign n2271 = /* LUT   13 25  1 */ n850;
assign n2272 = /* LUT    3 21  3 */ (n276 ? (io_33_1_1 ? 1'b0 : (n317 ? 1'b1 : n301)) : (io_33_1_1 ? 1'b0 : n317));
assign n2273 = /* LUT   13 22  5 */ (n708 ? (n790 ? (n1290 ? 1'b1 : n512) : n1290) : (n790 ? n512 : 1'b0));
assign n2274 = /* LUT    7 28  0 */ (n666 ? n731 : n725);
assign n2278 = /* LUT    7 18  3 */ (n678 ? (n684 ? (n118 ? 1'b1 : n675) : 1'b1) : (n684 ? (n118 ? 1'b1 : n675) : n118));
assign n2279 = /* LUT    9 27  3 */ (n964 ? (n779 ? 1'b1 : !n130) : (n779 ? n130 : 1'b0));
assign n2280 = /* LUT   12 16  5 */ (io_33_1_1 ? 1'b0 : io_33_13_0);
assign n2281 = /* LUT   11 24  2 */ (n780 ? (n234 ? 1'b1 : n130) : (n234 ? !n130 : 1'b0));
assign n2282 = /* LUT    4 26  1 */ (\wb_dat_i[19]  ? !n118 : 1'b0);
assign n2283 = /* LUT   21 22  6 */ (n1137 ? (n1004 ? 1'b0 : n1285) : (n1004 ? n1338 : (n1285 ? 1'b1 : n1338)));
assign n2284 = /* LUT   13 26  0 */ (n130 ? \dd_pad_i[15]  : \dd_pad_i[5] );
assign n2285 = /* LUT    3 18  2 */ (n33 ? (n359 ? (n168 ? 1'b1 : io_33_1_1) : 1'b1) : (n359 ? (n168 ? 1'b1 : io_33_1_1) : 1'b0));
assign n2286 = /* LUT    2 22  0 */ (n169 ? n107 : n92);
assign n2287 = /* LUT   11 22  1 */ (n1052 ? 1'b0 : (n1149 ? 1'b0 : (n1146 ? 1'b0 : !n817)));
assign n2288 = /* LUT    5 16  4 */ (n472 ? (io_33_1_1 ? 1'b0 : n447) : (n449 ? (io_33_1_1 ? 1'b0 : n447) : 1'b0));
assign n2289 = /* LUT   10 18  0 */ (n460 ? (io_33_1_1 ? 1'b0 : n996) : n786);
assign n2290 = /* LUT    6 26  7 */ (n632 ? 1'b0 : (n222 ? 1'b1 : (n376 ? !n130 : 1'b1)));
assign n2291 = /* LUT    5 29  2 */ (n648 ? (n660 ? !io_33_1_1 : (io_33_1_1 ? 1'b0 : !n287)) : (n660 ? (io_33_1_1 ? 1'b0 : n287) : 1'b0));
assign n2292 = /* LUT    7 19  0 */ \dd_pad_i[5] ;
assign n2293 = /* LUT    9 20  2 */ io_33_8_0;
assign n2294 = /* LUT   12 23  4 */ (n1154 ? (n1244 ? 1'b1 : n675) : (n1244 ? !n675 : 1'b0));
assign n2295 = /* LUT    4 25  0 */ \wb_dat_i[5] ;
assign n2296 = /* LUT   10 22  5 */ (n639 ? (n1055 ? !io_33_1_1 : (io_33_1_1 ? 1'b0 : !n287)) : (n1055 ? (io_33_1_1 ? 1'b0 : n287) : 1'b0));
assign n2297 = /* LUT    9 25  4 */ (n720 ? (n764 ? 1'b1 : !n130) : (n764 ? n130 : 1'b0));
assign n2298 = /* LUT   13 27  7 */ (n130 ? n874 : n872);
assign n2299 = /* LUT    3 19  1 */ (n260 ? n67 : n367);
assign n1162 = /* LUT   11 23  2 */ (n1056 ? (n1161 ? (n286 ? 1'b1 : \wb_adr_i[5] ) : \wb_adr_i[5] ) : (n1161 ? n286 : 1'b0));
assign n2301 = /* LUT   10 21  1 */ (n1045 ? !n1047 : (n1047 ? 1'b0 : !n798));
assign n2302 = /* LUT   15 19  3 */ (n758 ? (n1390 ? 1'b1 : (n1333 ? 1'b1 : n993)) : (n1390 ? 1'b1 : n1333));
assign n2303 = /* LUT   12 27  3 */ (n130 ? n635 : n538);
assign n2304 = /* LUT   15 28  7 */ (n1271 ? (n1382 ? 1'b1 : !n675) : (n1382 ? n675 : 1'b0));
assign n2305 = /* LUT    9 21  1 */ (n758 ? (n685 ? 1'b1 : (n701 ? n650 : 1'b0)) : (n701 ? n650 : 1'b0));
assign n2306 = /* LUT   13 31  4 */ (n677 ? n1332 : n1279);
assign n2307 = /* LUT   18 22  7 */ (n92 ? (n1517 ? (n1302 ? 1'b1 : n708) : n708) : (n1517 ? n1302 : 1'b0));
assign n2308 = /* LUT    6 24  0 */ (n130 ? n414 : n315);
assign n2309 = /* LUT    4 24  7 */ (n118 ? 1'b0 : io_33_9_0);
assign n2310 = /* LUT    9 26  5 */ (n130 ? (n621 ? 1'b0 : !n376) : (n621 ? (n376 ? !n418 : 1'b0) : (n376 ? !n418 : 1'b1)));
assign n2311 = /* LUT   13 28  6 */ (n634 ? (n636 ? 1'b1 : n130) : (n636 ? !n130 : 1'b0));
assign n1515 = /* LUT   18 21  3 */ (\wb_dat_i[2]  ? 1'b0 : (n1514 ? (io_33_8_0 ? 1'b0 : !io_33_7_0) : 1'b0));
assign n2312 = /* LUT    2 24  2 */ (n322 ? (n206 ? n67 : !n67) : (n206 ? !n67 : n67));
assign n2313 = /* LUT   11 20  3 */ (n798 ? (n1140 ? 1'b0 : n1040) : !n1140);
assign n2314 = /* LUT    5 18  6 */ (n264 ? !n344 : 1'b0);
assign n2315 = /* LUT   12 26  0 */ (n969 ? (n1179 ? 1'b1 : n666) : (n1179 ? !n666 : 1'b0));
assign n2316 = /* LUT   17 21  7 */ (\wb_dat_i[2]  ? 1'b0 : (io_33_8_0 ? (io_33_7_0 ? n1486 : 1'b0) : 1'b0));
assign n2320 = /* LUT   17 24  4 */ (n286 ? (n1503 ? (n1409 ? 1'b1 : !n675) : (n1409 ? n675 : 1'b0)) : 1'b0);
assign n2321 = /* LUT    4 28  4 */ (n437 ? (io_33_1_1 ? 1'b0 : (n287 ? 1'b1 : n233)) : (io_33_1_1 ? 1'b0 : (n287 ? 1'b0 : n233)));
assign n2322 = /* LUT    7 17  6 */ (n744 ? (n67 ? n572 : !n572) : (n67 ? !n572 : n572));
assign n922  = /* LUT    9 22  0 */ (n514 ? (\wb_adr_i[5]  ? (n96 ? 1'b1 : n813) : n96) : (\wb_adr_i[5]  ? n813 : 1'b0));
assign n2324 = /* LUT   14 26  0 */ (n130 ? wb_cyc_i : \wb_sel_i[1] );
assign n722  = /* LUT    6 27  1 */ (n430 ? (n376 ? 1'b0 : !n623) : (n376 ? !n130 : !n623));
assign n2326 = /* LUT    9 32  6 */ (n279 ? 1'b1 : (n809 ? 1'b1 : (n808 ? 1'b1 : n988)));
assign n1511 = /* LUT   18 20  0 */ (io_33_7_0 ? 1'b0 : (io_33_8_0 ? 1'b0 : (n1478 ? n1486 : 1'b0)));
assign n2328 = /* LUT    6 21  0 */ (n603 ? (n697 ? (n701 ? 1'b1 : n512) : n512) : (n697 ? n701 : 1'b0));
assign n2329 = /* LUT   11 21  4 */ (n907 ? (n991 ? (n104 ? 1'b1 : n96) : n96) : (n991 ? n104 : 1'b0));
assign n2330 = /* LUT    5 19  1 */ (n587 ? (n270 ? 1'b1 : n75) : (n270 ? !n75 : 1'b0));
assign n1058 = /* LUT   10 23  3 */ (n666 ? n858 : n920);
assign n2332 = /* LUT   15 26  4 */ (io_33_1_1 ? 1'b0 : \wb_dat_i[18] );
assign n2333 = /* LUT    7 21  3 */ (io_33_1_1 ? 1'b0 : \dd_pad_i[2] );
assign n2334 = /* LUT   12 25  1 */ (n131 ? (n337 ? 1'b1 : !n130) : (n337 ? n130 : 1'b0));
assign n481  = /* LUT    4 19  5 */ (n452 ? (n480 ? (n458 ? 1'b1 : n273) : 1'b1) : 1'b1);
assign n2336 = /* LUT    9 28  6 */ (n130 ? n720 : n764);
assign n2337 = /* LUT   18 24  5 */ (n1461 ? (n1521 ? (n286 ? 1'b1 : \wb_adr_i[5] ) : \wb_adr_i[5] ) : (n1521 ? n286 : 1'b0));
assign n2338 = /* LUT   14 21  1 */ (\wb_dat_i[25]  ? !io_33_1_1 : 1'b0);
assign n2339 = /* LUT   11 17  1 */ (n798 ? (n1116 ? 1'b0 : n789) : !n1116);
assign n2340 = /* LUT   13 19  3 */ (\wb_dat_i[22]  ? !io_33_1_1 : 1'b0);
assign n2341 = /* LUT   15 21  2 */ (n1045 ? (n1046 ? 1'b0 : n1338) : (n1046 ? n1285 : (n1285 ? 1'b1 : n1338)));
assign n1329 = /* LUT   13 30  4 */ (n677 ? n1274 : n1328);
assign n2343 = /* LUT    2 17  5 */ (n251 ? (n67 ? n243 : !n243) : (n67 ? !n243 : n243));
assign n1518 = /* LUT   18 23  1 */ (n286 ? (n708 ? (n738 ? 1'b1 : n95) : n738) : (n708 ? n95 : 1'b0));
assign n2345 = /* LUT    6 20  3 */ (n387 ? (n319 ? (n104 ? 1'b1 : n465) : n104) : (n319 ? n465 : 1'b0));
assign n2346 = /* LUT   11 18  5 */ (n892 ? (n1007 ? !n992 : (n893 ? 1'b1 : !n992)) : (n1007 ? 1'b0 : n893));
assign n2347 = /* LUT    5 20  0 */ (n320 ? (n473 ? (n465 ? n474 : 1'b0) : 1'b0) : (n473 ? n465 : 1'b0));
assign n2348 = /* LUT   15 22  4 */ (\dd_pad_i[12]  ? !io_33_1_1 : 1'b0);
assign n2349 = /* LUT    9 19  4 */ (n794 ? (n898 ? 1'b1 : n793) : (n898 ? !n793 : 1'b0));
assign n2350 = /* LUT   12 19  7 */ (n1023 ? 1'b0 : (n798 ? n1114 : 1'b1));
assign n2351 = /* LUT   12 24  6 */ (n836 ? (n1251 ? 1'b1 : !n677) : (n1251 ? n677 : 1'b0));
assign n2352 = /* LUT   17 23  1 */ (n1498 ? 1'b1 : (n1499 ? 1'b1 : (n1231 ? 1'b1 : n1036)));
assign n2353 = /* LUT    4 18  6 */ (n239 ? 1'b0 : (n242 ? 1'b0 : !n243));
assign n2354 = /* LUT    9 29  5 */ (n636 ? (n634 ? 1'b1 : n130) : (n634 ? !n130 : 1'b0));
assign n2355 = /* LUT    7 23  4 */ (io_33_1_1 ? 1'b0 : \wb_dat_i[4] );
assign n2356 = /* LUT   11 30  0 */ (n847 ? (n966 ? 1'b1 : n130) : (n966 ? !n130 : 1'b0));
assign n2357 = /* LUT   16 23  5 */ (n700 ? (n96 ? 1'b1 : n192) : n192);
assign n2358 = /* LUT   16 28  4 */ (n1431 ? (n1477 ? n286 : (n286 ? n675 : 1'b0)) : (n1477 ? (n286 ? !n675 : 1'b0) : 1'b0));
assign n2359 = /* LUT   13 20  2 */ (wb_clk_i ? !io_33_1_1 : 1'b0);
assign n2360 = /* LUT    6 23  2 */ (n609 ? (io_33_1_1 ? 1'b0 : (n287 ? 1'b1 : n627)) : (io_33_1_1 ? 1'b0 : (n287 ? 1'b0 : n627)));
assign n2361 = /* LUT   12 28  3 */ (n130 ? n850 : n849);
assign n2362 = /* LUT   11 19  6 */ (n1025 ? 1'b0 : (n798 ? n900 : 1'b1));
assign n2363 = /* LUT    5 21  3 */ (n75 ? (n320 ? !n456 : 1'b1) : (n320 ? !n49 : 1'b1));
assign n2364 = /* LUT   15 24  6 */ (n915 ? (n746 ? !n1351 : 1'b0) : (n762 ? 1'b1 : (n746 ? !n1351 : 1'b0)));
assign n2365 = /* LUT    7 27  1 */ (n130 ? (n770 ? 1'b0 : (n223 ? 1'b1 : !n376)) : !n770);
assign n2366 = /* LUT   12 18  4 */ (n1223 ? (n67 ? n52 : !n52) : (n67 ? !n52 : n52));
assign n2367 = /* LUT   12 31  7 */ (n130 ? n526 : n633);
assign n2368 = /* LUT   16 24  1 */ (n677 ? n1416 : n1172);
assign n2369 = /* LUT    9 30  4 */ (n130 ? n780 : n234);
assign n2370 = /* LUT    7 20  5 */ (\wb_dat_i[21]  ? !io_33_1_1 : 1'b0);
assign n2371 = /* LUT    9 17  5 */ (io_33_8_0 ? 1'b0 : !io_33_7_0);
assign n2372 = /* LUT   14 23  3 */ (\wb_dat_i[23]  ? !io_33_1_1 : 1'b0);
assign n2373 = /* LUT   16 27  5 */ (n130 ? n962 : n547);
assign n2374 = /* LUT   13 21  1 */ (n1017 ? (n398 ? (n701 ? 1'b1 : n758) : n758) : (n398 ? n701 : 1'b0));
assign n2375 = /* LUT    6 22  5 */ (n75 ? n618 : n581);
assign n2376 = /* LUT   11 16  7 */ (io_33_14_0 ? !io_33_1_1 : 1'b0);
assign n2377 = /* LUT    5 22  2 */ (n596 ? 1'b0 : (n509 ? 1'b0 : (n595 ? 1'b0 : !n473)));
assign n2378 = /* LUT   15 25  1 */ (n1360 ? 1'b1 : (n1417 ? 1'b1 : (n1362 ? 1'b1 : n1335)));
assign n2379 = /* LUT   15 20  6 */ (io_33_1_1 ? 1'b0 : \wb_dat_i[30] );
assign n2380 = /* LUT    7 24  0 */ (n686 ? 1'b0 : (n408 ? (n709 ? 1'b0 : !n710) : 1'b0));
assign n2381 = /* LUT   12 17  5 */ (io_33_1_1 ? 1'b1 : \wb_dat_i[21] );
assign n2382 = /* LUT   12 30  4 */ (n966 ? (n847 ? 1'b1 : n130) : (n847 ? !n130 : 1'b0));
assign n2383 = /* LUT    5 24  1 */ (\wb_dat_i[20]  ? !n118 : 1'b0);
assign n2384 = /* LUT    4 16  0 */ n342;
assign n2385 = /* LUT    9 18  4 */ (n475 ? 1'b1 : (n887 ? 1'b1 : (n573 ? 1'b1 : n886)));
assign n2386 = /* LUT   14 29  5 */ (n130 ? n547 : n962);
assign n2387 = /* LUT   14 22  4 */ (n1286 ? 1'b1 : (n1345 ? 1'b1 : (n1232 ? 1'b1 : n1034)));
assign n2388 = /* LUT    6 18  2 */ (n51 ? 1'b1 : (n459 ? io_33_1_1 : 1'b1));
assign n2389 = /* LUT   11 28  2 */ (n1105 ? (n978 ? 1'b1 : !n130) : (n978 ? n130 : 1'b0));
assign n2390 = /* LUT   16 26  6 */ (n677 ? n876 : n1415);
assign n2391 = /* LUT   13 22  0 */ (n925 ? (n1175 ? 1'b1 : n677) : (n1175 ? !n677 : 1'b0));
assign n404  = /* LUT    3 22  2 */ (n299 ? (n403 ? (n402 ? !n185 : 1'b0) : 1'b0) : 1'b0);
assign n2392 = /* LUT    6 17  4 */ (n671 ? (io_33_1_1 ? !n450 : (n450 ? n464 : 1'b1)) : (io_33_1_1 ? 1'b0 : (n450 ? n464 : 1'b0)));
assign n2393 = /* LUT   10 30  0 */ (n130 ? n1105 : n978);
assign n2394 = /* LUT    4 20  5 */ (n495 ? (n67 ? n381 : !n381) : (n67 ? !n381 : n381));
assign n2395 = /* LUT    7 18  6 */ (n51 ? (io_33_1_1 ? 1'b0 : (n459 ? n53 : 1'b1)) : (io_33_1_1 ? 1'b0 : !n459));
assign n2396 = /* LUT    7 25  7 */ (n643 ? (n130 ? n719 : 1'b1) : (n130 ? n719 : 1'b0));
assign n2397 = /* LUT   12 16  2 */ (io_33_1_1 ? 1'b0 : \wb_dat_i[0] );
assign n2398 = /* LUT   14 18  1 */ (\wb_dat_o[5]  ? 1'b1 : io_33_1_1);
assign n2399 = /* LUT   12 29  5 */ (n547 ? (n962 ? 1'b1 : !n130) : (n962 ? n130 : 1'b0));
assign n2400 = /* LUT    1 20  2 */ (n183 ? (io_33_1_1 ? !n163 : (n164 ? 1'b1 : !n163)) : (io_33_1_1 ? 1'b0 : (n164 ? n163 : 1'b0)));
assign n2401 = /* LUT   17 18  2 */ (\wb_dat_i[19]  ? !io_33_1_1 : 1'b0);
assign n2402 = /* LUT    5 25  2 */ (n474 ? !io_33_1_1 : 1'b0);
assign n2403 = /* LUT    4 23  1 */ (n238 ? !io_33_1_1 : 1'b0);
assign n2404 = /* LUT    9 24  2 */ (n130 ? \dd_pad_i[0]  : \dd_pad_i[6] );
assign n1379 = /* LUT   14 28  6 */ (n1315 ? (n1182 ? 1'b1 : !n666) : (n1182 ? n666 : 1'b0));
assign n2406 = /* LUT    2 22  5 */ (n285 ? (n305 ? 1'b1 : !n169) : (n305 ? n169 : 1'b0));
assign n2407 = /* LUT   11 22  4 */ (n1147 ? (n1150 ? 1'b1 : n677) : (n1150 ? !n677 : 1'b0));
assign n2408 = /* LUT   11 29  5 */ (n130 ? n966 : n847);
assign n2409 = /* LUT   10 15  5 */ (n273 ? !n67 : n67);
assign n1448 = /* LUT   16 20  0 */ (n1037 ? n512 : 1'b0);
assign n2411 = /* LUT   15 18  7 */ (io_33_1_1 ? 1'b1 : \wb_dat_i[20] );
assign n411  = /* LUT    3 23  1 */ (n319 ? (n287 ? n308 : 1'b1) : (n287 ? n308 : 1'b0));
assign n2413 = /* LUT    2 21  1 */ (n289 ? (n67 ? n266 : !n266) : (n67 ? !n266 : n266));
assign n2414 = /* LUT   12 20  7 */ (io_33_1_1 ? 1'b0 : \wb_dat_i[16] );
assign n2415 = /* LUT   10 17  1 */ (n893 ? (n999 ? 1'b0 : n747) : !n999);
assign n2416 = /* LUT    7 19  5 */ (n487 ? 1'b0 : (n754 ? 1'b1 : (n666 ? !n686 : n686)));
assign n2417 = /* LUT    3 24  5 */ (\wb_dat_o[5]  ? !n118 : 1'b0);
assign n1244 = /* LUT   12 23  3 */ (n870 ? (n1163 ? 1'b1 : n677) : (n1163 ? !n677 : 1'b0));
assign n2419 = /* LUT    5 26  3 */ \wb_dat_i[5] ;
assign n2420 = /* LUT   11 25  2 */ (n827 ? (n828 ? 1'b1 : n130) : (n828 ? !n130 : 1'b0));
assign n2421 = /* LUT    4 22  2 */ (n280 ? (n181 ? io_33_1_1 : (io_33_1_1 ? 1'b1 : !n173)) : io_33_1_1);
assign n2422 = /* LUT    9 25  1 */ (n130 ? n828 : n827);
assign n2423 = /* LUT   11 26  4 */ (n130 ? n827 : n828);
assign n2424 = /* LUT   16 19  1 */ (n1113 ? (n1442 ? 1'b1 : (n1439 ? 1'b1 : n758)) : (n1442 ? 1'b1 : n1439));
assign n2425 = /* LUT    3 20  0 */ (n379 ? io_33_1_1 : (io_33_1_1 ? 1'b1 : (n182 ? 1'b0 : n202)));
assign n2426 = /* LUT    2 20  2 */ (n181 ? !io_33_1_1 : (n278 ? (io_33_1_1 ? 1'b0 : n173) : 1'b0));
assign n2427 = /* LUT   12 27  6 */ (n547 ? (n962 ? 1'b1 : n130) : (n962 ? !n130 : 1'b0));
assign n2428 = /* LUT    6 19  6 */ io_33_15_1;
assign n1433 = /* LUT   15 28  2 */ (n666 ? n775 : n1080);
assign n1238 = /* LUT   12 22  0 */ (n1143 ? (n1121 ? (n96 ? 1'b1 : n104) : n96) : (n1121 ? n104 : 1'b0));
assign n2431 = /* LUT    1 22  0 */ (io_33_1_1 ? 1'b0 : io_33_5_0);
assign n2432 = /* LUT    5 27  4 */ (n130 ? n418 : n335);
assign n2433 = /* LUT    4 21  3 */ (n300 ? (io_33_1_1 ? 1'b0 : n507) : n373);
assign n2434 = /* LUT    9 26  0 */ (n840 ? 1'b0 : (n335 ? 1'b1 : (n376 ? !n130 : 1'b1)));
assign n2435 = /* LUT    2 24  7 */ (n327 ? n220 : !n220);
assign n2436 = /* LUT   14 19  7 */ (\wb_dat_i[14]  ? !io_33_1_1 : 1'b0);
assign n2437 = /* LUT   11 20  6 */ (n892 ? (n1039 ? !n1134 : (n893 ? 1'b1 : !n1134)) : (n1039 ? 1'b0 : n893));
assign n2438 = /* LUT   11 27  7 */ (n636 ? (n634 ? 1'b1 : n130) : (n634 ? !n130 : 1'b0));
assign n2439 = /* LUT    3 21  7 */ (n276 ? (n301 ? !io_33_1_1 : 1'b0) : 1'b0);
assign n2440 = /* LUT    2 23  3 */ (n212 ? (io_33_1_1 ? 1'b1 : (n197 ? 1'b1 : !n205)) : (io_33_1_1 ? n205 : (n197 ? n205 : 1'b0)));
assign n2441 = /* LUT   20 22  3 */ (n903 ? (n1285 ? !n1040 : 1'b0) : (n1285 ? (n1338 ? 1'b1 : !n1040) : n1338));
assign n2442 = /* LUT   12 26  5 */ (n872 ? (n874 ? 1'b1 : n130) : (n874 ? !n130 : 1'b0));
assign n1503 = /* LUT   17 24  3 */ (n677 ? n983 : n837);
assign n1019 = /* LUT   10 19  3 */ (n587 ? (n270 ? 1'b1 : n75) : (n270 ? (n75 ? n801 : 1'b1) : (n75 ? n801 : 1'b0)));
assign n2445 = /* LUT    7 17  3 */ (n741 ? (n67 ? n569 : !n569) : (n67 ? !n569 : n569));
assign n2446 = /* LUT    7 28  4 */ (n666 ? n658 : n728);
assign n2447 = /* LUT   14 26  5 */ n764;
assign n2448 = /* LUT   12 21  1 */ (\wb_dat_i[25]  ? !io_33_1_1 : 1'b0);
assign n2449 = /* LUT    5 28  5 */ (n438 ? (io_33_1_1 ? 1'b0 : (n287 ? 1'b1 : n657)) : (io_33_1_1 ? 1'b0 : (n287 ? 1'b0 : n657)));
assign n2450 = /* LUT   14 25  1 */ (n130 ? n779 : n964);
assign n2451 = /* LUT    3 17  4 */ (n147 ? (io_33_1_1 ? 1'b1 : (n254 ? n341 : 1'b1)) : (io_33_1_1 ? n254 : (n254 ? n341 : 1'b0)));
assign n2452 = /* LUT    6 21  7 */ (n90 ? (n611 ? 1'b1 : !n169) : (n611 ? n169 : 1'b0));
assign n2453 = /* LUT   11 24  6 */ (n781 ? (n130 ? n338 : 1'b1) : (n130 ? n338 : 1'b0));
assign n2454 = /* LUT   15 17  2 */ (io_33_1_1 ? 1'b0 : \wb_dat_i[8] );
assign n2455 = /* LUT    3 18  6 */ (n254 ? (io_33_1_1 ? 1'b0 : n343) : n35);
assign n2456 = /* LUT   12 25  4 */ (n666 ? n839 : n224);
assign n564  = /* LUT    5 16  0 */ (n240 ? 1'b1 : (n245 ? 1'b1 : (n243 ? 1'b1 : n244)));
assign n2458 = /* LUT   10 25  5 */ (n130 ? n780 : n234);
assign n2459 = /* LUT   10 18  4 */ (n460 ? (io_33_1_1 ? 1'b1 : n1001) : n586);
assign n2460 = /* LUT    7 22  2 */ (n474 ? !io_33_1_1 : 1'b0);
assign n2461 = /* LUT   14 21  4 */ (io_33_1_1 ? 1'b0 : \wb_dat_i[24] );
assign n2462 = /* LUT    6 26  3 */ (n718 ? 1'b0 : (n315 ? 1'b1 : (n376 ? !n130 : 1'b1)));
assign n1118 = /* LUT   11 17  6 */ (n892 ? (n1112 ? !n1005 : (n893 ? 1'b1 : !n1005)) : (n1112 ? 1'b0 : n893));
assign n1356 = /* LUT   14 24  2 */ (n1076 ? (n712 ? 1'b1 : n677) : (n712 ? !n677 : 1'b0));
assign n2465 = /* LUT    6 20  4 */ !n594;
assign n2466 = /* LUT    6 25  7 */ (n130 ? (n545 ? 1'b0 : !n376) : (n545 ? (n376 ? !n310 : 1'b0) : (n376 ? !n310 : 1'b1)));
assign n1122 = /* LUT   11 18  0 */ (n798 ? (n892 ? (n1113 ? !n796 : 1'b1) : !n1113) : (n892 ? !n796 : 1'b0));
assign n1054 = /* LUT   10 22  1 */ (n75 ? n802 : n793);
assign n2468 = /* LUT   15 22  3 */ (\wb_dat_i[30]  ? !io_33_1_1 : 1'b0);
assign n2469 = /* LUT   18 18  6 */ (io_33_16_1 ? !io_33_1_1 : 1'b0);
assign n2470 = /* LUT    3 19  5 */ (n254 ? (io_33_1_1 ? 1'b0 : n271) : n70);
assign n2471 = /* LUT   12 24  3 */ (n1250 ? (n1215 ? 1'b1 : !n677) : (n1215 ? n677 : 1'b0));
assign n2472 = /* LUT    5 17  3 */ io_33_13_0;
assign n2473 = /* LUT   10 24  6 */ (n941 ? (n943 ? 1'b1 : !n666) : (n943 ? n666 : 1'b0));
assign n2474 = /* LUT   10 21  5 */ (n919 ? !n1049 : (n1049 ? 1'b0 : !n893));
assign n2475 = /* LUT    7 23  1 */ (io_33_1_1 ? 1'b0 : io_33_15_1);
assign n2476 = /* LUT   14 20  7 */ (n1128 ? (io_33_7_0 ? (io_33_8_0 ? 1'b0 : n1337) : 1'b0) : 1'b0);
assign n2477 = /* LUT   17 20  0 */ (n708 ? (n755 ? (n512 ? 1'b1 : n86) : n86) : (n755 ? n512 : 1'b0));
assign n2478 = /* LUT   11 30  7 */ (n130 ? n1105 : n978);
assign n2479 = /* LUT   16 28  1 */ (n1430 ? 1'b1 : (n1476 ? 1'b1 : (n1336 ? 1'b1 : n1429)));
assign n1330 = /* LUT   13 31  0 */ (n666 ? n860 : n967);
assign n2481 = /* LUT   18 22  3 */ (n758 ? (n1516 ? 1'b1 : (n1495 ? 1'b1 : n40)) : (n1516 ? 1'b1 : n1495));
assign n2482 = /* LUT   14 27  3 */ (n1307 ? (n666 ? n1256 : 1'b1) : (n666 ? n1256 : 1'b0));
assign n2483 = /* LUT    6 24  4 */ (n130 ? n310 : n222);
assign n2484 = /* LUT   11 19  3 */ (n1128 ? !n1132 : (n1132 ? 1'b0 : !n798));
assign n2485 = /* LUT   13 17  1 */ (\dd_pad_i[12]  ? !io_33_1_1 : 1'b0);
assign n1407 = /* LUT   15 23  0 */ (n96 ? (n1347 ? 1'b1 : (n104 ? n1125 : 1'b0)) : (n104 ? n1125 : 1'b0));
assign n2487 = /* LUT   18 21  7 */ (\wb_dat_i[2]  ? !io_33_8_0 : 1'b1);
assign n1282 = /* LUT   12 31  2 */ (n855 ? (n871 ? 1'b1 : !n666) : (n871 ? n666 : 1'b0));
assign n578  = /* LUT    5 18  2 */ (n275 ? io_33_1_1 : (n452 ? (io_33_1_1 ? 1'b1 : !n273) : io_33_1_1));
assign n2490 = /* LUT   10 27  7 */ (n169 ? n707 : n228);
assign n1032 = /* LUT   10 20  6 */ (n792 ? 1'b0 : (n169 ? (n896 ? 1'b0 : n700) : 1'b0));
assign n2491 = /* LUT    7 20  0 */ (n517 ? (io_33_1_1 ? 1'b1 : n708) : io_33_1_1);
assign n2492 = /* LUT   14 23  6 */ (io_33_1_1 ? 1'b0 : \wb_dat_i[4] );
assign n1490 = /* LUT   17 21  3 */ (n1041 ? !io_33_8_0 : 1'b0);
assign n2494 = /* LUT    1 18  4 */ (n159 ? (n67 ? n60 : !n60) : (n67 ? !n60 : n60));
assign n1217 = /* LUT   11 31  4 */ (n1184 ? (n854 ? 1'b1 : !n666) : (n854 ? n666 : 1'b0));
assign n2496 = /* LUT   16 27  0 */ (n1105 ? (n978 ? 1'b1 : !n130) : (n978 ? n130 : 1'b0));
assign n705  = /* LUT    6 22  2 */ (n388 ? (n704 ? (n498 ? 1'b0 : \wb_adr_i[5] ) : 1'b1) : !n704);
assign n724  = /* LUT    6 27  5 */ (n425 ? (n376 ? 1'b0 : !n625) : (n376 ? !n130 : !n625));
assign n2499 = /* LUT   11 16  2 */ (io_33_1_1 ? 1'b1 : io_33_16_1);
assign n2500 = /* LUT   13 18  0 */ (n701 ? (n891 ? (n512 ? 1'b1 : n612) : n612) : (n891 ? n512 : 1'b0));
assign n2501 = /* LUT   15 20  1 */ (\wb_dat_i[18]  ? !io_33_1_1 : 1'b0);
assign n1512 = /* LUT   18 20  4 */ (io_33_7_0 ? 1'b0 : (io_33_8_0 ? 1'b0 : n1337));
assign n2502 = /* LUT   12 30  1 */ (n130 ? n964 : n779);
assign n2503 = /* LUT    5 24  4 */ (n118 ? 1'b0 : \dd_pad_i[7] );
assign n2504 = /* LUT    5 19  5 */ (n390 ? 1'b0 : (n590 ? (io_33_1_1 ? 1'b0 : !n77) : 1'b0));
assign n2505 = /* LUT   10 26  0 */ (n130 ? n780 : n234);
assign n2506 = /* LUT   10 23  7 */ (n675 ? n927 : n1059);
assign n2507 = /* LUT   15 26  0 */ (n677 ? n560 : n834);
assign n1344 = /* LUT   14 22  1 */ (n675 ? n1289 : n1343);
assign n2509 = /* LUT    6 18  7 */ (n50 ? (n682 ? (io_33_1_1 ? !n460 : 1'b1) : (io_33_1_1 ? 1'b0 : n460)) : (n682 ? !n460 : 1'b0));
assign n2510 = /* LUT   17 22  2 */ (n905 ? (n1494 ? 1'b1 : (n1456 ? 1'b1 : n512)) : (n1494 ? 1'b1 : n1456));
assign n2511 = /* LUT   11 28  5 */ (n130 ? n966 : n847);
assign n2512 = /* LUT    4 19  1 */ (n466 ? (n479 ? (io_33_1_1 ? 1'b0 : n360) : !io_33_1_1) : (n479 ? 1'b0 : !io_33_1_1));
assign n2513 = /* LUT    9 28  2 */ (n130 ? n827 : n828);
assign n1520 = /* LUT   18 24  1 */ (io_33_7_0 ? (\wb_adr_i[5]  ? 1'b1 : n1488) : (\wb_adr_i[5]  ? 1'b1 : (n1488 ? 1'b1 : \wb_dat_i[2] )));
assign n2514 = /* LUT    6 17  3 */ (n670 ? (io_33_1_1 ? 1'b1 : (n574 ? 1'b1 : !n450)) : (io_33_1_1 ? n450 : (n574 ? n450 : 1'b0)));
assign n2515 = /* LUT   10 30  5 */ (n964 ? (n779 ? 1'b1 : !n130) : (n779 ? n130 : 1'b0));
assign n2516 = /* LUT    9 14  5 */ (\wb_dat_o[5]  ? 1'b1 : io_33_1_1);
assign n2517 = /* LUT   13 19  7 */ (io_33_1_1 ? 1'b0 : wb_clk_i);
assign n2518 = /* LUT    3 27  1 */ (n130 ? \dd_pad_i[5]  : \dd_pad_i[15] );
assign n2519 = /* LUT    2 17  1 */ (n247 ? (n67 ? n239 : !n239) : (n67 ? !n239 : n239));
assign n2520 = /* LUT   14 18  6 */ (io_33_1_1 ? 1'b1 : \dd_pad_i[2] );
assign n2521 = /* LUT   12 29  0 */ (n1094 ? (n1197 ? 1'b1 : n666) : (n1197 ? !n666 : 1'b0));
assign n2522 = /* LUT    5 20  4 */ (n388 ? (n598 ? (n505 ? 1'b0 : n509) : 1'b0) : 1'b0);
assign n2523 = /* LUT   10 29  1 */ (n962 ? (n547 ? 1'b1 : n130) : (n547 ? !n130 : 1'b0));
assign n2524 = /* LUT   12 19  3 */ (n1015 ? 1'b0 : (n798 ? n1027 : 1'b1));
assign n2525 = /* LUT   17 23  5 */ iordy_pad_i;
assign n2526 = /* LUT   11 29  2 */ (n538 ? (n635 ? 1'b1 : n130) : (n635 ? !n130 : 1'b0));
assign n2527 = /* LUT   16 25  2 */ (io_33_1_1 ? 1'b0 : \dd_pad_i[7] );
assign n467  = /* LUT    4 18  2 */ (n240 ? 1'b0 : (n244 ? 1'b0 : (n245 ? 1'b0 : !n241)));
assign n2529 = /* LUT    9 29  1 */ (n780 ? (n234 ? 1'b1 : n130) : (n234 ? !n130 : 1'b0));
assign n2530 = /* LUT   13 23  4 */ (n1295 ? (n1168 ? 1'b1 : !n169) : (n1168 ? n169 : 1'b0));
assign n2531 = /* LUT   16 23  1 */ (n1168 ? (n1463 ? 1'b1 : (n1406 ? 1'b1 : n701)) : (n1463 ? 1'b1 : n1406));
assign n2532 = /* LUT   13 20  6 */ (\wb_dat_i[17]  ? !io_33_1_1 : 1'b0);
assign n2533 = /* LUT    3 24  0 */ (n118 ? 1'b0 : \wb_dat_i[30] );
assign n2534 = /* LUT   11 12  3 */ (\wb_dat_i[8]  ? !io_33_1_1 : 1'b0);
assign n2535 = /* LUT    5 26  6 */ \wb_dat_i[8] ;
assign n2536 = /* LUT   11 25  7 */ (n130 ? n764 : n720);
assign n2537 = /* LUT    5 21  7 */ (n75 ? n474 : n473);
assign n2538 = /* LUT   10 28  2 */ (n130 ? n337 : n131);
assign n2539 = /* LUT   15 24  2 */ (\wb_dat_i[14]  ? !io_33_1_1 : 1'b0);
assign n2543 = /* LUT   14 16  3 */ (io_33_1_1 ? 1'b0 : io_33_9_0);
assign n2544 = /* LUT    6 28  5 */ (n75 ? n531 : n585);
assign n2545 = /* LUT   11 26  3 */ (n719 ? (n643 ? 1'b1 : !n130) : (n643 ? n130 : 1'b0));
assign n2546 = /* LUT   12 32  6 */ (n1187 ? (n1183 ? 1'b1 : n666) : (n1183 ? !n666 : 1'b0));
assign n2547 = /* LUT    9 30  0 */ (n973 ? (n865 ? 1'b1 : n666) : (n865 ? !n666 : 1'b0));
assign n2548 = /* LUT   13 24  5 */ (n720 ? (n764 ? 1'b1 : !n130) : (n764 ? n130 : 1'b0));
assign n2549 = /* LUT    6 19  1 */ io_33_5_0;
assign n2550 = /* LUT   10 16  7 */ (n892 ? (n603 ? !n885 : (n893 ? 1'b1 : !n885)) : (n603 ? 1'b0 : n893));
assign n2551 = /* LUT   13 21  5 */ (n1167 ? (n1011 ? (n701 ? 1'b1 : n758) : n701) : (n1011 ? n758 : 1'b0));
assign n2552 = /* LUT    2 19  3 */ (n265 ? (n79 ? io_33_1_1 : 1'b1) : (n79 ? io_33_1_1 : 1'b0));
assign n2553 = /* LUT   20 18  3 */ (io_33_5_0 ? !io_33_1_1 : 1'b0);
assign n1508 = /* LUT   17 28  3 */ (n677 ? n1104 : n1303);
assign n2555 = /* LUT    5 27  1 */ (n316 ? (n223 ? 1'b1 : n130) : (n223 ? !n130 : 1'b0));
assign n2556 = /* LUT    5 22  6 */ (n317 ? (n181 ? !io_33_1_1 : 1'b0) : 1'b0);
assign n2557 = /* LUT   10 31  3 */ (n666 ? n965 : n982);
assign n2558 = /* LUT   15 25  5 */ (n1385 ? n708 : 1'b0);
assign n2559 = /* LUT   14 19  2 */ (io_33_1_1 ? 1'b1 : io_33_16_1);
assign n2560 = /* LUT   11 27  0 */ (n130 ? n968 : n769);
assign n2561 = /* LUT    4 27  5 */ (n75 ? n532 : n421);
assign n2562 = /* LUT   13 25  6 */ (n130 ? wb_inta_o : \dd_pad_i[1] );
assign n2563 = /* LUT   18 16  5 */ (\wb_dat_i[4]  ? !io_33_1_1 : 1'b0);
assign n2564 = /* LUT   14 29  1 */ (n130 ? n1105 : n978);
assign n2565 = /* LUT   18 29  6 */ (n778 ? (n1421 ? 1'b1 : !n677) : (n1421 ? n677 : 1'b0));
assign n2566 = /* LUT   16 21  3 */ (n504 ? n512 : 1'b0);
assign n2567 = /* LUT   10 19  6 */ (n792 ? n67 : n1021);
assign n2568 = /* LUT   15 29  2 */ (n1190 ? (n1206 ? 1'b1 : n666) : (n1206 ? !n666 : 1'b0));
assign n2569 = /* LUT   13 22  4 */ (n1233 ? 1'b1 : (n1293 ? 1'b1 : (n917 ? 1'b1 : n1235)));
assign n2570 = /* LUT    2 18  4 */ (n163 ? (io_33_1_1 ? 1'b1 : n196) : n170);
assign n2571 = /* LUT    4 20  1 */ (n491 ? (n67 ? n384 : !n384) : (n67 ? !n384 : n384));
assign n2572 = /* LUT    7 18  2 */ (n684 ? (n677 ? !n118 : 1'b0) : (n675 ? !n118 : 1'b0));
assign n2573 = /* LUT    9 27  4 */ (n130 ? n849 : n850);
assign n2574 = /* LUT   11 24  1 */ (n130 ? n234 : n780);
assign n2575 = /* LUT    4 26  6 */ (n118 ? 1'b0 : wb_clk_i);
assign n2576 = /* LUT    4 23  5 */ (n276 ? (io_33_1_1 ? 1'b0 : (n297 ? 1'b1 : n202)) : (io_33_1_1 ? 1'b0 : n297));
assign n2577 = /* LUT    9 24  6 */ (n130 ? \dd_pad_i[13]  : \dd_pad_i[8] );
assign n2578 = /* LUT   13 26  7 */ n769;
assign n1378 = /* LUT   14 28  2 */ (n677 ? n1377 : n1312);
assign n2580 = /* LUT    2 22  1 */ (n93 ? (n106 ? 1'b1 : !n169) : (n106 ? n169 : 1'b0));
assign n1149 = /* LUT   11 22  0 */ (n330 ? (n762 ? !n1043 : 1'b0) : (n762 ? (n746 ? 1'b1 : !n1043) : n746));
assign n2582 = /* LUT    5 16  7 */ (n447 ? io_33_1_1 : (io_33_1_1 ? 1'b1 : (n449 ? 1'b1 : n472)));
assign n2583 = /* LUT   16 20  4 */ (\wb_dat_i[20]  ? !io_33_1_1 : 1'b0);
assign n2584 = /* LUT   10 18  1 */ (io_33_1_1 ? (n1008 ? !n460 : 1'b0) : (n1012 ? (n1008 ? 1'b1 : n460) : (n1008 ? !n460 : 1'b0)));
assign n2585 = /* LUT   15 18  3 */ (io_33_1_1 ? 1'b1 : \wb_dat_i[22] );
assign n2586 = /* LUT    2 21  5 */ (n293 ? (n67 ? n268 : !n268) : (n67 ? !n268 : n268));
assign n2587 = /* LUT   12 20  3 */ (io_33_1_1 ? 1'b0 : io_33_15_1);
assign n2588 = /* LUT    5 29  3 */ (n75 ? n453 : n332);
assign n752  = /* LUT    7 19  1 */ (n693 ? (n677 ? (n698 ? !n675 : n675) : 1'b1) : (n677 ? 1'b1 : (n698 ? !n675 : n675)));
assign n2590 = /* LUT    9 20  5 */ \wb_adr_i[4] ;
assign n2591 = /* LUT    6 25  2 */ (n376 ? (n518 ? 1'b0 : !n130) : !n540);
assign n2592 = /* LUT    4 25  7 */ io_33_9_0;
assign n2593 = /* LUT   10 22  6 */ (n911 ? (n287 ? io_33_1_1 : 1'b1) : 1'b1);
assign n2594 = /* LUT    4 22  6 */ (io_33_1_1 ? 1'b0 : (n514 ? !io_31_0_1 : 1'b0));
assign n2595 = /* LUT    9 25  5 */ (n130 ? n720 : n764);
assign n2596 = /* LUT   13 27  0 */ (n547 ? (n962 ? 1'b1 : !n130) : (n962 ? n130 : 1'b0));
assign n2597 = /* LUT   11 23  3 */ (n1033 ? 1'b1 : (n1162 ? 1'b1 : (n989 ? 1'b1 : n1158)));
assign n2598 = /* LUT    5 17  4 */ wb_we_i;
assign n2599 = /* LUT   16 19  5 */ (n1387 ? 1'b1 : (n1443 ? 1'b1 : (n73 ? 1'b1 : n561)));
assign n1047 = /* LUT   10 21  0 */ (n892 ? (n1046 ? !n814 : (n893 ? 1'b1 : !n814)) : (n1046 ? 1'b0 : n893));
assign n2601 = /* LUT   15 19  0 */ (n990 ? (n701 ? (n303 ? 1'b1 : n104) : n104) : (n701 ? n303 : 1'b0));
assign n2602 = /* LUT    2 20  6 */ (n181 ? !io_33_1_1 : (io_33_1_1 ? 1'b0 : (n177 ? !n173 : 1'b0)));
assign n2603 = /* LUT   12 27  2 */ (n538 ? (n635 ? 1'b1 : n130) : (n635 ? !n130 : 1'b0));
assign n2604 = /* LUT   13 31  5 */ (\wb_adr_i[5]  ? (n286 ? (n1280 ? 1'b1 : n1277) : n1280) : (n286 ? n1277 : 1'b0));
assign n1239 = /* LUT   12 22  4 */ (n1156 ? (n1165 ? 1'b1 : !n675) : (n1165 ? n675 : 1'b0));
assign n2606 = /* LUT    6 24  1 */ (n416 ? (n431 ? 1'b1 : n130) : (n431 ? !n130 : 1'b0));
assign n2607 = /* LUT    4 24  0 */ (\wb_dat_i[27]  ? !n118 : 1'b0);
assign n2608 = /* LUT    4 21  7 */ (n300 ? (n508 ? !io_33_1_1 : 1'b0) : n370);
assign n2609 = /* LUT    9 26  4 */ (n376 ? (n957 ? 1'b0 : (n126 ? 1'b1 : !n130)) : !n957);
assign n1318 = /* LUT   13 28  1 */ (n666 ? n1093 : n525);
assign n1514 = /* LUT   18 21  2 */ (\wb_adr_i[5]  ? 1'b0 : !\wb_adr_i[3] );
assign n2611 = /* LUT   14 30  4 */ n643;
assign n2612 = /* LUT    2 24  3 */ (n323 ? (n67 ? n207 : !n207) : (n67 ? !n207 : n207));
assign n1140 = /* LUT   11 20  2 */ (n892 ? (n903 ? !n1053 : (n893 ? 1'b1 : !n1053)) : (n903 ? 1'b0 : n893));
assign n2614 = /* LUT   17 27  3 */ (io_33_1_1 ? 1'b0 : \wb_dat_i[24] );
assign n2615 = /* LUT    5 18  5 */ (n465 ? (n84 ? 1'b1 : (n477 ? 1'b1 : n54)) : (n477 ? 1'b1 : n54));
assign n1031 = /* LUT   10 20  3 */ (n892 ? (n1029 ? !n783 : (n783 ? n893 : 1'b1)) : (n1029 ? 1'b0 : n893));
assign n2617 = /* LUT    2 23  7 */ (n216 ? (io_33_1_1 ? !n205 : (n111 ? 1'b1 : !n205)) : (io_33_1_1 ? 1'b0 : (n111 ? n205 : 1'b0)));
assign n2618 = /* LUT   12 26  1 */ (n964 ? (n779 ? 1'b1 : n130) : (n779 ? !n130 : 1'b0));
assign n1491 = /* LUT   17 21  4 */ (n1119 ? (n1490 ? (n1337 ? 1'b1 : n512) : n512) : (n1490 ? n1337 : 1'b0));
assign n2620 = /* LUT    7 17  7 */ (n745 ? n476 : !n476);
assign n2621 = /* LUT   14 26  1 */ n978;
assign n2622 = /* LUT   12 21  5 */ (\wb_dat_i[23]  ? !io_33_1_1 : 1'b0);
assign n2623 = /* LUT    6 27  0 */ (n130 ? (n622 ? 1'b0 : !n376) : (n622 ? (n376 ? !n313 : 1'b0) : (n376 ? !n313 : 1'b1)));
assign n2624 = /* LUT   13 29  2 */ (n666 ? n1254 : n1305);
assign n2625 = /* LUT   18 20  1 */ (io_33_8_0 ? n1511 : (n1511 ? 1'b1 : (n1337 ? n805 : 1'b0)));
assign n2626 = /* LUT    3 17  0 */ (n71 ? (io_33_1_1 ? 1'b1 : (n254 ? n45 : 1'b1)) : (io_33_1_1 ? n254 : (n254 ? n45 : 1'b0)));
assign n1365 = /* LUT   14 25  5 */ (n666 ? n1089 : n1355);
assign n2628 = /* LUT   11 21  5 */ (n320 ? (n879 ? (n96 ? 1'b1 : n104) : n96) : (n879 ? n104 : 1'b0));
assign n589  = /* LUT    5 19  2 */ (n588 ? (n263 ? n356 : 1'b1) : (n263 ? n356 : (n165 ? 1'b1 : n356)));
assign n2629 = /* LUT   10 23  2 */ (n130 ? n234 : n780);
assign n2630 = /* LUT   15 17  6 */ (io_33_1_1 ? 1'b0 : io_33_9_0);
assign n2631 = /* LUT    7 21  4 */ (\wb_dat_i[27]  ? !io_33_1_1 : 1'b0);
assign n2632 = /* LUT   12 25  0 */ (n666 ? n963 : n1170);
assign n2633 = /* LUT   17 22  5 */ (n286 ? (n94 ? (n1195 ? 1'b1 : n708) : n1195) : (n94 ? n708 : 1'b0));
assign n2634 = /* LUT    1 19  0 */ io_33_13_0;
assign n2635 = /* LUT   10 25  1 */ (n130 ? n849 : n850);
assign n480  = /* LUT    4 19  4 */ (n75 ? n456 : n49);
assign n2636 = /* LUT    7 22  6 */ (n698 ? (n408 ? (n118 ? 1'b0 : n709) : !n118) : (n408 ? (n118 ? 1'b0 : n709) : 1'b0));
assign n934  = /* LUT    9 23  0 */ (n820 ? (n730 ? 1'b1 : !n677) : (n730 ? n677 : 1'b0));
assign n2638 = /* LUT   14 21  0 */ (io_33_1_1 ? 1'b0 : \wb_dat_i[17] );
assign n2639 = /* LUT   11 17  2 */ (n1002 ? 1'b0 : (n893 ? n881 : 1'b1));
assign n2640 = /* LUT    1 13  4 */ arst_i;
assign n1328 = /* LUT   13 30  3 */ (n666 ? n1091 : n1082);
assign n2642 = /* LUT    2 17  4 */ (n250 ? (n67 ? n242 : !n242) : (n67 ? !n242 : n242));
assign n2643 = /* LUT   18 23  0 */ (n889 ? (n104 ? 1'b1 : (n96 ? n1497 : 1'b0)) : (n96 ? n1497 : 1'b0));
assign n2644 = /* LUT   14 24  6 */ (io_33_1_1 ? 1'b0 : \wb_dat_i[16] );
assign n694  = /* LUT    6 20  0 */ (n84 ? (io_33_1_1 ? 1'b0 : (n78 ? 1'b0 : n514)) : 1'b0);
assign n2646 = /* LUT   11 15  7 */ (n883 ? (n221 ? (n512 ? 1'b1 : n708) : n512) : (n221 ? n708 : 1'b0));
assign n2647 = /* LUT   11 18  4 */ (n798 ? (n892 ? (n1121 ? !n880 : 1'b1) : !n880) : (n892 ? !n1121 : 1'b0));
assign n598  = /* LUT    5 20  3 */ (n319 ? 1'b0 : (n595 ? 1'b0 : (n483 ? 1'b0 : !io_33_1_1)));
assign n2648 = /* LUT   15 27  4 */ (n666 ? n861 : n1372);
assign n2649 = /* LUT   15 22  7 */ (\wb_dat_i[0]  ? !io_33_1_1 : 1'b0);
assign n2650 = /* LUT    7 26  5 */ (n169 ? n650 : n601);
assign n2651 = /* LUT    9 19  5 */ \wb_adr_i[3] ;
assign n2652 = /* LUT   12 19  6 */ (n1022 ? 1'b0 : (n1227 ? 1'b1 : !n798));
assign n2653 = /* LUT   12 24  7 */ (n677 ? n961 : n841);
assign n2654 = /* LUT   17 26  5 */ (\wb_dat_i[11]  ? !io_33_1_1 : 1'b0);
assign n2655 = /* LUT   10 24  2 */ (n337 ? (n131 ? 1'b1 : !n130) : (n131 ? n130 : 1'b0));
assign n2656 = /* LUT    4 18  7 */ (n466 ? (n350 ? 1'b0 : (io_33_1_1 ? 1'b0 : n352)) : !io_33_1_1);
assign n2657 = /* LUT    7 23  5 */ (io_33_1_1 ? 1'b0 : \wb_dat_i[0] );
assign n2658 = /* LUT    9 16  1 */ (n882 ? 1'b0 : (n798 ? n784 : 1'b1));
assign n2659 = /* LUT   11 30  3 */ (n130 ? n633 : n526);
assign n2660 = /* LUT   16 23  4 */ \dd_pad_i[9] ;
assign n2661 = /* LUT   16 28  5 */ (n706 ? (\wb_adr_i[5]  ? (n1428 ? 1'b1 : n96) : n96) : (\wb_adr_i[5]  ? n1428 : 1'b0));
assign n2662 = /* LUT   20 19  7 */ (io_33_1_1 ? 1'b0 : io_33_19_0);
assign n2663 = /* LUT   14 27  7 */ (n872 ? (n874 ? 1'b1 : n130) : (n874 ? !n130 : 1'b0));
assign n1267 = /* LUT   12 28  4 */ (n666 ? n1092 : n1083);
assign n2665 = /* LUT   11 19  7 */ (n892 ? (n420 ? !n1125 : (n893 ? 1'b1 : !n1125)) : (n420 ? 1'b0 : n893));
assign n604  = /* LUT    5 21  0 */ (n401 ? (n474 ? (n510 ? 1'b0 : !n75) : (n510 ? n75 : 1'b1)) : (n510 ? 1'b0 : !n75));
assign n2667 = /* LUT   15 24  5 */ (n677 ? n926 : n832);
assign n2668 = /* LUT   15 23  4 */ (n512 ? n420 : 1'b0);
assign n2669 = /* LUT    7 27  6 */ (n686 ? 1'b0 : (n408 ? (n709 ? !n710 : 1'b0) : 1'b0));
assign n2670 = /* LUT   12 18  5 */ (n1224 ? (n67 ? n573 : !n573) : (n67 ? !n573 : n573));
assign n2671 = /* LUT   12 31  6 */ (n526 ? (n633 ? 1'b1 : !n130) : (n633 ? n130 : 1'b0));
assign n2672 = /* LUT    7 20  4 */ (\wb_dat_i[19]  ? !io_33_1_1 : 1'b0);
assign n2673 = /* LUT   14 23  2 */ (io_33_1_1 ? 1'b0 : io_33_17_0);
assign n2674 = /* LUT   11 31  0 */ (n1067 ? (n1108 ? 1'b1 : n666) : (n1108 ? !n666 : 1'b0));
assign n2675 = /* LUT   16 27  4 */ (n547 ? (n962 ? 1'b1 : n130) : (n962 ? !n130 : 1'b0));
assign n2676 = /* LUT    6 22  6 */ (n169 ? n612 : n687);
assign n2677 = /* LUT    5 22  1 */ (n498 ? (n613 ? 1'b0 : (wb_we_i ? !n509 : n509)) : (n613 ? 1'b0 : n509));
assign n2678 = /* LUT   15 25  2 */ \dd_pad_i[1] ;
assign n2679 = /* LUT   15 20  5 */ (\wb_dat_i[27]  ? 1'b1 : io_33_1_1);
assign n2680 = /* LUT    7 24  7 */ (n408 ? (n118 ? 1'b0 : n686) : (n693 ? !n118 : 1'b0));
assign n1276 = /* LUT   12 30  5 */ (n666 ? n1258 : n1208);
assign n2682 = /* LUT    5 24  0 */ (n118 ? 1'b0 : \wb_dat_i[24] );
assign n2683 = /* LUT   10 26  4 */ (n130 ? n526 : n633);
assign n2684 = /* LUT    4 16  1 */ (io_0_6_0 ? (n17 ? 1'b0 : wb_stb_i) : 1'b0);
assign n2685 = /* LUT    7 14  2 */ (io_0_3_1 ? (n237 ? (io_0_4_0 ? !n606 : 1'b1) : 1'b0) : n237);
assign n2686 = /* LUT    9 18  3 */ (n67 ? !n166 : n166);
assign n2687 = /* LUT   14 29  4 */ (n1323 ? (n735 ? 1'b1 : !n666) : (n735 ? n666 : 1'b0));
assign n2688 = /* LUT   14 22  5 */ \dd_pad_i[3] ;
assign n2689 = /* LUT    6 18  3 */ (n567 ? 1'b1 : (n569 ? 1'b1 : n570));
assign n2690 = /* LUT   11 28  1 */ (n130 ? n781 : n338);
assign n406  = /* LUT    3 22  5 */ (n185 ? io_33_1_1 : (n405 ? (io_33_1_1 ? 1'b1 : n402) : io_33_1_1));
assign n2692 = /* LUT    6 17  7 */ (n674 ? (io_33_1_1 ? !n450 : (n676 ? 1'b1 : !n450)) : (io_33_1_1 ? 1'b0 : (n676 ? n450 : 1'b0)));
assign n2693 = /* LUT   10 30  1 */ (n872 ? (n874 ? 1'b1 : n130) : (n874 ? !n130 : 1'b0));
assign n2694 = /* LUT    4 20  6 */ (n496 ? (n382 ? n67 : !n67) : (n382 ? !n67 : n67));
assign n2695 = /* LUT   15 30  3 */ (n1316 ? (n1435 ? 1'b1 : !n675) : (n1435 ? n675 : 1'b0));
assign n2696 = /* LUT    7 25  0 */ (n737 ? (n123 ? 1'b1 : n666) : (n123 ? !n666 : 1'b0));
assign n2697 = /* LUT   12 16  3 */ (io_33_1_1 ? 1'b0 : io_33_14_0);
assign n2698 = /* LUT   14 18  2 */ (io_33_1_1 ? 1'b1 : \wb_dat_i[22] );
assign n2699 = /* LUT   12 29  4 */ (n130 ? n547 : n962);
assign n2700 = /* LUT    1 20  5 */ (n163 ? (io_33_1_1 ? 1'b1 : n184) : n83);
assign n2701 = /* LUT   17 18  1 */ (n807 ? 1'b1 : (n1479 ? 1'b1 : (n1474 ? 1'b1 : n1438)));
assign n2702 = /* LUT    4 23  0 */ (n407 ? (n318 ? 1'b0 : dmarq_pad_i) : (n318 ? 1'b0 : (dmarq_pad_i ? 1'b1 : n238)));
assign n2703 = /* LUT   14 28  7 */ (n1199 ? (n1379 ? 1'b1 : n677) : (n1379 ? !n677 : 1'b0));
assign n2704 = /* LUT    2 22  6 */ (n169 ? n105 : n95);
assign n2705 = /* LUT    6 29  2 */ (n652 ? (io_33_1_1 ? 1'b0 : (n287 ? 1'b1 : n641)) : (io_33_1_1 ? 1'b0 : (n287 ? 1'b0 : n641)));
assign n2706 = /* LUT   11 22  7 */ (n675 ? (n1151 ? 1'b0 : \wb_adr_i[3] ) : (n1051 ? 1'b0 : \wb_adr_i[3] ));
assign n2707 = /* LUT   11 29  6 */ (n234 ? (n780 ? 1'b1 : !n130) : (n780 ? n130 : 1'b0));
assign n2708 = /* LUT   16 20  1 */ (n1114 ? (n1448 ? 1'b1 : (n758 ? 1'b1 : n1393)) : (n1448 ? 1'b1 : n1393));
assign n2709 = /* LUT   15 18  6 */ (\wb_dat_i[11]  ? 1'b1 : io_33_1_1);
assign n2710 = /* LUT    3 23  6 */ (n115 ? (n413 ? !io_33_1_1 : (io_33_1_1 ? 1'b0 : !n287)) : (n413 ? (io_33_1_1 ? 1'b0 : n287) : 1'b0));
assign n999  = /* LUT   10 17  0 */ (n798 ? (n892 ? (n40 ? !n889 : 1'b1) : !n40) : (n892 ? !n889 : 1'b0));
assign n2715 = /* LUT    3 24  4 */ (n118 ? 1'b0 : \wb_dat_i[0] );
assign n2716 = /* LUT    7 30  1 */ (io_33_1_1 ? 1'b1 : \wb_dat_i[19] );
assign n2717 = /* LUT   12 23  2 */ (n708 ? (n1242 ? 1'b1 : (n512 ? n799 : 1'b0)) : (n512 ? n799 : 1'b0));
assign n2718 = /* LUT    5 26  2 */ wb_clk_i;
assign n2719 = /* LUT   11 25  3 */ (n130 ? n828 : n827);
assign n2720 = /* LUT   10 28  6 */ (n130 ? n338 : n781);
assign n2721 = /* LUT    4 22  3 */ (n317 ? !n173 : (n173 ? 1'b0 : !n84));
assign n732  = /* LUT    6 28  1 */ (n75 ? n703 : n582);
assign n2723 = /* LUT   11 23  4 */ \dd_pad_i[15] ;
assign n2724 = /* LUT   11 26  7 */ (n849 ? (n850 ? 1'b1 : !n130) : (n850 ? n130 : 1'b0));
assign n1442 = /* LUT   16 19  0 */ (n1388 ? (n96 ? 1'b1 : (n104 ? n796 : 1'b0)) : (n104 ? n796 : 1'b0));
assign n1391 = /* LUT   15 19  5 */ (n758 ? (n885 ? (n104 ? 1'b1 : n784) : n784) : (n885 ? n104 : 1'b0));
assign n2727 = /* LUT   13 24  1 */ (n526 ? (n633 ? 1'b1 : !n130) : (n633 ? n130 : 1'b0));
assign n2728 = /* LUT    3 20  7 */ (n191 ? (io_33_1_1 ? !n163 : (n200 ? 1'b1 : !n163)) : (io_33_1_1 ? 1'b0 : (n200 ? n163 : 1'b0)));
assign n2729 = /* LUT    2 20  3 */ (n276 ? (io_33_1_1 ? 1'b0 : (n171 ? n174 : 1'b0)) : !io_33_1_1);
assign n2730 = /* LUT    6 19  5 */ \wb_dat_i[21] ;
assign n2731 = /* LUT   10 16  3 */ (\wb_dat_i[21]  ? 1'b1 : io_33_1_1);
assign n2732 = /* LUT   15 28  1 */ (n844 ? (n1371 ? 1'b1 : n666) : (n1371 ? !n666 : 1'b0));
assign n2733 = /* LUT   12 22  1 */ (n1145 ? 1'b1 : (n1238 ? 1'b1 : (n1144 ? 1'b1 : n785)));
assign n2734 = /* LUT    1 22  7 */ (io_33_1_1 ? 1'b0 : \wb_dat_i[30] );
assign n2735 = /* LUT    5 27  5 */ (n125 ? (n313 ? 1'b1 : !n130) : (n313 ? n130 : 1'b0));
assign n2736 = /* LUT   10 31  7 */ (n666 ? n971 : n1103);
assign n2737 = /* LUT    4 21  2 */ (n372 ? (io_33_1_1 ? !n300 : (n399 ? 1'b1 : !n300)) : (io_33_1_1 ? 1'b0 : (n399 ? n300 : 1'b0)));
assign n2738 = /* LUT    2 24  4 */ (n324 ? (n208 ? n67 : !n67) : (n208 ? !n67 : n67));
assign n2739 = /* LUT   14 19  6 */ (io_33_1_1 ? 1'b0 : \dd_pad_i[7] );
assign n2740 = /* LUT   11 20  5 */ (n798 ? (n1141 ? 1'b0 : n1041) : !n1141);
assign n2741 = /* LUT   11 27  4 */ (n130 ? n872 : n874);
assign n549  = /* LUT    4 27  1 */ (n75 ? n533 : n124);
assign n2743 = /* LUT   13 25  2 */ (n130 ? \dd_pad_i[14]  : \dd_pad_i[9] );
assign n2744 = /* LUT   15 15  5 */ (n169 ? n1386 : n1385);
assign n2745 = /* LUT    3 21  0 */ (n363 ? (n96 ? (n104 ? 1'b1 : n317) : n104) : (n96 ? n317 : 1'b0));
assign n2746 = /* LUT    2 23  2 */ (n65 ? (n312 ? (n311 ? !io_33_1_1 : 1'b0) : 1'b1) : (n312 ? (n311 ? !io_33_1_1 : 1'b0) : 1'b0));
assign n2747 = /* LUT   17 24  2 */ wb_cyc_i;
assign n2748 = /* LUT   10 19  2 */ (n587 ? 1'b1 : (n801 ? 1'b1 : !n75));
assign n2749 = /* LUT    7 28  3 */ (n726 ? (n773 ? 1'b1 : !n666) : (n773 ? n666 : 1'b0));
assign n2750 = /* LUT   14 26  6 */ (n130 ? iordy_pad_i : DMA_req);
assign n2751 = /* LUT   12 21  0 */ (io_33_1_1 ? 1'b0 : \wb_dat_i[17] );
assign n2752 = /* LUT    9 27  0 */ (n130 ? n828 : n827);
assign n2753 = /* LUT   14 25  0 */ (n964 ? (n779 ? 1'b1 : n130) : (n779 ? !n130 : 1'b0));
assign n2754 = /* LUT    3 17  5 */ (n148 ? (io_33_1_1 ? !n254 : (n348 ? 1'b1 : !n254)) : (io_33_1_1 ? 1'b0 : (n348 ? n254 : 1'b0)));
assign n2755 = /* LUT    6 21  6 */ (n169 ? n610 : n600);
assign n2756 = /* LUT   11 21  2 */ (n169 ? n1028 : n1042);
assign n2757 = /* LUT   11 24  5 */ (n338 ? (n130 ? n781 : 1'b1) : (n130 ? n781 : 1'b0));
assign n2758 = /* LUT    4 26  2 */ (n118 ? 1'b0 : \wb_dat_i[22] );
assign n2759 = /* LUT   18 19  0 */ (io_33_7_0 ? 1'b0 : (n1486 ? (n1510 ? !io_33_8_0 : 1'b0) : 1'b0));
assign n359  = /* LUT    3 18  1 */ (io_33_1_1 ? 1'b1 : (n358 ? (n356 ? 1'b0 : n263) : !n356));
assign n2760 = /* LUT    5 16  3 */ (n447 ? io_33_1_1 : (io_33_1_1 ? 1'b1 : (n449 ? 1'b0 : !n472)));
assign n2761 = /* LUT   10 25  4 */ (n234 ? (n780 ? 1'b1 : n130) : (n780 ? !n130 : 1'b0));
assign n1014 = /* LUT   10 18  5 */ (n792 ? 1'b0 : (n169 ? 1'b0 : (n896 ? 1'b0 : n692)));
assign n2762 = /* LUT    6 26  4 */ (n130 ? (n415 ? !n630 : (n630 ? 1'b0 : !n376)) : !n630);
assign n2763 = /* LUT   11 17  7 */ (n798 ? (n1118 ? 1'b0 : n462) : !n1118);
assign n2764 = /* LUT    5 29  7 */ (n75 ? n454 : n333);
assign n2765 = /* LUT   16 29  5 */ (n130 ? n962 : n547);
assign n2766 = /* LUT    9 20  1 */ io_33_7_0;
assign n2767 = /* LUT   14 24  3 */ (\wb_adr_i[3]  ? (n1356 ? (n1296 ? 1'b0 : !n675) : (n1296 ? n675 : 1'b1)) : 1'b0);
assign n2768 = /* LUT   11 18  3 */ (n262 ? !n1123 : (n1123 ? 1'b0 : !n798));
assign n2769 = /* LUT    4 25  3 */ \wb_dat_i[8] ;
assign n2770 = /* LUT   10 22  2 */ (n287 ? (n1054 ? 1'b1 : io_33_1_1) : 1'b1);
assign n2771 = /* LUT   15 22  2 */ (io_33_17_0 ? !io_33_1_1 : 1'b0);
assign n2772 = /* LUT   13 27  4 */ (n636 ? (n634 ? 1'b1 : n130) : (n634 ? !n130 : 1'b0));
assign n2773 = /* LUT    3 19  2 */ (n59 ? 1'b1 : (n61 ? 1'b1 : (n60 ? 1'b1 : n57)));
assign n2774 = /* LUT   17 26  0 */ (n1136 ? (n746 ? !n1469 : 1'b0) : (n762 ? 1'b1 : (n746 ? !n1469 : 1'b0)));
assign n2775 = /* LUT    1  7  5 */ !\wb_sel_i[0] ;
assign n2776 = /* LUT    5 17  0 */ \wb_dat_i[0] ;
assign n2777 = /* LUT   10 24  7 */ (n130 ? n526 : n633);
assign n1049 = /* LUT   10 21  4 */ (n892 ? (n916 ? !n1043 : (n798 ? 1'b1 : !n1043)) : (n916 ? 1'b0 : n798));
assign n2779 = /* LUT   14 20  4 */ (n758 ? (n1249 ? (n701 ? 1'b1 : n788) : n788) : (n1249 ? n701 : 1'b0));
assign n2780 = /* LUT   17 20  3 */ (n1129 ? (n96 ? (n104 ? 1'b1 : n1445) : n104) : (n96 ? n1445 : 1'b0));
assign n2781 = /* LUT   11 30  6 */ (n827 ? (n828 ? 1'b1 : n130) : (n828 ? !n130 : 1'b0));
assign n2782 = /* LUT    5 30  6 */ (n555 ? (io_33_1_1 ? 1'b0 : (n287 ? 1'b1 : n645)) : (io_33_1_1 ? 1'b0 : (n287 ? 1'b0 : n645)));
assign n2783 = /* LUT   16 28  2 */ \wb_sel_i[1] ;
assign n1331 = /* LUT   13 31  1 */ (n1265 ? (n1330 ? 1'b1 : n677) : (n1330 ? !n677 : 1'b0));
assign n2785 = /* LUT   14 27  2 */ (n130 ? n769 : n968);
assign n2786 = /* LUT    6 24  5 */ (n119 ? (n417 ? 1'b1 : n130) : (n417 ? !n130 : 1'b0));
assign n1131 = /* LUT   11 19  0 */ (n1129 ? (n755 ? 1'b0 : n893) : (n892 ? 1'b1 : (n755 ? 1'b0 : n893)));
assign n2788 = /* LUT    4 24  4 */ (io_33_14_0 ? !n118 : 1'b0);
assign n1408 = /* LUT   15 23  1 */ (n1027 ? (n1407 ? 1'b1 : (n758 ? 1'b1 : n1348)) : (n1407 ? 1'b1 : n1348));
assign n2790 = /* LUT   13 28  5 */ (n1320 ? (n1261 ? 1'b1 : !n677) : (n1261 ? n677 : 1'b0));
assign n2791 = /* LUT   18 21  6 */ (\wb_adr_i[5]  ? 1'b0 : (\wb_adr_i[3]  ? 1'b0 : \wb_dat_i[2] ));
assign n2792 = /* LUT    5 18  1 */ (n273 ? 1'b1 : (n577 ? 1'b1 : (n452 ? n275 : 1'b1)));
assign n2793 = /* LUT   16 24  7 */ (n1405 ? 1'b1 : (n1402 ? 1'b1 : (n1403 ? 1'b1 : n733)));
assign n2794 = /* LUT   10 20  7 */ (n892 ? (n1032 ? (n1018 ? !n504 : 1'b1) : !n1018) : (n1032 ? !n504 : 1'b0));
assign n2795 = /* LUT   14 23  5 */ (\wb_dat_i[8]  ? !io_33_1_1 : 1'b0);
assign n2796 = /* LUT   17 21  0 */ (n1450 ? 1'b1 : (n305 ? (n465 ? 1'b1 : n701) : n465));
assign n2797 = /* LUT    1 18  3 */ (n158 ? (n155 ? n67 : !n67) : (n155 ? !n67 : n67));
assign n2798 = /* LUT   11 31  5 */ (n677 ? n1217 : n1106);
assign n2799 = /* LUT   16 27  3 */ (n130 ? n874 : n872);
assign n924  = /* LUT    9 22  3 */ (n677 ? n921 : n759);
assign n2801 = /* LUT    6 22  3 */ (n596 ? (n705 ? 1'b0 : (\wb_adr_i[5]  ? 1'b0 : !n17)) : (n705 ? 1'b0 : !n17));
assign n2802 = /* LUT    6 27  4 */ (n130 ? (n723 ? 1'b0 : (n376 ? n229 : 1'b1)) : !n723);
assign n2803 = /* LUT   15 20  0 */ (io_33_1_1 ? 1'b0 : \wb_dat_i[14] );
assign n1513 = /* LUT   18 20  5 */ (n512 ? (n1512 ? 1'b1 : (n1334 ? 1'b1 : n1228)) : (n1512 ? 1'b1 : n1334));
assign n2805 = /* LUT    5 24  7 */ (io_33_19_0 ? !n118 : 1'b0);
assign n2806 = /* LUT    5 19  6 */ (n486 ? (n75 ? 1'b1 : n471) : (n490 ? (n75 ? 1'b1 : n471) : 1'b0));
assign n2807 = /* LUT   10 26  1 */ (n968 ? (n769 ? 1'b1 : n130) : (n769 ? !n130 : 1'b0));
assign n1059 = /* LUT   10 23  6 */ (n677 ? n867 : n112);
assign n2809 = /* LUT    7 21  0 */ (\wb_adr_i[4]  ? !io_33_1_1 : 1'b0);
assign n2810 = /* LUT   14 22  2 */ (\wb_adr_i[5]  ? (n1344 ? (n286 ? 1'b1 : n1288) : n1288) : (n1344 ? n286 : 1'b0));
assign n1494 = /* LUT   17 22  1 */ (n900 ? (n1493 ? 1'b1 : (n1487 ? 1'b1 : n758)) : (n1493 ? 1'b1 : n1487));
assign n2812 = /* LUT   11 28  4 */ (n847 ? (n966 ? 1'b1 : n130) : (n966 ? !n130 : 1'b0));
assign n479  = /* LUT    4 19  0 */ (n275 ? n67 : n361);
assign n2814 = /* LUT    9 28  5 */ (n849 ? (n850 ? 1'b1 : !n130) : (n850 ? n130 : 1'b0));
assign n2815 = /* LUT    9 23  4 */ (n331 ? (n829 ? 1'b1 : !n677) : (n829 ? n677 : 1'b0));
assign n2816 = /* LUT   18 24  6 */ (n817 ? 1'b0 : (n1074 ? 1'b0 : (n1340 ? 1'b0 : !n765)));
assign n2817 = /* LUT    6 17  2 */ (n669 ? (io_33_1_1 ? 1'b1 : (n450 ? n576 : 1'b1)) : (io_33_1_1 ? n450 : (n450 ? n576 : 1'b0)));
assign n2818 = /* LUT   10 30  6 */ (n130 ? n633 : n526);
assign n2819 = /* LUT   13 19  0 */ (n701 ? (n517 ? 1'b1 : io_33_1_1) : io_33_1_1);
assign n2820 = /* LUT   13 30  7 */ (n847 ? (n966 ? 1'b1 : !n130) : (n966 ? n130 : 1'b0));
assign n2824 = /* LUT   18 23  4 */ (io_33_1_1 ? 1'b0 : \wb_dat_i[30] );
assign n2825 = /* LUT   14 18  7 */ (io_33_1_1 ? 1'b0 : io_33_17_0);
assign n2826 = /* LUT   11 15  3 */ (n512 ? (n517 ? 1'b1 : io_33_1_1) : io_33_1_1);
assign n2827 = /* LUT    5 20  7 */ (n509 ? (n474 ? 1'b0 : (n596 ? 1'b0 : !n595)) : 1'b0);
assign n2828 = /* LUT   10 29  0 */ (n130 ? n547 : n962);
assign n2829 = /* LUT   15 27  0 */ (n666 ? n859 : n1370);
assign n2830 = /* LUT    7 26  1 */ (n651 ? (n434 ? 1'b1 : n666) : (n434 ? !n666 : 1'b0));
assign n2831 = /* LUT    9 19  1 */ io_33_7_0;
assign n2832 = /* LUT   12 19  2 */ (n893 ? (n1229 ? 1'b0 : n1137) : !n1229);
assign n2833 = /* LUT   11 29  3 */ (n130 ? n234 : n780);
assign n2834 = /* LUT    4 18  3 */ (n152 ? 1'b0 : (n467 ? (n351 ? n352 : 1'b0) : 1'b0));
assign n2835 = /* LUT    9 29  6 */ (n130 ? n338 : n781);
assign n2836 = /* LUT    9 16  5 */ (n356 ? 1'b0 : (n53 ? n263 : 1'b1));
assign n2837 = /* LUT   18 27  7 */ (n817 ? 1'b0 : (n1413 ? 1'b0 : (n1339 ? 1'b0 : !n1504)));
assign n1463 = /* LUT   16 23  0 */ (n708 ? (n1111 ? (n512 ? 1'b1 : n1295) : n1295) : (n1111 ? n512 : 1'b0));
assign n2839 = /* LUT   10 17  7 */ (n892 ? (n883 ? !n782 : (n893 ? 1'b1 : !n782)) : (n883 ? 1'b0 : n893));
assign n2840 = /* LUT   13 20  1 */ (io_33_1_1 ? 1'b0 : io_33_15_1);
assign n1266 = /* LUT   12 28  0 */ (n666 ? n231 : n1194);
assign n1482 = /* LUT   17 19  3 */ (n1026 ? (n1126 ? (n701 ? 1'b1 : n758) : n701) : (n1126 ? n758 : 1'b0));
assign n2843 = /* LUT    5 26  5 */ io_33_17_0;
assign n2844 = /* LUT    5 21  4 */ (n401 ? 1'b0 : (wb_we_i ? (n509 ? n474 : 1'b0) : 1'b0));
assign n2845 = /* LUT   10 28  3 */ (n337 ? (n131 ? 1'b1 : !n130) : (n131 ? n130 : 1'b0));
assign n2846 = /* LUT   15 24  1 */ (n1341 ? 1'b0 : (n1411 ? 1'b0 : (n1354 ? 1'b0 : !n817)));
assign n2847 = /* LUT    7 27  2 */ (n686 ? (n408 ? (n709 ? 1'b0 : n710) : 1'b0) : 1'b0);
assign n2848 = /* LUT   12 18  1 */ (n1220 ? (n67 ? n357 : !n357) : (n67 ? !n357 : n357));
assign n2849 = /* LUT   11 26  2 */ (n130 ? n719 : n643);
assign n2850 = /* LUT   10 14  0 */ (\wb_adr_i[4]  ? 1'b1 : io_33_1_1);
assign n2851 = /* LUT    9 30  7 */ (n666 ? n852 : n979);
assign n2852 = /* LUT   13 24  4 */ (n130 ? n720 : n764);
assign n2853 = /* LUT    6 19  0 */ io_33_8_0;
assign n2854 = /* LUT   16 22  3 */ (n1039 ? n512 : 1'b0);
assign n2855 = /* LUT   13 21  2 */ (n102 ? (n664 ? (n758 ? 1'b1 : n701) : n701) : (n664 ? n758 : 1'b0));
assign n2856 = /* LUT    2 19  2 */ (n78 ? 1'b1 : n258);
assign n2857 = /* LUT   17 28  2 */ (n446 ? (n1384 ? (n286 ? 1'b1 : \wb_adr_i[5] ) : \wb_adr_i[5] ) : (n1384 ? n286 : 1'b0));
assign n2858 = /* LUT    5 27  2 */ (n130 ? n519 : n415);
assign n2859 = /* LUT    5 22  5 */ (n591 ? (n409 ? 1'b1 : (n410 ? !n317 : 1'b0)) : 1'b0);
assign n2860 = /* LUT   10 31  2 */ (n338 ? (n781 ? 1'b1 : n130) : (n781 ? !n130 : 1'b0));
assign n2861 = /* LUT   15 25  6 */ (n1298 ? (n1364 ? 1'b1 : n677) : (n1364 ? !n677 : 1'b0));
assign n2862 = /* LUT    7 24  3 */ (n118 ? 1'b0 : (n763 ? (n408 ? 1'b0 : n686) : (n408 ? 1'b1 : n686)));
assign n2863 = /* LUT   12 17  0 */ (\wb_adr_i[4]  ? 1'b1 : io_33_1_1);
assign n2864 = /* LUT   14 19  1 */ (io_33_1_1 ? 1'b1 : \wb_dat_i[27] );
assign n2865 = /* LUT   11 27  1 */ (n968 ? (n769 ? 1'b1 : !n130) : (n769 ? n130 : 1'b0));
assign n2866 = /* LUT    4 27  4 */ (n287 ? (n550 ? !io_33_1_1 : 1'b0) : (n548 ? !io_33_1_1 : 1'b0));
assign n2867 = /* LUT    7 14  6 */ (n687 ? n708 : 1'b0);
assign n2868 = /* LUT   13 25  7 */ n779;
assign n2869 = /* LUT   16 21  2 */ (n103 ? (n1452 ? 1'b1 : (n701 ? 1'b1 : n1398)) : (n1452 ? 1'b1 : n1398));
assign n1021 = /* LUT   10 19  5 */ (n692 ? (n1020 ? 1'b1 : (n700 ? 1'b0 : n169)) : (n1020 ? 1'b1 : (n700 ? !n169 : 1'b1)));
assign n1434 = /* LUT   15 29  3 */ (n1081 ? (n666 ? n970 : 1'b1) : (n666 ? n970 : 1'b0));
assign n1293 = /* LUT   13 22  3 */ (\wb_adr_i[5]  ? (n1292 ? (n286 ? 1'b1 : n1236) : n1236) : (n1292 ? n286 : 1'b0));
assign n403  = /* LUT    3 22  1 */ (n204 ? 1'b0 : (n208 ? 1'b0 : (n206 ? 1'b0 : !n207)));
assign n2873 = /* LUT    4 20  2 */ (n492 ? (n380 ? n67 : !n67) : (n380 ? !n67 : n67));
assign n2874 = /* LUT    7 18  5 */ (n452 ? (io_33_1_1 ? 1'b0 : (n219 ? n459 : 1'b1)) : (io_33_1_1 ? 1'b0 : !n219));
assign n2875 = /* LUT    9 27  5 */ (n849 ? (n850 ? 1'b1 : !n130) : (n850 ? n130 : 1'b0));
assign n2876 = /* LUT    7 25  4 */ (n719 ? (n130 ? n643 : 1'b1) : (n130 ? n643 : 1'b0));
assign n2877 = /* LUT    1 20  1 */ (n185 ? !n67 : n67);
assign n2878 = /* LUT   17 18  5 */ (n749 ? (n104 ? 1'b1 : (n1437 ? n96 : 1'b0)) : (n1437 ? n96 : 1'b0));
assign n2879 = /* LUT   11 24  0 */ (n666 ? n1071 : n1060);
assign n2880 = /* LUT    4 26  7 */ (\wb_dat_i[5]  ? !n118 : 1'b0);
assign n2881 = /* LUT    4 23  4 */ (n402 ? 1'b1 : (n176 ? 1'b1 : io_33_1_1));
assign n2882 = /* LUT    9 24  1 */ n633;
assign n2883 = /* LUT   13 26  6 */ (n130 ? \dd_pad_i[10]  : \dd_pad_i[3] );
assign n2884 = /* LUT   14 28  3 */ (n675 ? n1376 : n1378);
assign n2885 = /* LUT    2 22  2 */ (n169 ? n97 : n94);
assign n1150 = /* LUT   11 22  3 */ (n1070 ? (n1148 ? 1'b1 : n666) : (n1148 ? !n666 : 1'b0));
assign n2887 = /* LUT    5 16  6 */ (n452 ? 1'b1 : (n566 ? io_33_1_1 : 1'b1));
assign n2888 = /* LUT   10 18  2 */ (n460 ? (io_33_1_1 ? 1'b0 : n1013) : n1009);
assign n2889 = /* LUT    3 23  2 */ (n317 ? (n411 ? !io_33_1_1 : 1'b0) : (n411 ? (io_33_1_1 ? 1'b0 : n287) : 1'b0));
assign n2890 = /* LUT    2 21  4 */ (n292 ? (n267 ? n67 : !n67) : (n267 ? !n67 : n67));
assign n2891 = /* LUT   12 20  4 */ (wb_clk_i ? !io_33_1_1 : 1'b0);
assign n2892 = /* LUT    3 14  6 */ n141;
assign n2893 = /* LUT    7 19  6 */ (n678 ? (n698 ? (n675 ? !n693 : n693) : 1'b1) : (n698 ? 1'b1 : (n675 ? !n693 : n693)));
assign n2894 = /* LUT    9 20  4 */ io_33_5_0;
assign n2895 = /* LUT   12 23  6 */ (n677 ? n1077 : n1174);
assign n321  = /* CARRY  2 24  0 */ (n185 & 1'b0) | ((n185 | 1'b0) & n1547);
assign n739  = /* CARRY  7 17  0 */ (n273 & 1'b0) | ((n273 | 1'b0) & n1556);
assign n292  = /* CARRY  2 21  3 */ (n193 & n67) | ((n193 | n67) & n291);
assign n326  = /* CARRY  2 24  5 */ (n209 & n67) | ((n209 | n67) & n325);
assign n158  = /* CARRY  1 18  2 */ (n59 & n67) | ((n59 | n67) & n157);
assign n743  = /* CARRY  7 17  4 */ (n570 & n67) | ((n570 | n67) & n742);
assign n250  = /* CARRY  2 17  3 */ (n241 & n67) | ((n241 | n67) & n249);
assign n1226 = /* CARRY 12 18  6 */ (n886 & n67) | ((n886 | n67) & n1225);
assign n494  = /* CARRY  4 20  3 */ (n385 & n67) | ((n385 | n67) & n493);
assign n322  = /* CARRY  2 24  1 */ (n204 & n67) | ((n204 | n67) & n321);
assign n740  = /* CARRY  7 17  1 */ (n567 & n67) | ((n567 | n67) & n739);
assign n253  = /* CARRY  2 17  6 */ (n244 & n67) | ((n244 | n67) & n252);
assign n162  = /* CARRY  1 18  6 */ (n61 & n67) | ((n61 | n67) & n161);
assign n291  = /* CARRY  2 21  2 */ (n151 & n67) | ((n151 | n67) & n290);
assign n1222 = /* CARRY 12 18  2 */ (n475 & n67) | ((n475 | n67) & n1221);
assign n157  = /* CARRY  1 18  1 */ (n56 & n67) | ((n56 | n67) & n156);
assign n744  = /* CARRY  7 17  5 */ (n571 & n67) | ((n571 | n67) & n743);
assign n249  = /* CARRY  2 17  2 */ (n240 & n67) | ((n240 | n67) & n248);
assign n495  = /* CARRY  4 20  4 */ (n67 & n391) | ((n67 | n391) & n494);
assign n295  = /* CARRY  2 21  6 */ (n269 & n67) | ((n269 | n67) & n294);
assign n327  = /* CARRY  2 24  6 */ (n67 & n210) | ((n67 | n210) & n326);
assign n741  = /* CARRY  7 17  2 */ (n568 & n67) | ((n568 | n67) & n740);
assign n161  = /* CARRY  1 18  5 */ (n57 & n67) | ((n57 | n67) & n160);
assign n1223 = /* CARRY 12 18  3 */ (n261 & n67) | ((n261 | n67) & n1222);
assign n491  = /* CARRY  4 20  0 */ (n182 & 1'b0) | ((n182 | 1'b0) & n2277);
assign n323  = /* CARRY  2 24  2 */ (n67 & n206) | ((n67 | n206) & n322);
assign n156  = /* CARRY  1 18  0 */ (n58 & 1'b0) | ((n58 | 1'b0) & n2319);
assign n745  = /* CARRY  7 17  6 */ (n572 & n67) | ((n572 | n67) & n744);
assign n252  = /* CARRY  2 17  5 */ (n243 & n67) | ((n243 | n67) & n251);
assign n1224 = /* CARRY 12 18  4 */ (n52 & n67) | ((n52 | n67) & n1223);
assign n496  = /* CARRY  4 20  5 */ (n381 & n67) | ((n381 | n67) & n495);
assign n290  = /* CARRY  2 21  1 */ (n266 & n67) | ((n266 | n67) & n289);
assign n742  = /* CARRY  7 17  3 */ (n569 & n67) | ((n569 | n67) & n741);
assign n160  = /* CARRY  1 18  4 */ (n60 & n67) | ((n60 | n67) & n159);
assign n248  = /* CARRY  2 17  1 */ (n239 & n67) | ((n239 | n67) & n247);
assign n1220 = /* CARRY 12 18  0 */ (n166 & 1'b0) | ((n166 | 1'b0) & n2542);
assign n492  = /* CARRY  4 20  1 */ (n384 & n67) | ((n384 | n67) & n491);
assign n294  = /* CARRY  2 21  5 */ (n268 & n67) | ((n268 | n67) & n293);
assign n324  = /* CARRY  2 24  3 */ (n207 & n67) | ((n207 | n67) & n323);
assign n251  = /* CARRY  2 17  4 */ (n242 & n67) | ((n242 | n67) & n250);
assign n1225 = /* CARRY 12 18  5 */ (n573 & n67) | ((n573 | n67) & n1224);
assign n497  = /* CARRY  4 20  6 */ (n67 & n382) | ((n67 | n382) & n496);
assign n289  = /* CARRY  2 21  0 */ (n69 & 1'b0) | ((n69 | 1'b0) & n2713);
assign n325  = /* CARRY  2 24  4 */ (n67 & n208) | ((n67 | n208) & n324);
assign n159  = /* CARRY  1 18  3 */ (n67 & n155) | ((n67 | n155) & n158);
assign n247  = /* CARRY  2 17  0 */ (n152 & 1'b0) | ((n152 | 1'b0) & n2823);
assign n1221 = /* CARRY 12 18  1 */ (n357 & n67) | ((n357 | n67) & n1220);
assign n493  = /* CARRY  4 20  2 */ (n67 & n380) | ((n67 | n380) & n492);
assign n293  = /* CARRY  2 21  4 */ (n67 & n267) | ((n67 | n267) & n292);
/* FF  4 25  6 */ always @(posedge \dd_pad_i[11] ) if (n172) n333 <= 1'b0 ? 1'b0 : n1527;
/* FF  4 22  7 */ assign n390 = n1528;
/* FF  9 25  2 */ always @(posedge \dd_pad_i[11] ) if (n429) n433 <= 1'b0 ? 1'b0 : n1529;
/* FF 13 27  1 */ always @(posedge \dd_pad_i[11] ) if (n552) n1254 <= 1'b0 ? 1'b0 : n1530;
/* FF 11 23  0 */ assign n1531 = n1160;
/* FF 16 19  4 */ assign n1532 = n1443;
/* FF 10 21  3 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n343 <= 1'b0 ? 1'b0 : n1533;
/* FF  2 20  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n177 <= 1'b0; else if (1'b1) n177 <= n1534;
/* FF 20 23  7 */ assign wb_err_o = n1535;
/* FF 12 27  5 */ always @(posedge \dd_pad_i[11] ) if (n552) n1190 <= 1'b0 ? 1'b0 : n1536;
/* FF 15 28  5 */ assign n1375 = n1537;
/* FF 13 31  6 */ assign n1279 = n1538;
/* FF 12 22  5 */ assign n1145 = n1539;
/* FF  1 22  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n91 <= 1'b0; else if (n194) n91 <= n1540;
/* FF  4 24  1 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n415 <= 1'b0; else if (n2) n415 <= n1541;
/* FF  4 21  6 */ assign n379 = n1542;
/* FF  9 26  3 */ assign n1543 = n957;
/* FF 13 28  0 */ assign n1261 = n1544;
/* FF  2 24  0 */ assign n1545 = n1546;
/* FF 11 20  1 */ assign n1023 = n1548;
/* FF 16 18  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1228 <= 1'b1; else if (n451) n1228 <= n1549;
/* FF 10 20  0 */ assign n1550 = n1030;
/* FF  3 21  4 */ assign n276 = n393;
/* FF  2 23  6 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n209 <= 1'b0; else if (n113) n209 <= n1551;
/* FF 12 26  6 */ assign n1086 = n1552;
/* FF 17 21  5 */ assign \wb_dat_o[9]  = n1553;
/* FF  7 17  0 */ assign n1554 = n1555;
/* FF  9 22  6 */ always @(posedge \dd_pad_i[11] ) if (n31) n813 <= 1'b0 ? 1'b0 : n1557;
/* FF  7 28  7 */ assign n730 = n1558;
/* FF 14 26  2 */ always @(posedge \dd_pad_i[11] ) if (n1) n781 <= 1'b0 ? 1'b0 : n1559;
/* FF 12 21  4 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1053 <= 1'b0; else if (n4) n1053 <= n1560;
/* FF 13 29  3 */ assign n1561 = n1326;
/* FF  3 17  1 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n239 <= 1'b1; else if (n44) n239 <= n1562;
/* FF 14 25  4 */ assign n1301 = n1563;
/* FF  6 21  2 */ assign n596 = n1564;
/* FF 11 21  6 */ assign n917 = n1565;
/* FF  5 19  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n180 <= 1'b0; else if (1'b1) n180 <= n1566;
/* FF 10 23  1 */ always @(posedge \dd_pad_i[11] ) if (n656) n926 <= 1'b0 ? 1'b0 : n1567;
/* FF 15 26  6 */ assign io_33_28_0 = n1568;
/* FF 15 17  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n462 <= 1'b0; else if (n6) n462 <= n1569;
/* FF  7 21  5 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n303 <= 1'b0; else if (n756) n303 <= n1570;
/* FF  3 18  5 */ assign n255 = n1571;
/* FF 12 25  7 */ assign n1175 = n1572;
/* FF  1 19  1 */ always @(posedge \dd_pad_i[11] ) if (n172) n49 <= 1'b0 ? 1'b0 : n1573;
/* FF 10 25  0 */ assign n841 = n1574;
/* FF  4 19  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n288 <= 1'b0; else if (1'b1) n288 <= n1575;
/* FF  7 22  1 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) resetn_pad_o <= 1'b0; else if (1'b1) resetn_pad_o <= n1576;
/* FF  9 23  1 */ assign n818 = n1577;
/* FF 12 15  2 */ assign n762 = n1578;
/* FF 14 21  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1227 <= 1'b0; else if (n6) n1227 <= n1579;
/* FF  6 26  0 */ always @(posedge \dd_pad_i[11] ) if (n638) n637 <= 1'b0 ? 1'b0 : n1580;
/* FF 11 17  3 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n797 <= 1'b0 ? 1'b0 : n1581;
/* FF 15 21  4 */ assign n1146 = n1582;
/* FF 13 30  2 */ assign n1273 = n1583;
/* FF  2 17  7 */ assign n150 = n1584;
/* FF  6 20  1 */ assign n591 = n695;
/* FF 11 18  7 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n50 <= 1'b0 ? 1'b0 : n1585;
/* FF  5 20  2 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n483 <= 1'b0 ? 1'b0 : n1586;
/* FF 15 27  5 */ always @(posedge \dd_pad_i[11] ) if (n429) n1372 <= 1'b0 ? 1'b0 : n1587;
/* FF 11 32  5 */ always @(posedge \dd_pad_i[11] ) if (n227) n1109 <= 1'b0 ? 1'b0 : n1588;
/* FF 15 22  6 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1167 <= 1'b0; else if (n756) n1167 <= n1589;
/* FF  9 19  6 */ assign n794 = n1590;
/* FF  3 19  6 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n57 <= 1'b0; else if (n62) n57 <= n1591;
/* FF 12 24  0 */ assign n1163 = n1592;
/* FF 17 23  3 */ assign n1460 = n1593;
/* FF 10 24  3 */ assign n939 = n1594;
/* FF  4 18  4 */ assign n1595 = n468;
/* FF  7 23  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n514 <= 1'b0; else if (n329) n514 <= n1596;
/* FF 14 20  0 */ assign n932 = n1597;
/* FF 11 30  2 */ always @(posedge \dd_pad_i[11] ) if (n721) n1100 <= 1'b0 ? 1'b0 : n1598;
/* FF 16 28  6 */ assign n1431 = n1599;
/* FF 14 27  6 */ assign n1309 = n1600;
/* FF 12 28  5 */ assign n1601 = n1268;
/* FF 11 19  4 */ assign n1602 = n1133;
/* FF  5 21  1 */ assign n1603 = n605;
/* FF 15 24  4 */ assign n1352 = n1604;
/* FF 15 23  5 */ assign n1349 = n1605;
/* FF  7 27  7 */ assign n552 = n1606;
/* FF 12 31  1 */ assign n1211 = n1607;
/* FF 17 16  2 */ assign n4 = n1608;
/* FF 22 20  6 */ assign n1285 = n1609;
/* FF  7 20  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n689 <= 1'b0; else if (n194) n689 <= n1610;
/* FF  9 17  3 */ assign n256 = n1611;
/* FF 14 23  1 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n285 <= 1'b0; else if (n194) n285 <= n1612;
/* FF  1 18  7 */ assign n39 = n1613;
/* FF 11 31  1 */ assign n1614 = n1216;
/* FF 16 22  4 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1400 <= 1'b0; else if (n329) n1400 <= n1615;
/* FF 16 27  7 */ assign n1376 = n1616;
/* FF  6 22  7 */ assign n517 = n1617;
/* FF  5 22  0 */ assign n506 = n613;
/* FF 15 25  3 */ assign n1360 = n1618;
/* FF 13 18  3 */ assign n1016 = n1619;
/* FF 15 20  4 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1119 <= 1'b0; else if (n451) n1119 <= n1620;
/* FF  3 26  1 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n330 <= 1'b0; else if (n329) n330 <= n1621;
/* FF 12 30  2 */ always @(posedge \dd_pad_i[11] ) if (n424) n1206 <= 1'b0 ? 1'b0 : n1622;
/* FF  5 24  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n519 <= 1'b0; else if (n2) n519 <= n1623;
/* FF 10 26  5 */ always @(posedge \dd_pad_i[11] ) if (n552) n848 <= 1'b0 ? 1'b0 : n1624;
/* FF  9 18  2 */ assign n588 = n1625;
/* FF 14 29  7 */ assign n1324 = n1626;
/* FF 14 22  6 */ assign n1289 = n1627;
/* FF 11 28  0 */ always @(posedge \dd_pad_i[11] ) if (n227) n775 <= 1'b0 ? 1'b0 : n1628;
/* FF 16 21  5 */ assign n1398 = n1629;
/* FF 16 26  4 */ assign n1630 = n1471;
/* FF  9 28  1 */ always @(posedge \dd_pad_i[11] ) if (n655) n851 <= 1'b0 ? 1'b0 : n1631;
/* FF  3 22  4 */ assign n299 = n405;
/* FF 18 24  2 */ assign \wb_dat_o[11]  = n1632;
/* FF  6 17  6 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n571 <= 1'b0; else if (n346) n571 <= n1633;
/* FF 10 30  2 */ always @(posedge \dd_pad_i[11] ) if (n655) n972 <= 1'b0 ? 1'b0 : n1634;
/* FF  4 20  7 */ assign n374 = n1635;
/* FF 13 19  4 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n699 <= 1'b0; else if (n756) n699 <= n1636;
/* FF 15 30  2 */ assign n1637 = n1435;
/* FF 14 18  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n750 <= 1'b1; else if (n451) n750 <= n1638;
/* FF 12 29  3 */ assign n1199 = n1639;
/* FF  1 20  4 */ assign n68 = n1640;
/* FF 19 25  6 */ assign io_33_27_0 = n1641;
/* FF 17 18  0 */ assign n1642 = n1479;
/* FF  5 25  0 */ always @(posedge \dd_pad_i[11] ) if (n429) n525 <= 1'b0 ? 1'b0 : n1643;
/* FF 10 29  4 */ always @(posedge \dd_pad_i[11] ) if (n227) n970 <= 1'b0 ? 1'b0 : n1644;
/* FF  4 23  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n402 <= 1'b0; else if (1'b1) n402 <= n1645;
/* FF 14 28  4 */ always @(posedge \dd_pad_i[11] ) if (n424) n1314 <= 1'b0 ? 1'b0 : n1646;
/* FF  6 29  5 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) \wb_dat_i[12]  <= 1'b0; else if (1'b1) \wb_dat_i[12]  <= n1647;
/* FF 11 22  6 */ assign n1648 = n1151;
/* FF 11 29  7 */ always @(posedge \dd_pad_i[11] ) if (n655) n977 <= 1'b0 ? 1'b0 : n1649;
/* FF  9 29  2 */ always @(posedge \dd_pad_i[11] ) if (n227) n651 <= 1'b0 ? 1'b0 : n1650;
/* FF 13 23  1 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n114 <= 1'b0 ? 1'b0 : n1651;
/* FF  3 23  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n258 <= 1'b0; else if (1'b1) n258 <= n1652;
/* FF  2 21  3 */ assign n188 = n1653;
/* FF  7 29  6 */ always @(posedge \dd_pad_i[11] ) if (n656) n734 <= 1'b0 ? 1'b0 : n1654;
/* FF 18 27  3 */ assign n1507 = n1655;
/* FF 10 17  3 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n347 <= 1'b0 ? 1'b0 : n1656;
/* FF 13 20  5 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1046 <= 1'b0; else if (n451) n1046 <= n1657;
/* FF  3 24  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n314 <= 1'b0; else if (n2) n314 <= n1658;
/* FF  5 15  6 */ always @(posedge \dd_pad_i[11] ) if (n31) n446 <= 1'b0 ? 1'b0 : n1659;
/* FF  5 26  1 */ always @(posedge \dd_pad_i[11] ) if (n478) n530 <= 1'b0 ? 1'b0 : n1660;
/* FF 11 25  4 */ always @(posedge \dd_pad_i[11] ) if (n552) n953 <= 1'b0 ? 1'b0 : n1661;
/* FF 16 16  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n789 <= 1'b0; else if (n6) n789 <= n1662;
/* FF 10 28  7 */ always @(posedge \dd_pad_i[11] ) if (n655) n774 <= 1'b0 ? 1'b0 : n1663;
/* FF  4 22  0 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n182 <= 1'b1; else if (n298) n182 <= n1664;
/* FF 11 26  6 */ always @(posedge \dd_pad_i[11] ) if (n656) n961 <= 1'b0 ? 1'b0 : n1665;
/* FF 16 19  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1388 <= 1'b0; else if (n329) n1388 <= n1666;
/* FF  9 30  3 */ assign n867 = n1667;
/* FF 13 24  0 */ always @(posedge \dd_pad_i[11] ) if (n424) n1245 <= 1'b0 ? 1'b0 : n1668;
/* FF 15 14  1 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n993 <= 1'b0; else if (n6) n993 <= n1669;
/* FF  3 20  6 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n268 <= 1'b0; else if (n153) n268 <= n1670;
/* FF  2 20  0 */ assign n1671 = n277;
/* FF  6 19  4 */ always @(posedge \dd_pad_i[11] ) if (n172) n582 <= 1'b0 ? 1'b0 : n1672;
/* FF  4 10  6 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n342 <= 1'b0 ? 1'b0 : n1673;
/* FF 10 16  0 */ assign n785 = n1674;
/* FF 15 28  0 */ assign n1325 = n1675;
/* FF 13 21  6 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n507 <= 1'b0 ? 1'b0 : n1676;
/* FF  1 22  6 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n94 <= 1'b0; else if (n194) n94 <= n1677;
/* FF  5 27  6 */ always @(posedge \dd_pad_i[11] ) if (n376) n545 <= 1'b0 ? 1'b0 : n1678;
/* FF 22 16  2 */ assign n6 = n1679;
/* FF 16 31  6 */ assign n738 = n1680;
/* FF  4 21  1 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n380 <= 1'b1; else if (n298) n380 <= n1681;
/* FF  2 24  5 */ assign n215 = n1682;
/* FF 14 19  5 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1128 <= 1'b0; else if (n6) n1128 <= n1683;
/* FF 11 20  4 */ assign n1684 = n1141;
/* FF 11 27  5 */ always @(posedge \dd_pad_i[11] ) if (n429) n1085 <= 1'b0 ? 1'b0 : n1685;
/* FF 13 25  3 */ always @(posedge \dd_pad_i[11] ) if (n1) n538 <= 1'b0 ? 1'b0 : n1686;
/* FF  3 21  1 */ assign n1 = n1687;
/* FF  2 23  1 */ assign n205 = n312;
/* FF 10 19  1 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n75 <= 1'b0; else if (1'b1) n75 <= n1688;
/* FF  7 28  2 */ always @(posedge \dd_pad_i[11] ) if (n721) n726 <= 1'b0 ? 1'b0 : n1689;
/* FF 14 26  7 */ always @(posedge \dd_pad_i[11] ) if (n1) n872 <= 1'b0 ? 1'b0 : n1690;
/* FF 14 15  0 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1005 <= 1'b0; else if (n4) n1005 <= n1691;
/* FF  1 23  1 */ always @(posedge \dd_pad_i[11] ) if (n31) n100 <= 1'b0 ? 1'b0 : n1692;
/* FF  7 18  1 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n677 <= 1'b0; else if (1'b1) n677 <= n1693;
/* FF  9 27  1 */ always @(posedge \dd_pad_i[11] ) if (n227) n839 <= 1'b0 ? 1'b0 : n1694;
/* FF  3 17  6 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n244 <= 1'b0; else if (n44) n244 <= n1695;
/* FF 14 25  3 */ always @(posedge \dd_pad_i[11] ) if (n656) n1300 <= 1'b0 ? 1'b0 : n1696;
/* FF  6 30  0 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) \dd_pad_o[6]  <= 1'b0; else if (1'b1) \dd_pad_o[6]  <= n1697;
/* FF 11 21  3 */ assign n1033 = n1698;
/* FF 11 24  4 */ assign n1062 = n1699;
/* FF  4 26  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n432 <= 1'b0; else if (n2) n432 <= n1700;
/* FF  9 24  5 */ always @(posedge \dd_pad_i[11] ) if (n1) n636 <= 1'b0 ? 1'b0 : n1701;
/* FF  3 18  0 */ assign n53 = n358;
/* FF 18 28  6 */ assign n1702 = n1523;
/* FF 16 15  0 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1386 <= 1'b0; else if (n756) n1386 <= n1703;
/* FF  5 16  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n447 <= 1'b0; else if (1'b1) n447 <= n1704;
/* FF 10 25  7 */ always @(posedge \dd_pad_i[11] ) if (n429) n947 <= 1'b0 ? 1'b0 : n1705;
/* FF 10 18  6 */ assign n888 = n1706;
/* FF 20 27  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n228 <= 1'b0; else if (n329) n228 <= n1707;
/* FF 14 21  6 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1041 <= 1'b0; else if (n6) n1041 <= n1708;
/* FF 12 20  0 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1134 <= 1'b1; else if (n4) n1134 <= n1709;
/* FF  6 26  5 */ always @(posedge \dd_pad_i[11] ) if (n638) n641 <= 1'b0 ? 1'b0 : n1710;
/* FF  7 19  2 */ assign n389 = n753;
/* FF  9 20  0 */ always @(posedge \dd_pad_i[11] ) if (n478) n800 <= 1'b0 ? 1'b0 : n1711;
/* FF 14 24  0 */ assign n1074 = n1712;
/* FF  2  7  4 */ assign n17 = n1713;
/* FF  6 25  1 */ assign n628 = n1714;
/* FF 11 18  2 */ assign n1715 = n1123;
/* FF  4 25  2 */ always @(posedge \dd_pad_i[11] ) if (n172) n422 <= 1'b0 ? 1'b0 : n1716;
/* FF 10 22  3 */ assign n913 = n1717;
/* FF  9 25  6 */ assign n834 = n1718;
/* FF 13 27  5 */ always @(posedge \dd_pad_i[11] ) if (n552) n1258 <= 1'b0 ? 1'b0 : n1719;
/* FF  3 19  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n59 <= 1'b0; else if (n62) n59 <= n1720;
/* FF  5 17  1 */ always @(posedge \dd_pad_i[11] ) if (n478) n454 <= 1'b0 ? 1'b0 : n1721;
/* FF 10 24  4 */ always @(posedge \dd_pad_i[11] ) if (n424) n940 <= 1'b0 ? 1'b0 : n1722;
/* FF 10 21  7 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n365 <= 1'b0 ? 1'b0 : n1723;
/* FF 12 27  1 */ always @(posedge \dd_pad_i[11] ) if (n552) n1186 <= 1'b0 ? 1'b0 : n1724;
/* FF 17 20  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1445 <= 1'b0; else if (n329) n1445 <= n1725;
/* FF 16 28  3 */ assign n1726 = n1477;
/* FF  7 16  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n664 <= 1'b1; else if (n6) n664 <= n1727;
/* FF  9 21  3 */ assign n809 = n1728;
/* FF 13 31  2 */ assign n1277 = n1729;
/* FF 18 22  5 */ assign n1484 = n1730;
/* FF 14 27  1 */ always @(posedge \dd_pad_i[11] ) if (n424) n1304 <= 1'b0 ? 1'b0 : n1731;
/* FF  6 24  2 */ always @(posedge \dd_pad_i[11] ) if (n376) n621 <= 1'b0 ? 1'b0 : n1732;
/* FF 11 19  1 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n1012 <= 1'b0 ? 1'b0 : n1733;
/* FF  4 24  5 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n418 <= 1'b0; else if (n2) n418 <= n1734;
/* FF  9 26  7 */ always @(posedge \dd_pad_i[11] ) if (n638) n233 <= 1'b0 ? 1'b0 : n1735;
/* FF 13 28  4 */ assign n1736 = n1320;
/* FF 18 21  1 */ assign n708 = n1737;
/* FF 17 27  0 */ assign n1470 = n1738;
/* FF  5 18  0 */ assign n458 = n577;
/* FF 10 27  5 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n907 <= 1'b0; else if (n329) n907 <= n1739;
/* FF 10 20  4 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n576 <= 1'b0 ? 1'b0 : n1740;
/* FF 12 26  2 */ always @(posedge \dd_pad_i[11] ) if (n721) n960 <= 1'b0 ? 1'b0 : n1741;
/* FF 17 21  1 */ assign n104 = n1742;
/* FF  1 18  2 */ assign n34 = n1743;
/* FF 16 27  2 */ always @(posedge \dd_pad_i[11] ) if (n656) n1416 <= 1'b0 ? 1'b0 : n1744;
/* FF  7 17  4 */ assign n672 = n1745;
/* FF  9 22  2 */ assign \wb_dat_o[8]  = n1746;
/* FF  6 27  3 */ assign n1747 = n723;
/* FF 13 18  6 */ assign n824 = n1748;
/* FF  5 24  6 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n522 <= 1'b0; else if (n2) n522 <= n1749;
/* FF  5 19  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n474 <= 1'b0; else if (1'b1) n474 <= n1750;
/* FF 10 26  2 */ always @(posedge \dd_pad_i[11] ) if (n552) n942 <= 1'b0 ? 1'b0 : n1751;
/* FF 10 23  5 */ always @(posedge \dd_pad_i[11] ) if (n656) n928 <= 1'b0 ? 1'b0 : n1752;
/* FF  7 21  1 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n102 <= 1'b0; else if (n756) n102 <= n1753;
/* FF 14 22  3 */ assign n1754 = n1345;
/* FF 12 25  3 */ assign n1172 = n1755;
/* FF 17 22  0 */ assign n1756 = n1493;
/* FF  4 19  3 */ assign n361 = n1757;
/* FF  9 28  4 */ always @(posedge \dd_pad_i[11] ) if (n655) n231 <= 1'b0 ? 1'b0 : n1758;
/* FF  9 23  5 */ assign n1759 = n935;
/* FF 10 30  7 */ always @(posedge \dd_pad_i[11] ) if (n655) n731 <= 1'b0 ? 1'b0 : n1760;
/* FF 13 19  1 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n612 <= 1'b0; else if (n756) n612 <= n1761;
/* FF 15 21  0 */ assign n1339 = n1762;
/* FF 13 30  6 */ always @(posedge \dd_pad_i[11] ) if (n656) n1274 <= 1'b0 ? 1'b0 : n1763;
/* FF  2 17  3 */ assign n146 = n1764;
/* FF 10 32  5 */ always @(posedge \dd_pad_i[11] ) if (n655) n987 <= 1'b0 ? 1'b0 : n1765;
/* FF  5 20  6 */ assign n487 = n1766;
/* FF 15 27  1 */ always @(posedge \dd_pad_i[11] ) if (n429) n1370 <= 1'b0 ? 1'b0 : n1767;
/* FF  7 26  0 */ assign n716 = n1768;
/* FF  9 19  2 */ assign n616 = n1769;
/* FF 12 19  5 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n341 <= 1'b0 ? 1'b0 : n1770;
/* FF 12 24  4 */ always @(posedge \dd_pad_i[11] ) if (n424) n1148 <= 1'b0 ? 1'b0 : n1771;
/* FF 16 25  0 */ assign n1413 = n1772;
/* FF  4 18  0 */ assign n349 = n1773;
/* FF 13 23  6 */ assign n1240 = n1774;
/* FF  7 23  6 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n388 <= 1'b0; else if (n329) n388 <= n1775;
/* FF 16 23  3 */ assign n1403 = n1776;
/* FF 10 17  6 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n464 <= 1'b0 ? 1'b0 : n1777;
/* FF 12 28  1 */ assign n1193 = n1778;
/* FF 17 19  4 */ assign \wb_dat_i[3]  = n1779;
/* FF  5 26  4 */ always @(posedge \dd_pad_i[11] ) if (n478) n533 <= 1'b0 ? 1'b0 : n1780;
/* FF  5 21  5 */ assign n501 = n1781;
/* FF 10 28  0 */ always @(posedge \dd_pad_i[11] ) if (n655) n863 <= 1'b0 ? 1'b0 : n1782;
/* FF 15 24  0 */ assign n1783 = n1411;
/* FF  7 27  3 */ assign n429 = n1784;
/* FF 12 18  6 */ assign n1008 = n1785;
/* FF 12 31  5 */ assign n1213 = n1786;
/* FF 12 32  0 */ assign n1787 = n1284;
/* FF  9 30  6 */ assign n825 = n1788;
/* FF 13 24  7 */ always @(posedge \dd_pad_i[11] ) if (n424) n1248 <= 1'b0 ? 1'b0 : n1789;
/* FF  7 20  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n86 <= 1'b0; else if (n194) n86 <= n1790;
/* FF 16 22  0 */ assign n1791 = n1458;
/* FF 10 16  5 */ assign n318 = n1792;
/* FF 13 21  3 */ assign n1232 = n1793;
/* FF  3 25  1 */ always @(posedge \dd_pad_i[11] ) if (n429) n123 <= 1'b0 ? 1'b0 : n1794;
/* FF  5 27  3 */ always @(posedge \dd_pad_i[11] ) if (n376) n542 <= 1'b0 ? 1'b0 : n1795;
/* FF  5 22  4 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n510 <= 1'b0; else if (1'b1) n510 <= n1796;
/* FF 10 31  1 */ always @(posedge \dd_pad_i[11] ) if (n721) n981 <= 1'b0 ? 1'b0 : n1797;
/* FF  7 24  2 */ assign n1798 = n763;
/* FF 12 17  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1114 <= 1'b1; else if (n6) n1114 <= n1799;
/* FF 14 19  0 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1115 <= 1'b1; else if (n6) n1115 <= n1800;
/* FF 12 30  6 */ assign n1203 = n1801;
/* FF  4 27  7 */ assign n438 = n1802;
/* FF 13 25  4 */ always @(posedge \dd_pad_i[11] ) if (n1) n780 <= 1'b0 ? 1'b0 : n1803;
/* FF  9 18  6 */ assign n787 = n1804;
/* FF 14 29  3 */ assign n778 = n1805;
/* FF 16 21  1 */ assign n1806 = n1452;
/* FF 10 19  4 */ assign n896 = n1020;
/* FF 15 29  4 */ assign n1382 = n1807;
/* FF 13 22  2 */ assign n1808 = n1292;
/* FF  3 22  0 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) io_0_6_1 <= 1'b1; else if (1'b1) io_0_6_1 <= n1809;
/* FF  4 20  3 */ assign n370 = n1810;
/* FF  7 18  4 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n377 <= 1'b0; else if (1'b1) n377 <= n1811;
/* FF  9 27  6 */ always @(posedge \dd_pad_i[11] ) if (n227) n826 <= 1'b0 ? 1'b0 : n1812;
/* FF  7 25  5 */ assign n714 = n766;
/* FF 12 16  0 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n799 <= 1'b0; else if (n451) n799 <= n1813;
/* FF 12 29  7 */ always @(posedge \dd_pad_i[11] ) if (n721) n1202 <= 1'b0 ? 1'b0 : n1814;
/* FF  4 26  4 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n335 <= 1'b0; else if (n2) n335 <= n1815;
/* FF  4 23  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) diown_pad_o <= 1'b0; else if (1'b1) diown_pad_o <= n1816;
/* FF  9 24  0 */ always @(posedge \dd_pad_i[11] ) if (n1) n633 <= 1'b0 ? 1'b0 : n1817;
/* FF 13 26  5 */ always @(posedge \dd_pad_i[11] ) if (n1) n547 <= 1'b0 ? 1'b0 : n1818;
/* FF 14 28  0 */ assign n1312 = n1819;
/* FF  2 22  3 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n197 <= 1'b0 ? 1'b0 : n1820;
/* FF 10 18  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n357 <= 1'b0; else if (n563) n357 <= n1821;
/* FF 15 18  5 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1121 <= 1'b1; else if (n4) n1121 <= n1822;
/* FF  3 23  3 */ assign n307 = n412;
/* FF  2 21  7 */ assign n183 = n1823;
/* FF  7 29  2 */ assign n1824 = n777;
/* FF 12 20  5 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n387 <= 1'b0; else if (n4) n387 <= n1825;
/* FF  5 29  1 */ assign n1826 = n660;
/* FF  7 19  7 */ assign n409 = n1827;
/* FF  9 20  7 */ always @(posedge \dd_pad_i[11] ) if (n478) n703 <= 1'b0 ? 1'b0 : n1828;
/* FF  3 24  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n316 <= 1'b0; else if (n2) n316 <= n1829;
/* FF 12 23  1 */ assign io_33_21_0 = n1830;
/* FF 11 25  0 */ always @(posedge \dd_pad_i[11] ) if (n552) n1067 <= 1'b0 ? 1'b0 : n1831;
/* FF  4 25  5 */ always @(posedge \dd_pad_i[11] ) if (n172) n332 <= 1'b0 ? 1'b0 : n1832;
/* FF  4 22  4 */ assign n1833 = n516;
/* FF  9 25  3 */ assign n832 = n1834;
/* FF 13 27  2 */ always @(posedge \dd_pad_i[11] ) if (n552) n1255 <= 1'b0 ? 1'b0 : n1835;
/* FF  6 28  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) \dd_pad_o[14]  <= 1'b0; else if (1'b1) \dd_pad_o[14]  <= n1836;
/* FF 11 23  1 */ assign n1837 = n1161;
/* FF 10 21  2 */ assign n1838 = n1048;
/* FF 15 19  6 */ assign n1336 = n1839;
/* FF  3 20  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n266 <= 1'b0; else if (n153) n266 <= n1840;
/* FF  2 20  4 */ assign n175 = n1841;
/* FF 12 27  4 */ always @(posedge \dd_pad_i[11] ) if (n552) n1189 <= 1'b0 ? 1'b0 : n1842;
/* FF  5 30  0 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) \dd_pad_o[5]  <= 1'b0; else if (1'b1) \dd_pad_o[5]  <= n1843;
/* FF  9 21  4 */ assign n1844 = n909;
/* FF 13 31  7 */ always @(posedge \dd_pad_i[11] ) if (n31) n1280 <= 1'b0 ? 1'b0 : n1845;
/* FF 12 22  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1143 <= 1'b0; else if (n329) n1143 <= n1846;
/* FF  1 22  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n90 <= 1'b0; else if (n194) n90 <= n1847;
/* FF  4 24  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n416 <= 1'b0; else if (n2) n416 <= n1848;
/* FF  4 21  5 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n384 <= 1'b0; else if (n298) n384 <= n1849;
/* FF  9 26  2 */ always @(posedge \dd_pad_i[11] ) if (n638) n230 <= 1'b0 ? 1'b0 : n1850;
/* FF 13 28  3 */ assign n1262 = n1851;
/* FF  2 24  1 */ assign n211 = n1852;
/* FF 11 20  0 */ assign n1022 = n1853;
/* FF 10 20  1 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n264 <= 1'b0 ? 1'b0 : n1854;
/* FF 15 15  6 */ assign n1333 = n1855;
/* FF  3 21  5 */ assign n282 = n1856;
/* FF  2 23  5 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n208 <= 1'b0; else if (n113) n208 <= n1857;
/* FF 20 22  5 */ assign \wb_dat_o[26]  = n1858;
/* FF 12 26  7 */ assign n1087 = n1859;
/* FF 17 24  1 */ assign \wb_dat_i[28]  = n1860;
/* FF  7 17  1 */ assign n669 = n1861;
/* FF  9 22  5 */ assign n812 = n1862;
/* FF  7 28  6 */ always @(posedge \dd_pad_i[11] ) if (n721) n729 <= 1'b0 ? 1'b0 : n1863;
/* FF 14 26  3 */ always @(posedge \dd_pad_i[11] ) if (n1) n338 <= 1'b0 ? 1'b0 : n1864;
/* FF 12 21  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1138 <= 1'b0; else if (n4) n1138 <= n1865;
/* FF 13 29  0 */ always @(posedge \dd_pad_i[11] ) if (n656) n1210 <= 1'b0 ? 1'b0 : n1866;
/* FF 14 25  7 */ assign n1302 = n1867;
/* FF  3 17  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n240 <= 1'b1; else if (n44) n240 <= n1868;
/* FF  6 21  5 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n508 <= 1'b0 ? 1'b0 : n1869;
/* FF 11 21  7 */ assign n1036 = n1870;
/* FF 16 17  5 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n906 <= 1'b0; else if (n329) n906 <= n1871;
/* FF 10 23  0 */ always @(posedge \dd_pad_i[11] ) if (n656) n925 <= 1'b0 ? 1'b0 : n1872;
/* FF 13 15  1 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n221 <= 1'b0; else if (n194) n221 <= n1873;
/* FF 15 17  0 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n40 <= 1'b0; else if (n6) n40 <= n1874;
/* FF  7 21  6 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n697 <= 1'b0; else if (n756) n697 <= n1875;
/* FF 18 19  3 */ assign n1481 = n1876;
/* FF  3 18  4 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n154 <= 1'b0; else if (n62) n154 <= n1877;
/* FF 12 25  6 */ assign n1174 = n1878;
/* FF 17 25  2 */ always @(posedge \dd_pad_i[11] ) if (n31) n1467 <= 1'b0 ? 1'b0 : n1879;
/* FF 10 25  3 */ assign n759 = n1880;
/* FF  4 19  6 */ assign n1881 = n482;
/* FF  7 22  0 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) dd_padoe_o <= 1'b0; else if (1'b1) dd_padoe_o <= n1882;
/* FF  9 23  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n819 <= 1'b0; else if (n329) n819 <= n1883;
/* FF 14 21  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1045 <= 1'b0; else if (n6) n1045 <= n1884;
/* FF  6 26  1 */ assign n638 = n1885;
/* FF 11 17  4 */ assign n1886 = n1117;
/* FF 15 21  5 */ assign n1341 = n1887;
/* FF 13 30  1 */ assign n1888 = n1327;
/* FF  2 17  6 */ assign n149 = n1889;
/* FF 14 24  4 */ assign n1890 = n1357;
/* FF  6 20  6 */ assign n594 = n696;
/* FF  6 25  5 */ assign n631 = n1891;
/* FF 11 18  6 */ assign n1892 = n1124;
/* FF 13 16  0 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n885 <= 1'b0; else if (n4) n885 <= n1893;
/* FF 15 22  1 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n305 <= 1'b0; else if (n756) n305 <= n1894;
/* FF  9 19  7 */ always @(posedge \dd_pad_i[11] ) if (n172) n795 <= 1'b0 ? 1'b0 : n1895;
/* FF 12 24  1 */ always @(posedge \dd_pad_i[11] ) if (n424) n1164 <= 1'b0 ? 1'b0 : n1896;
/* FF 17 26  3 */ assign n1468 = n1897;
/* FF 10 24  0 */ assign n936 = n1898;
/* FF  4 18  5 */ assign n44 = n1899;
/* FF  7 23  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n320 <= 1'b0; else if (n329) n320 <= n1900;
/* FF 11 30  5 */ always @(posedge \dd_pad_i[11] ) if (n721) n1102 <= 1'b0 ? 1'b0 : n1901;
/* FF 16 23  6 */ assign n1406 = n1902;
/* FF 14 27  5 */ always @(posedge \dd_pad_i[11] ) if (n424) n1308 <= 1'b0 ? 1'b0 : n1903;
/* FF 12 28  6 */ assign n1195 = n1904;
/* FF  6 24  6 */ always @(posedge \dd_pad_i[11] ) if (n376) n625 <= 1'b0 ? 1'b0 : n1905;
/* FF 11 19  5 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n271 <= 1'b0 ? 1'b0 : n1906;
/* FF 13 17  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n897 <= 1'b0; else if (n4) n897 <= n1907;
/* FF 15 23  2 */ assign diorn_pad_o = n1908;
/* FF  7 27  4 */ assign n655 = n1909;
/* FF 18 21  5 */ assign n1488 = n1910;
/* FF 12 31  0 */ assign n1911 = n1281;
/* FF  4 17  4 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n78 <= 1'b0; else if (1'b1) n78 <= n1912;
/* FF  7 20  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n688 <= 1'b0; else if (n194) n688 <= n1913;
/* FF  9 17  0 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n574 <= 1'b0 ? 1'b0 : n1914;
/* FF 14 23  0 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n272 <= 1'b0; else if (n194) n272 <= n1915;
/* FF  1 18  6 */ assign n38 = n1916;
/* FF 11 31  6 */ always @(posedge \dd_pad_i[11] ) if (n424) n1108 <= 1'b0 ? 1'b0 : n1917;
/* FF 16 22  5 */ assign n1401 = n1918;
/* FF  2 19  4 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n164 <= 1'b0 ? 1'b0 : n1919;
/* FF  6 22  0 */ assign n595 = n1920;
/* FF  6 27  7 */ always @(posedge \dd_pad_i[11] ) if (n638) n648 <= 1'b0 ? 1'b0 : n1921;
/* FF 13 18  2 */ assign n477 = n1922;
/* FF  7 24  5 */ assign n118 = n1923;
/* FF 18 20  6 */ assign \wb_dat_o[27]  = n1924;
/* FF 12 30  3 */ assign n1207 = n1925;
/* FF  5 24  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n518 <= 1'b0; else if (n2) n518 <= n1926;
/* FF 10 26  6 */ always @(posedge \dd_pad_i[11] ) if (n552) n952 <= 1'b0 ? 1'b0 : n1927;
/* FF  9 18  1 */ assign n1928 = n894;
/* FF 11 28  7 */ always @(posedge \dd_pad_i[11] ) if (n227) n1093 <= 1'b0 ? 1'b0 : n1929;
/* FF 16 21  4 */ assign n1930 = n1453;
/* FF 16 26  5 */ assign n1418 = n1931;
/* FF  9 28  0 */ always @(posedge \dd_pad_i[11] ) if (n655) n658 <= 1'b0 ? 1'b0 : n1932;
/* FF  3 22  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n301 <= 1'b0; else if (1'b1) n301 <= n1933;
/* FF 10 30  3 */ always @(posedge \dd_pad_i[11] ) if (n655) n973 <= 1'b0 ? 1'b0 : n1934;
/* FF 13 19  5 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n610 <= 1'b0; else if (n756) n610 <= n1935;
/* FF  7 25  2 */ always @(posedge \dd_pad_i[11] ) if (n429) n224 <= 1'b0 ? 1'b0 : n1936;
/* FF 14 18  4 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1137 <= 1'b1; else if (n451) n1137 <= n1937;
/* FF 12 29  2 */ always @(posedge \dd_pad_i[11] ) if (n721) n1198 <= 1'b0 ? 1'b0 : n1938;
/* FF  1 20  7 */ assign n71 = n1939;
/* FF  5 25  1 */ always @(posedge \dd_pad_i[11] ) if (n429) n434 <= 1'b0 ? 1'b0 : n1940;
/* FF 10 29  7 */ always @(posedge \dd_pad_i[11] ) if (n227) n537 <= 1'b0 ? 1'b0 : n1941;
/* FF  4 23  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n392 <= 1'b0; else if (1'b1) n392 <= n1942;
/* FF 14 28  5 */ always @(posedge \dd_pad_i[11] ) if (n424) n1315 <= 1'b0 ? 1'b0 : n1943;
/* FF 12 19  1 */ assign n1944 = n1229;
/* FF 11 29  0 */ always @(posedge \dd_pad_i[11] ) if (n655) n1094 <= 1'b0 ? 1'b0 : n1945;
/* FF 16 20  3 */ assign n1393 = n1946;
/* FF 21 19  4 */ assign n1338 = n1947;
/* FF  9 29  3 */ always @(posedge \dd_pad_i[11] ) if (n227) n843 <= 1'b0 ? 1'b0 : n1948;
/* FF 13 23  2 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n109 <= 1'b0 ? 1'b0 : n1949;
/* FF  3 23  4 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n308 <= 1'b0; else if (1'b1) n308 <= n1950;
/* FF  2 21  2 */ assign n170 = n1951;
/* FF  7 29  7 */ always @(posedge \dd_pad_i[11] ) if (n656) n560 <= 1'b0 ? 1'b0 : n1952;
/* FF 18 27  2 */ assign n1953 = n1522;
/* FF  6 16  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n273 <= 1'b0; else if (n346) n273 <= n1954;
/* FF 10 17  2 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n575 <= 1'b0 ? 1'b0 : n1955;
/* FF 13 20  4 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n901 <= 1'b0; else if (n451) n901 <= n1956;
/* FF  3 24  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n119 <= 1'b0; else if (n2) n119 <= n1957;
/* FF  1 21  4 */ assign n83 = n1958;
/* FF  5 26  0 */ always @(posedge \dd_pad_i[11] ) if (n478) n529 <= 1'b0 ? 1'b0 : n1959;
/* FF 11 25  5 */ always @(posedge \dd_pad_i[11] ) if (n552) n1071 <= 1'b0 ? 1'b0 : n1960;
/* FF 10 28  4 */ always @(posedge \dd_pad_i[11] ) if (n655) n955 <= 1'b0 ? 1'b0 : n1961;
/* FF  4 22  1 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n391 <= 1'b1; else if (n298) n391 <= n1962;
/* FF 12 18  2 */ assign n680 = n1963;
/* FF  6 28  7 */ assign n654 = n1964;
/* FF 11 26  1 */ always @(posedge \dd_pad_i[11] ) if (n656) n1076 <= 1'b0 ? 1'b0 : n1965;
/* FF  9 30  2 */ always @(posedge \dd_pad_i[11] ) if (n721) n866 <= 1'b0 ? 1'b0 : n1966;
/* FF 13 24  3 */ always @(posedge \dd_pad_i[11] ) if (n424) n1237 <= 1'b0 ? 1'b0 : n1967;
/* FF  3 20  5 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n267 <= 1'b1; else if (n153) n267 <= n1968;
/* FF  2 20  1 */ assign n171 = n278;
/* FF 18 26  5 */ assign n1504 = n1969;
/* FF  6 19  3 */ always @(posedge \dd_pad_i[11] ) if (n172) n581 <= 1'b0 ? 1'b0 : n1970;
/* FF  1 22  5 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n93 <= 1'b0; else if (n194) n93 <= n1971;
/* FF  5 27  7 */ always @(posedge \dd_pad_i[11] ) if (n376) n546 <= 1'b0 ? 1'b0 : n1972;
/* FF 10 31  5 */ always @(posedge \dd_pad_i[11] ) if (n721) n984 <= 1'b0 ? 1'b0 : n1973;
/* FF  4 21  0 */ assign n79 = n1974;
/* FF 12 17  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1113 <= 1'b1; else if (n6) n1113 <= n1975;
/* FF 14 19  4 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1126 <= 1'b0; else if (n6) n1126 <= n1976;
/* FF 11 27  2 */ always @(posedge \dd_pad_i[11] ) if (n429) n1082 <= 1'b0 ? 1'b0 : n1977;
/* FF  4 27  3 */ assign n1978 = n550;
/* FF 13 25  0 */ always @(posedge \dd_pad_i[11] ) if (n1) n850 <= 1'b0 ? 1'b0 : n1979;
/* FF  3 21  2 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n280 <= 1'b0 ? 1'b0 : n1980;
/* FF  2 23  0 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n204 <= 1'b0; else if (n113) n204 <= n1981;
/* FF 10 19  0 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) \wb_dat_i[29]  <= 1'b0; else if (1'b1) \wb_dat_i[29]  <= n1982;
/* FF 15 29  0 */ assign n1380 = n1983;
/* FF 13 22  6 */ always @(posedge \dd_pad_i[11] ) if (n31) n1236 <= 1'b0 ? 1'b0 : n1984;
/* FF  7 28  1 */ always @(posedge \dd_pad_i[11] ) if (n721) n725 <= 1'b0 ? 1'b0 : n1985;
/* FF  1 23  2 */ always @(posedge \dd_pad_i[11] ) if (n31) n101 <= 1'b0 ? 1'b0 : n1986;
/* FF  7 18  0 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n666 <= 1'b0; else if (1'b1) n666 <= n1987;
/* FF  9 27  2 */ always @(posedge \dd_pad_i[11] ) if (n227) n440 <= 1'b0 ? 1'b0 : n1988;
/* FF 14 25  2 */ always @(posedge \dd_pad_i[11] ) if (n656) n1299 <= 1'b0 ? 1'b0 : n1989;
/* FF  3 17  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n245 <= 1'b0; else if (n44) n245 <= n1990;
/* FF 11 24  3 */ assign n112 = n1991;
/* FF  4 26  0 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n430 <= 1'b0; else if (n2) n430 <= n1992;
/* FF  9 24  4 */ always @(posedge \dd_pad_i[11] ) if (n1) n634 <= 1'b0 ? 1'b0 : n1993;
/* FF 13 26  1 */ always @(posedge \dd_pad_i[11] ) if (n1) n847 <= 1'b0 ? 1'b0 : n1994;
/* FF  3 18  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n61 <= 1'b0; else if (n62) n61 <= n1995;
/* FF 18 28  7 */ assign \wb_dat_o[19]  = n1996;
/* FF  5 16  5 */ assign n219 = n566;
/* FF 10 25  6 */ assign n768 = n1997;
/* FF 10 18  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n52 <= 1'b1; else if (n563) n52 <= n1998;
/* FF 12 20  1 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1135 <= 1'b1; else if (n4) n1135 <= n1999;
/* FF  6 26  6 */ always @(posedge \dd_pad_i[11] ) if (n638) n553 <= 1'b0 ? 1'b0 : n2000;
/* FF  5 29  5 */ assign n556 = n2001;
/* FF  7 19  3 */ assign n73 = n2002;
/* FF  9 20  3 */ always @(posedge \dd_pad_i[11] ) if (n478) n802 <= 1'b0 ? 1'b0 : n2003;
/* FF 12 23  5 */ always @(posedge \dd_pad_i[11] ) if (n31) n1153 <= 1'b0 ? 1'b0 : n2004;
/* FF  6 25  0 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n220 <= 1'b0; else if (n113) n220 <= n2005;
/* FF 10 22  4 */ assign n2006 = n1055;
/* FF  9 25  7 */ always @(posedge \dd_pad_i[11] ) if (n429) n835 <= 1'b0 ? 1'b0 : n2007;
/* FF 13 27  6 */ always @(posedge \dd_pad_i[11] ) if (n552) n1259 <= 1'b0 ? 1'b0 : n2008;
/* FF  3 19  0 */ assign n2009 = n367;
/* FF 16 14  0 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1385 <= 1'b0; else if (n194) n1385 <= n2010;
/* FF 10 24  5 */ always @(posedge \dd_pad_i[11] ) if (n424) n933 <= 1'b0 ? 1'b0 : n2011;
/* FF 10 21  6 */ assign n2012 = n1050;
/* FF 15 19  2 */ assign n2013 = n1390;
/* FF 12 27  0 */ always @(posedge \dd_pad_i[11] ) if (n552) n1185 <= 1'b0 ? 1'b0 : n2014;
/* FF 17 20  5 */ assign n1447 = n2015;
/* FF  2 11  6 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n141 <= 1'b0 ? 1'b0 : n2016;
/* FF  9 21  0 */ assign n807 = n2017;
/* FF 13 31  3 */ assign n2018 = n1332;
/* FF 18 22  6 */ assign n286 = n1517;
/* FF 14 27  0 */ assign n1303 = n2019;
/* FF  6 24  3 */ always @(posedge \dd_pad_i[11] ) if (n376) n622 <= 1'b0 ? 1'b0 : n2020;
/* FF  4 24  6 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n328 <= 1'b0; else if (n2) n328 <= n2021;
/* FF  9 26  6 */ assign n2022 = n958;
/* FF 13 28  7 */ always @(posedge \dd_pad_i[11] ) if (n656) n1265 <= 1'b0 ? 1'b0 : n2023;
/* FF 18 21  0 */ assign n1485 = n2024;
/* FF 10 27  4 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n959 <= 1'b0; else if (n329) n959 <= n2025;
/* FF 10 20  5 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n85 <= 1'b0 ? 1'b0 : n2026;
/* FF  3 30  0 */ always @(posedge \dd_pad_i[11] ) if (n1) n337 <= 1'b0 ? 1'b0 : n2027;
/* FF 12 26  3 */ assign n649 = n2028;
/* FF 17 21  6 */ assign n512 = n2029;
/* FF  1 18  1 */ assign n33 = n2030;
/* FF  7 17  5 */ assign n673 = n2031;
/* FF  9 22  1 */ assign n2032 = n923;
/* FF  6 27  2 */ always @(posedge \dd_pad_i[11] ) if (n638) n645 <= 1'b0 ? 1'b0 : n2033;
/* FF 13 18  5 */ assign n1219 = n2034;
/* FF 13 29  4 */ assign n1271 = n2035;
/* FF  6 21  1 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n311 <= 1'b0 ? 1'b0 : n2036;
/* FF  5 19  0 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) \da_pad_o[2]  <= 1'b0; else if (1'b1) \da_pad_o[2]  <= n2037;
/* FF 10 26  3 */ always @(posedge \dd_pad_i[11] ) if (n552) n951 <= 1'b0 ? 1'b0 : n2038;
/* FF 10 23  4 */ assign n927 = n2039;
/* FF 15 26  5 */ assign n2040 = n1420;
/* FF  7 21  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n107 <= 1'b0; else if (n756) n107 <= n2041;
/* FF 12 25  2 */ always @(posedge \dd_pad_i[11] ) if (n721) n1171 <= 1'b0 ? 1'b0 : n2042;
/* FF  4 19  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) dmackn_pad_o <= 1'b1; else if (1'b1) dmackn_pad_o <= n2043;
/* FF  9 23  6 */ assign \wb_dat_o[18]  = n2044;
/* FF 18 24  4 */ assign n2045 = n1521;
/* FF 11 17  0 */ assign n2046 = n1116;
/* FF  5 23  5 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n420 <= 1'b0; else if (n451) n420 <= n2047;
/* FF 13 19  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n904 <= 1'b0; else if (n756) n904 <= n2048;
/* FF 13 30  5 */ assign n561 = n2049;
/* FF  2 17  2 */ assign n145 = n2050;
/* FF 18 23  2 */ assign \wb_dat_o[31]  = n2051;
/* FF  6 20  2 */ assign n257 = n2052;
/* FF  5 20  1 */ assign n2053 = n597;
/* FF 10 29  2 */ always @(posedge \dd_pad_i[11] ) if (n227) n954 <= 1'b0 ? 1'b0 : n2054;
/* FF 15 27  6 */ always @(posedge \dd_pad_i[11] ) if (n429) n1355 <= 1'b0 ? 1'b0 : n2055;
/* FF 15 22  5 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1249 <= 1'b0; else if (n756) n1249 <= n2056;
/* FF  7 26  3 */ assign n718 = n2057;
/* FF  9 19  3 */ assign n2058 = n898;
/* FF 12 19  4 */ assign n2059 = n1230;
/* FF 12 24  5 */ assign n2060 = n1251;
/* FF 17 23  0 */ assign n2061 = n1499;
/* FF  4 18  1 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n263 <= 1'b0; else if (1'b1) n263 <= n2062;
/* FF  9 29  4 */ always @(posedge \dd_pad_i[11] ) if (n227) n859 <= 1'b0 ? 1'b0 : n2063;
/* FF 13 23  7 */ assign n1241 = n2064;
/* FF  7 23  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n707 <= 1'b0; else if (n329) n707 <= n2065;
/* FF 11 30  1 */ always @(posedge \dd_pad_i[11] ) if (n721) n1099 <= 1'b0 ? 1'b0 : n2066;
/* FF 13 20  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n902 <= 1'b0; else if (n451) n902 <= n2067;
/* FF 12 28  2 */ always @(posedge \dd_pad_i[11] ) if (n721) n1194 <= 1'b0 ? 1'b0 : n2068;
/* FF 17 19  5 */ assign n1441 = n2069;
/* FF  5 21  2 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n498 <= 1'b0 ? 1'b0 : n2070;
/* FF 10 28  1 */ always @(posedge \dd_pad_i[11] ) if (n655) n659 <= 1'b0 ? 1'b0 : n2071;
/* FF  7 27  0 */ assign n2072 = n770;
/* FF 12 18  7 */ assign n1009 = n2073;
/* FF 12 31  4 */ assign n1212 = n2074;
/* FF 12 32  1 */ assign n136 = n2075;
/* FF 16 24  0 */ assign n1409 = n2076;
/* FF  9 30  5 */ always @(posedge \dd_pad_i[11] ) if (n721) n869 <= 1'b0 ? 1'b0 : n2077;
/* FF 13 24  6 */ always @(posedge \dd_pad_i[11] ) if (n424) n1183 <= 1'b0 ? 1'b0 : n2078;
/* FF  7 20  6 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n601 <= 1'b0; else if (n194) n601 <= n2079;
/* FF 11 31  2 */ assign n663 = n2080;
/* FF 16 22  1 */ assign n1155 = n2081;
/* FF  6 22  4 */ assign wb_rty_o = n2082;
/* FF 17 28  4 */ assign n1475 = n2083;
/* FF  5 22  3 */ assign n490 = n2084;
/* FF 10 31  0 */ assign n980 = n2085;
/* FF 15 25  0 */ assign n2086 = n1417;
/* FF  3  7  7 */ assign n237 = n2087;
/* FF 15 20  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n504 <= 1'b0; else if (n451) n504 <= n2088;
/* FF  7 24  1 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n709 <= 1'b0; else if (1'b1) n709 <= n2089;
/* FF 12 17  6 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1004 <= 1'b1; else if (n6) n1004 <= n2090;
/* FF 12 30  7 */ always @(posedge \dd_pad_i[11] ) if (n424) n1209 <= 1'b0 ? 1'b0 : n2091;
/* FF 13 25  5 */ always @(posedge \dd_pad_i[11] ) if (n1) n234 <= 1'b0 ? 1'b0 : n2092;
/* FF 14 29  2 */ always @(posedge \dd_pad_i[11] ) if (n429) n1321 <= 1'b0 ? 1'b0 : n2093;
/* FF 11 28  3 */ always @(posedge \dd_pad_i[11] ) if (n227) n862 <= 1'b0 ? 1'b0 : n2094;
/* FF 16 21  0 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1395 <= 1'b0; else if (n329) n1395 <= n2095;
/* FF 13 22  1 */ assign n2096 = n1291;
/* FF  3 22  3 */ assign n298 = n2097;
/* FF  6 17  5 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n570 <= 1'b0; else if (n346) n570 <= n2098;
/* FF  4 20  4 */ assign n371 = n2099;
/* FF  7 18  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n505 <= 1'b0; else if (1'b1) n505 <= n2100;
/* FF  9 27  7 */ always @(posedge \dd_pad_i[11] ) if (n227) n846 <= 1'b0 ? 1'b0 : n2101;
/* FF  7 25  6 */ assign n2 = n2102;
/* FF 12 16  1 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n790 <= 1'b0; else if (n451) n790 <= n2103;
/* FF 14 18  0 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1029 <= 1'b1; else if (n451) n1029 <= n2104;
/* FF 12 29  6 */ assign n1147 = n2105;
/* FF  1 20  3 */ assign n67 = n186;
/* FF  4 26  5 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n125 <= 1'b0; else if (n2) n125 <= n2106;
/* FF  4 23  6 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n408 <= 1'b0; else if (1'b1) n408 <= n2107;
/* FF  9 24  3 */ always @(posedge \dd_pad_i[11] ) if (n1) n827 <= 1'b0 ? 1'b0 : n2108;
/* FF 13 26  4 */ always @(posedge \dd_pad_i[11] ) if (n1) n962 <= 1'b0 ? 1'b0 : n2109;
/* FF 14 28  1 */ assign n2110 = n1377;
/* FF  2 22  4 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n198 <= 1'b0 ? 1'b0 : n2111;
/* FF 11 22  5 */ assign n748 = n2112;
/* FF 11 29  4 */ always @(posedge \dd_pad_i[11] ) if (n655) n976 <= 1'b0 ? 1'b0 : n2113;
/* FF 15 18  4 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n749 <= 1'b1; else if (n4) n749 <= n2114;
/* FF  3 23  0 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n287 <= 1'b0; else if (1'b1) n287 <= n2115;
/* FF  2 21  6 */ assign n191 = n2116;
/* FF  7 29  3 */ assign n733 = n2117;
/* FF 12 20  6 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1130 <= 1'b0; else if (n4) n1130 <= n2118;
/* FF  7 19  4 */ assign n2119 = n754;
/* FF  9 20  6 */ always @(posedge \dd_pad_i[11] ) if (n478) n618 <= 1'b0 ? 1'b0 : n2120;
/* FF  3 24  6 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n223 <= 1'b0; else if (n2) n223 <= n2121;
/* FF 12 23  0 */ assign n2122 = n1243;
/* FF 11 25  1 */ always @(posedge \dd_pad_i[11] ) if (n552) n1068 <= 1'b0 ? 1'b0 : n2123;
/* FF  4 25  4 */ always @(posedge \dd_pad_i[11] ) if (n172) n225 <= 1'b0 ? 1'b0 : n2124;
/* FF  4 22  5 */ assign n396 = n2125;
/* FF  9 25  0 */ assign n767 = n2126;
/* FF 13 27  3 */ always @(posedge \dd_pad_i[11] ) if (n552) n1256 <= 1'b0 ? 1'b0 : n2127;
/* FF  6 28  3 */ assign n652 = n2128;
/* FF 11 23  6 */ assign n1057 = n2129;
/* FF 11 26  5 */ always @(posedge \dd_pad_i[11] ) if (n656) n1078 <= 1'b0 ? 1'b0 : n2130;
/* FF  2 20  5 */ assign n153 = n2131;
/* FF 12 27  7 */ always @(posedge \dd_pad_i[11] ) if (n552) n1191 <= 1'b0 ? 1'b0 : n2132;
/* FF  6 19  7 */ always @(posedge \dd_pad_i[11] ) if (n172) n585 <= 1'b0 ? 1'b0 : n2133;
/* FF 15 28  3 */ assign n1374 = n2134;
/* FF  9 21  5 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n169 <= 1'b0 ? 1'b0 : n2135;
/* FF  7 31  4 */ always @(posedge \dd_pad_i[11] ) if (n227) n737 <= 1'b0 ? 1'b0 : n2136;
/* FF 12 22  3 */ assign n1144 = n2137;
/* FF  4 24  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n129 <= 1'b0; else if (n2) n129 <= n2138;
/* FF  4 21  4 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n383 <= 1'b0; else if (n298) n383 <= n2139;
/* FF  9 26  1 */ assign n2140 = n956;
/* FF 13 28  2 */ assign n2141 = n1319;
/* FF  2 24  6 */ assign n216 = n2142;
/* FF 11 20  7 */ assign n1025 = n2143;
/* FF 17 27  6 */ assign n1432 = n2144;
/* FF 11 27  6 */ always @(posedge \dd_pad_i[11] ) if (n429) n855 <= 1'b0 ? 1'b0 : n2145;
/* FF  3 21  6 */ assign n283 = n2146;
/* FF  2 23  4 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n207 <= 1'b0; else if (n113) n207 <= n2147;
/* FF 12 26  4 */ always @(posedge \dd_pad_i[11] ) if (n721) n1180 <= 1'b0 ? 1'b0 : n2148;
/* FF 17 24  0 */ assign n2149 = n1502;
/* FF  7 17  2 */ assign n670 = n2150;
/* FF  9 22  4 */ assign n811 = n2151;
/* FF  7 28  5 */ always @(posedge \dd_pad_i[11] ) if (n721) n728 <= 1'b0 ? 1'b0 : n2152;
/* FF 14 26  4 */ always @(posedge \dd_pad_i[11] ) if (n1) n874 <= 1'b0 ? 1'b0 : n2153;
/* FF 12 21  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n915 <= 1'b0; else if (n4) n915 <= n2154;
/* FF 19 20  0 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n386 <= 1'b0; else if (n4) n386 <= n2155;
/* FF 13 29  1 */ always @(posedge \dd_pad_i[11] ) if (n656) n1269 <= 1'b0 ? 1'b0 : n2156;
/* FF 12 11  1 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1110 <= 1'b0; else if (n4) n1110 <= n2157;
/* FF 14 25  6 */ assign n2158 = n1366;
/* FF  3 17  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n241 <= 1'b0; else if (n44) n241 <= n2159;
/* FF  6 21  4 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n302 <= 1'b0 ? 1'b0 : n2160;
/* FF 11 24  7 */ assign n837 = n2161;
/* FF 15 17  1 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n998 <= 1'b0; else if (n6) n998 <= n2162;
/* FF  7 21  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n611 <= 1'b0; else if (n756) n611 <= n2163;
/* FF  3 18  7 */ assign n62 = n2164;
/* FF 12 25  5 */ assign n1173 = n2165;
/* FF  5 16  1 */ assign n2166 = n565;
/* FF 10 25  2 */ always @(posedge \dd_pad_i[11] ) if (n429) n945 <= 1'b0 ? 1'b0 : n2167;
/* FF  9 23  3 */ assign n820 = n2168;
/* FF 14 21  5 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1027 <= 1'b0; else if (n6) n1027 <= n2169;
/* FF  6 26  2 */ always @(posedge \dd_pad_i[11] ) if (n638) n639 <= 1'b0 ? 1'b0 : n2170;
/* FF 11 17  5 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n996 <= 1'b0 ? 1'b0 : n2171;
/* FF 15 21  6 */ assign n1342 = n2172;
/* FF 13 30  0 */ assign n1272 = n2173;
/* FF 14 24  5 */ assign n1296 = n2174;
/* FF  6 20  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n319 <= 1'b0; else if (1'b1) n319 <= n2175;
/* FF  6 25  4 */ assign n630 = n2176;
/* FF 11 18  1 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n681 <= 1'b0 ? 1'b0 : n2177;
/* FF 10 22  0 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) \wb_dat_o[24]  <= 1'b0; else if (1'b1) \wb_dat_o[24]  <= n2178;
/* FF 15 22  0 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1028 <= 1'b0; else if (n756) n1028 <= n2179;
/* FF  3 19  4 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n60 <= 1'b0; else if (n62) n60 <= n2180;
/* FF 12 24  2 */ assign n2181 = n1250;
/* FF  5 17  2 */ always @(posedge \dd_pad_i[11] ) if (n478) n455 <= 1'b0 ? 1'b0 : n2182;
/* FF 10 24  1 */ always @(posedge \dd_pad_i[11] ) if (n424) n937 <= 1'b0 ? 1'b0 : n2183;
/* FF  7 23  0 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n706 <= 1'b1; else if (n329) n706 <= n2184;
/* FF 11 30  4 */ always @(posedge \dd_pad_i[11] ) if (n721) n986 <= 1'b0 ? 1'b0 : n2185;
/* FF 16 28  0 */ assign n2186 = n1476;
/* FF 18 22  2 */ assign n2187 = n1516;
/* FF 14 27  4 */ always @(posedge \dd_pad_i[11] ) if (n424) n1307 <= 1'b0 ? 1'b0 : n2188;
/* FF 12 28  7 */ assign n1192 = n2189;
/* FF  6 24  7 */ always @(posedge \dd_pad_i[11] ) if (n376) n626 <= 1'b0 ? 1'b0 : n2190;
/* FF 11 19  2 */ assign n2191 = n1132;
/* FF 13 17  0 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n889 <= 1'b0; else if (n4) n889 <= n2192;
/* FF 15 23  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1347 <= 1'b0; else if (n329) n1347 <= n2193;
/* FF  7 27  5 */ assign n656 = n2194;
/* FF 18 21  4 */ assign n1487 = n2195;
/* FF 12 31  3 */ assign n2196 = n1283;
/* FF  5 18  3 */ assign n460 = n2197;
/* FF 10 27  0 */ assign n329 = n2198;
/* FF  7 20  1 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n687 <= 1'b0; else if (n194) n687 <= n2199;
/* FF  9 17  1 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n353 <= 1'b0 ? 1'b0 : n2200;
/* FF 14 23  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1295 <= 1'b0; else if (n194) n1295 <= n2201;
/* FF 17 21  2 */ assign n1450 = n2202;
/* FF  1 18  5 */ assign n37 = n2203;
/* FF 11 31  7 */ always @(posedge \dd_pad_i[11] ) if (n424) n948 <= 1'b0 ? 1'b0 : n2204;
/* FF 16 27  1 */ always @(posedge \dd_pad_i[11] ) if (n656) n1422 <= 1'b0 ? 1'b0 : n2205;
/* FF  6 22  1 */ assign n606 = n704;
/* FF  6 27  6 */ always @(posedge \dd_pad_i[11] ) if (n638) n647 <= 1'b0 ? 1'b0 : n2206;
/* FF 11 16  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n991 <= 1'b0; else if (n4) n991 <= n2207;
/* FF  9 13  7 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n203 <= 1'b0 ? 1'b0 : n2208;
/* FF 15 20  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n903 <= 1'b0; else if (n451) n903 <= n2209;
/* FF  7 24  4 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n710 <= 1'b0; else if (1'b1) n710 <= n2210;
/* FF 18 20  7 */ assign n758 = n2211;
/* FF 12 30  0 */ assign n1204 = n2212;
/* FF  5 24  5 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n521 <= 1'b0; else if (n2) n521 <= n2213;
/* FF  5 19  4 */ assign n471 = n590;
/* FF 10 26  7 */ always @(posedge \dd_pad_i[11] ) if (n552) n830 <= 1'b0 ? 1'b0 : n2214;
/* FF 15 26  1 */ assign n1368 = n2215;
/* FF  9 18  0 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n476 <= 1'b0; else if (n346) n476 <= n2216;
/* FF 14 22  0 */ assign n2217 = n1343;
/* FF  6 18  6 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n475 <= 1'b1; else if (n563) n475 <= n2218;
/* FF 17 22  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1455 <= 1'b0; else if (n329) n1455 <= n2219;
/* FF 11 28  6 */ always @(posedge \dd_pad_i[11] ) if (n227) n1088 <= 1'b0 ? 1'b0 : n2220;
/* FF  9 28  3 */ always @(posedge \dd_pad_i[11] ) if (n655) n853 <= 1'b0 ? 1'b0 : n2221;
/* FF  3 22  6 */ assign n300 = n2222;
/* FF 10 30  4 */ always @(posedge \dd_pad_i[11] ) if (n655) n969 <= 1'b0 ? 1'b0 : n2223;
/* FF 13 19  6 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n650 <= 1'b0; else if (n756) n650 <= n2224;
/* FF  7 25  3 */ assign n331 = n2225;
/* FF 14 18  5 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1037 <= 1'b1; else if (n451) n1037 <= n2226;
/* FF 12 29  1 */ always @(posedge \dd_pad_i[11] ) if (n721) n1197 <= 1'b0 ? 1'b0 : n2227;
/* FF  1 20  6 */ assign n70 = n2228;
/* FF  5 20  5 */ assign n486 = n2229;
/* FF 10 29  6 */ always @(posedge \dd_pad_i[11] ) if (n227) n135 <= 1'b0 ? 1'b0 : n2230;
/* FF 15 27  2 */ always @(posedge \dd_pad_i[11] ) if (n429) n1371 <= 1'b0 ? 1'b0 : n2231;
/* FF 12 19  0 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n43 <= 1'b0 ? 1'b0 : n2232;
/* FF 14 17  1 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n891 <= 1'b0; else if (n451) n891 <= n2233;
/* FF  6 29  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) \dd_pad_o[8]  <= 1'b0; else if (1'b1) \dd_pad_o[8]  <= n2234;
/* FF 11 29  1 */ always @(posedge \dd_pad_i[11] ) if (n655) n1095 <= 1'b0 ? 1'b0 : n2235;
/* FF 16 25  3 */ assign n1415 = n2236;
/* FF  9 29  0 */ always @(posedge \dd_pad_i[11] ) if (n227) n857 <= 1'b0 ? 1'b0 : n2237;
/* FF 13 23  3 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n110 <= 1'b0 ? 1'b0 : n2238;
/* FF  3 23  5 */ assign n2239 = n413;
/* FF  1 27  4 */ always @(posedge \dd_pad_i[11] ) if (n172) n124 <= 1'b0 ? 1'b0 : n2240;
/* FF 10 17  5 */ assign n2241 = n1000;
/* FF 13 20  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n919 <= 1'b0; else if (n451) n919 <= n2242;
/* FF  3 24  1 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n313 <= 1'b0; else if (n2) n313 <= n2243;
/* FF  1 21  5 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n84 <= 1'b0 ? 1'b0 : n2244;
/* FF 17 19  1 */ assign n1439 = n2245;
/* FF  5 26  7 */ always @(posedge \dd_pad_i[11] ) if (n478) n536 <= 1'b0 ? 1'b0 : n2246;
/* FF 11 25  6 */ always @(posedge \dd_pad_i[11] ) if (n552) n1072 <= 1'b0 ? 1'b0 : n2247;
/* FF  5 21  6 */ assign n488 = n2248;
/* FF 10 28  5 */ always @(posedge \dd_pad_i[11] ) if (n655) n232 <= 1'b0 ? 1'b0 : n2249;
/* FF 15 24  3 */ assign n2250 = n1412;
/* FF 12 18  3 */ assign n586 = n2251;
/* FF 11 26  0 */ always @(posedge \dd_pad_i[11] ) if (n656) n1075 <= 1'b0 ? 1'b0 : n2252;
/* FF  9 30  1 */ always @(posedge \dd_pad_i[11] ) if (n721) n865 <= 1'b0 ? 1'b0 : n2253;
/* FF 13 24  2 */ always @(posedge \dd_pad_i[11] ) if (n424) n1246 <= 1'b0 ? 1'b0 : n2254;
/* FF  3 20  4 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n193 <= 1'b0; else if (n153) n193 <= n2255;
/* FF 12 13  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n877 <= 1'b0; else if (n194) n877 <= n2256;
/* FF 18 26  6 */ assign n1505 = n2257;
/* FF  6 19  2 */ always @(posedge \dd_pad_i[11] ) if (n172) n580 <= 1'b0 ? 1'b0 : n2258;
/* FF 10 16  6 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n603 <= 1'b0; else if (n451) n603 <= n2259;
/* FF  1 22  4 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n92 <= 1'b0; else if (n194) n92 <= n2260;
/* FF 17 28  0 */ assign n1473 = n2261;
/* FF  5 27  0 */ always @(posedge \dd_pad_i[11] ) if (n376) n539 <= 1'b0 ? 1'b0 : n2262;
/* FF  5 22  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n511 <= 1'b0; else if (1'b1) n511 <= n2263;
/* FF 10 31  4 */ assign n876 = n2264;
/* FF 15 25  4 */ assign n1361 = n2265;
/* FF 12 17  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n679 <= 1'b0; else if (n6) n679 <= n2266;
/* FF 14 19  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n685 <= 1'b0; else if (n6) n685 <= n2267;
/* FF 11 27  3 */ always @(posedge \dd_pad_i[11] ) if (n429) n1083 <= 1'b0 ? 1'b0 : n2268;
/* FF  4 27  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) \da_pad_o[1]  <= 1'b0; else if (1'b1) \da_pad_o[1]  <= n2269;
/* FF  9 31  6 */ always @(posedge \dd_pad_i[11] ) if (n227) n871 <= 1'b0 ? 1'b0 : n2270;
/* FF 13 25  1 */ always @(posedge \dd_pad_i[11] ) if (n1) n849 <= 1'b0 ? 1'b0 : n2271;
/* FF  3 21  3 */ assign n281 = n2272;
/* FF 13 22  5 */ assign n1235 = n2273;
/* FF  7 28  0 */ assign n441 = n2274;
/* FF  4 20  0 */ assign n2275 = n2276;
/* FF  7 18  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n678 <= 1'b1; else if (1'b1) n678 <= n2278;
/* FF  9 27  3 */ always @(posedge \dd_pad_i[11] ) if (n227) n844 <= 1'b0 ? 1'b0 : n2279;
/* FF 12 16  5 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1112 <= 1'b0; else if (n451) n1112 <= n2280;
/* FF 11 24  2 */ always @(posedge \dd_pad_i[11] ) if (n424) n1061 <= 1'b0 ? 1'b0 : n2281;
/* FF  4 26  1 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n126 <= 1'b0; else if (n2) n126 <= n2282;
/* FF 21 22  6 */ assign n1526 = n2283;
/* FF 13 26  0 */ always @(posedge \dd_pad_i[11] ) if (n1) n966 <= 1'b0 ? 1'b0 : n2284;
/* FF  3 18  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n56 <= 1'b1; else if (n62) n56 <= n2285;
/* FF  2 22  0 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n184 <= 1'b0 ? 1'b0 : n2286;
/* FF 11 22  1 */ assign \wb_dat_o[15]  = n2287;
/* FF  5 16  4 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n449 <= 1'b0; else if (1'b1) n449 <= n2288;
/* FF 10 18  0 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n166 <= 1'b0; else if (n563) n166 <= n2289;
/* FF  6 26  7 */ always @(posedge \dd_pad_i[11] ) if (n638) n642 <= 1'b0 ? 1'b0 : n2290;
/* FF  5 29  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) \dd_pad_o[13]  <= 1'b0; else if (1'b1) \dd_pad_o[13]  <= n2291;
/* FF  7 19  0 */ always @(posedge \dd_pad_i[11] ) if (n31) n683 <= 1'b0 ? 1'b0 : n2292;
/* FF  9 20  2 */ always @(posedge \dd_pad_i[11] ) if (n478) n587 <= 1'b0 ? 1'b0 : n2293;
/* FF 12 23  4 */ assign n1152 = n2294;
/* FF  4 25  0 */ always @(posedge \dd_pad_i[11] ) if (n172) n421 <= 1'b0 ? 1'b0 : n2295;
/* FF 10 22  5 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) io_21_33_0 <= 1'b0; else if (1'b1) io_21_33_0 <= n2296;
/* FF  9 25  4 */ always @(posedge \dd_pad_i[11] ) if (n429) n833 <= 1'b0 ? 1'b0 : n2297;
/* FF 13 27  7 */ always @(posedge \dd_pad_i[11] ) if (n552) n1260 <= 1'b0 ? 1'b0 : n2298;
/* FF  3 19  1 */ assign n259 = n2299;
/* FF 11 23  2 */ assign n2300 = n1162;
/* FF 10 21  1 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n274 <= 1'b0 ? 1'b0 : n2301;
/* FF 15 19  3 */ assign n1335 = n2302;
/* FF 12 27  3 */ always @(posedge \dd_pad_i[11] ) if (n552) n1188 <= 1'b0 ? 1'b0 : n2303;
/* FF 15 28  7 */ assign n558 = n2304;
/* FF  9 21  1 */ assign n808 = n2305;
/* FF 13 31  4 */ assign n1278 = n2306;
/* FF 18 22  7 */ assign n1462 = n2307;
/* FF  6 24  0 */ always @(posedge \dd_pad_i[11] ) if (n376) n619 <= 1'b0 ? 1'b0 : n2308;
/* FF  4 24  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n419 <= 1'b0; else if (n2) n419 <= n2309;
/* FF  9 26  5 */ assign n840 = n2310;
/* FF 13 28  6 */ always @(posedge \dd_pad_i[11] ) if (n656) n1264 <= 1'b0 ? 1'b0 : n2311;
/* FF 18 21  3 */ assign n96 = n1515;
/* FF  2 24  2 */ assign n212 = n2312;
/* FF 11 20  3 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n355 <= 1'b0 ? 1'b0 : n2313;
/* FF  5 18  6 */ assign n356 = n2314;
/* FF 12 26  0 */ assign n1178 = n2315;
/* FF 17 21  7 */ assign n701 = n2316;
/* FF  1 18  0 */ assign n2317 = n2318;
/* FF 17 24  4 */ assign n1466 = n2320;
/* FF  4 28  4 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) \dd_pad_o[2]  <= 1'b0; else if (1'b1) \dd_pad_o[2]  <= n2321;
/* FF  7 17  6 */ assign n674 = n2322;
/* FF  9 22  0 */ assign n2323 = n922;
/* FF 14 26  0 */ always @(posedge \dd_pad_i[11] ) if (n1) n978 <= 1'b0 ? 1'b0 : n2324;
/* FF  6 27  1 */ assign n2325 = n722;
/* FF  9 32  6 */ assign \dd_pad_o[15]  = n2326;
/* FF 18 20  0 */ assign n2327 = n1511;
/* FF  6 21  0 */ assign n513 = n2328;
/* FF 11 21  4 */ assign n1034 = n2329;
/* FF  5 19  1 */ assign n470 = n2330;
/* FF 10 23  3 */ assign n2331 = n1058;
/* FF 15 26  4 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1369 <= 1'b0; else if (n329) n1369 <= n2332;
/* FF  7 21  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n106 <= 1'b0; else if (n756) n106 <= n2333;
/* FF 12 25  1 */ always @(posedge \dd_pad_i[11] ) if (n721) n1170 <= 1'b0 ? 1'b0 : n2334;
/* FF  4 19  5 */ assign n2335 = n481;
/* FF  9 28  6 */ always @(posedge \dd_pad_i[11] ) if (n655) n773 <= 1'b0 ? 1'b0 : n2336;
/* FF 18 24  5 */ assign n1498 = n2337;
/* FF 14 21  1 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n916 <= 1'b0; else if (n6) n916 <= n2338;
/* FF 11 17  1 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n676 <= 1'b0 ? 1'b0 : n2339;
/* FF 13 19  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n691 <= 1'b0; else if (n756) n691 <= n2340;
/* FF 15 21  2 */ assign n1340 = n2341;
/* FF 13 30  4 */ assign n2342 = n1329;
/* FF  2 17  5 */ assign n148 = n2343;
/* FF 18 23  1 */ assign n2344 = n1518;
/* FF  6 20  3 */ assign n592 = n2345;
/* FF 11 18  5 */ assign n1003 = n2346;
/* FF  5 20  0 */ assign n192 = n2347;
/* FF 15 22  4 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n103 <= 1'b0; else if (n756) n103 <= n2348;
/* FF  9 19  4 */ assign n792 = n2349;
/* FF 12 19  7 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n45 <= 1'b0 ? 1'b0 : n2350;
/* FF 12 24  6 */ assign n1156 = n2351;
/* FF 17 23  1 */ assign \wb_dat_o[1]  = n2352;
/* FF  4 18  6 */ assign n351 = n2353;
/* FF  9 29  5 */ always @(posedge \dd_pad_i[11] ) if (n227) n860 <= 1'b0 ? 1'b0 : n2354;
/* FF  7 23  4 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n692 <= 1'b0; else if (n329) n692 <= n2355;
/* FF 11 30  0 */ always @(posedge \dd_pad_i[11] ) if (n721) n1098 <= 1'b0 ? 1'b0 : n2356;
/* FF 16 23  5 */ assign n1405 = n2357;
/* FF 16 28  4 */ assign n1429 = n2358;
/* FF 13 20  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n755 <= 1'b0; else if (n451) n755 <= n2359;
/* FF  6 23  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) \wb_dat_o[30]  <= 1'b0; else if (1'b1) \wb_dat_o[30]  <= n2360;
/* FF 12 28  3 */ always @(posedge \dd_pad_i[11] ) if (n721) n1184 <= 1'b0 ? 1'b0 : n2361;
/* FF 11 19  6 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n42 <= 1'b0 ? 1'b0 : n2362;
/* FF  5 21  3 */ assign n499 = n2363;
/* FF 15 24  6 */ assign n1354 = n2364;
/* FF  7 27  1 */ always @(posedge \dd_pad_i[11] ) if (n638) n115 <= 1'b0 ? 1'b0 : n2365;
/* FF 12 18  4 */ assign n1010 = n2366;
/* FF 12 31  7 */ always @(posedge \dd_pad_i[11] ) if (n656) n1215 <= 1'b0 ? 1'b0 : n2367;
/* FF 16 24  1 */ assign n1176 = n2368;
/* FF  9 30  4 */ always @(posedge \dd_pad_i[11] ) if (n721) n868 <= 1'b0 ? 1'b0 : n2369;
/* FF  7 20  5 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n600 <= 1'b0; else if (n194) n600 <= n2370;
/* FF  9 17  5 */ assign n746 = n2371;
/* FF 14 23  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1042 <= 1'b0; else if (n194) n1042 <= n2372;
/* FF 16 27  5 */ always @(posedge \dd_pad_i[11] ) if (n656) n1425 <= 1'b0 ? 1'b0 : n2373;
/* FF 13 21  1 */ assign n1231 = n2374;
/* FF  6 22  5 */ assign n609 = n2375;
/* FF 11 16  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n992 <= 1'b0; else if (n4) n992 <= n2376;
/* FF  5 22  2 */ assign n172 = n2377;
/* FF 15 25  1 */ assign \wb_dat_o[16]  = n2378;
/* FF 15 20  6 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n747 <= 1'b0; else if (n451) n747 <= n2379;
/* FF  7 24  0 */ assign n424 = n2380;
/* FF 12 17  5 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n880 <= 1'b1; else if (n6) n880 <= n2381;
/* FF 12 30  4 */ always @(posedge \dd_pad_i[11] ) if (n424) n1208 <= 1'b0 ? 1'b0 : n2382;
/* FF  5 24  1 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n425 <= 1'b0; else if (n2) n425 <= n2383;
/* FF  4 16  0 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n344 <= 1'b0 ? 1'b0 : n2384;
/* FF  9 18  4 */ assign n165 = n2385;
/* FF 14 29  5 */ always @(posedge \dd_pad_i[11] ) if (n429) n1323 <= 1'b0 ? 1'b0 : n2386;
/* FF 14 22  4 */ assign \wb_dat_o[3]  = n2387;
/* FF  6 18  2 */ assign n563 = n2388;
/* FF 11 28  2 */ always @(posedge \dd_pad_i[11] ) if (n227) n1090 <= 1'b0 ? 1'b0 : n2389;
/* FF 16 26  6 */ assign n1419 = n2390;
/* FF 13 22  0 */ assign n1234 = n2391;
/* FF  3 22  2 */ assign n297 = n404;
/* FF  6 17  4 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n569 <= 1'b0; else if (n346) n569 <= n2392;
/* FF 10 30  0 */ always @(posedge \dd_pad_i[11] ) if (n655) n971 <= 1'b0 ? 1'b0 : n2393;
/* FF  4 20  5 */ assign n372 = n2394;
/* FF  7 18  6 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n51 <= 1'b0; else if (1'b1) n51 <= n2395;
/* FF  7 25  7 */ always @(posedge \dd_pad_i[11] ) if (n429) n715 <= 1'b0 ? 1'b0 : n2396;
/* FF 12 16  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1111 <= 1'b0; else if (n451) n1111 <= n2397;
/* FF 14 18  1 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n883 <= 1'b1; else if (n451) n883 <= n2398;
/* FF 12 29  5 */ always @(posedge \dd_pad_i[11] ) if (n721) n1201 <= 1'b0 ? 1'b0 : n2399;
/* FF  1 20  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n66 <= 1'b0; else if (n153) n66 <= n2400;
/* FF 17 18  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1437 <= 1'b0; else if (n329) n1437 <= n2401;
/* FF  5 25  2 */ assign n489 = n2402;
/* FF  4 23  1 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n407 <= 1'b0; else if (1'b1) n407 <= n2403;
/* FF  9 24  2 */ always @(posedge \dd_pad_i[11] ) if (n1) n828 <= 1'b0 ? 1'b0 : n2404;
/* FF 14 28  6 */ assign n2405 = n1379;
/* FF  2 22  5 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n199 <= 1'b0 ? 1'b0 : n2406;
/* FF 11 22  4 */ assign n1051 = n2407;
/* FF 11 29  5 */ always @(posedge \dd_pad_i[11] ) if (n655) n1097 <= 1'b0 ? 1'b0 : n2408;
/* FF 10 15  5 */ assign n668 = n2409;
/* FF 16 20  0 */ assign n2410 = n1448;
/* FF 15 18  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1139 <= 1'b1; else if (n4) n1139 <= n2411;
/* FF  3 23  1 */ assign n2412 = n411;
/* FF  2 21  1 */ assign n187 = n2413;
/* FF 12 20  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n814 <= 1'b0; else if (n4) n814 <= n2414;
/* FF 10 17  1 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n41 <= 1'b0 ? 1'b0 : n2415;
/* FF  7 19  5 */ assign n684 = n2416;
/* FF  3 24  5 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n315 <= 1'b0; else if (n2) n315 <= n2417;
/* FF 12 23  3 */ assign n2418 = n1244;
/* FF  5 26  3 */ always @(posedge \dd_pad_i[11] ) if (n478) n532 <= 1'b0 ? 1'b0 : n2419;
/* FF 11 25  2 */ always @(posedge \dd_pad_i[11] ) if (n552) n1069 <= 1'b0 ? 1'b0 : n2420;
/* FF  4 22  2 */ assign n394 = n2421;
/* FF  9 25  1 */ always @(posedge \dd_pad_i[11] ) if (n429) n831 <= 1'b0 ? 1'b0 : n2422;
/* FF 11 26  4 */ always @(posedge \dd_pad_i[11] ) if (n656) n1077 <= 1'b0 ? 1'b0 : n2423;
/* FF 16 19  1 */ assign n1387 = n2424;
/* FF  3 20  0 */ assign n265 = n2425;
/* FF  2 20  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n173 <= 1'b0; else if (1'b1) n173 <= n2426;
/* FF 12 27  6 */ always @(posedge \dd_pad_i[11] ) if (n552) n1182 <= 1'b0 ? 1'b0 : n2427;
/* FF  6 19  6 */ always @(posedge \dd_pad_i[11] ) if (n172) n584 <= 1'b0 ? 1'b0 : n2428;
/* FF 15 28  2 */ assign n2429 = n1433;
/* FF 12 22  0 */ assign n2430 = n1238;
/* FF  1 22  0 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n89 <= 1'b0; else if (n194) n89 <= n2431;
/* FF  5 27  4 */ always @(posedge \dd_pad_i[11] ) if (n376) n543 <= 1'b0 ? 1'b0 : n2432;
/* FF  4 21  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n382 <= 1'b0; else if (n298) n382 <= n2433;
/* FF  9 26  0 */ always @(posedge \dd_pad_i[11] ) if (n638) n657 <= 1'b0 ? 1'b0 : n2434;
/* FF  2 24  7 */ assign n217 = n2435;
/* FF 14 19  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1044 <= 1'b0; else if (n6) n1044 <= n2436;
/* FF 11 20  6 */ assign n1024 = n2437;
/* FF 11 27  7 */ always @(posedge \dd_pad_i[11] ) if (n429) n967 <= 1'b0 ? 1'b0 : n2438;
/* FF  3 21  7 */ assign n284 = n2439;
/* FF  2 23  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n206 <= 1'b1; else if (n113) n206 <= n2440;
/* FF 20 22  3 */ assign n1519 = n2441;
/* FF 12 26  5 */ always @(posedge \dd_pad_i[11] ) if (n721) n1181 <= 1'b0 ? 1'b0 : n2442;
/* FF 17 24  3 */ assign n2443 = n1503;
/* FF 10 19  3 */ assign n2444 = n1019;
/* FF  7 17  3 */ assign n671 = n2445;
/* FF  7 28  4 */ assign n727 = n2446;
/* FF 14 26  5 */ always @(posedge \dd_pad_i[11] ) if (n1) n720 <= 1'b0 ? 1'b0 : n2447;
/* FF 12 21  1 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1043 <= 1'b0; else if (n4) n1043 <= n2448;
/* FF  5 28  5 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) \dd_pad_o[3]  <= 1'b0; else if (1'b1) \dd_pad_o[3]  <= n2449;
/* FF 14 25  1 */ always @(posedge \dd_pad_i[11] ) if (n656) n1252 <= 1'b0 ? 1'b0 : n2450;
/* FF  3 17  4 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n242 <= 1'b1; else if (n44) n242 <= n2451;
/* FF  6 21  7 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n400 <= 1'b0 ? 1'b0 : n2452;
/* FF 11 24  6 */ always @(posedge \dd_pad_i[11] ) if (n424) n1064 <= 1'b0 ? 1'b0 : n2453;
/* FF 15 17  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n788 <= 1'b0; else if (n6) n788 <= n2454;
/* FF  3 18  6 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n155 <= 1'b0; else if (n62) n155 <= n2455;
/* FF 12 25  4 */ assign n1159 = n2456;
/* FF  5 16  0 */ assign n2457 = n564;
/* FF 10 25  5 */ always @(posedge \dd_pad_i[11] ) if (n429) n920 <= 1'b0 ? 1'b0 : n2458;
/* FF 10 18  4 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n261 <= 1'b1; else if (n563) n261 <= n2459;
/* FF  7 22  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n401 <= 1'b0; else if (1'b1) n401 <= n2460;
/* FF 14 21  4 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1040 <= 1'b0; else if (n6) n1040 <= n2461;
/* FF  6 26  3 */ always @(posedge \dd_pad_i[11] ) if (n638) n627 <= 1'b0 ? 1'b0 : n2462;
/* FF 11 17  6 */ assign n2463 = n1118;
/* FF 14 24  2 */ assign n2464 = n1356;
/* FF  6 20  4 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) io_27_33_1 <= 1'b1; else if (1'b1) io_27_33_1 <= n2465;
/* FF  6 25  7 */ assign n632 = n2466;
/* FF 11 18  0 */ assign n2467 = n1122;
/* FF 10 22  1 */ assign n911 = n1054;
/* FF 15 22  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n105 <= 1'b0; else if (n756) n105 <= n2468;
/* FF 18 18  6 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1478 <= 1'b0; else if (n329) n1478 <= n2469;
/* FF  3 19  5 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n58 <= 1'b0; else if (n62) n58 <= n2470;
/* FF 12 24  3 */ assign n1165 = n2471;
/* FF  5 17  3 */ always @(posedge \dd_pad_i[11] ) if (n478) n364 <= 1'b0 ? 1'b0 : n2472;
/* FF 10 24  6 */ assign n836 = n2473;
/* FF 10 21  5 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n366 <= 1'b0 ? 1'b0 : n2474;
/* FF  7 23  1 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n317 <= 1'b0; else if (n329) n317 <= n2475;
/* FF 14 20  7 */ assign n816 = n2476;
/* FF 17 20  0 */ assign n1444 = n2477;
/* FF 11 30  7 */ always @(posedge \dd_pad_i[11] ) if (n721) n1103 <= 1'b0 ? 1'b0 : n2478;
/* FF 16 28  1 */ assign \wb_dat_o[23]  = n2479;
/* FF 13 31  0 */ assign n2480 = n1330;
/* FF 18 22  3 */ assign n1492 = n2481;
/* FF 14 27  3 */ assign n1306 = n2482;
/* FF  6 24  4 */ always @(posedge \dd_pad_i[11] ) if (n376) n623 <= 1'b0 ? 1'b0 : n2483;
/* FF 11 19  3 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n1013 <= 1'b0 ? 1'b0 : n2484;
/* FF 13 17  1 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1018 <= 1'b0; else if (n4) n1018 <= n2485;
/* FF 15 23  0 */ assign n2486 = n1407;
/* FF 18 21  7 */ assign n1489 = n2487;
/* FF 12 31  2 */ assign n2488 = n1282;
/* FF  5 18  2 */ assign n2489 = n578;
/* FF 10 27  7 */ assign n130 = n2490;
/* FF 10 20  6 */ assign n893 = n1032;
/* FF  7 20  0 */ assign n194 = n2491;
/* FF 14 23  6 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1290 <= 1'b0; else if (n194) n1290 <= n2492;
/* FF 17 21  3 */ assign n2493 = n1490;
/* FF  1 18  4 */ assign n36 = n2494;
/* FF 11 31  4 */ assign n2495 = n1217;
/* FF 16 27  0 */ always @(posedge \dd_pad_i[11] ) if (n656) n1421 <= 1'b0 ? 1'b0 : n2496;
/* FF  6 22  2 */ assign n2497 = n705;
/* FF  6 27  5 */ assign n2498 = n724;
/* FF 11 16  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n990 <= 1'b1; else if (n4) n990 <= n2499;
/* FF 13 18  0 */ assign n54 = n2500;
/* FF 15 20  1 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1038 <= 1'b0; else if (n451) n1038 <= n2501;
/* FF 18 20  4 */ assign n465 = n1512;
/* FF 12 30  1 */ always @(posedge \dd_pad_i[11] ) if (n424) n1205 <= 1'b0 ? 1'b0 : n2502;
/* FF  5 24  4 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n520 <= 1'b0; else if (n2) n520 <= n2503;
/* FF  5 19  5 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n472 <= 1'b0; else if (1'b1) n472 <= n2504;
/* FF 10 26  0 */ always @(posedge \dd_pad_i[11] ) if (n552) n949 <= 1'b0 ? 1'b0 : n2505;
/* FF 10 23  7 */ assign n929 = n2506;
/* FF 15 26  0 */ assign n1367 = n2507;
/* FF 14 22  1 */ assign n2508 = n1344;
/* FF  6 18  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n573 <= 1'b0; else if (n563) n573 <= n2509;
/* FF 17 22  2 */ assign \wb_dat_o[25]  = n2510;
/* FF 11 28  5 */ always @(posedge \dd_pad_i[11] ) if (n227) n1092 <= 1'b0 ? 1'b0 : n2511;
/* FF  4 19  1 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n360 <= 1'b0; else if (1'b1) n360 <= n2512;
/* FF  9 28  2 */ always @(posedge \dd_pad_i[11] ) if (n655) n852 <= 1'b0 ? 1'b0 : n2513;
/* FF 18 24  1 */ assign n817 = n1520;
/* FF  6 17  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n568 <= 1'b1; else if (n346) n568 <= n2514;
/* FF 10 30  5 */ always @(posedge \dd_pad_i[11] ) if (n655) n974 <= 1'b0 ? 1'b0 : n2515;
/* FF  9 14  5 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n782 <= 1'b1; else if (n4) n782 <= n2516;
/* FF 13 19  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1026 <= 1'b0; else if (n756) n1026 <= n2517;
/* FF  3 27  1 */ always @(posedge \dd_pad_i[11] ) if (n1) n131 <= 1'b0 ? 1'b0 : n2518;
/* FF  2 17  1 */ assign n144 = n2519;
/* FF 14 18  6 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1039 <= 1'b1; else if (n451) n1039 <= n2520;
/* FF 12 29  0 */ assign n1104 = n2521;
/* FF  5 20  4 */ assign n485 = n2522;
/* FF 10 29  1 */ always @(posedge \dd_pad_i[11] ) if (n227) n662 <= 1'b0 ? 1'b0 : n2523;
/* FF 12 19  3 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n246 <= 1'b0 ? 1'b0 : n2524;
/* FF 17 23  5 */ always @(posedge \dd_pad_i[11] ) if (n31) n1461 <= 1'b0 ? 1'b0 : n2525;
/* FF 11 29  2 */ always @(posedge \dd_pad_i[11] ) if (n655) n1096 <= 1'b0 ? 1'b0 : n2526;
/* FF 16 25  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1414 <= 1'b0; else if (n329) n1414 <= n2527;
/* FF  4 18  2 */ assign n2528 = n467;
/* FF  9 29  1 */ always @(posedge \dd_pad_i[11] ) if (n227) n858 <= 1'b0 ? 1'b0 : n2529;
/* FF 13 23  4 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n111 <= 1'b0 ? 1'b0 : n2530;
/* FF 16 23  1 */ assign n1402 = n2531;
/* FF 13 20  6 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n918 <= 1'b0; else if (n451) n918 <= n2532;
/* FF  3 24  0 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n310 <= 1'b0; else if (n2) n310 <= n2533;
/* FF 11 12  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n879 <= 1'b0; else if (n4) n879 <= n2534;
/* FF  5 26  6 */ always @(posedge \dd_pad_i[11] ) if (n478) n535 <= 1'b0 ? 1'b0 : n2535;
/* FF 11 25  7 */ always @(posedge \dd_pad_i[11] ) if (n552) n1073 <= 1'b0 ? 1'b0 : n2536;
/* FF  5 21  7 */ assign n502 = n2537;
/* FF 10 28  2 */ always @(posedge \dd_pad_i[11] ) if (n655) n963 <= 1'b0 ? 1'b0 : n2538;
/* FF 15 24  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1351 <= 1'b0; else if (n329) n1351 <= n2539;
/* FF 12 18  0 */ assign n2540 = n2541;
/* FF 14 16  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1006 <= 1'b0; else if (n4) n1006 <= n2543;
/* FF  6 28  5 */ assign n653 = n2544;
/* FF 11 26  3 */ always @(posedge \dd_pad_i[11] ) if (n656) n829 <= 1'b0 ? 1'b0 : n2545;
/* FF 12 32  6 */ assign n1218 = n2546;
/* FF  9 30  0 */ assign n864 = n2547;
/* FF 13 24  5 */ always @(posedge \dd_pad_i[11] ) if (n424) n1177 <= 1'b0 ? 1'b0 : n2548;
/* FF  6 19  1 */ always @(posedge \dd_pad_i[11] ) if (n172) n579 <= 1'b0 ? 1'b0 : n2549;
/* FF 10 16  7 */ assign n882 = n2550;
/* FF 13 21  5 */ assign n1233 = n2551;
/* FF  2 19  3 */ assign n163 = n2552;
/* FF 20 18  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n784 <= 1'b0; else if (n6) n784 <= n2553;
/* FF 17 28  3 */ assign n2554 = n1508;
/* FF  5 27  1 */ always @(posedge \dd_pad_i[11] ) if (n376) n540 <= 1'b0 ? 1'b0 : n2555;
/* FF  5 22  6 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n376 <= 1'b0; else if (1'b1) n376 <= n2556;
/* FF 10 31  3 */ assign n983 = n2557;
/* FF 15 25  5 */ assign n1362 = n2558;
/* FF 14 19  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n805 <= 1'b1; else if (n6) n805 <= n2559;
/* FF 11 27  0 */ always @(posedge \dd_pad_i[11] ) if (n429) n1080 <= 1'b0 ? 1'b0 : n2560;
/* FF  4 27  5 */ assign n437 = n2561;
/* FF 13 25  6 */ always @(posedge \dd_pad_i[11] ) if (n1) n779 <= 1'b0 ? 1'b0 : n2562;
/* FF 18 16  5 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1011 <= 1'b0; else if (n6) n1011 <= n2563;
/* FF 14 29  1 */ always @(posedge \dd_pad_i[11] ) if (n429) n1275 <= 1'b0 ? 1'b0 : n2564;
/* FF 18 29  6 */ assign n1509 = n2565;
/* FF 16 21  3 */ assign n1397 = n2566;
/* FF 10 19  6 */ assign n892 = n2567;
/* FF 15 29  2 */ assign n1381 = n2568;
/* FF 13 22  4 */ assign \wb_dat_i[1]  = n2569;
/* FF  2 18  4 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n151 <= 1'b1; else if (n153) n151 <= n2570;
/* FF  4 20  1 */ assign n368 = n2571;
/* FF  7 18  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n675 <= 1'b0; else if (1'b1) n675 <= n2572;
/* FF  9 27  4 */ always @(posedge \dd_pad_i[11] ) if (n227) n845 <= 1'b0 ? 1'b0 : n2573;
/* FF 11 24  1 */ always @(posedge \dd_pad_i[11] ) if (n424) n1060 <= 1'b0 ? 1'b0 : n2574;
/* FF  4 26  6 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n428 <= 1'b0; else if (n2) n428 <= n2575;
/* FF  4 23  5 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n202 <= 1'b0; else if (1'b1) n202 <= n2576;
/* FF  9 24  6 */ always @(posedge \dd_pad_i[11] ) if (n1) n764 <= 1'b0 ? 1'b0 : n2577;
/* FF 13 26  7 */ always @(posedge \dd_pad_i[11] ) if (n1) n968 <= 1'b0 ? 1'b0 : n2578;
/* FF 14 28  2 */ assign n2579 = n1378;
/* FF  2 22  1 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n195 <= 1'b0 ? 1'b0 : n2580;
/* FF 11 22  0 */ assign n2581 = n1149;
/* FF  5 16  7 */ assign n450 = n2582;
/* FF 16 20  4 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1394 <= 1'b0; else if (n329) n1394 <= n2583;
/* FF 10 18  1 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n886 <= 1'b0; else if (n563) n886 <= n2584;
/* FF 15 18  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n796 <= 1'b1; else if (n4) n796 <= n2585;
/* FF  2 21  5 */ assign n190 = n2586;
/* FF 12 20  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n363 <= 1'b0; else if (n4) n363 <= n2587;
/* FF  5 29  3 */ assign n555 = n2588;
/* FF  7 19  1 */ assign n2589 = n752;
/* FF  9 20  5 */ always @(posedge \dd_pad_i[11] ) if (n478) n804 <= 1'b0 ? 1'b0 : n2590;
/* FF  6 25  2 */ assign n629 = n2591;
/* FF  4 25  7 */ always @(posedge \dd_pad_i[11] ) if (n172) n334 <= 1'b0 ? 1'b0 : n2592;
/* FF 10 22  6 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) \wb_dat_o[28]  <= 1'b1; else if (1'b1) \wb_dat_o[28]  <= n2593;
/* FF  4 22  6 */ assign n397 = n2594;
/* FF  9 25  5 */ always @(posedge \dd_pad_i[11] ) if (n429) n122 <= 1'b0 ? 1'b0 : n2595;
/* FF 13 27  0 */ always @(posedge \dd_pad_i[11] ) if (n552) n1253 <= 1'b0 ? 1'b0 : n2596;
/* FF 11 23  3 */ assign io_33_23_0 = n2597;
/* FF  5 17  4 */ always @(posedge \dd_pad_i[11] ) if (n478) n456 <= 1'b0 ? 1'b0 : n2598;
/* FF 16 19  5 */ assign \dd_pad_o[0]  = n2599;
/* FF 10 21  0 */ assign n2600 = n1047;
/* FF 15 19  0 */ assign n1334 = n2601;
/* FF  2 20  6 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n176 <= 1'b0; else if (1'b1) n176 <= n2602;
/* FF 12 27  2 */ always @(posedge \dd_pad_i[11] ) if (n552) n1187 <= 1'b0 ? 1'b0 : n2603;
/* FF 13 31  5 */ assign n988 = n2604;
/* FF 12 22  4 */ assign n2605 = n1239;
/* FF  6 24  1 */ always @(posedge \dd_pad_i[11] ) if (n376) n620 <= 1'b0 ? 1'b0 : n2606;
/* FF  4 24  0 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n414 <= 1'b0; else if (n2) n414 <= n2607;
/* FF  4 21  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n385 <= 1'b0; else if (n298) n385 <= n2608;
/* FF  9 26  4 */ always @(posedge \dd_pad_i[11] ) if (n638) n548 <= 1'b0 ? 1'b0 : n2609;
/* FF 13 28  1 */ assign n2610 = n1318;
/* FF 18 21  2 */ assign n1486 = n1514;
/* FF 14 30  4 */ always @(posedge \dd_pad_i[11] ) if (n1) n719 <= 1'b0 ? 1'b0 : n2611;
/* FF  2 24  3 */ assign n213 = n2612;
/* FF 11 20  2 */ assign n2613 = n1140;
/* FF 17 27  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1472 <= 1'b0; else if (n329) n1472 <= n2614;
/* FF  5 18  5 */ assign n461 = n2615;
/* FF 10 20  3 */ assign n2616 = n1031;
/* FF  2 23  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n210 <= 1'b0; else if (n113) n210 <= n2617;
/* FF 12 26  1 */ always @(posedge \dd_pad_i[11] ) if (n721) n1179 <= 1'b0 ? 1'b0 : n2618;
/* FF 17 21  4 */ assign n2619 = n1491;
/* FF  7 17  7 */ assign n667 = n2620;
/* FF 14 26  1 */ always @(posedge \dd_pad_i[11] ) if (n1) n1105 <= 1'b0 ? 1'b0 : n2621;
/* FF 12 21  5 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1125 <= 1'b0; else if (n4) n1125 <= n2622;
/* FF  6 27  0 */ assign n644 = n2623;
/* FF 13 29  2 */ assign n1270 = n2624;
/* FF 18 20  1 */ assign n1483 = n2625;
/* FF  3 17  0 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n152 <= 1'b1; else if (n44) n152 <= n2626;
/* FF 14 25  5 */ assign n2627 = n1365;
/* FF 11 21  5 */ assign n1035 = n2628;
/* FF  5 19  2 */ assign n466 = n589;
/* FF 10 23  2 */ always @(posedge \dd_pad_i[11] ) if (n656) n921 <= 1'b0 ? 1'b0 : n2629;
/* FF 15 17  6 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n890 <= 1'b0; else if (n6) n890 <= n2630;
/* FF  7 21  4 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n97 <= 1'b0; else if (n756) n97 <= n2631;
/* FF 12 25  0 */ assign n1157 = n2632;
/* FF 17 22  5 */ assign n1456 = n2633;
/* FF  1 19  0 */ always @(posedge \dd_pad_i[11] ) if (n172) n48 <= 1'b0 ? 1'b0 : n2634;
/* FF 10 25  1 */ always @(posedge \dd_pad_i[11] ) if (n429) n944 <= 1'b0 ? 1'b0 : n2635;
/* FF  4 19  4 */ assign n362 = n480;
/* FF  7 22  6 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n698 <= 1'b0; else if (1'b1) n698 <= n2636;
/* FF  9 23  0 */ assign n2637 = n934;
/* FF 14 21  0 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n815 <= 1'b0; else if (n6) n815 <= n2638;
/* FF 11 17  2 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n995 <= 1'b0 ? 1'b0 : n2639;
/* FF  1 13  4 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n24 <= 1'b0 ? 1'b0 : n2640;
/* FF 13 30  3 */ assign n2641 = n1328;
/* FF  2 17  4 */ assign n147 = n2642;
/* FF 18 23  0 */ assign n1495 = n2643;
/* FF 14 24  6 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1297 <= 1'b0; else if (n329) n1297 <= n2644;
/* FF  6 20  0 */ assign n2645 = n694;
/* FF 11 15  7 */ assign n989 = n2646;
/* FF 11 18  4 */ assign n1002 = n2647;
/* FF  5 20  3 */ assign n484 = n598;
/* FF 15 27  4 */ assign n1317 = n2648;
/* FF 15 22  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1168 <= 1'b0; else if (n756) n1168 <= n2649;
/* FF  7 26  5 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n399 <= 1'b0 ? 1'b0 : n2650;
/* FF  9 19  5 */ always @(posedge \dd_pad_i[11] ) if (n172) n793 <= 1'b0 ? 1'b0 : n2651;
/* FF 12 19  6 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n55 <= 1'b0 ? 1'b0 : n2652;
/* FF 12 24  7 */ assign n1166 = n2653;
/* FF 17 26  5 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1469 <= 1'b0; else if (n329) n1469 <= n2654;
/* FF 10 24  2 */ always @(posedge \dd_pad_i[11] ) if (n424) n938 <= 1'b0 ? 1'b0 : n2655;
/* FF  4 18  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n352 <= 1'b0; else if (1'b1) n352 <= n2656;
/* FF  7 23  5 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n700 <= 1'b0; else if (n329) n700 <= n2657;
/* FF  9 16  1 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n457 <= 1'b0 ? 1'b0 : n2658;
/* FF 11 30  3 */ always @(posedge \dd_pad_i[11] ) if (n721) n1101 <= 1'b0 ? 1'b0 : n2659;
/* FF 16 23  4 */ always @(posedge \dd_pad_i[11] ) if (n31) n1404 <= 1'b0 ? 1'b0 : n2660;
/* FF 16 28  5 */ assign n1430 = n2661;
/* FF 20 19  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1510 <= 1'b0; else if (n329) n1510 <= n2662;
/* FF 14 27  7 */ always @(posedge \dd_pad_i[11] ) if (n424) n1310 <= 1'b0 ? 1'b0 : n2663;
/* FF 12 28  4 */ assign n2664 = n1267;
/* FF 11 19  7 */ assign n1015 = n2665;
/* FF  5 21  0 */ assign n2666 = n604;
/* FF 15 24  5 */ assign n1353 = n2667;
/* FF 15 23  4 */ assign n1348 = n2668;
/* FF  7 27  6 */ assign n721 = n2669;
/* FF 12 18  5 */ assign n682 = n2670;
/* FF 12 31  6 */ always @(posedge \dd_pad_i[11] ) if (n656) n1214 <= 1'b0 ? 1'b0 : n2671;
/* FF  7 20  4 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n599 <= 1'b0; else if (n194) n599 <= n2672;
/* FF 14 23  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1294 <= 1'b0; else if (n194) n1294 <= n2673;
/* FF 11 31  0 */ assign n1106 = n2674;
/* FF 16 27  4 */ always @(posedge \dd_pad_i[11] ) if (n656) n1424 <= 1'b0 ? 1'b0 : n2675;
/* FF  6 22  6 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n515 <= 1'b0 ? 1'b0 : n2676;
/* FF  5 22  1 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n509 <= 1'b0; else if (1'b1) n509 <= n2677;
/* FF 15 25  2 */ always @(posedge \dd_pad_i[11] ) if (n31) n1359 <= 1'b0 ? 1'b0 : n2678;
/* FF 15 20  5 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n905 <= 1'b1; else if (n451) n905 <= n2679;
/* FF  7 24  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n693 <= 1'b0; else if (1'b1) n693 <= n2680;
/* FF 12 30  5 */ assign n2681 = n1276;
/* FF  5 24  0 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n427 <= 1'b0; else if (n2) n427 <= n2682;
/* FF 10 26  4 */ always @(posedge \dd_pad_i[11] ) if (n552) n943 <= 1'b0 ? 1'b0 : n2683;
/* FF  4 16  1 */ assign n345 = n2684;
/* FF  7 14  2 */ assign \wb_dat_o[7]  = n2685;
/* FF  9 18  3 */ assign n786 = n2686;
/* FF 14 29  4 */ assign n1322 = n2687;
/* FF 14 22  5 */ always @(posedge \dd_pad_i[11] ) if (n31) n1288 <= 1'b0 ? 1'b0 : n2688;
/* FF  6 18  3 */ assign n275 = n2689;
/* FF 11 28  1 */ always @(posedge \dd_pad_i[11] ) if (n227) n1089 <= 1'b0 ? 1'b0 : n2690;
/* FF  3 22  5 */ assign n2691 = n406;
/* FF  6 17  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n572 <= 1'b0; else if (n346) n572 <= n2692;
/* FF 10 30  1 */ always @(posedge \dd_pad_i[11] ) if (n655) n856 <= 1'b0 ? 1'b0 : n2693;
/* FF  4 20  6 */ assign n373 = n2694;
/* FF 15 30  3 */ assign n1384 = n2695;
/* FF  7 25  0 */ assign n712 = n2696;
/* FF 12 16  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1007 <= 1'b0; else if (n451) n1007 <= n2697;
/* FF 14 18  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1120 <= 1'b1; else if (n451) n1120 <= n2698;
/* FF 12 29  4 */ always @(posedge \dd_pad_i[11] ) if (n721) n1200 <= 1'b0 ? 1'b0 : n2699;
/* FF  1 20  5 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n69 <= 1'b1; else if (n153) n69 <= n2700;
/* FF 17 18  1 */ assign io_33_24_0 = n2701;
/* FF  4 23  0 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) dmarq_pad_i <= 1'b0; else if (1'b1) dmarq_pad_i <= n2702;
/* FF 14 28  7 */ assign n1316 = n2703;
/* FF  2 22  6 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n200 <= 1'b0 ? 1'b0 : n2704;
/* FF  6 29  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) \dd_pad_o[11]  <= 1'b0; else if (1'b1) \dd_pad_o[11]  <= n2705;
/* FF 11 22  7 */ assign n1052 = n2706;
/* FF 11 29  6 */ always @(posedge \dd_pad_i[11] ) if (n655) n736 <= 1'b0 ? 1'b0 : n2707;
/* FF 16 20  1 */ assign n1392 = n2708;
/* FF 15 18  6 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1136 <= 1'b1; else if (n4) n1136 <= n2709;
/* FF  3 23  6 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) cs0n_pad_o <= 1'b0; else if (1'b1) cs0n_pad_o <= n2710;
/* FF  2 21  0 */ assign n2711 = n2712;
/* FF 10 17  0 */ assign n2714 = n999;
/* FF  3 24  4 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n222 <= 1'b0; else if (n2) n222 <= n2715;
/* FF  7 30  1 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n262 <= 1'b1; else if (n6) n262 <= n2716;
/* FF 12 23  2 */ assign n711 = n2717;
/* FF  5 26  2 */ always @(posedge \dd_pad_i[11] ) if (n478) n531 <= 1'b0 ? 1'b0 : n2718;
/* FF 11 25  3 */ always @(posedge \dd_pad_i[11] ) if (n552) n1070 <= 1'b0 ? 1'b0 : n2719;
/* FF 10 28  6 */ always @(posedge \dd_pad_i[11] ) if (n655) n965 <= 1'b0 ? 1'b0 : n2720;
/* FF  4 22  3 */ assign n395 = n2721;
/* FF  6 28  1 */ assign n2722 = n732;
/* FF 11 23  4 */ always @(posedge \dd_pad_i[11] ) if (n31) n1056 <= 1'b0 ? 1'b0 : n2723;
/* FF 11 26  7 */ always @(posedge \dd_pad_i[11] ) if (n656) n1079 <= 1'b0 ? 1'b0 : n2724;
/* FF 16 19  0 */ assign n2725 = n1442;
/* FF 15 19  5 */ assign n2726 = n1391;
/* FF 13 24  1 */ always @(posedge \dd_pad_i[11] ) if (n424) n838 <= 1'b0 ? 1'b0 : n2727;
/* FF  3 20  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n269 <= 1'b0; else if (n153) n269 <= n2728;
/* FF  2 20  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n174 <= 1'b0; else if (1'b1) n174 <= n2729;
/* FF  6 19  5 */ always @(posedge \dd_pad_i[11] ) if (n172) n583 <= 1'b0 ? 1'b0 : n2730;
/* FF 10 16  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n881 <= 1'b1; else if (n451) n881 <= n2731;
/* FF 15 28  1 */ assign n1373 = n2732;
/* FF 12 22  1 */ assign \wb_dat_o[0]  = n2733;
/* FF  1 22  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n95 <= 1'b0; else if (n194) n95 <= n2734;
/* FF  5 27  5 */ always @(posedge \dd_pad_i[11] ) if (n376) n544 <= 1'b0 ? 1'b0 : n2735;
/* FF 10 31  7 */ assign n985 = n2736;
/* FF  4 21  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n381 <= 1'b0; else if (n298) n381 <= n2737;
/* FF  2 24  4 */ assign n214 = n2738;
/* FF 14 19  6 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1127 <= 1'b0; else if (n6) n1127 <= n2739;
/* FF 11 20  5 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n348 <= 1'b0 ? 1'b0 : n2740;
/* FF 11 27  4 */ always @(posedge \dd_pad_i[11] ) if (n429) n1084 <= 1'b0 ? 1'b0 : n2741;
/* FF  4 27  1 */ assign n2742 = n549;
/* FF 13 25  2 */ always @(posedge \dd_pad_i[11] ) if (n1) n635 <= 1'b0 ? 1'b0 : n2743;
/* FF 15 15  5 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n665 <= 1'b0 ? 1'b0 : n2744;
/* FF  3 21  0 */ assign n279 = n2745;
/* FF  2 23  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n185 <= 1'b0; else if (n113) n185 <= n2746;
/* FF 17 24  2 */ always @(posedge \dd_pad_i[11] ) if (n31) n1465 <= 1'b0 ? 1'b0 : n2747;
/* FF 10 19  2 */ assign n895 = n2748;
/* FF  7 28  3 */ assign n134 = n2749;
/* FF 14 26  6 */ always @(posedge \dd_pad_i[11] ) if (n1) n769 <= 1'b0 ? 1'b0 : n2750;
/* FF 12 21  0 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n931 <= 1'b0; else if (n4) n931 <= n2751;
/* FF  9 27  0 */ always @(posedge \dd_pad_i[11] ) if (n227) n842 <= 1'b0 ? 1'b0 : n2752;
/* FF 14 25  0 */ always @(posedge \dd_pad_i[11] ) if (n656) n1298 <= 1'b0 ? 1'b0 : n2753;
/* FF  3 17  5 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n243 <= 1'b0; else if (n44) n243 <= n2754;
/* FF  6 21  6 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n309 <= 1'b0 ? 1'b0 : n2755;
/* FF 11 21  2 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n378 <= 1'b0 ? 1'b0 : n2756;
/* FF 11 24  5 */ always @(posedge \dd_pad_i[11] ) if (n424) n1063 <= 1'b0 ? 1'b0 : n2757;
/* FF  4 26  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n431 <= 1'b0; else if (n2) n431 <= n2758;
/* FF 18 19  0 */ assign n1480 = n2759;
/* FF  3 18  1 */ assign n254 = n359;
/* FF  5 16  3 */ assign n448 = n2760;
/* FF 10 25  4 */ always @(posedge \dd_pad_i[11] ) if (n429) n946 <= 1'b0 ? 1'b0 : n2761;
/* FF 10 18  5 */ assign n798 = n1014;
/* FF  6 26  4 */ always @(posedge \dd_pad_i[11] ) if (n638) n640 <= 1'b0 ? 1'b0 : n2762;
/* FF 11 17  7 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n997 <= 1'b0 ? 1'b0 : n2763;
/* FF  5 29  7 */ assign n557 = n2764;
/* FF 16 29  5 */ always @(posedge \dd_pad_i[11] ) if (n429) n1383 <= 1'b0 ? 1'b0 : n2765;
/* FF  9 20  1 */ always @(posedge \dd_pad_i[11] ) if (n478) n801 <= 1'b0 ? 1'b0 : n2766;
/* FF 14 24  3 */ assign n765 = n2767;
/* FF 11 18  3 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n1001 <= 1'b0 ? 1'b0 : n2768;
/* FF  4 25  3 */ always @(posedge \dd_pad_i[11] ) if (n172) n423 <= 1'b0 ? 1'b0 : n2769;
/* FF 10 22  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) \wb_dat_o[6]  <= 1'b1; else if (1'b1) \wb_dat_o[6]  <= n2770;
/* FF 15 22  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1169 <= 1'b0; else if (n756) n1169 <= n2771;
/* FF 13 27  4 */ always @(posedge \dd_pad_i[11] ) if (n552) n1257 <= 1'b0 ? 1'b0 : n2772;
/* FF  3 19  2 */ assign n260 = n2773;
/* FF 17 26  0 */ assign n1426 = n2774;
/* FF  1  7  5 */ assign n5 = n2775;
/* FF  5 17  0 */ always @(posedge \dd_pad_i[11] ) if (n478) n453 <= 1'b0 ? 1'b0 : n2776;
/* FF 10 24  7 */ always @(posedge \dd_pad_i[11] ) if (n424) n941 <= 1'b0 ? 1'b0 : n2777;
/* FF 10 21  4 */ assign n2778 = n1049;
/* FF 14 20  4 */ assign n1065 = n2779;
/* FF 17 20  3 */ assign n1446 = n2780;
/* FF 11 30  6 */ always @(posedge \dd_pad_i[11] ) if (n721) n979 <= 1'b0 ? 1'b0 : n2781;
/* FF  5 30  6 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) \dd_pad_o[12]  <= 1'b0; else if (1'b1) \dd_pad_o[12]  <= n2782;
/* FF 16 28  2 */ always @(posedge \dd_pad_i[11] ) if (n31) n1428 <= 1'b0 ? 1'b0 : n2783;
/* FF 13 31  1 */ assign n2784 = n1331;
/* FF 14 27  2 */ always @(posedge \dd_pad_i[11] ) if (n424) n1305 <= 1'b0 ? 1'b0 : n2785;
/* FF  6 24  5 */ always @(posedge \dd_pad_i[11] ) if (n376) n624 <= 1'b0 ? 1'b0 : n2786;
/* FF 11 19  0 */ assign n2787 = n1131;
/* FF  4 24  4 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n417 <= 1'b0; else if (n2) n417 <= n2788;
/* FF 15 23  1 */ assign n2789 = n1408;
/* FF 13 28  5 */ assign n1263 = n2790;
/* FF 18 21  6 */ assign n1337 = n2791;
/* FF  5 18  1 */ assign n459 = n2792;
/* FF 16 24  7 */ assign \wb_dat_o[29]  = n2793;
/* FF 10 20  7 */ assign n899 = n2794;
/* FF 14 23  5 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1242 <= 1'b0; else if (n194) n1242 <= n2795;
/* FF 17 21  0 */ assign n1449 = n2796;
/* FF  1 18  3 */ assign n35 = n2797;
/* FF 11 31  5 */ assign n1107 = n2798;
/* FF 16 27  3 */ always @(posedge \dd_pad_i[11] ) if (n656) n1423 <= 1'b0 ? 1'b0 : n2799;
/* FF  9 22  3 */ assign n2800 = n924;
/* FF  6 22  3 */ assign io_18_33_0 = n2801;
/* FF  6 27  4 */ always @(posedge \dd_pad_i[11] ) if (n638) n646 <= 1'b0 ? 1'b0 : n2802;
/* FF 15 20  0 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n757 <= 1'b0; else if (n451) n757 <= n2803;
/* FF 18 20  5 */ assign n2804 = n1513;
/* FF  5 24  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n523 <= 1'b0; else if (n2) n523 <= n2805;
/* FF  5 19  6 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n473 <= 1'b0; else if (1'b1) n473 <= n2806;
/* FF 10 26  1 */ always @(posedge \dd_pad_i[11] ) if (n552) n950 <= 1'b0 ? 1'b0 : n2807;
/* FF 10 23  6 */ assign n2808 = n1059;
/* FF  7 21  0 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n398 <= 1'b0; else if (n756) n398 <= n2809;
/* FF 14 22  2 */ assign n1286 = n2810;
/* FF 17 22  1 */ assign n2811 = n1494;
/* FF 11 28  4 */ always @(posedge \dd_pad_i[11] ) if (n227) n1091 <= 1'b0 ? 1'b0 : n2812;
/* FF  4 19  0 */ assign n2813 = n479;
/* FF  9 28  5 */ always @(posedge \dd_pad_i[11] ) if (n655) n854 <= 1'b0 ? 1'b0 : n2814;
/* FF  9 23  4 */ assign n821 = n2815;
/* FF 18 24  6 */ assign \wb_dat_o[4]  = n2816;
/* FF  6 17  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n567 <= 1'b1; else if (n346) n567 <= n2817;
/* FF 10 30  6 */ always @(posedge \dd_pad_i[11] ) if (n655) n975 <= 1'b0 ? 1'b0 : n2818;
/* FF 13 19  0 */ assign n756 = n2819;
/* FF 13 30  7 */ always @(posedge \dd_pad_i[11] ) if (n656) n1196 <= 1'b0 ? 1'b0 : n2820;
/* FF  2 17  0 */ assign n2821 = n2822;
/* FF 18 23  4 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1497 <= 1'b0; else if (n329) n1497 <= n2824;
/* FF 14 18  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n994 <= 1'b0; else if (n451) n994 <= n2825;
/* FF 11 15  3 */ assign n451 = n2826;
/* FF  5 20  7 */ assign n478 = n2827;
/* FF 10 29  0 */ always @(posedge \dd_pad_i[11] ) if (n227) n735 <= 1'b0 ? 1'b0 : n2828;
/* FF 15 27  0 */ assign n1364 = n2829;
/* FF  7 26  1 */ assign n717 = n2830;
/* FF  9 19  1 */ always @(posedge \dd_pad_i[11] ) if (n172) n791 <= 1'b0 ? 1'b0 : n2831;
/* FF 12 19  2 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n168 <= 1'b0 ? 1'b0 : n2832;
/* FF 11 29  3 */ always @(posedge \dd_pad_i[11] ) if (n655) n873 <= 1'b0 ? 1'b0 : n2833;
/* FF  4 18  3 */ assign n350 = n2834;
/* FF  9 29  6 */ always @(posedge \dd_pad_i[11] ) if (n227) n861 <= 1'b0 ? 1'b0 : n2835;
/* FF  9 16  5 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n31 <= 1'b0 ? 1'b0 : n2836;
/* FF 18 27  7 */ assign \wb_dat_o[21]  = n2837;
/* FF 16 23  0 */ assign n2838 = n1463;
/* FF 10 17  7 */ assign n884 = n2839;
/* FF 13 20  1 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n908 <= 1'b0; else if (n451) n908 <= n2840;
/* FF 12 28  0 */ assign n2841 = n1266;
/* FF 17 19  3 */ assign n2842 = n1482;
/* FF  5 26  5 */ always @(posedge \dd_pad_i[11] ) if (n478) n534 <= 1'b0 ? 1'b0 : n2843;
/* FF  5 21  4 */ assign n500 = n2844;
/* FF 10 28  3 */ always @(posedge \dd_pad_i[11] ) if (n655) n442 <= 1'b0 ? 1'b0 : n2845;
/* FF 15 24  1 */ assign io_33_30_0 = n2846;
/* FF  7 27  2 */ assign n227 = n2847;
/* FF 12 18  1 */ assign n751 = n2848;
/* FF 11 26  2 */ always @(posedge \dd_pad_i[11] ) if (n656) n1066 <= 1'b0 ? 1'b0 : n2849;
/* FF 10 14  0 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n783 <= 1'b1; else if (n4) n783 <= n2850;
/* FF  9 30  7 */ assign n870 = n2851;
/* FF 13 24  4 */ always @(posedge \dd_pad_i[11] ) if (n424) n1247 <= 1'b0 ? 1'b0 : n2852;
/* FF  6 19  0 */ always @(posedge \dd_pad_i[11] ) if (n172) n270 <= 1'b0 ? 1'b0 : n2853;
/* FF 16 22  3 */ assign n1399 = n2854;
/* FF 13 21  2 */ assign n1158 = n2855;
/* FF  2 19  2 */ assign n77 = n2856;
/* FF 17 28  2 */ assign n1474 = n2857;
/* FF  5 27  2 */ always @(posedge \dd_pad_i[11] ) if (n376) n541 <= 1'b0 ? 1'b0 : n2858;
/* FF  5 22  5 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n181 <= 1'b0; else if (1'b1) n181 <= n2859;
/* FF 10 31  2 */ always @(posedge \dd_pad_i[11] ) if (n721) n982 <= 1'b0 ? 1'b0 : n2860;
/* FF 15 25  6 */ assign n1363 = n2861;
/* FF  7 24  3 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n686 <= 1'b0; else if (1'b1) n686 <= n2862;
/* FF 12 17  0 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1017 <= 1'b1; else if (n6) n1017 <= n2863;
/* FF 14 19  1 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n900 <= 1'b1; else if (n6) n900 <= n2864;
/* FF 11 27  1 */ always @(posedge \dd_pad_i[11] ) if (n429) n1081 <= 1'b0 ? 1'b0 : n2865;
/* FF  4 27  4 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) \dd_pad_o[9]  <= 1'b0; else if (1'b1) \dd_pad_o[9]  <= n2866;
/* FF  7 14  6 */ assign n562 = n2867;
/* FF 13 25  7 */ always @(posedge \dd_pad_i[11] ) if (n1) n964 <= 1'b0 ? 1'b0 : n2868;
/* FF 16 21  2 */ assign cs1n_pad_o = n2869;
/* FF 10 19  5 */ assign n2870 = n1021;
/* FF 15 29  3 */ assign n2871 = n1434;
/* FF 13 22  3 */ assign n2872 = n1293;
/* FF  3 22  1 */ assign n296 = n403;
/* FF  4 20  2 */ assign n369 = n2873;
/* FF  7 18  5 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n452 <= 1'b0; else if (1'b1) n452 <= n2874;
/* FF  9 27  5 */ always @(posedge \dd_pad_i[11] ) if (n227) n772 <= 1'b0 ? 1'b0 : n2875;
/* FF  7 25  4 */ always @(posedge \dd_pad_i[11] ) if (n429) n713 <= 1'b0 ? 1'b0 : n2876;
/* FF  1 20  1 */ assign n65 = n2877;
/* FF 17 18  5 */ assign n1438 = n2878;
/* FF 11 24  0 */ assign n760 = n2879;
/* FF  4 26  7 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n229 <= 1'b0; else if (n2) n229 <= n2880;
/* FF  4 23  4 */ assign n113 = n2881;
/* FF  9 24  1 */ always @(posedge \dd_pad_i[11] ) if (n1) n526 <= 1'b0 ? 1'b0 : n2882;
/* FF 13 26  6 */ always @(posedge \dd_pad_i[11] ) if (n1) n643 <= 1'b0 ? 1'b0 : n2883;
/* FF 14 28  3 */ assign n1313 = n2884;
/* FF  2 22  2 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n196 <= 1'b0 ? 1'b0 : n2885;
/* FF 11 22  3 */ assign n2886 = n1150;
/* FF  5 16  6 */ assign n346 = n2887;
/* FF 10 18  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n887 <= 1'b0; else if (n563) n887 <= n2888;
/* FF  3 23  2 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) io_14_33_0 <= 1'b0; else if (1'b1) io_14_33_0 <= n2889;
/* FF  2 21  4 */ assign n189 = n2890;
/* FF 12 20  4 */ always @(posedge \dd_pad_i[11] , posedge n5) if (n5) n1129 <= 1'b0; else if (n4) n1129 <= n2891;
/* FF  3 14  6 */ always @(posedge \dd_pad_i[11] ) if (1'b1) n238 <= 1'b0 ? 1'b0 : n2892;
/* FF  7 19  6 */ assign n410 = n2893;
/* FF  9 20  4 */ always @(posedge \dd_pad_i[11] ) if (n478) n803 <= 1'b0 ? 1'b0 : n2894;
/* FF 12 23  6 */ assign n1154 = n2895;

// Warning: unmatched port '\dd_pad_i[4] '
// Warning: unmatched port '\wb_dat_o[20] '
// Warning: unmatched port 'wb_ack_o'
// Warning: unmatched port '\da_pad_o[0] '
// Warning: unmatched port '\wb_dat_i[31] '
// Warning: unmatched port 'DMA_Ack'
// Warning: unmatched port '\dd_pad_o[4] '
// Warning: unmatched port 'wb_rst_i'
// Warning: unmatched port '\wb_dat_i[13] '
// Warning: unmatched port '\wb_dat_i[10] '
// Warning: unmatched port '\wb_dat_o[10] '
// Warning: unmatched port '\wb_dat_i[7] '
// Warning: unmatched port '\dd_pad_o[7] '
// Warning: unmatched port '\wb_dat_i[9] '
// Warning: unmatched port 'intrq_pad_i'
// Warning: unmatched port '\wb_dat_o[13] '
// Warning: unmatched port '\wb_adr_i[6] '
// Warning: unmatched port '\wb_adr_i[2] '
// Warning: unmatched port '\wb_sel_i[2] '
// Warning: unmatched port '\wb_dat_o[22] '
// Warning: unmatched port '\wb_dat_i[26] '
// Warning: unmatched port '\dd_pad_o[1] '
// Warning: unmatched port '\wb_dat_i[6] '
// Warning: unmatched port '\wb_dat_o[2] '
// Warning: unmatched port '\wb_dat_o[17] '
// Warning: unmatched port '\wb_dat_o[14] '
// Warning: unmatched port '\wb_dat_i[15] '
// Warning: unmatched port '\dd_pad_o[10] '
// Warning: unmatched port '\wb_dat_o[12] '

endmodule

