
module chip (input clk, output \rco[191] , output \rco[22] , output \rco[184] , output \rco[187] , output \rco[193] , output \rco[194] , output \rco[195] , output \rco[154] , output \rco[156] , output \rco[155] , output \rco[21] , output \rco[159] , output \rco[160] , output \rco[131] , output \rco[161] , output \rco[123] , output \rco[10] , output \rco[130] , output \rco[3] , output \rco[12] , output \rco[24] , output \rco[11] , output \rco[0] , output \rco[13] , output \rco[16] , output \rco[19] , output \rco[7] , output \rco[8] , output \rco[5] , output \rco[4] , output \rco[27] , output \rco[28] , output \rco[29] , output \rco[6] , output \rco[2] , output \rco[18] , output \rco[14] , output \rco[20] , output \rco[17] , output \rco[23] , output \rco[15] , output \rco[26] , output \rco[25] , output \rco[127] , output \rco[9] , output \rco[125] , output \rco[124] , output \rco[126] , output \rco[148] , output \rco[147] , output \rco[134] , output \rco[153] , output \rco[103] , output \rco[158] , output \rco[157] , output \rco[110] , output \rco[135] , output \rco[136] , output \rco[99] , output \rco[137] , output \rco[122] , output \rco[199] , output \rco[67] , input en_in, output \rco[166] , output \rco[132] , output \rco[113] , output \rco[42] , output \rco[43] , output \rco[107] , output \rco[145] , output \rco[108] , output \rco[109] , output \rco[165] , output \rco[164] , output \rco[152] , output \rco[112] , output \rco[68] , output \rco[162] , output \rco[172] , output \rco[151] , output \rco[69] , output \rco[102] , output \rco[54] , output \rco[97] , output \rco[93] , output \rco[60] , output \rco[143] , output \rco[120] , output \rco[106] , output \rco[105] , output \rco[61] , output \rco[104] , output \rco[62] , output \rco[53] , output \rco[65] , output \rco[40] , output \rco[1] , output \rco[101] , output \rco[100] , output \rco[88] , output \rco[39] , output \rco[149] , output \rco[83] , output \rco[118] , output \rco[119] , output \rco[115] , output \rco[87] , output \rco[142] , output \rco[138] , output \rco[116] , output \rco[111] , output \rco[198] , output \rco[58] , output \rco[86] , output \rco[90] , output \rco[114] , output \rco[173] , output \rco[182] , output \rco[98] , output \rco[192] , output \rco[30] , output \rco[179] , output \rco[91] , output \rco[85] , output \rco[144] , output \rco[141] , output \rco[41] , output \rco[183] , output \rco[117] , output \rco[133] , output \rco[180] , output \rco[176] , output \rco[150] , output \rco[37] , output \rco[51] , output \rco[181] , output \rco[34] , output \rco[84] , output \rco[89] , output \rco[92] , output \rco[96] , output \rco[52] , output \rco[56] , output \rco[197] , output \rco[174] , output \rco[146] , output \rco[47] , output \rco[74] , output \rco[57] , output \rco[31] , output \rco[196] , output \rco[169] , output \rco[168] , output \rco[94] , output \rco[95] , output \rco[44] , output \rco[48] , output \rco[59] , output \rco[175] , output \rco[46] , output \rco[177] , output \rco[45] , output \rco[55] , output \rco[121] , output \rco[66] , output \rco[38] , output \rco[188] , output \rco[178] , output \rco[82] , output \rco[64] , output \rco[63] , output \rco[33] , output \rco[36] , output \rco[35] , output \rco[79] , output \rco[78] , output \rco[32] , output \rco[81] , output \rco[70] , output \rco[171] , output \rco[170] , output \rco[167] , output \rco[163] , output \rco[139] , output \rco[50] , output \rco[75] , output \rco[76] , output \rco[77] , output \rco[80] , output \rco[72] , output \rco[140] , output \rco[73] , output \rco[71] , output \rco[186] , output \rco[185] , output \rco[190] , output \rco[189] , output \rco[129] , output \rco[128] , output \rco[49] );

wire n1, n2, clk, \rco[191] , \rco[22] , \rco[184] , \rco[187] , \rco[193] , \rco[194] , \rco[195] ;
wire \rco[154] , \rco[156] , \rco[155] , \rco[21] , n21, \rco[159] , \rco[160] , \rco[131] , \rco[161] , \rco[123] ;
wire \rco[10] , \rco[130] , n37, \rco[3] , n39, \rco[12] , \rco[24] , \rco[11] , n54, n56;
wire \rco[13] , \rco[16] , n59, \rco[19] , n76, n77, n78, n79, \rco[7] , \rco[8] ;
wire \rco[5] , n83, \rco[4] , n85, \rco[27] , \rco[28] , \rco[29] , \rco[6] , n115, n116;
wire n117, n118, n119, n121, \rco[2] , \rco[18] , n126, \rco[14] , \rco[20] , \rco[17] ;
wire \rco[23] , \rco[15] , \rco[26] , \rco[25] , \rco[127] , \rco[9] , \rco[125] , \rco[124] , \rco[126] , \rco[148] ;
wire \rco[147] , \rco[134] , \rco[153] , \rco[103] , \rco[158] , \rco[157] , n153, n168, n175, n184;
wire n195, n197, n202, n203, n207, n215, n216, n224, \rco[110] , n246;
wire \rco[135] , \rco[136] , n251, n260, n277, n285, n286, n288, n290, n302;
wire n325, n328, n329, n335, \rco[99] , n338, n339, n340, n341, n349;
wire n350, n351, n352, n360, n363, \rco[137] , \rco[122] , \rco[199] , \rco[67] , en_in;
wire \rco[166] , n402, n403, n404, n405, n406, n407, n410, n411, n438;
wire n439, n440, n454, n455, n456, n458, n459, n460, n461, n462;
wire \rco[132] , \rco[113] , \rco[42] , n501, n502, n503, n511, n512, n513, n514;
wire n545, n546, n547, n549, n552, n553, n554, n562, n563, n564;
wire n567, \rco[43] , \rco[107] , n570, n588, n589, n629, n630, \rco[145] , n645;
wire n657, n658, n659, n660, n670, n671, n672, n673, n675, n676;
wire n677, n695, n697, \rco[108] , \rco[109] , \rco[165] , \rco[164] , \rco[152] , n718, n726;
wire n727, n728, n732, n733, n736, n739, n750, n765, n766, n767;
wire n768, n777, n778, n779, n780, n781, n782, \rco[112] , n796, n804;
wire \rco[68] , \rco[162] , n807, \rco[172] , n809, n814, n815, n816, n817, n818;
wire n819, n820, n821, \rco[151] , n823, n850, \rco[69] , n891, n900, n912;
wire n922, n954, \rco[102] , n961, n962, \rco[54] , \rco[97] , \rco[93] , n977, n982;
wire n983, n988, n990, n996, n1015, n1030, \rco[60] , \rco[143] , n1056, n1057;
wire n1065, n1069, \rco[120] , \rco[106] , n1089, n1090, n1091, \rco[105] , \rco[61] , \rco[104] ;
wire \rco[62] , n1115, \rco[53] , \rco[65] , \rco[40] , n1131, \rco[1] , n1136, n1137, n1154;
wire n1155, n1176, n1177, n1178, n1187, n1188, n1196, n1197, n1205, n1213;
wire n1222, n1243, n1245, n1246, \rco[101] , \rco[100] , n1271, \rco[88] , \rco[39] , \rco[149] ;
wire \rco[83] , n1335, n1336, n1337, \rco[118] , n1339, n1340, n1347, n1355, n1356;
wire n1357, \rco[119] , \rco[115] , n1375, n1383, n1384, n1393, n1394, n1402, \rco[87] ;
wire n1460, n1461, n1491, n1500, n1501, \rco[142] , \rco[138] , n1511, n1512, n1520;
wire n1521, n1532, \rco[116] , \rco[111] , n1541, n1542, \rco[198] , n1557, n1559, n1560;
wire \rco[58] , \rco[86] , \rco[90] , n1577, n1584, n1592, n1601, n1602, n1620, n1621;
wire n1622, n1623, n1624, n1625, n1666, n1671, n1672, n1673, n1674, n1675;
wire n1683, n1685, \rco[114] , n1697, n1698, n1699, n1700, n1710, \rco[173] , \rco[182] ;
wire \rco[98] , n1741, n1742, n1743, n1744, n1752, n1761, n1771, n1773, n1774;
wire n1775, n1776, n1791, n1792, n1825, n1826, n1835, n1843, n1844, n1845;
wire n1860, n1861, n1862, n1863, n1871, n1873, n1874, n1876, n1877, n1878;
wire \rco[192] , n1881, \rco[30] , \rco[179] , \rco[91] , \rco[85] , n1887, \rco[144] , \rco[141] , n1914;
wire n1933, n1936, \rco[41] , n1951, n1952, n1953, n1954, n1982, n1998, n1999;
wire n2000, n2003, \rco[183] , n2017, n2020, \rco[117] , \rco[133] , \rco[180] , \rco[176] , \rco[150] ;
wire n2037, n2045, n2054, n2055, n2056, n2057, \rco[37] , \rco[51] , n2076, n2085;
wire n2094, n2109, n2110, n2111, n2112, n2113, n2123, n2164, n2174, n2175;
wire \rco[181] , n2195, n2196, \rco[34] , n2207, \rco[84] , \rco[89] , \rco[92] , n2229, n2230;
wire n2240, n2241, \rco[96] , n2247, n2257, n2258, n2259, n2260, n2270, n2271;
wire n2272, n2282, n2283, \rco[52] , \rco[56] , n2303, n2304, n2306, n2307, n2308;
wire n2322, n2323, n2324, n2325, n2347, n2348, n2358, n2384, \rco[197] , \rco[174] ;
wire \rco[146] , n2451, n2460, \rco[47] , n2470, \rco[74] , n2495, n2496, \rco[57] , n2511;
wire n2519, n2520, \rco[31] , n2523, n2524, n2534, n2535, n2536, n2538, n2540;
wire n2551, n2553, n2562, n2564, n2573, n2574, n2575, n2590, n2591, n2592;
wire n2593, n2602, n2612, n2613, n2614, n2615, n2628, \rco[196] , \rco[169] , \rco[168] ;
wire \rco[94] , \rco[95] , n2670, n2671, \rco[44] , n2678, n2679, n2680, n2682, \rco[48] ;
wire n2697, n2707, n2708, n2715, n2725, n2726, n2727, n2728, n2730, n2731;
wire \rco[59] , n2757, n2760, n2775, n2785, n2786, n2787, n2812, n2813, \rco[175] ;
wire \rco[46] , n2841, n2844, n2852, n2853, n2854, n2855, n2856, n2859, n2865;
wire n2866, n2881, n2886, n2896, n2897, n2910, n2952, n2953, n2961, n2970;
wire n2971, \rco[177] , \rco[45] , n2989, n3006, n3007, n3008, n3009, n3029, n3030;
wire n3031, \rco[55] , n3033, n3034, n3045, n3065, n3067, n3068, n3069, n3087;
wire n3104, n3112, n3113, n3114, n3124, n3141, n3142, \rco[121] , n3158, n3175;
wire n3198, n3199, \rco[66] , n3216, \rco[38] , n3233, n3249, n3258, n3259, n3260;
wire n3261, n3262, n3295, \rco[188] , \rco[178] , \rco[82] , n3330, n3331, \rco[64] , \rco[63] ;
wire n3351, n3352, n3368, n3376, \rco[33] , n3393, \rco[36] , n3411, n3421, n3422;
wire n3424, n3432, n3457, n3458, n3459, n3460, n3462, n3464, n3465, n3466;
wire n3467, n3468, \rco[35] , n3470, \rco[79] , n3488, \rco[78] , n3525, n3526, n3527;
wire n3553, \rco[32] , n3555, \rco[81] , n3593, n3594, n3603, n3604, n3605, \rco[70] ;
wire n3621, n3639, n3640, n3664, n3665, n3666, n3683, n3684, n3685, n3686;
wire n3703, n3704, n3718, n3733, n3749, n3750, n3751, n3752, n3765, \rco[171] ;
wire n3785, n3786, \rco[170] , n3788, \rco[167] , \rco[163] , n3814, n3815, \rco[139] , \rco[50] ;
wire \rco[75] , \rco[76] , \rco[77] , \rco[80] , n3848, n3876, \rco[72] , n3892, \rco[140] , \rco[73] ;
wire \rco[71] , \rco[186] , \rco[185] , \rco[190] , \rco[189] , \rco[129] , \rco[128] , \rco[49] , n3911, n3912;
wire n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922;
wire n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932;
wire n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942;
wire n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952;
wire n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962;
wire n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972;
wire n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982;
wire n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992;
wire n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002;
wire n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012;
wire n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022;
wire n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032;
wire n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042;
wire n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052;
wire n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062;
wire n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072;
wire n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082;
wire n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092;
wire n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102;
wire n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112;
wire n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122;
wire n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132;
wire n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142;
wire n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152;
wire n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162;
wire n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172;
wire n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182;
wire n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192;
wire n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202;
wire n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212;
wire n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222;
wire n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232;
wire n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242;
wire n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252;
wire n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262;
wire n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272;
wire n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282;
wire n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292;
wire n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302;
wire n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312;
wire n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322;
wire n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332;
wire n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342;
wire n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352;
wire n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362;
wire n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372;
wire n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382;
wire n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392;
wire n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402;
wire n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412;
wire n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422;
wire n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432;
wire n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442;
wire n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452;
wire n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462;
wire n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472;
wire n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482;
wire n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492;
wire n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502;
wire n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512;
wire n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522;
wire n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532;
wire n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542;
wire n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552;
wire n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562;
wire n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572;
wire n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582;
wire n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592;
wire n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602;
wire n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612;
wire n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622;
wire n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632;
wire n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642;
wire n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652;
wire n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662;
wire n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672;
wire n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682;
wire n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692;
wire n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702;
wire n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712;
wire n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722;
wire n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732;
wire n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742;
wire n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752;
wire n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762;
wire n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772;
wire n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782;
wire n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792;
wire n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802;
wire n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812;
wire n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822;
wire n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832;
wire n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842;
wire n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852;
wire n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862;
wire n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872;
wire n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882;
wire n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892;
wire n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902;
wire n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912;
wire n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922;
wire n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932;
wire n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942;
wire n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952;
wire n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962;
wire n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972;
wire n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982;
wire n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992;
wire n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002;
wire n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012;
wire n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022;
wire n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032;
wire n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042;
wire n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052;
wire n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062;
wire n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072;
wire n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082;
wire n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092;
wire n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102;
wire n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112;
wire n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122;
wire n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132;
wire n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142;
wire n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152;
wire n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162;
wire n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172;
wire n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182;
wire n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192;
wire n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202;
wire n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212;
wire n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222;
wire n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232;
wire n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242;
wire n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252;
wire n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262;
wire n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272;
wire n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282;
wire n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292;
wire n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302;
wire n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312;
wire n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322;
wire n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332;
wire n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342;
wire n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352;
wire n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362;
wire n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372;
wire n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382;
wire n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392;
wire n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402;
wire n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412;
wire n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422;
wire n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432;
wire n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442;
wire n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452;
wire n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462;
wire n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472;
wire n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482;
wire n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492;
wire n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502;
wire n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512;
wire n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522;
wire n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532;
wire n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542;
wire n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552;
wire n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562;
wire n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572;
wire n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582;
wire n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592;
wire n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602;
wire n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612;
wire n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622;
wire n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632;
wire n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642;
wire n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652;
wire n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662;
wire n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672;
wire n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682;
wire n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692;
wire n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702;
wire n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712;
wire n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722;
wire n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732;
wire n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742;
wire n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752;
wire n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762;
wire n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772;
wire n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782;
wire n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792;
wire n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802;
wire n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812;
wire n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822;
wire n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832;
wire n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842;
wire n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852;
wire n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862;
wire n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872;
wire n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882;
wire n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892;
wire n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902;
wire n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912;
wire n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922;
wire n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932;
wire n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942;
wire n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952;
wire n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962;
wire n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972;
wire n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982;
wire n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992;
wire n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002;
wire n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012;
wire n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022;
wire n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032;
wire n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042;
wire n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052;
wire n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062;
wire n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072;
wire n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082;
wire n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092;
wire n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102;
wire n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112;
wire n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122;
wire n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132;
wire n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142;
wire n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152;
wire n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162;
wire n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172;
wire n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182;
wire n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192;
wire n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202;
wire n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212;
wire n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222;
wire n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232;
wire n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242;
wire n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252;
wire n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262;
wire n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272;
wire n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282;
wire n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292;
wire n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302;
wire n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312;
wire n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322;
wire n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332;
wire n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342;
wire n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352;
wire n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362;
wire n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372;
wire n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382;
wire n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392;
wire n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402;
wire n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412;
wire n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422;
wire n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432;
wire n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442;
wire n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452;
wire n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462;
wire n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472;
wire n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482;
wire n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492;
wire n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502;
wire n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512;
wire n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522;
wire n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532;
wire n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542;
wire n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552;
wire n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562;
wire n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572;
wire n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582;
wire n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592;
wire n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602;
wire n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612;
wire n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622;
wire n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632;
wire n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642;
wire n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652;
wire n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662;
wire n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672;
wire n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682;
wire n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692;
wire n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702;
wire n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712;
wire n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722;
wire n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732;
wire n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742;
wire n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752;
wire n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762;
wire n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772;
wire n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782;
wire n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792;
wire n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802;
wire n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812;
wire n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822;
wire n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832;
wire n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842;
wire n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852;
wire n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862;
wire n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872;
wire n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882;
wire n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892;
wire n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902;
wire n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912;
wire n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922;
wire n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932;
wire n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942;
wire n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952;
wire n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962;
wire n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972;
wire n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982;
wire n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992;
wire n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002;
wire n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012;
wire n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022;
wire n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032;
wire n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042;
wire n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052;
wire n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062;
wire n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072;
wire n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082;
wire n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092;
wire n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102;
wire n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112;
wire n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122;
wire n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132;
wire n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142;
wire n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152;
wire n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162;
wire n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172;
wire n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182;
wire n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192;
wire n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202;
wire n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212;
wire n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222;
wire n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232;
wire n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242;
wire n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252;
wire n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262;
wire n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272;
wire n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282;
wire n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292;
wire n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302;
wire n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312;
wire n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322;
wire n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332;
wire n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342;
wire n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352;
wire n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362;
wire n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372;
wire n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382;
wire n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392;
wire n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402;
wire n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412;
wire n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422;
wire n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432;
wire n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442;
wire n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452;
wire n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462;
wire n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472;
wire n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482;
wire n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492;
wire n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502;
wire n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512;
wire n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522;
wire n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532;
wire n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542;
wire n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552;
wire n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562;
wire n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572;
wire n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582;
wire n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592;
wire n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602;
wire n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612;
wire n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622;
wire n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632;
wire n7633, n7634, n7635, n7636, n7637, n7638;
reg n14 = 0, n15 = 0, n16 = 0, n17 = 0, n18 = 0, n19 = 0, n24 = 0, n28 = 0, n29 = 0, n30 = 0;
reg n31 = 0, n32 = 0, n33 = 0, n34 = 0, n40 = 0, n41 = 0, n42 = 0, n46 = 0, n47 = 0, n48 = 0;
reg n49 = 0, n50 = 0, n51 = 0, n52 = 0, n53 = 0, \rco[0]  = 0, n60 = 0, n61 = 0, n62 = 0, n63 = 0;
reg n64 = 0, n65 = 0, n66 = 0, n68 = 0, n69 = 0, n70 = 0, n71 = 0, n72 = 0, n73 = 0, n74 = 0;
reg n75 = 0, n86 = 0, n87 = 0, n88 = 0, n89 = 0, n90 = 0, n91 = 0, n92 = 0, n93 = 0, n94 = 0;
reg n98 = 0, n99 = 0, n100 = 0, n101 = 0, n102 = 0, n103 = 0, n104 = 0, n105 = 0, n106 = 0, n107 = 0;
reg n108 = 0, n109 = 0, n110 = 0, n111 = 0, n113 = 0, n114 = 0, n120 = 0, n122 = 0, n123 = 0, n129 = 0;
reg n137 = 0, n148 = 0, n149 = 0, n150 = 0, n151 = 0, n152 = 0, n154 = 0, n155 = 0, n156 = 0, n157 = 0;
reg n158 = 0, n159 = 0, n160 = 0, n161 = 0, n162 = 0, n163 = 0, n164 = 0, n165 = 0, n166 = 0, n167 = 0;
reg n169 = 0, n170 = 0, n171 = 0, n172 = 0, n173 = 0, n174 = 0, n176 = 0, n177 = 0, n178 = 0, n179 = 0;
reg n180 = 0, n181 = 0, n182 = 0, n183 = 0, n185 = 0, n186 = 0, n187 = 0, n188 = 0, n189 = 0, n190 = 0;
reg n191 = 0, n192 = 0, n193 = 0, n194 = 0, n196 = 0, n198 = 0, n199 = 0, n200 = 0, n201 = 0, n204 = 0;
reg n205 = 0, n206 = 0, n208 = 0, n209 = 0, n210 = 0, n211 = 0, n212 = 0, n213 = 0, n214 = 0, n217 = 0;
reg n218 = 0, n219 = 0, n220 = 0, n221 = 0, n222 = 0, n223 = 0, n225 = 0, n226 = 0, n227 = 0, n228 = 0;
reg n229 = 0, n230 = 0, n231 = 0, n232 = 0, n233 = 0, n234 = 0, n235 = 0, n236 = 0, n237 = 0, n238 = 0;
reg n239 = 0, n240 = 0, n241 = 0, n242 = 0, n243 = 0, n244 = 0, n247 = 0, n250 = 0, n252 = 0, n253 = 0;
reg n254 = 0, n255 = 0, n256 = 0, n257 = 0, n258 = 0, n259 = 0, n261 = 0, n262 = 0, n263 = 0, n264 = 0;
reg n265 = 0, n266 = 0, n267 = 0, n268 = 0, n269 = 0, n270 = 0, n271 = 0, n272 = 0, n273 = 0, n274 = 0;
reg n275 = 0, n276 = 0, n278 = 0, n279 = 0, n280 = 0, n281 = 0, n282 = 0, n283 = 0, n284 = 0, n287 = 0;
reg n289 = 0, n291 = 0, n292 = 0, n293 = 0, n294 = 0, n295 = 0, n296 = 0, n297 = 0, n298 = 0, n299 = 0;
reg n300 = 0, n301 = 0, n303 = 0, n304 = 0, n305 = 0, n306 = 0, n307 = 0, n308 = 0, n309 = 0, n310 = 0;
reg n311 = 0, n312 = 0, n313 = 0, n314 = 0, n315 = 0, n316 = 0, n317 = 0, n318 = 0, n319 = 0, n320 = 0;
reg n321 = 0, n322 = 0, n323 = 0, n324 = 0, n326 = 0, n327 = 0, n330 = 0, n331 = 0, n332 = 0, n333 = 0;
reg n334 = 0, n336 = 0, n342 = 0, n343 = 0, n344 = 0, n345 = 0, n346 = 0, n347 = 0, n348 = 0, n353 = 0;
reg n354 = 0, n355 = 0, n356 = 0, n357 = 0, n358 = 0, n359 = 0, n361 = 0, n362 = 0, n365 = 0, n371 = 0;
reg n372 = 0, n373 = 0, n374 = 0, n375 = 0, n376 = 0, n377 = 0, n378 = 0, n379 = 0, n380 = 0, n381 = 0;
reg n382 = 0, n383 = 0, n384 = 0, n385 = 0, n386 = 0, n387 = 0, n388 = 0, n389 = 0, n390 = 0, n391 = 0;
reg n392 = 0, n393 = 0, n394 = 0, n395 = 0, n396 = 0, n397 = 0, n398 = 0, n399 = 0, n400 = 0, n401 = 0;
reg n408 = 0, n409 = 0, n412 = 0, n413 = 0, n414 = 0, n415 = 0, n416 = 0, n417 = 0, n418 = 0, n419 = 0;
reg n420 = 0, n421 = 0, n422 = 0, n423 = 0, n424 = 0, n425 = 0, n426 = 0, n427 = 0, n428 = 0, n429 = 0;
reg n430 = 0, n431 = 0, n432 = 0, n433 = 0, n434 = 0, n435 = 0, n436 = 0, n437 = 0, n441 = 0, n442 = 0;
reg n443 = 0, n444 = 0, n445 = 0, n446 = 0, n447 = 0, n448 = 0, n449 = 0, n450 = 0, n451 = 0, n452 = 0;
reg n453 = 0, n457 = 0, n463 = 0, n465 = 0, n468 = 0, n469 = 0, n470 = 0, n471 = 0, n472 = 0, n473 = 0;
reg n474 = 0, n475 = 0, n476 = 0, n477 = 0, n478 = 0, n479 = 0, n480 = 0, n481 = 0, n482 = 0, n483 = 0;
reg n484 = 0, n485 = 0, n486 = 0, n487 = 0, n488 = 0, n489 = 0, n490 = 0, n491 = 0, n492 = 0, n493 = 0;
reg n494 = 0, n495 = 0, n496 = 0, n497 = 0, n498 = 0, n499 = 0, n500 = 0, n504 = 0, n505 = 0, n506 = 0;
reg n507 = 0, n508 = 0, n509 = 0, n510 = 0, n515 = 0, n516 = 0, n517 = 0, n518 = 0, n519 = 0, n520 = 0;
reg n521 = 0, n522 = 0, n523 = 0, n524 = 0, n525 = 0, n526 = 0, n527 = 0, n528 = 0, n529 = 0, n530 = 0;
reg n531 = 0, n532 = 0, n533 = 0, n534 = 0, n535 = 0, n536 = 0, n537 = 0, n538 = 0, n539 = 0, n540 = 0;
reg n541 = 0, n542 = 0, n543 = 0, n544 = 0, n548 = 0, n550 = 0, n551 = 0, n555 = 0, n556 = 0, n557 = 0;
reg n558 = 0, n559 = 0, n560 = 0, n561 = 0, n565 = 0, n566 = 0, n571 = 0, n572 = 0, n573 = 0, n574 = 0;
reg n575 = 0, n576 = 0, n577 = 0, n578 = 0, n579 = 0, n580 = 0, n581 = 0, n582 = 0, n583 = 0, n584 = 0;
reg n585 = 0, n586 = 0, n587 = 0, n590 = 0, n591 = 0, n592 = 0, n593 = 0, n594 = 0, n595 = 0, n596 = 0;
reg n597 = 0, n598 = 0, n599 = 0, n600 = 0, n601 = 0, n602 = 0, n603 = 0, n604 = 0, n605 = 0, n606 = 0;
reg n607 = 0, n608 = 0, n609 = 0, n610 = 0, n611 = 0, n612 = 0, n613 = 0, n614 = 0, n615 = 0, n616 = 0;
reg n617 = 0, n618 = 0, n619 = 0, n620 = 0, n621 = 0, n622 = 0, n623 = 0, n624 = 0, n625 = 0, n626 = 0;
reg n627 = 0, n628 = 0, n631 = 0, n632 = 0, n633 = 0, n634 = 0, n635 = 0, n636 = 0, n637 = 0, n638 = 0;
reg n639 = 0, n640 = 0, n641 = 0, n642 = 0, n643 = 0, n646 = 0, n647 = 0, n648 = 0, n649 = 0, n650 = 0;
reg n651 = 0, n652 = 0, n653 = 0, n654 = 0, n655 = 0, n656 = 0, n661 = 0, n662 = 0, n663 = 0, n664 = 0;
reg n665 = 0, n666 = 0, n667 = 0, n668 = 0, n669 = 0, n674 = 0, n678 = 0, n679 = 0, n680 = 0, n681 = 0;
reg n682 = 0, n683 = 0, n684 = 0, n685 = 0, n686 = 0, n687 = 0, n688 = 0, n689 = 0, n690 = 0, n691 = 0;
reg n692 = 0, n693 = 0, n694 = 0, n696 = 0, n698 = 0, n699 = 0, n700 = 0, n706 = 0, n707 = 0, n708 = 0;
reg n709 = 0, n710 = 0, n711 = 0, n712 = 0, n713 = 0, n714 = 0, n715 = 0, n716 = 0, n717 = 0, n719 = 0;
reg n720 = 0, n721 = 0, n722 = 0, n723 = 0, n724 = 0, n725 = 0, n729 = 0, n730 = 0, n731 = 0, n734 = 0;
reg n735 = 0, n737 = 0, n738 = 0, n740 = 0, n741 = 0, n742 = 0, n743 = 0, n744 = 0, n745 = 0, n746 = 0;
reg n747 = 0, n748 = 0, n749 = 0, n751 = 0, n752 = 0, n753 = 0, n754 = 0, n755 = 0, n756 = 0, n757 = 0;
reg n758 = 0, n759 = 0, n760 = 0, n761 = 0, n762 = 0, n763 = 0, n764 = 0, n769 = 0, n770 = 0, n771 = 0;
reg n772 = 0, n773 = 0, n774 = 0, n775 = 0, n776 = 0, n783 = 0, n784 = 0, n785 = 0, n786 = 0, n787 = 0;
reg n788 = 0, n789 = 0, n790 = 0, n791 = 0, n792 = 0, n793 = 0, n795 = 0, n797 = 0, n798 = 0, n799 = 0;
reg n800 = 0, n801 = 0, n802 = 0, n803 = 0, n810 = 0, n811 = 0, n812 = 0, n813 = 0, n824 = 0, n825 = 0;
reg n826 = 0, n827 = 0, n828 = 0, n829 = 0, n830 = 0, n831 = 0, n832 = 0, n833 = 0, n834 = 0, n835 = 0;
reg n836 = 0, n837 = 0, n838 = 0, n839 = 0, n840 = 0, n841 = 0, n842 = 0, n843 = 0, n844 = 0, n845 = 0;
reg n846 = 0, n847 = 0, n848 = 0, n849 = 0, n851 = 0, n852 = 0, n853 = 0, n855 = 0, n856 = 0, n857 = 0;
reg n858 = 0, n859 = 0, n860 = 0, n861 = 0, n862 = 0, n863 = 0, n864 = 0, n865 = 0, n866 = 0, n867 = 0;
reg n868 = 0, n869 = 0, n870 = 0, n871 = 0, n872 = 0, n873 = 0, n874 = 0, n875 = 0, n876 = 0, n877 = 0;
reg n878 = 0, n879 = 0, n880 = 0, n881 = 0, n882 = 0, n883 = 0, n884 = 0, n885 = 0, n886 = 0, n887 = 0;
reg n888 = 0, n889 = 0, n890 = 0, n892 = 0, n893 = 0, n894 = 0, n895 = 0, n896 = 0, n897 = 0, n898 = 0;
reg n899 = 0, n901 = 0, n902 = 0, n903 = 0, n904 = 0, n905 = 0, n906 = 0, n907 = 0, n908 = 0, n909 = 0;
reg n910 = 0, n911 = 0, n913 = 0, n914 = 0, n915 = 0, n916 = 0, n917 = 0, n918 = 0, n919 = 0, n920 = 0;
reg n921 = 0, n923 = 0, n924 = 0, n925 = 0, n926 = 0, n927 = 0, n928 = 0, n929 = 0, n930 = 0, n931 = 0;
reg n932 = 0, n933 = 0, n934 = 0, n935 = 0, n936 = 0, n937 = 0, n938 = 0, n939 = 0, n940 = 0, n941 = 0;
reg n942 = 0, n943 = 0, n944 = 0, n945 = 0, n946 = 0, n947 = 0, n948 = 0, n949 = 0, n950 = 0, n951 = 0;
reg n952 = 0, n953 = 0, n955 = 0, n956 = 0, n957 = 0, n958 = 0, n959 = 0, n966 = 0, n967 = 0, n968 = 0;
reg n969 = 0, n970 = 0, n971 = 0, n972 = 0, n973 = 0, n974 = 0, n975 = 0, n976 = 0, n978 = 0, n979 = 0;
reg n980 = 0, n981 = 0, n984 = 0, n985 = 0, n986 = 0, n987 = 0, n989 = 0, n991 = 0, n992 = 0, n993 = 0;
reg n994 = 0, n995 = 0, n997 = 0, n998 = 0, n999 = 0, n1000 = 0, n1001 = 0, n1002 = 0, n1003 = 0, n1004 = 0;
reg n1005 = 0, n1006 = 0, n1007 = 0, n1008 = 0, n1009 = 0, n1010 = 0, n1011 = 0, n1012 = 0, n1013 = 0, n1014 = 0;
reg n1016 = 0, n1017 = 0, n1018 = 0, n1019 = 0, n1020 = 0, n1021 = 0, n1022 = 0, n1023 = 0, n1024 = 0, n1025 = 0;
reg n1026 = 0, n1027 = 0, n1028 = 0, n1029 = 0, n1031 = 0, n1032 = 0, n1033 = 0, n1034 = 0, n1035 = 0, n1036 = 0;
reg n1037 = 0, n1038 = 0, n1039 = 0, n1040 = 0, n1042 = 0, n1043 = 0, n1044 = 0, n1045 = 0, n1046 = 0, n1047 = 0;
reg n1048 = 0, n1049 = 0, n1050 = 0, n1051 = 0, n1052 = 0, n1053 = 0, n1054 = 0, n1058 = 0, n1059 = 0, n1060 = 0;
reg n1061 = 0, n1062 = 0, n1063 = 0, n1064 = 0, n1066 = 0, n1067 = 0, n1068 = 0, n1070 = 0, n1072 = 0, n1073 = 0;
reg n1074 = 0, n1075 = 0, n1076 = 0, n1077 = 0, n1078 = 0, n1079 = 0, n1080 = 0, n1081 = 0, n1082 = 0, n1083 = 0;
reg n1084 = 0, n1085 = 0, n1086 = 0, n1087 = 0, n1093 = 0, n1094 = 0, n1095 = 0, n1096 = 0, n1097 = 0, n1098 = 0;
reg n1099 = 0, n1101 = 0, n1102 = 0, n1103 = 0, n1104 = 0, n1105 = 0, n1106 = 0, n1107 = 0, n1108 = 0, n1109 = 0;
reg n1110 = 0, n1111 = 0, n1113 = 0, n1119 = 0, n1120 = 0, n1121 = 0, n1122 = 0, n1123 = 0, n1124 = 0, n1125 = 0;
reg n1126 = 0, n1127 = 0, n1128 = 0, n1129 = 0, n1130 = 0, n1132 = 0, n1133 = 0, n1134 = 0, n1138 = 0, n1139 = 0;
reg n1140 = 0, n1141 = 0, n1142 = 0, n1143 = 0, n1144 = 0, n1145 = 0, n1146 = 0, n1147 = 0, n1148 = 0, n1149 = 0;
reg n1150 = 0, n1151 = 0, n1152 = 0, n1153 = 0, n1156 = 0, n1157 = 0, n1158 = 0, n1159 = 0, n1160 = 0, n1161 = 0;
reg n1162 = 0, n1163 = 0, n1164 = 0, n1165 = 0, n1166 = 0, n1167 = 0, n1168 = 0, n1169 = 0, n1170 = 0, n1171 = 0;
reg n1172 = 0, n1173 = 0, n1174 = 0, n1175 = 0, n1179 = 0, n1180 = 0, n1181 = 0, n1182 = 0, n1183 = 0, n1184 = 0;
reg n1185 = 0, n1186 = 0, n1189 = 0, n1190 = 0, n1191 = 0, n1192 = 0, n1193 = 0, n1194 = 0, n1195 = 0, n1198 = 0;
reg n1199 = 0, n1200 = 0, n1201 = 0, n1202 = 0, n1203 = 0, n1204 = 0, n1206 = 0, n1207 = 0, n1208 = 0, n1209 = 0;
reg n1210 = 0, n1211 = 0, n1212 = 0, n1214 = 0, n1215 = 0, n1216 = 0, n1217 = 0, n1218 = 0, n1219 = 0, n1220 = 0;
reg n1221 = 0, n1223 = 0, n1224 = 0, n1225 = 0, n1226 = 0, n1227 = 0, n1228 = 0, n1229 = 0, n1230 = 0, n1231 = 0;
reg n1232 = 0, n1233 = 0, n1234 = 0, n1235 = 0, n1236 = 0, n1237 = 0, n1238 = 0, n1239 = 0, n1240 = 0, n1241 = 0;
reg n1242 = 0, n1244 = 0, n1247 = 0, n1248 = 0, n1249 = 0, n1250 = 0, n1251 = 0, n1252 = 0, n1253 = 0, n1254 = 0;
reg n1255 = 0, n1256 = 0, n1257 = 0, n1258 = 0, n1259 = 0, n1260 = 0, n1261 = 0, n1262 = 0, n1264 = 0, n1265 = 0;
reg n1266 = 0, n1267 = 0, n1268 = 0, n1269 = 0, n1272 = 0, n1273 = 0, n1278 = 0, n1279 = 0, n1280 = 0, n1281 = 0;
reg n1282 = 0, n1283 = 0, n1284 = 0, n1285 = 0, n1286 = 0, n1287 = 0, n1288 = 0, n1289 = 0, n1290 = 0, n1291 = 0;
reg n1292 = 0, n1293 = 0, n1294 = 0, n1295 = 0, n1296 = 0, n1297 = 0, n1298 = 0, n1299 = 0, n1300 = 0, n1301 = 0;
reg n1302 = 0, n1303 = 0, n1304 = 0, n1305 = 0, n1306 = 0, n1307 = 0, n1308 = 0, n1309 = 0, n1310 = 0, n1311 = 0;
reg n1312 = 0, n1313 = 0, n1314 = 0, n1315 = 0, n1316 = 0, n1317 = 0, n1318 = 0, n1319 = 0, n1320 = 0, n1321 = 0;
reg n1322 = 0, n1323 = 0, n1324 = 0, n1325 = 0, n1326 = 0, n1327 = 0, n1328 = 0, n1329 = 0, n1330 = 0, n1331 = 0;
reg n1332 = 0, n1333 = 0, n1334 = 0, n1341 = 0, n1342 = 0, n1343 = 0, n1344 = 0, n1345 = 0, n1346 = 0, n1348 = 0;
reg n1349 = 0, n1350 = 0, n1351 = 0, n1352 = 0, n1353 = 0, n1354 = 0, n1358 = 0, n1359 = 0, n1360 = 0, n1361 = 0;
reg n1362 = 0, n1363 = 0, n1364 = 0, n1365 = 0, n1367 = 0, n1368 = 0, n1369 = 0, n1370 = 0, n1371 = 0, n1372 = 0;
reg n1373 = 0, n1376 = 0, n1377 = 0, n1378 = 0, n1379 = 0, n1380 = 0, n1381 = 0, n1382 = 0, n1385 = 0, n1386 = 0;
reg n1387 = 0, n1388 = 0, n1389 = 0, n1390 = 0, n1391 = 0, n1392 = 0, n1395 = 0, n1396 = 0, n1397 = 0, n1398 = 0;
reg n1399 = 0, n1400 = 0, n1401 = 0, n1403 = 0, n1404 = 0, n1405 = 0, n1406 = 0, n1407 = 0, n1409 = 0, n1410 = 0;
reg n1411 = 0, n1412 = 0, n1413 = 0, n1414 = 0, n1415 = 0, n1416 = 0, n1417 = 0, n1418 = 0, n1419 = 0, n1420 = 0;
reg n1421 = 0, n1422 = 0, n1423 = 0, n1424 = 0, n1425 = 0, n1426 = 0, n1427 = 0, n1428 = 0, n1429 = 0, n1430 = 0;
reg n1431 = 0, n1432 = 0, n1433 = 0, n1434 = 0, n1435 = 0, n1436 = 0, n1437 = 0, n1438 = 0, n1439 = 0, n1440 = 0;
reg n1441 = 0, n1442 = 0, n1443 = 0, n1444 = 0, n1445 = 0, n1446 = 0, n1447 = 0, n1448 = 0, n1449 = 0, n1450 = 0;
reg n1451 = 0, n1452 = 0, n1453 = 0, n1454 = 0, n1455 = 0, n1456 = 0, n1457 = 0, n1458 = 0, n1459 = 0, n1462 = 0;
reg n1463 = 0, n1464 = 0, n1465 = 0, n1466 = 0, n1467 = 0, n1468 = 0, n1469 = 0, n1470 = 0, n1471 = 0, n1472 = 0;
reg n1473 = 0, n1474 = 0, n1475 = 0, n1476 = 0, n1477 = 0, n1478 = 0, n1479 = 0, n1480 = 0, n1481 = 0, n1482 = 0;
reg n1483 = 0, n1484 = 0, n1485 = 0, n1486 = 0, n1487 = 0, n1488 = 0, n1489 = 0, n1490 = 0, n1492 = 0, n1493 = 0;
reg n1494 = 0, n1495 = 0, n1496 = 0, n1497 = 0, n1498 = 0, n1499 = 0, n1503 = 0, n1504 = 0, n1505 = 0, n1506 = 0;
reg n1507 = 0, n1508 = 0, n1509 = 0, n1513 = 0, n1514 = 0, n1515 = 0, n1516 = 0, n1517 = 0, n1518 = 0, n1519 = 0;
reg n1522 = 0, n1523 = 0, n1524 = 0, n1525 = 0, n1526 = 0, n1527 = 0, n1528 = 0, n1529 = 0, n1530 = 0, n1531 = 0;
reg n1535 = 0, n1536 = 0, n1537 = 0, n1538 = 0, n1539 = 0, n1540 = 0, n1543 = 0, n1544 = 0, n1545 = 0, n1546 = 0;
reg n1547 = 0, n1548 = 0, n1549 = 0, n1550 = 0, n1551 = 0, n1553 = 0, n1554 = 0, n1555 = 0, n1556 = 0, n1558 = 0;
reg n1561 = 0, n1562 = 0, n1563 = 0, n1564 = 0, n1565 = 0, n1566 = 0, n1567 = 0, n1571 = 0, n1572 = 0, n1573 = 0;
reg n1574 = 0, n1575 = 0, n1576 = 0, n1578 = 0, n1579 = 0, n1580 = 0, n1581 = 0, n1582 = 0, n1583 = 0, n1585 = 0;
reg n1586 = 0, n1587 = 0, n1588 = 0, n1589 = 0, n1590 = 0, n1591 = 0, n1593 = 0, n1594 = 0, n1595 = 0, n1596 = 0;
reg n1597 = 0, n1598 = 0, n1599 = 0, n1600 = 0, n1603 = 0, n1604 = 0, n1605 = 0, n1606 = 0, n1607 = 0, n1608 = 0;
reg n1609 = 0, n1610 = 0, n1611 = 0, n1612 = 0, n1613 = 0, n1614 = 0, n1615 = 0, n1616 = 0, n1617 = 0, n1618 = 0;
reg n1619 = 0, n1626 = 0, n1627 = 0, n1628 = 0, n1629 = 0, n1630 = 0, n1631 = 0, n1632 = 0, n1633 = 0, n1634 = 0;
reg n1635 = 0, n1636 = 0, n1637 = 0, n1638 = 0, n1639 = 0, n1640 = 0, n1641 = 0, n1642 = 0, n1643 = 0, n1644 = 0;
reg n1645 = 0, n1646 = 0, n1647 = 0, n1648 = 0, n1649 = 0, n1650 = 0, n1651 = 0, n1652 = 0, n1653 = 0, n1654 = 0;
reg n1655 = 0, n1656 = 0, n1657 = 0, n1658 = 0, n1659 = 0, n1660 = 0, n1661 = 0, n1662 = 0, n1663 = 0, n1664 = 0;
reg n1665 = 0, n1667 = 0, n1668 = 0, n1669 = 0, n1670 = 0, n1676 = 0, n1677 = 0, n1678 = 0, n1679 = 0, n1680 = 0;
reg n1681 = 0, n1682 = 0, n1684 = 0, n1686 = 0, n1687 = 0, n1688 = 0, n1689 = 0, n1690 = 0, n1691 = 0, n1692 = 0;
reg n1693 = 0, n1694 = 0, n1695 = 0, n1701 = 0, n1702 = 0, n1703 = 0, n1704 = 0, n1705 = 0, n1706 = 0, n1707 = 0;
reg n1708 = 0, n1709 = 0, n1711 = 0, n1712 = 0, n1713 = 0, n1714 = 0, n1715 = 0, n1716 = 0, n1717 = 0, n1718 = 0;
reg n1719 = 0, n1720 = 0, n1721 = 0, n1722 = 0, n1725 = 0, n1726 = 0, n1727 = 0, n1728 = 0, n1729 = 0, n1730 = 0;
reg n1731 = 0, n1733 = 0, n1734 = 0, n1735 = 0, n1736 = 0, n1737 = 0, n1738 = 0, n1739 = 0, n1740 = 0, n1745 = 0;
reg n1746 = 0, n1747 = 0, n1748 = 0, n1749 = 0, n1750 = 0, n1751 = 0, n1753 = 0, n1754 = 0, n1755 = 0, n1756 = 0;
reg n1757 = 0, n1758 = 0, n1759 = 0, n1760 = 0, n1762 = 0, n1763 = 0, n1764 = 0, n1765 = 0, n1766 = 0, n1767 = 0;
reg n1768 = 0, n1769 = 0, n1770 = 0, n1772 = 0, n1777 = 0, n1778 = 0, n1779 = 0, n1780 = 0, n1781 = 0, n1782 = 0;
reg n1783 = 0, n1784 = 0, n1785 = 0, n1786 = 0, n1787 = 0, n1788 = 0, n1789 = 0, n1790 = 0, n1793 = 0, n1794 = 0;
reg n1795 = 0, n1796 = 0, n1797 = 0, n1798 = 0, n1799 = 0, n1800 = 0, n1801 = 0, n1802 = 0, n1803 = 0, n1804 = 0;
reg n1805 = 0, n1806 = 0, n1807 = 0, n1808 = 0, n1809 = 0, n1810 = 0, n1811 = 0, n1812 = 0, n1813 = 0, n1814 = 0;
reg n1815 = 0, n1816 = 0, n1817 = 0, n1818 = 0, n1819 = 0, n1820 = 0, n1821 = 0, n1822 = 0, n1823 = 0, n1824 = 0;
reg n1827 = 0, n1828 = 0, n1829 = 0, n1830 = 0, n1831 = 0, n1832 = 0, n1833 = 0, n1834 = 0, n1836 = 0, n1837 = 0;
reg n1838 = 0, n1839 = 0, n1840 = 0, n1841 = 0, n1842 = 0, n1846 = 0, n1847 = 0, n1848 = 0, n1849 = 0, n1850 = 0;
reg n1851 = 0, n1852 = 0, n1853 = 0, n1854 = 0, n1855 = 0, n1856 = 0, n1857 = 0, n1858 = 0, n1859 = 0, n1864 = 0;
reg n1865 = 0, n1866 = 0, n1867 = 0, n1868 = 0, n1869 = 0, n1870 = 0, n1872 = 0, n1875 = 0, n1879 = 0, n1886 = 0;
reg n1888 = 0, n1889 = 0, n1890 = 0, n1891 = 0, n1892 = 0, n1893 = 0, n1894 = 0, n1895 = 0, n1896 = 0, n1897 = 0;
reg n1898 = 0, n1899 = 0, n1900 = 0, n1901 = 0, n1902 = 0, n1903 = 0, n1904 = 0, n1907 = 0, n1908 = 0, n1909 = 0;
reg n1910 = 0, n1911 = 0, n1912 = 0, n1913 = 0, n1915 = 0, n1916 = 0, n1917 = 0, n1918 = 0, n1919 = 0, n1920 = 0;
reg n1921 = 0, n1922 = 0, n1923 = 0, n1924 = 0, n1925 = 0, n1926 = 0, n1927 = 0, n1928 = 0, n1929 = 0, n1930 = 0;
reg n1931 = 0, n1932 = 0, n1934 = 0, n1935 = 0, n1937 = 0, n1938 = 0, n1939 = 0, n1940 = 0, n1941 = 0, n1943 = 0;
reg n1944 = 0, n1945 = 0, n1946 = 0, n1947 = 0, n1948 = 0, n1949 = 0, n1950 = 0, n1955 = 0, n1956 = 0, n1957 = 0;
reg n1958 = 0, n1959 = 0, n1960 = 0, n1961 = 0, n1962 = 0, n1963 = 0, n1964 = 0, n1965 = 0, n1966 = 0, n1967 = 0;
reg n1968 = 0, n1969 = 0, n1970 = 0, n1971 = 0, n1972 = 0, n1973 = 0, n1974 = 0, n1975 = 0, n1976 = 0, n1977 = 0;
reg n1978 = 0, n1979 = 0, n1980 = 0, n1981 = 0, n1983 = 0, n1984 = 0, n1985 = 0, n1986 = 0, n1987 = 0, n1988 = 0;
reg n1989 = 0, n1990 = 0, n1991 = 0, n1992 = 0, n1993 = 0, n1994 = 0, n1995 = 0, n1996 = 0, n1997 = 0, n2001 = 0;
reg n2002 = 0, n2004 = 0, n2005 = 0, n2006 = 0, n2007 = 0, n2008 = 0, n2010 = 0, n2011 = 0, n2012 = 0, n2013 = 0;
reg n2014 = 0, n2015 = 0, n2016 = 0, n2018 = 0, n2019 = 0, n2025 = 0, n2026 = 0, n2027 = 0, n2028 = 0, n2029 = 0;
reg n2030 = 0, n2031 = 0, n2032 = 0, n2033 = 0, n2034 = 0, n2035 = 0, n2038 = 0, n2039 = 0, n2040 = 0, n2041 = 0;
reg n2042 = 0, n2043 = 0, n2044 = 0, n2046 = 0, n2047 = 0, n2048 = 0, n2049 = 0, n2050 = 0, n2051 = 0, n2052 = 0;
reg n2053 = 0, n2059 = 0, n2060 = 0, n2061 = 0, n2062 = 0, n2063 = 0, n2064 = 0, n2065 = 0, n2066 = 0, n2067 = 0;
reg n2068 = 0, n2069 = 0, n2070 = 0, n2071 = 0, n2072 = 0, n2073 = 0, n2075 = 0, n2077 = 0, n2078 = 0, n2079 = 0;
reg n2080 = 0, n2081 = 0, n2082 = 0, n2083 = 0, n2084 = 0, n2086 = 0, n2087 = 0, n2088 = 0, n2089 = 0, n2090 = 0;
reg n2091 = 0, n2092 = 0, n2093 = 0, n2095 = 0, n2096 = 0, n2097 = 0, n2098 = 0, n2099 = 0, n2100 = 0, n2101 = 0;
reg n2102 = 0, n2103 = 0, n2104 = 0, n2105 = 0, n2106 = 0, n2107 = 0, n2108 = 0, n2114 = 0, n2115 = 0, n2116 = 0;
reg n2117 = 0, n2118 = 0, n2119 = 0, n2120 = 0, n2121 = 0, n2122 = 0, n2124 = 0, n2125 = 0, n2126 = 0, n2127 = 0;
reg n2128 = 0, n2129 = 0, n2130 = 0, n2131 = 0, n2132 = 0, n2133 = 0, n2134 = 0, n2135 = 0, n2136 = 0, n2137 = 0;
reg n2138 = 0, n2139 = 0, n2140 = 0, n2141 = 0, n2142 = 0, n2143 = 0, n2144 = 0, n2145 = 0, n2146 = 0, n2147 = 0;
reg n2148 = 0, n2149 = 0, n2150 = 0, n2151 = 0, n2152 = 0, n2153 = 0, n2154 = 0, n2155 = 0, n2156 = 0, n2157 = 0;
reg n2158 = 0, n2159 = 0, n2160 = 0, n2161 = 0, n2162 = 0, n2163 = 0, n2165 = 0, n2166 = 0, n2167 = 0, n2168 = 0;
reg n2169 = 0, n2170 = 0, n2171 = 0, n2172 = 0, n2173 = 0, n2176 = 0, n2177 = 0, n2178 = 0, n2179 = 0, n2180 = 0;
reg n2181 = 0, n2182 = 0, n2183 = 0, n2185 = 0, n2186 = 0, n2187 = 0, n2188 = 0, n2189 = 0, n2190 = 0, n2191 = 0;
reg n2192 = 0, n2193 = 0, n2194 = 0, n2197 = 0, n2198 = 0, n2199 = 0, n2200 = 0, n2201 = 0, n2202 = 0, n2203 = 0;
reg n2204 = 0, n2205 = 0, n2211 = 0, n2212 = 0, n2213 = 0, n2214 = 0, n2215 = 0, n2216 = 0, n2217 = 0, n2218 = 0;
reg n2219 = 0, n2220 = 0, n2221 = 0, n2222 = 0, n2223 = 0, n2224 = 0, n2225 = 0, n2226 = 0, n2227 = 0, n2228 = 0;
reg n2231 = 0, n2232 = 0, n2233 = 0, n2234 = 0, n2235 = 0, n2236 = 0, n2237 = 0, n2238 = 0, n2239 = 0, n2243 = 0;
reg n2244 = 0, n2245 = 0, n2246 = 0, n2248 = 0, n2249 = 0, n2250 = 0, n2251 = 0, n2252 = 0, n2253 = 0, n2254 = 0;
reg n2255 = 0, n2256 = 0, n2261 = 0, n2262 = 0, n2263 = 0, n2264 = 0, n2265 = 0, n2266 = 0, n2267 = 0, n2268 = 0;
reg n2269 = 0, n2273 = 0, n2274 = 0, n2275 = 0, n2276 = 0, n2277 = 0, n2278 = 0, n2279 = 0, n2280 = 0, n2281 = 0;
reg n2285 = 0, n2286 = 0, n2287 = 0, n2288 = 0, n2289 = 0, n2290 = 0, n2291 = 0, n2292 = 0, n2293 = 0, n2295 = 0;
reg n2296 = 0, n2297 = 0, n2298 = 0, n2299 = 0, n2300 = 0, n2301 = 0, n2302 = 0, n2305 = 0, n2309 = 0, n2310 = 0;
reg n2311 = 0, n2312 = 0, n2313 = 0, n2314 = 0, n2315 = 0, n2316 = 0, n2317 = 0, n2318 = 0, n2319 = 0, n2320 = 0;
reg n2321 = 0, n2326 = 0, n2327 = 0, n2328 = 0, n2329 = 0, n2330 = 0, n2331 = 0, n2332 = 0, n2333 = 0, n2334 = 0;
reg n2335 = 0, n2336 = 0, n2337 = 0, n2338 = 0, n2339 = 0, n2340 = 0, n2341 = 0, n2342 = 0, n2343 = 0, n2344 = 0;
reg n2345 = 0, n2346 = 0, n2349 = 0, n2350 = 0, n2351 = 0, n2352 = 0, n2353 = 0, n2354 = 0, n2355 = 0, n2356 = 0;
reg n2357 = 0, n2359 = 0, n2360 = 0, n2361 = 0, n2362 = 0, n2363 = 0, n2364 = 0, n2365 = 0, n2366 = 0, n2367 = 0;
reg n2368 = 0, n2369 = 0, n2370 = 0, n2371 = 0, n2372 = 0, n2373 = 0, n2374 = 0, n2375 = 0, n2376 = 0, n2377 = 0;
reg n2378 = 0, n2379 = 0, n2380 = 0, n2381 = 0, n2382 = 0, n2383 = 0, n2385 = 0, n2386 = 0, n2387 = 0, n2388 = 0;
reg n2389 = 0, n2390 = 0, n2391 = 0, n2392 = 0, n2393 = 0, n2394 = 0, n2395 = 0, n2396 = 0, n2397 = 0, n2398 = 0;
reg n2399 = 0, n2400 = 0, n2402 = 0, n2403 = 0, n2404 = 0, n2405 = 0, n2406 = 0, n2407 = 0, n2408 = 0, n2409 = 0;
reg n2410 = 0, n2411 = 0, n2412 = 0, n2413 = 0, n2414 = 0, n2415 = 0, n2416 = 0, n2417 = 0, n2418 = 0, n2419 = 0;
reg n2420 = 0, n2421 = 0, n2422 = 0, n2423 = 0, n2425 = 0, n2426 = 0, n2427 = 0, n2428 = 0, n2429 = 0, n2430 = 0;
reg n2431 = 0, n2432 = 0, n2433 = 0, n2435 = 0, n2436 = 0, n2437 = 0, n2438 = 0, n2439 = 0, n2440 = 0, n2441 = 0;
reg n2442 = 0, n2443 = 0, n2444 = 0, n2445 = 0, n2446 = 0, n2447 = 0, n2448 = 0, n2449 = 0, n2450 = 0, n2452 = 0;
reg n2453 = 0, n2454 = 0, n2455 = 0, n2456 = 0, n2457 = 0, n2458 = 0, n2459 = 0, n2461 = 0, n2462 = 0, n2463 = 0;
reg n2464 = 0, n2465 = 0, n2466 = 0, n2467 = 0, n2468 = 0, n2471 = 0, n2472 = 0, n2473 = 0, n2474 = 0, n2475 = 0;
reg n2476 = 0, n2477 = 0, n2478 = 0, n2479 = 0, n2480 = 0, n2481 = 0, n2482 = 0, n2483 = 0, n2484 = 0, n2485 = 0;
reg n2486 = 0, n2487 = 0, n2488 = 0, n2489 = 0, n2490 = 0, n2491 = 0, n2492 = 0, n2494 = 0, n2497 = 0, n2498 = 0;
reg n2499 = 0, n2500 = 0, n2501 = 0, n2502 = 0, n2503 = 0, n2504 = 0, n2506 = 0, n2507 = 0, n2508 = 0, n2509 = 0;
reg n2510 = 0, n2512 = 0, n2513 = 0, n2514 = 0, n2515 = 0, n2516 = 0, n2517 = 0, n2518 = 0, n2521 = 0, n2525 = 0;
reg n2526 = 0, n2527 = 0, n2528 = 0, n2529 = 0, n2530 = 0, n2531 = 0, n2532 = 0, n2533 = 0, n2537 = 0, n2539 = 0;
reg n2541 = 0, n2542 = 0, n2543 = 0, n2544 = 0, n2545 = 0, n2546 = 0, n2547 = 0, n2548 = 0, n2549 = 0, n2550 = 0;
reg n2552 = 0, n2554 = 0, n2555 = 0, n2556 = 0, n2557 = 0, n2558 = 0, n2559 = 0, n2560 = 0, n2561 = 0, n2563 = 0;
reg n2565 = 0, n2566 = 0, n2567 = 0, n2568 = 0, n2569 = 0, n2570 = 0, n2571 = 0, n2572 = 0, n2576 = 0, n2577 = 0;
reg n2578 = 0, n2579 = 0, n2580 = 0, n2581 = 0, n2582 = 0, n2583 = 0, n2584 = 0, n2585 = 0, n2586 = 0, n2587 = 0;
reg n2588 = 0, n2589 = 0, n2594 = 0, n2595 = 0, n2596 = 0, n2597 = 0, n2598 = 0, n2599 = 0, n2600 = 0, n2601 = 0;
reg n2603 = 0, n2604 = 0, n2605 = 0, n2606 = 0, n2607 = 0, n2608 = 0, n2609 = 0, n2610 = 0, n2611 = 0, n2616 = 0;
reg n2617 = 0, n2618 = 0, n2619 = 0, n2620 = 0, n2621 = 0, n2622 = 0, n2623 = 0, n2624 = 0, n2625 = 0, n2626 = 0;
reg n2627 = 0, n2630 = 0, n2631 = 0, n2632 = 0, n2633 = 0, n2634 = 0, n2635 = 0, n2636 = 0, n2637 = 0, n2638 = 0;
reg n2639 = 0, n2640 = 0, n2641 = 0, n2642 = 0, n2643 = 0, n2644 = 0, n2645 = 0, n2646 = 0, n2647 = 0, n2648 = 0;
reg n2653 = 0, n2654 = 0, n2655 = 0, n2656 = 0, n2657 = 0, n2658 = 0, n2659 = 0, n2660 = 0, n2661 = 0, n2662 = 0;
reg n2663 = 0, n2664 = 0, n2665 = 0, n2666 = 0, n2667 = 0, n2668 = 0, n2669 = 0, n2672 = 0, n2673 = 0, n2674 = 0;
reg n2675 = 0, n2676 = 0, n2681 = 0, n2683 = 0, n2684 = 0, n2685 = 0, n2686 = 0, n2687 = 0, n2688 = 0, n2689 = 0;
reg n2690 = 0, n2691 = 0, n2692 = 0, n2693 = 0, n2694 = 0, n2695 = 0, n2698 = 0, n2699 = 0, n2700 = 0, n2701 = 0;
reg n2702 = 0, n2703 = 0, n2704 = 0, n2705 = 0, n2706 = 0, n2709 = 0, n2710 = 0, n2711 = 0, n2712 = 0, n2713 = 0;
reg n2714 = 0, n2716 = 0, n2717 = 0, n2718 = 0, n2719 = 0, n2720 = 0, n2721 = 0, n2722 = 0, n2723 = 0, n2724 = 0;
reg n2729 = 0, n2732 = 0, n2733 = 0, n2734 = 0, n2735 = 0, n2736 = 0, n2737 = 0, n2738 = 0, n2739 = 0, n2740 = 0;
reg n2741 = 0, n2742 = 0, n2743 = 0, n2744 = 0, n2745 = 0, n2746 = 0, n2747 = 0, n2749 = 0, n2750 = 0, n2751 = 0;
reg n2752 = 0, n2753 = 0, n2754 = 0, n2755 = 0, n2756 = 0, n2758 = 0, n2759 = 0, n2761 = 0, n2762 = 0, n2763 = 0;
reg n2764 = 0, n2765 = 0, n2766 = 0, n2767 = 0, n2768 = 0, n2769 = 0, n2770 = 0, n2771 = 0, n2772 = 0, n2773 = 0;
reg n2774 = 0, n2776 = 0, n2777 = 0, n2778 = 0, n2779 = 0, n2780 = 0, n2781 = 0, n2782 = 0, n2783 = 0, n2784 = 0;
reg n2788 = 0, n2789 = 0, n2790 = 0, n2791 = 0, n2792 = 0, n2793 = 0, n2794 = 0, n2795 = 0, n2796 = 0, n2797 = 0;
reg n2798 = 0, n2799 = 0, n2800 = 0, n2801 = 0, n2802 = 0, n2803 = 0, n2804 = 0, n2805 = 0, n2806 = 0, n2807 = 0;
reg n2808 = 0, n2809 = 0, n2810 = 0, n2811 = 0, n2814 = 0, n2815 = 0, n2816 = 0, n2817 = 0, n2818 = 0, n2819 = 0;
reg n2820 = 0, n2821 = 0, n2822 = 0, n2823 = 0, n2824 = 0, n2825 = 0, n2826 = 0, n2827 = 0, n2828 = 0, n2830 = 0;
reg n2832 = 0, n2833 = 0, n2834 = 0, n2835 = 0, n2836 = 0, n2837 = 0, n2838 = 0, n2839 = 0, n2840 = 0, n2842 = 0;
reg n2843 = 0, n2845 = 0, n2846 = 0, n2847 = 0, n2848 = 0, n2849 = 0, n2850 = 0, n2851 = 0, n2857 = 0, n2858 = 0;
reg n2860 = 0, n2861 = 0, n2862 = 0, n2863 = 0, n2864 = 0, n2867 = 0, n2868 = 0, n2869 = 0, n2870 = 0, n2871 = 0;
reg n2872 = 0, n2873 = 0, n2874 = 0, n2875 = 0, n2876 = 0, n2877 = 0, n2878 = 0, n2879 = 0, n2880 = 0, n2882 = 0;
reg n2883 = 0, n2884 = 0, n2885 = 0, n2887 = 0, n2888 = 0, n2889 = 0, n2890 = 0, n2891 = 0, n2892 = 0, n2893 = 0;
reg n2894 = 0, n2895 = 0, n2898 = 0, n2899 = 0, n2900 = 0, n2901 = 0, n2902 = 0, n2903 = 0, n2904 = 0, n2905 = 0;
reg n2906 = 0, n2907 = 0, n2908 = 0, n2909 = 0, n2911 = 0, n2912 = 0, n2913 = 0, n2914 = 0, n2915 = 0, n2916 = 0;
reg n2917 = 0, n2918 = 0, n2919 = 0, n2920 = 0, n2921 = 0, n2922 = 0, n2923 = 0, n2924 = 0, n2925 = 0, n2926 = 0;
reg n2927 = 0, n2928 = 0, n2929 = 0, n2930 = 0, n2931 = 0, n2932 = 0, n2933 = 0, n2934 = 0, n2935 = 0, n2936 = 0;
reg n2937 = 0, n2938 = 0, n2939 = 0, n2940 = 0, n2941 = 0, n2942 = 0, n2943 = 0, n2944 = 0, n2945 = 0, n2946 = 0;
reg n2947 = 0, n2948 = 0, n2949 = 0, n2950 = 0, n2951 = 0, n2954 = 0, n2955 = 0, n2956 = 0, n2957 = 0, n2958 = 0;
reg n2959 = 0, n2960 = 0, n2962 = 0, n2963 = 0, n2964 = 0, n2965 = 0, n2966 = 0, n2967 = 0, n2968 = 0, n2969 = 0;
reg n2972 = 0, n2973 = 0, n2974 = 0, n2975 = 0, n2976 = 0, n2977 = 0, n2978 = 0, n2979 = 0, n2980 = 0, n2981 = 0;
reg n2982 = 0, n2983 = 0, n2984 = 0, n2985 = 0, n2986 = 0, n2990 = 0, n2991 = 0, n2992 = 0, n2993 = 0, n2994 = 0;
reg n2995 = 0, n2996 = 0, n2997 = 0, n2998 = 0, n2999 = 0, n3000 = 0, n3001 = 0, n3002 = 0, n3003 = 0, n3004 = 0;
reg n3005 = 0, n3010 = 0, n3011 = 0, n3012 = 0, n3013 = 0, n3014 = 0, n3015 = 0, n3016 = 0, n3017 = 0, n3018 = 0;
reg n3019 = 0, n3020 = 0, n3021 = 0, n3022 = 0, n3023 = 0, n3024 = 0, n3025 = 0, n3026 = 0, n3027 = 0, n3028 = 0;
reg n3035 = 0, n3036 = 0, n3037 = 0, n3038 = 0, n3039 = 0, n3040 = 0, n3041 = 0, n3042 = 0, n3043 = 0, n3044 = 0;
reg n3046 = 0, n3047 = 0, n3048 = 0, n3049 = 0, n3050 = 0, n3051 = 0, n3052 = 0, n3053 = 0, n3054 = 0, n3055 = 0;
reg n3056 = 0, n3057 = 0, n3058 = 0, n3059 = 0, n3060 = 0, n3061 = 0, n3062 = 0, n3063 = 0, n3064 = 0, n3066 = 0;
reg n3070 = 0, n3071 = 0, n3072 = 0, n3073 = 0, n3074 = 0, n3075 = 0, n3076 = 0, n3077 = 0, n3078 = 0, n3079 = 0;
reg n3080 = 0, n3081 = 0, n3082 = 0, n3083 = 0, n3084 = 0, n3085 = 0, n3086 = 0, n3088 = 0, n3089 = 0, n3090 = 0;
reg n3091 = 0, n3092 = 0, n3093 = 0, n3094 = 0, n3095 = 0, n3096 = 0, n3097 = 0, n3098 = 0, n3099 = 0, n3100 = 0;
reg n3101 = 0, n3102 = 0, n3103 = 0, n3105 = 0, n3106 = 0, n3107 = 0, n3108 = 0, n3109 = 0, n3110 = 0, n3111 = 0;
reg n3115 = 0, n3116 = 0, n3117 = 0, n3118 = 0, n3119 = 0, n3120 = 0, n3121 = 0, n3122 = 0, n3123 = 0, n3125 = 0;
reg n3126 = 0, n3127 = 0, n3128 = 0, n3129 = 0, n3130 = 0, n3131 = 0, n3132 = 0, n3133 = 0, n3134 = 0, n3135 = 0;
reg n3136 = 0, n3137 = 0, n3138 = 0, n3139 = 0, n3140 = 0, n3143 = 0, n3144 = 0, n3145 = 0, n3146 = 0, n3147 = 0;
reg n3148 = 0, n3149 = 0, n3151 = 0, n3152 = 0, n3153 = 0, n3154 = 0, n3155 = 0, n3156 = 0, n3157 = 0, n3159 = 0;
reg n3160 = 0, n3161 = 0, n3162 = 0, n3163 = 0, n3164 = 0, n3165 = 0, n3166 = 0, n3167 = 0, n3168 = 0, n3169 = 0;
reg n3170 = 0, n3171 = 0, n3172 = 0, n3173 = 0, n3174 = 0, n3176 = 0, n3177 = 0, n3178 = 0, n3179 = 0, n3180 = 0;
reg n3181 = 0, n3182 = 0, n3183 = 0, n3184 = 0, n3185 = 0, n3186 = 0, n3187 = 0, n3188 = 0, n3189 = 0, n3190 = 0;
reg n3191 = 0, n3192 = 0, n3193 = 0, n3194 = 0, n3195 = 0, n3196 = 0, n3197 = 0, n3200 = 0, n3201 = 0, n3202 = 0;
reg n3203 = 0, n3204 = 0, n3205 = 0, n3206 = 0, n3208 = 0, n3209 = 0, n3210 = 0, n3211 = 0, n3212 = 0, n3213 = 0;
reg n3214 = 0, n3215 = 0, n3217 = 0, n3218 = 0, n3219 = 0, n3220 = 0, n3221 = 0, n3222 = 0, n3223 = 0, n3224 = 0;
reg n3225 = 0, n3226 = 0, n3227 = 0, n3228 = 0, n3229 = 0, n3230 = 0, n3232 = 0, n3234 = 0, n3235 = 0, n3236 = 0;
reg n3237 = 0, n3238 = 0, n3239 = 0, n3240 = 0, n3241 = 0, n3242 = 0, n3243 = 0, n3244 = 0, n3245 = 0, n3246 = 0;
reg n3247 = 0, n3248 = 0, n3250 = 0, n3251 = 0, n3252 = 0, n3253 = 0, n3254 = 0, n3255 = 0, n3256 = 0, n3257 = 0;
reg n3263 = 0, n3264 = 0, n3265 = 0, n3266 = 0, n3267 = 0, n3268 = 0, n3269 = 0, n3270 = 0, n3271 = 0, n3272 = 0;
reg n3273 = 0, n3274 = 0, n3275 = 0, n3276 = 0, n3277 = 0, n3278 = 0, n3279 = 0, n3280 = 0, n3281 = 0, n3282 = 0;
reg n3283 = 0, n3284 = 0, n3285 = 0, n3286 = 0, n3287 = 0, n3288 = 0, n3289 = 0, n3290 = 0, n3291 = 0, n3292 = 0;
reg n3293 = 0, n3294 = 0, n3296 = 0, n3297 = 0, n3298 = 0, n3299 = 0, n3300 = 0, n3301 = 0, n3302 = 0, n3303 = 0;
reg n3305 = 0, n3306 = 0, n3307 = 0, n3308 = 0, n3309 = 0, n3310 = 0, n3311 = 0, n3312 = 0, n3313 = 0, n3314 = 0;
reg n3315 = 0, n3316 = 0, n3317 = 0, n3319 = 0, n3320 = 0, n3321 = 0, n3322 = 0, n3323 = 0, n3324 = 0, n3325 = 0;
reg n3326 = 0, n3327 = 0, n3328 = 0, n3332 = 0, n3333 = 0, n3334 = 0, n3335 = 0, n3336 = 0, n3337 = 0, n3338 = 0;
reg n3339 = 0, n3340 = 0, n3341 = 0, n3342 = 0, n3343 = 0, n3344 = 0, n3345 = 0, n3346 = 0, n3347 = 0, n3348 = 0;
reg n3353 = 0, n3354 = 0, n3355 = 0, n3356 = 0, n3357 = 0, n3358 = 0, n3359 = 0, n3360 = 0, n3361 = 0, n3362 = 0;
reg n3363 = 0, n3364 = 0, n3365 = 0, n3366 = 0, n3367 = 0, n3369 = 0, n3370 = 0, n3371 = 0, n3372 = 0, n3373 = 0;
reg n3374 = 0, n3375 = 0, n3377 = 0, n3378 = 0, n3379 = 0, n3380 = 0, n3381 = 0, n3382 = 0, n3383 = 0, n3384 = 0;
reg n3385 = 0, n3386 = 0, n3387 = 0, n3388 = 0, n3389 = 0, n3390 = 0, n3391 = 0, n3394 = 0, n3395 = 0, n3396 = 0;
reg n3397 = 0, n3398 = 0, n3399 = 0, n3400 = 0, n3401 = 0, n3402 = 0, n3403 = 0, n3404 = 0, n3405 = 0, n3406 = 0;
reg n3407 = 0, n3408 = 0, n3410 = 0, n3412 = 0, n3413 = 0, n3414 = 0, n3415 = 0, n3416 = 0, n3417 = 0, n3418 = 0;
reg n3419 = 0, n3420 = 0, n3423 = 0, n3425 = 0, n3426 = 0, n3427 = 0, n3428 = 0, n3429 = 0, n3430 = 0, n3431 = 0;
reg n3433 = 0, n3434 = 0, n3435 = 0, n3436 = 0, n3437 = 0, n3438 = 0, n3439 = 0, n3440 = 0, n3441 = 0, n3442 = 0;
reg n3443 = 0, n3444 = 0, n3445 = 0, n3446 = 0, n3447 = 0, n3448 = 0, n3449 = 0, n3450 = 0, n3451 = 0, n3452 = 0;
reg n3453 = 0, n3454 = 0, n3455 = 0, n3456 = 0, n3461 = 0, n3463 = 0, n3472 = 0, n3473 = 0, n3474 = 0, n3475 = 0;
reg n3476 = 0, n3477 = 0, n3478 = 0, n3479 = 0, n3480 = 0, n3481 = 0, n3482 = 0, n3483 = 0, n3484 = 0, n3485 = 0;
reg n3486 = 0, n3487 = 0, n3490 = 0, n3491 = 0, n3492 = 0, n3493 = 0, n3494 = 0, n3495 = 0, n3496 = 0, n3497 = 0;
reg n3498 = 0, n3499 = 0, n3500 = 0, n3501 = 0, n3502 = 0, n3503 = 0, n3504 = 0, n3505 = 0, n3506 = 0, n3507 = 0;
reg n3508 = 0, n3509 = 0, n3510 = 0, n3511 = 0, n3512 = 0, n3513 = 0, n3514 = 0, n3515 = 0, n3516 = 0, n3517 = 0;
reg n3518 = 0, n3519 = 0, n3520 = 0, n3521 = 0, n3522 = 0, n3523 = 0, n3524 = 0, n3528 = 0, n3529 = 0, n3530 = 0;
reg n3531 = 0, n3532 = 0, n3533 = 0, n3534 = 0, n3535 = 0, n3536 = 0, n3537 = 0, n3538 = 0, n3539 = 0, n3540 = 0;
reg n3541 = 0, n3542 = 0, n3543 = 0, n3544 = 0, n3545 = 0, n3546 = 0, n3547 = 0, n3548 = 0, n3549 = 0, n3550 = 0;
reg n3551 = 0, n3552 = 0, n3556 = 0, n3557 = 0, n3558 = 0, n3559 = 0, n3560 = 0, n3561 = 0, n3562 = 0, n3563 = 0;
reg n3564 = 0, n3565 = 0, n3566 = 0, n3567 = 0, n3568 = 0, n3569 = 0, n3570 = 0, n3571 = 0, n3572 = 0, n3573 = 0;
reg n3574 = 0, n3575 = 0, n3576 = 0, n3577 = 0, n3578 = 0, n3579 = 0, n3580 = 0, n3581 = 0, n3582 = 0, n3583 = 0;
reg n3585 = 0, n3586 = 0, n3587 = 0, n3588 = 0, n3589 = 0, n3590 = 0, n3591 = 0, n3592 = 0, n3595 = 0, n3596 = 0;
reg n3597 = 0, n3598 = 0, n3599 = 0, n3600 = 0, n3601 = 0, n3602 = 0, n3606 = 0, n3607 = 0, n3608 = 0, n3609 = 0;
reg n3610 = 0, n3611 = 0, n3612 = 0, n3613 = 0, n3614 = 0, n3615 = 0, n3616 = 0, n3617 = 0, n3618 = 0, n3619 = 0;
reg n3622 = 0, n3623 = 0, n3624 = 0, n3625 = 0, n3626 = 0, n3627 = 0, n3628 = 0, n3629 = 0, n3630 = 0, n3631 = 0;
reg n3632 = 0, n3633 = 0, n3634 = 0, n3635 = 0, n3636 = 0, n3637 = 0, n3638 = 0, n3641 = 0, n3642 = 0, n3643 = 0;
reg n3644 = 0, n3645 = 0, n3646 = 0, n3647 = 0, n3648 = 0, n3649 = 0, n3650 = 0, n3651 = 0, n3652 = 0, n3653 = 0;
reg n3654 = 0, n3655 = 0, n3656 = 0, n3657 = 0, n3658 = 0, n3659 = 0, n3660 = 0, n3661 = 0, n3662 = 0, n3663 = 0;
reg n3667 = 0, n3668 = 0, n3669 = 0, n3670 = 0, n3671 = 0, n3672 = 0, n3673 = 0, n3674 = 0, n3675 = 0, n3676 = 0;
reg n3677 = 0, n3678 = 0, n3679 = 0, n3680 = 0, n3681 = 0, n3682 = 0, n3687 = 0, n3688 = 0, n3689 = 0, n3690 = 0;
reg n3691 = 0, n3692 = 0, n3693 = 0, n3694 = 0, n3695 = 0, n3696 = 0, n3697 = 0, n3698 = 0, n3699 = 0, n3700 = 0;
reg n3701 = 0, n3702 = 0, n3705 = 0, n3706 = 0, n3707 = 0, n3708 = 0, n3709 = 0, n3710 = 0, n3711 = 0, n3712 = 0;
reg n3713 = 0, n3714 = 0, n3715 = 0, n3716 = 0, n3717 = 0, n3719 = 0, n3720 = 0, n3721 = 0, n3722 = 0, n3723 = 0;
reg n3724 = 0, n3725 = 0, n3726 = 0, n3727 = 0, n3728 = 0, n3729 = 0, n3730 = 0, n3731 = 0, n3732 = 0, n3734 = 0;
reg n3735 = 0, n3736 = 0, n3737 = 0, n3738 = 0, n3739 = 0, n3740 = 0, n3741 = 0, n3742 = 0, n3743 = 0, n3744 = 0;
reg n3745 = 0, n3746 = 0, n3747 = 0, n3748 = 0, n3753 = 0, n3754 = 0, n3755 = 0, n3756 = 0, n3757 = 0, n3758 = 0;
reg n3759 = 0, n3760 = 0, n3761 = 0, n3762 = 0, n3763 = 0, n3764 = 0, n3766 = 0, n3767 = 0, n3768 = 0, n3769 = 0;
reg n3770 = 0, n3771 = 0, n3772 = 0, n3773 = 0, n3774 = 0, n3775 = 0, n3776 = 0, n3777 = 0, n3778 = 0, n3779 = 0;
reg n3780 = 0, n3781 = 0, n3782 = 0, n3783 = 0, n3791 = 0, n3792 = 0, n3793 = 0, n3794 = 0, n3795 = 0, n3796 = 0;
reg n3797 = 0, n3798 = 0, n3799 = 0, n3800 = 0, n3801 = 0, n3802 = 0, n3803 = 0, n3804 = 0, n3805 = 0, n3806 = 0;
reg n3807 = 0, n3808 = 0, n3809 = 0, n3810 = 0, n3811 = 0, n3812 = 0, n3813 = 0, n3818 = 0, n3819 = 0, n3820 = 0;
reg n3821 = 0, n3822 = 0, n3823 = 0, n3824 = 0, n3829 = 0, n3830 = 0, n3831 = 0, n3832 = 0, n3833 = 0, n3834 = 0;
reg n3835 = 0, n3836 = 0, n3837 = 0, n3838 = 0, n3839 = 0, n3840 = 0, n3841 = 0, n3842 = 0, n3843 = 0, n3844 = 0;
reg n3845 = 0, n3846 = 0, n3847 = 0, n3849 = 0, n3850 = 0, n3851 = 0, n3852 = 0, n3853 = 0, n3854 = 0, n3855 = 0;
reg n3856 = 0, n3857 = 0, n3858 = 0, n3859 = 0, n3860 = 0, n3861 = 0, n3862 = 0, n3863 = 0, n3864 = 0, n3865 = 0;
reg n3866 = 0, n3867 = 0, n3868 = 0, n3869 = 0, n3870 = 0, n3871 = 0, n3872 = 0, n3873 = 0, n3874 = 0, n3875 = 0;
reg n3877 = 0, n3878 = 0, n3879 = 0, n3880 = 0, n3881 = 0, n3882 = 0, n3883 = 0, n3885 = 0, n3886 = 0, n3887 = 0;
reg n3888 = 0, n3889 = 0, n3890 = 0, n3891 = 0, n3893 = 0, n3894 = 0, n3895 = 0, n3896 = 0, n3897 = 0, n3898 = 0;
reg n3899 = 0, n3900 = 0;

assign n3911 = /* LUT   24 20  4 */ n3415;
assign n3912 = /* LUT   16 16  2 */ n1956;
assign n3913 = /* LUT   22 12  4 */ n3039;
assign n3914 = /* LUT   10 22  7 */ (n696 ? (n114 ? (n551 ? n769 : 1'b0) : 1'b0) : 1'b0);
assign n3915 = /* LUT   21 28  2 */ n2980;
assign n3916 = /* LUT    4 22  7 */ (n120 ? (\rco[132]  ? n225 : 1'b0) : 1'b0);
assign n3917 = /* LUT   13 27  1 */ n1553;
assign n3918 = /* LUT   27 10  0 */ (n3646 ? (\rco[66]  ? (n3619 ? n3525 : 1'b0) : 1'b0) : 1'b0);
assign n3919 = /* LUT   15 13  0 */ n1782;
assign n3920 = /* LUT   20 20  3 */ n2763;
assign n3921 = /* LUT   23 18  4 */ n3245;
assign n3922 = /* LUT    5 12  5 */ n488;
assign n3923 = /* LUT   19 27  6 */ n2621;
assign n3924 = /* LUT   11 23  0 */ n1219;
assign n3925 = /* LUT   23 25  5 */ n3308;
assign n3926 = /* LUT   16 19  4 */ n1972;
assign n3927 = /* LUT    1 10  5 */ n42;
assign n3928 = /* LUT   10 21  3 */ n1060;
assign n3929 = /* LUT   15 19  1 */ n1817;
assign n3930 = /* LUT   20 26  4 */ n2808;
assign n3931 = /* LUT    3 20  3 */ n344;
assign n3932 = /* LUT    2 20  7 */ n234;
assign n3933 = /* LUT    6 14  6 */ n622;
assign n3934 = /* LUT   20 23  7 */ (n2785 ? 1'b0 : n1876);
assign n3935 = /* LUT   12 27  5 */ (\rco[99]  ? (n1543 ? \rco[0]  : 1'b0) : 1'b0);
assign n3936 = /* LUT   17 20  6 */ n1975;
assign n3937 = /* LUT   11  8  6 */ n1129;
assign n3938 = /* LUT   29  5  4 */ n3821;
assign n3939 = /* LUT   23 15  1 */ n3222;
assign n3940 = /* LUT   24 16  1 */ n3384;
assign n3941 = /* LUT   27 22  2 */ n3696;
assign n3942 = /* LUT    3 15  5 */ n297;
assign n3943 = /* LUT   18  3  1 */ (\rco[83]  ? n614 : 1'b0);
assign n3944 = /* LUT   21 11  0 */ (n2680 ? (\rco[0]  ? (n2416 ? \rco[48]  : 1'b0) : 1'b0) : 1'b0);
assign n3945 = /* LUT    7 16  7 */ n637;
assign n3946 = /* LUT    9 21  7 */ n920;
assign n3666 = /* LUT   26 18  3 */ (n2552 ? (n3665 ? (n2112 ? n2533 : 1'b0) : 1'b0) : 1'b0);
assign n3947 = /* LUT   12 22  5 */ n1352;
assign n3948 = /* LUT   26 15  4 */ n3543;
assign n3949 = /* LUT   17  9  0 */ (n2270 ? (\rco[23]  ? (n2269 ? n1933 : 1'b0) : 1'b0) : 1'b0);
assign n3950 = /* LUT   19 23  3 */ (n1340 ? (n2786 ? 1'b0 : (n912 ? !n2593 : 1'b0)) : 1'b0);
assign n3951 = /* LUT   28 20  5 */ (n3432 ? \rco[162]  : 1'b0);
assign n3952 = /* LUT   22 15  5 */ n3062;
assign n3953 = /* LUT    4 21  6 */ n453;
assign n3954 = /* LUT   13 28  0 */ n1566;
assign n3955 = /* LUT   27 11  3 */ n3625;
assign n3956 = /* LUT   20 11  2 */ (\rco[48]  ? (n2866 ? (\rco[0]  ? n2680 : 1'b0) : 1'b0) : 1'b0);
assign n3957 = /* LUT    6 10  3 */ n593;
assign n3958 = /* LUT   23 19  7 */ n3256;
assign n3959 = /* LUT    5 13  6 */ n497;
assign n3960 = /* LUT   19 24  7 */ n2795;
assign n3961 = /* LUT   11 20  1 */ n1189;
assign n3962 = /* LUT   29  9  1 */ (n3604 ? \rco[74]  : 1'b0);
assign n3963 = /* LUT   17 27  4 */ n2191;
assign n3964 = /* LUT   28 23  1 */ n3809;
assign n3965 = /* LUT    5 18  4 */ n534;
assign n3966 = /* LUT   19  5  3 */ n2437;
assign n3967 = /* LUT   10 20  0 */ n1053;
assign n3968 = /* LUT   15 16  0 */ n758;
assign n3069 = /* LUT   21 15  5 */ (n2470 ? (n3068 ? 1'b0 : (n2306 ? n2308 : 1'b0)) : 1'b0);
assign n3970 = /* LUT   20 25  5 */ n2802;
assign n3971 = /* LUT    3 21  4 */ (\rco[110]  ? (n460 ? (n363 ? n351 : 1'b0) : 1'b0) : 1'b0);
assign n3972 = /* LUT    6  9  7 */ (n717 ? (n590 ? en_in : 1'b0) : 1'b0);
assign n3973 = /* LUT   20 22  4 */ n2779;
assign n3974 = /* LUT   12 26  6 */ n1392;
assign n3975 = /* LUT   14  8  1 */ n1593;
assign n3976 = /* LUT   17 21  5 */ n2148;
assign n3977 = /* LUT   17 24  6 */ n2171;
assign n3978 = /* LUT   23 12  0 */ n3205;
assign n3979 = /* LUT   24 15  0 */ (n2122 ? (\rco[33]  ? \rco[0]  : 1'b0) : 1'b0);
assign n3980 = /* LUT   10  6  1 */ n975;
assign n3814 = /* LUT   27 23  1 */ (n2002 ? (n2361 ? (n2369 ? !n2589 : 1'b1) : 1'b1) : 1'b1);
assign n3982 = /* LUT    3 12  4 */ n282;
assign n3983 = /* LUT   31 24  3 */ (n116 ? \rco[127]  : 1'b0);
assign n3984 = /* LUT   18  2  6 */ n2204;
assign n3985 = /* LUT    7 17  0 */ n336;
assign n3986 = /* LUT   21 12  1 */ n2867;
assign n3987 = /* LUT   26 21  2 */ n3563;
assign n3988 = /* LUT   14 26  2 */ n1712;
assign n3989 = /* LUT   12 21  4 */ n1344;
assign n3990 = /* LUT   17 10  1 */ n2059;
assign n3991 = /* LUT   20  4  0 */ (\rco[93]  ? n2239 : 1'b0);
assign n3992 = /* LUT   19 20  2 */ n2566;
assign n3993 = /* LUT    1 12  6 */ n51;
assign n3994 = /* LUT   10  5  5 */ n970;
assign n3995 = /* LUT   22 14  2 */ n3052;
assign n3996 = /* LUT   27  8  2 */ (n3330 ? (\rco[0]  ? (n1752 ? \rco[66]  : 1'b0) : 1'b0) : 1'b0);
assign n3997 = /* LUT    3 17  1 */ n310;
assign n3998 = /* LUT   14 25  4 */ n1704;
assign n3999 = /* LUT    6 21  2 */ (n244 ? (n336 ? (n123 ? n326 : 1'b0) : 1'b0) : 1'b0);
assign n4000 = /* LUT   17  4  0 */ n2032;
assign n4001 = /* LUT   23 16  6 */ (\rco[99]  ? n1090 : 1'b0);
assign n4002 = /* LUT   11 14  7 */ n1295;
assign n4003 = /* LUT   20 10  1 */ n2683;
assign n4004 = /* LUT    5 14  7 */ n499;
assign n4005 = /* LUT   11 21  6 */ n1203;
assign n4006 = /* LUT   29 10  0 */ n3833;
assign n4007 = /* LUT   28 22  2 */ n3803;
assign n4008 = /* LUT   16 12  1 */ (n1772 ? \rco[41]  : 1'b0);
assign n4009 = /* LUT    5 19  3 */ n541;
assign n4010 = /* LUT   19  2  2 */ n2426;
assign n4011 = /* LUT   16 17  6 */ n1968;
assign n4012 = /* LUT   10 23  1 */ n1066;
assign n4013 = /* LUT   27  6  1 */ (\rco[0]  ? (n3718 ? (\rco[66]  ? n1752 : 1'b0) : 1'b0) : 1'b0);
assign n4014 = /* LUT   13 15  0 */ n812;
assign n4015 = /* LUT   30 12  0 */ n3463;
assign n4016 = /* LUT   15 17  7 */ n1800;
assign n4017 = /* LUT   18  6  3 */ n2233;
assign n4018 = /* LUT    7 21  5 */ n774;
assign n4019 = /* LUT    6  7  5 */ n575;
assign n4020 = /* LUT   20 24  2 */ n2789;
assign n4021 = /* LUT    3 18  5 */ n322;
assign n4022 = /* LUT    6  8  4 */ n577;
assign n4023 = /* LUT   20 21  5 */ n2774;
assign n4024 = /* LUT   14 11  0 */ n1617;
assign n4025 = /* LUT   17 22  4 */ n2155;
assign n4026 = /* LUT    1 19  1 */ n104;
assign n4027 = /* LUT   17 25  5 */ n2180;
assign n4028 = /* LUT   10 25  0 */ n1085;
assign n4029 = /* LUT   24 14  3 */ n3371;
assign n4030 = /* LUT   27 20  0 */ n3680;
assign n4031 = /* LUT    4 19  7 */ (\rco[123]  ? (\rco[0]  ? (n121 ? n336 : 1'b0) : 1'b0) : 1'b0);
assign n406  = /* LUT    3 13  3 */ (n56 ? 1'b0 : (n405 ? (n195 ? 1'b0 : n403) : 1'b0));
assign n4032 = /* LUT   22 10  7 */ n3028;
assign n4033 = /* LUT   18  5  7 */ n2222;
assign n4034 = /* LUT    7 22  1 */ n783;
assign n4035 = /* LUT    9 23  1 */ n769;
assign n4036 = /* LUT   21 13  2 */ n2875;
assign n4037 = /* LUT   26 20  1 */ (\rco[162]  ? (n2942 ? n3432 : 1'b0) : 1'b0);
assign n4038 = /* LUT   12 15  2 */ n1297;
assign n4039 = /* LUT   14 21  3 */ (n1671 ? (n1685 ? (\rco[0]  ? \rco[110]  : 1'b0) : 1'b0) : 1'b0);
assign n4040 = /* LUT   19 30  4 */ n2637;
assign n4041 = /* LUT   19 21  5 */ n2582;
assign n4042 = /* LUT   11 17  3 */ n1170;
assign n4043 = /* LUT   10 11  7 */ n1002;
assign n4044 = /* LUT   16  8  6 */ n1922;
assign n4045 = /* LUT    1 13  5 */ n65;
assign n4046 = /* LUT   24 17  7 */ n3400;
assign n4047 = /* LUT   28  7  4 */ n3722;
assign n4048 = /* LUT   22  9  3 */ n3016;
assign n4049 = /* LUT   15 21  4 */ n1839;
assign n4050 = /* LUT   20 28  7 */ n2830;
assign n4051 = /* LUT   17  5  3 */ (n823 ? \rco[145]  : 1'b0);
assign n4052 = /* LUT   20  9  0 */ (\rco[37]  ? (\rco[0]  ? (n1933 ? n2269 : 1'b0) : 1'b0) : 1'b0);
assign n4053 = /* LUT    6 20  1 */ n548;
assign n4054 = /* LUT   23 17  1 */ n3234;
assign n4055 = /* LUT   11 15  4 */ n1156;
assign n4056 = /* LUT   26  6  5 */ n3477;
assign n4057 = /* LUT   11 18  7 */ n1179;
assign n4058 = /* LUT   29 11  7 */ n3845;
assign n4059 = /* LUT   28 21  3 */ n3793;
assign n4060 = /* LUT   16 11  0 */ n2075;
assign n4061 = /* LUT   19  3  1 */ n2427;
assign n4062 = /* LUT    4 12  0 */ n491;
assign n4063 = /* LUT   13 16  1 */ n1477;
assign n4064 = /* LUT   27  7  2 */ n3598;
assign n4065 = /* LUT   15 22  6 */ n1852;
assign n4066 = /* LUT   18  9  2 */ n2253;
assign n4067 = /* LUT    7 26  4 */ n700;
assign n4068 = /* LUT    9 19  6 */ n908;
assign n4069 = /* LUT    3 19  6 */ n334;
assign n4070 = /* LUT    6 11  5 */ n603;
assign n4071 = /* LUT   12 24  0 */ n696;
assign n4072 = /* LUT   17 23  3 */ n2163;
assign n4073 = /* LUT   19 17  2 */ n2542;
assign n4074 = /* LUT   17 26  4 */ n2016;
assign n4075 = /* LUT   22 21  5 */ n3100;
assign n4076 = /* LUT   24 24  5 */ n3443;
assign n4077 = /* LUT   10 24  3 */ n1074;
assign n4078 = /* LUT   28 11  3 */ (n3033 ? (n3034 ? (n3463 ? n3636 : 1'b0) : 1'b0) : 1'b0);
assign n4079 = /* LUT   24 13  2 */ n3362;
assign n4080 = /* LUT   27 21  7 */ n3693;
assign n4081 = /* LUT    4 18  4 */ n433;
assign n4082 = /* LUT    3 10  2 */ n263;
assign n4083 = /* LUT   18  4  4 */ n2216;
assign n4084 = /* LUT    7 23  2 */ n791;
assign n4085 = /* LUT    9 16  0 */ n882;
assign n4086 = /* LUT   12 14  1 */ n1288;
assign n4087 = /* LUT   26 23  0 */ n3581;
assign n4088 = /* LUT   14 20  0 */ n1681;
assign n4089 = /* LUT    5  8  4 */ n472;
assign n4090 = /* LUT   19 31  7 */ n2647;
assign n4091 = /* LUT   23 21  6 */ n3276;
assign n4092 = /* LUT   19 18  4 */ n2557;
assign n4093 = /* LUT   10 10  0 */ (\rco[9]  ? \rco[0]  : 1'b0);
assign n4094 = /* LUT   16 23  7 */ n2165;
assign n4095 = /* LUT    1 14  4 */ n71;
assign n4096 = /* LUT   28  6  7 */ n3592;
assign n4097 = /* LUT   22  8  0 */ n3014;
assign n4098 = /* LUT   15 10  5 */ n1758;
assign n4099 = /* LUT    2 16  4 */ n201;
assign n4100 = /* LUT   20 19  6 */ n2754;
assign n4101 = /* LUT   18 22  0 */ (n2574 ? (n2357 ? (n2037 ? n817 : 1'b0) : 1'b0) : 1'b0);
assign n4102 = /* LUT   17  6  2 */ n2039;
assign n4103 = /* LUT    6 23  0 */ n361;
assign n4104 = /* LUT   20  8  7 */ n2657;
assign n4105 = /* LUT   12 28  5 */ n1398;
assign n4106 = /* LUT   23 22  0 */ n2934;
assign n4107 = /* LUT   11 19  4 */ n1172;
assign n4108 = /* LUT   29 12  6 */ n3855;
assign n4109 = /* LUT   16 10  3 */ n1928;
assign n676  = /* LUT    5 21  1 */ (n326 ? (n675 ? (n336 ? n562 : 1'b0) : 1'b0) : 1'b0);
assign n4111 = /* LUT   22 26  1 */ n3133;
assign n4112 = /* LUT   15 24  4 */ n1867;
assign n4113 = /* LUT   13 17  2 */ n1485;
assign n4114 = /* LUT   27  4  3 */ (\rco[74]  ? (n3175 ? n3456 : 1'b0) : 1'b0);
assign n4115 = /* LUT   15 23  5 */ n1856;
assign n4116 = /* LUT   18  8  1 */ n2254;
assign n4117 = /* LUT    3 16  7 */ n204;
assign n4118 = /* LUT   17 16  2 */ (\rco[0]  ? n2322 : 1'b0);
assign n4119 = /* LUT   19 14  3 */ n2515;
assign n4120 = /* LUT   22 20  6 */ n2924;
assign n4121 = /* LUT   10 14  5 */ n1011;
assign n4122 = /* LUT   24 23  4 */ n3438;
assign n4123 = /* LUT   22 25  5 */ n3129;
assign n4124 = /* LUT   10 27  2 */ n1094;
assign n4125 = /* LUT   24 12  5 */ n3357;
assign n2175 = /* LUT   16 24  3 */ (n117 ? (n2174 ? (n465 ? !\rco[0]  : 1'b1) : 1'b1) : 1'b1);
assign n4127 = /* LUT   28 10  0 */ n3636;
assign n4128 = /* LUT   27 18  6 */ n3662;
assign n4129 = /* LUT    4 17  5 */ n529;
assign n4130 = /* LUT    3 11  1 */ n270;
assign n4131 = /* LUT   18  7  5 */ n2245;
assign n4132 = /* LUT    9 17  3 */ n885;
assign n4133 = /* LUT   15  5  1 */ n1725;
assign n1860 = /* LUT   14 23  1 */ (n148 ? (n1113 ? n1231 : 1'b0) : 1'b0);
assign n4135 = /* LUT   20 12  4 */ n2701;
assign n4136 = /* LUT   19 19  7 */ (n1710 ? (n2760 ? (n2037 ? \rco[0]  : 1'b0) : 1'b0) : 1'b0);
assign n4137 = /* LUT   10 13  1 */ (\rco[99]  ? (n912 ? \rco[0]  : 1'b0) : 1'b0);
assign n4138 = /* LUT   16 22  4 */ n1989;
assign n4139 = /* LUT    1 15  3 */ (\rco[0]  ? n203 : 1'b0);
assign n4140 = /* LUT   16 27  7 */ n2194;
assign n4141 = /* LUT   22 11  1 */ (n2859 ? (n2494 ? \rco[53]  : 1'b0) : 1'b0);
assign n4142 = /* LUT   30 10  3 */ n3887;
assign n4143 = /* LUT   15 11  6 */ n1763;
assign n4144 = /* LUT    2 19  5 */ (\rco[99]  ? (n341 ? (n335 ? n216 : 1'b0) : 1'b0) : 1'b0);
assign n4145 = /* LUT    6 13  6 */ n620;
assign n4146 = /* LUT   15  6  5 */ n1737;
assign n4147 = /* LUT   17  7  5 */ n2050;
assign n4148 = /* LUT   18 25  1 */ n2377;
assign n4149 = /* LUT    6 22  7 */ n684;
assign n4150 = /* LUT   20 18  5 */ n2745;
assign n4151 = /* LUT   20 15  6 */ n2717;
assign n4152 = /* LUT   11 13  2 */ n1141;
assign n4153 = /* LUT   23 23  3 */ n3289;
assign n4154 = /* LUT   11 16  5 */ n1163;
assign n4155 = /* LUT    5 22  0 */ n682;
assign n4156 = /* LUT    9 13  1 */ n855;
assign n4157 = /* LUT   13  7  4 */ n1426;
assign n4158 = /* LUT   15 25  3 */ (\rco[183]  ? n1876 : 1'b0);
assign n4159 = /* LUT   13 18  3 */ n1494;
assign n4160 = /* LUT   27  5  4 */ n3588;
assign n4161 = /* LUT   18 11  0 */ (n2470 ? (\rco[41]  ? (\rco[0]  ? n2306 : 1'b0) : 1'b0) : 1'b0);
assign n4162 = /* LUT   15 20  4 */ n1830;
assign n4163 = /* LUT   26  7  3 */ n3483;
assign n4164 = /* LUT   17 17  1 */ n2114;
assign n4165 = /* LUT    2 14  0 */ n60;
assign n4166 = /* LUT   16  7  1 */ n1907;
assign n4167 = /* LUT   19 15  0 */ n2530;
assign n4168 = /* LUT   23  5  3 */ n3152;
assign n4169 = /* LUT   22 23  7 */ n3294;
assign n4170 = /* LUT   24 22  7 */ n3286;
assign n4171 = /* LUT   22 24  6 */ n3123;
assign n3466 = /* LUT   24 11  4 */ (n962 ? (n2680 ? n2067 : 1'b0) : 1'b0);
assign n1246 = /* LUT   10 26  5 */ (n1244 ? !n1243 : 1'b0);
assign n4172 = /* LUT   27 19  5 */ n3671;
assign n4173 = /* LUT   28  9  1 */ n3734;
assign n4174 = /* LUT    4 16  2 */ n421;
assign n4175 = /* LUT    9 18  2 */ n893;
assign n4176 = /* LUT   14 22  6 */ n1692;
assign n4177 = /* LUT   17  3  2 */ n2026;
assign n4178 = /* LUT    6 18  4 */ n652;
assign n4179 = /* LUT    5 10  6 */ n479;
assign n4180 = /* LUT   19 29  1 */ n2630;
assign n4181 = /* LUT   23 27  4 */ n3315;
assign n4182 = /* LUT   19 16  6 */ (n813 ? (n880 ? (n206 ? !n812 : 1'b1) : 1'b1) : 1'b1);
assign n4183 = /* LUT   11 28  0 */ n1260;
assign n4184 = /* LUT   10 12  2 */ n998;
assign n4185 = /* LUT   24 25  3 */ n3448;
assign n4186 = /* LUT   16 21  5 */ n1987;
assign n4187 = /* LUT    1  8  2 */ n15;
assign n4188 = /* LUT   16 26  4 */ n2015;
assign n4189 = /* LUT    9 28  1 */ n956;
assign n4190 = /* LUT    3 22  4 */ n356;
assign n4191 = /* LUT    2 18  2 */ n210;
assign n4192 = /* LUT    6 12  5 */ n610;
assign n4193 = /* LUT   15  7  6 */ (n587 ? (n1623 ? (\rco[0]  ? \rco[83]  : 1'b0) : 1'b0) : 1'b0);
assign n3009 = /* LUT   21  7  6 */ (n2440 ? (n2997 ? n2278 : 1'b0) : 1'b0);
assign n4194 = /* LUT   18 24  2 */ n2371;
assign n4195 = /* LUT   20 17  4 */ n2735;
assign n4196 = /* LUT   23 20  2 */ n3264;
assign n4197 = /* LUT   11 10  3 */ (n717 ? en_in : 1'b0);
assign n4198 = /* LUT   24  7  3 */ (n1491 ? (n3458 ? (n1752 ? \rco[59]  : 1'b0) : 1'b0) : 1'b0);
assign n4199 = /* LUT    9 14  0 */ n864;
assign n4200 = /* LUT    4 20  7 */ n102;
assign n1674 = /* LUT   13 19  4 */ (n777 ? (n667 ? (\rco[0]  ? !n335 : 1'b1) : 1'b1) : 1'b1);
assign n4202 = /* LUT   18 10  7 */ n2066;
assign n4203 = /* LUT   14 18  3 */ n1670;
assign n4204 = /* LUT   19 25  6 */ n2609;
assign n4205 = /* LUT   17 18  0 */ n2332;
assign n4206 = /* LUT   16  6  2 */ n1898;
assign n4207 = /* LUT   19 12  1 */ n2497;
assign n4208 = /* LUT   23 10  2 */ n3183;
assign n4209 = /* LUT   22 22  0 */ n2948;
assign n4210 = /* LUT   22 27  7 */ n3149;
assign n4211 = /* LUT   24 10  7 */ n3346;
assign n4212 = /* LUT   28  8  6 */ n3732;
assign n4213 = /* LUT   13  5  5 */ n1576;
assign n4214 = /* LUT    2 22  7 */ n353;
assign n4215 = /* LUT   17 12  3 */ n2079;
assign n4216 = /* LUT   19 26  0 */ (n2003 ? (\rco[172]  ? (n1998 ? \rco[0]  : 1'b0) : 1'b0) : 1'b0);
assign n4217 = /* LUT    5 11  1 */ n481;
assign n4218 = /* LUT   11 22  6 */ n565;
assign n4219 = /* LUT   23 24  5 */ n3303;
assign n4220 = /* LUT   23  7  4 */ n3169;
assign n4221 = /* LUT   11 29  7 */ n1268;
assign n4222 = /* LUT   10 15  3 */ n749;
assign n4223 = /* LUT   16 20  2 */ n2141;
assign n4224 = /* LUT    1  9  1 */ n160;
assign n4225 = /* LUT   16 25  5 */ n2007;
assign n4226 = /* LUT   21 24  2 */ n2954;
assign n4227 = /* LUT   13 23  1 */ n1524;
assign n4228 = /* LUT   27 14  0 */ n3647;
assign n4229 = /* LUT   18 14  4 */ (n2303 ? 1'b0 : (n2524 ? 1'b0 : (n2094 ? n1951 : 1'b0)));
assign n4230 = /* LUT    2 21  3 */ n229;
assign n4231 = /* LUT    6 15  4 */ n633;
assign n4232 = /* LUT   18 27  3 */ n2395;
assign n2897 = /* LUT   20 16  3 */ (n2550 ? (n2722 ? n2737 : 1'b0) : 1'b0);
assign n4233 = /* LUT    6 16  5 */ n642;
assign n4234 = /* LUT   20 13  4 */ n2709;
assign n4235 = /* LUT    4 11  5 */ n391;
assign n4236 = /* LUT   22 18  5 */ n3084;
assign n4237 = /* LUT   22  7  2 */ n2999;
assign n4238 = /* LUT   10 17  3 */ (\rco[99]  ? (n1176 ? 1'b0 : n912) : 1'b0);
assign n4239 = /* LUT    9 15  7 */ n873;
assign n4240 = /* LUT   24  6  0 */ n3327;
assign n4241 = /* LUT   28 12  3 */ n3755;
assign n4242 = /* LUT   13 20  5 */ n1507;
assign n4243 = /* LUT   18 13  6 */ n2300;
assign n4244 = /* LUT   16  5  3 */ n1890;
assign n4245 = /* LUT   23 11  1 */ n3190;
assign n4246 = /* LUT   11 25  4 */ n1234;
assign n4247 = /* LUT   22 17  1 */ n3072;
assign n4248 = /* LUT   24 20  1 */ n3414;
assign n4249 = /* LUT   16 16  7 */ n1957;
assign n4250 = /* LUT   10 28  7 */ n1107;
assign n4251 = /* LUT   24  9  6 */ n3339;
assign n4252 = /* LUT   13  6  4 */ n1418;
assign n4253 = /* LUT    4 22  0 */ (n113 ? (n462 ? (n122 ? \rco[132]  : 1'b0) : 1'b0) : 1'b0);
assign n4254 = /* LUT   21 23  0 */ n3066;
assign n4255 = /* LUT   15 13  5 */ n1781;
assign n4256 = /* LUT   29 19  5 */ n3865;
assign n4257 = /* LUT   14 16  4 */ n1649;
assign n4258 = /* LUT   17 13  0 */ n2092;
assign n4259 = /* LUT    5 12  0 */ n490;
assign n4260 = /* LUT   23 25  2 */ (\rco[183]  ? (n1876 ? n2797 : 1'b0) : 1'b0);
assign n4261 = /* LUT   11 23  5 */ n1218;
assign n4262 = /* LUT   19 27  3 */ n2618;
assign n4263 = /* LUT   11 26  6 */ n1242;
assign n4264 = /* LUT    1 10  0 */ n34;
assign n4265 = /* LUT   21 25  1 */ n2962;
assign n4266 = /* LUT    9 11  4 */ n845;
assign n4267 = /* LUT   13 24  0 */ (\rco[99]  ? \rco[0]  : 1'b0);
assign n4268 = /* LUT   15 14  1 */ n1783;
assign n4269 = /* LUT    3 20  6 */ n348;
assign n4270 = /* LUT    2 20  0 */ n222;
assign n4271 = /* LUT    6 14  3 */ n625;
assign n4272 = /* LUT   20 23  2 */ (n2002 ? (n2361 ? (n2369 ? n2589 : 1'b0) : 1'b0) : 1'b0);
assign n4273 = /* LUT   18 17  5 */ n2329;
assign n4274 = /* LUT   18 26  4 */ n2388;
assign n767  = /* LUT    6 19  4 */ (n336 ? n766 : 1'b0);
assign n4275 = /* LUT   11  8  1 */ n1123;
assign n4276 = /* LUT   29  5  1 */ n3818;
assign n4277 = /* LUT   28 19  1 */ n3777;
assign n4278 = /* LUT   19  9  3 */ n2473;
assign n4279 = /* LUT    4 10  6 */ n384;
assign n4280 = /* LUT   22 29  4 */ (n2539 ? (n982 ? \rco[172]  : 1'b0) : 1'b0);
assign n4281 = /* LUT   24 16  6 */ n3389;
assign n4282 = /* LUT   22  6  5 */ n2994;
assign n4283 = /* LUT   10 16  0 */ n1028;
assign n4284 = /* LUT   24  5  1 */ n3320;
assign n4285 = /* LUT   13 10  7 */ n1431;
assign n4286 = /* LUT   31 27  7 */ (\rco[138]  ? n1685 : 1'b0);
assign n4287 = /* LUT   18  3  4 */ (n1620 ? (\rco[0]  ? \rco[83]  : 1'b0) : 1'b0);
assign n4288 = /* LUT   13 21  6 */ n1519;
assign n4289 = /* LUT   18 12  5 */ n2290;
assign n4290 = /* LUT   21  6  2 */ n2834;
assign n4291 = /* LUT   29 23  2 */ n3882;
assign n1774 = /* LUT   14 12  1 */ (n1623 ? (n1773 ? 1'b0 : n1420) : 1'b0);
assign n4292 = /* LUT   19 23  4 */ (n1666 ? (n817 ? (\rco[23]  ? !n1620 : 1'b1) : 1'b1) : 1'b1);
assign n4293 = /* LUT   19 10  7 */ n2690;
assign n4294 = /* LUT   24 19  0 */ n3401;
assign n4295 = /* LUT   28 14  4 */ n3764;
assign n4296 = /* LUT    4 21  1 */ n447;
assign n4297 = /* LUT    7 13  0 */ (n811 ? (n737 ? \rco[153]  : 1'b0) : 1'b0);
assign n4298 = /* LUT   21  8  1 */ n2832;
assign n4299 = /* LUT   26 17  2 */ n3547;
assign n4300 = /* LUT   18 30  1 */ n2417;
assign n4301 = /* LUT   14 19  5 */ n1668;
assign n4302 = /* LUT   17 14  1 */ n1919;
assign n4303 = /* LUT   29 20  4 */ n3871;
assign n4304 = /* LUT    5 13  3 */ n500;
assign n4305 = /* LUT   19 24  2 */ n2595;
assign n4306 = /* LUT   11 20  4 */ n1192;
assign n4307 = /* LUT   11 27  5 */ n1251;
assign n4308 = /* LUT   16 18  0 */ n1499;
assign n4309 = /* LUT   21 26  0 */ (n2044 ? (\rco[172]  ? (n2563 ? n2400 : 1'b0) : 1'b0) : 1'b0);
assign n4310 = /* LUT   13 25  3 */ n1536;
assign n4311 = /* LUT   27 12  2 */ n3629;
assign n1952 = /* LUT   15 15  2 */ (n758 ? (n1130 ? (\rco[0]  ? !n823 : 1'b1) : 1'b1) : 1'b1);
assign n4313 = /* LUT    3 21  1 */ (n243 ? (n458 ? (n361 ? n439 : 1'b0) : 1'b0) : 1'b0);
assign n4314 = /* LUT   18 16  6 */ n2319;
assign n727  = /* LUT    6  9  2 */ (n76 ? (n726 ? (n54 ? n277 : 1'b0) : 1'b0) : 1'b0);
assign n4315 = /* LUT   18 29  5 */ n2412;
assign n4316 = /* LUT   20 22  1 */ n2776;
assign n4317 = /* LUT   28 18  2 */ n3774;
assign n4318 = /* LUT   19  6  2 */ n2444;
assign n4319 = /* LUT    4  9  7 */ n259;
assign n4320 = /* LUT   24 15  7 */ n3391;
assign n4321 = /* LUT   10 19  1 */ (\rco[99]  ? (n1188 ? 1'b0 : (n121 ? !n224 : 1'b0)) : 1'b0);
assign n4322 = /* LUT    9  9  5 */ n831;
assign n4323 = /* LUT   13 11  0 */ n1619;
assign n4324 = /* LUT   18  2  3 */ n2201;
assign n4325 = /* LUT   13 22  7 */ n1695;
assign n4326 = /* LUT   18 15  4 */ n2312;
assign n4327 = /* LUT   14 26  7 */ n1550;
assign n4328 = /* LUT   26 14  0 */ n3536;
assign n4329 = /* LUT   14 15  0 */ n1644;
assign n4330 = /* LUT    2  9  5 */ n24;
assign n4331 = /* LUT   20  4  5 */ n2654;
assign n4332 = /* LUT   19 20  5 */ n2569;
assign n4333 = /* LUT   19 11  4 */ n2489;
assign n4334 = /* LUT   23  9  7 */ n3182;
assign n4335 = /* LUT   22 19  3 */ (n3259 ? (n3261 ? (\rco[0]  ? \rco[153]  : 1'b0) : 1'b0) : 1'b0);
assign n4336 = /* LUT   10  5  0 */ \rco[0] ;
assign n4337 = /* LUT   24 18  3 */ n3404;
assign n4338 = /* LUT   28 13  5 */ n3650;
assign n4339 = /* LUT   21  9  2 */ n2846;
assign n4340 = /* LUT    9 27  1 */ n949;
assign n4341 = /* LUT    3 17  6 */ n316;
assign n4342 = /* LUT   14 25  3 */ n1703;
assign n4343 = /* LUT   29 21  7 */ n3798;
assign n4344 = /* LUT   17 15  6 */ n2106;
assign n4345 = /* LUT   20  7  1 */ n2661;
assign n4346 = /* LUT    5 14  2 */ n509;
assign n4347 = /* LUT   11 21  3 */ n1200;
assign n4348 = /* LUT   11 24  4 */ n1226;
assign n4349 = /* LUT   16 17  1 */ n1958;
assign n4350 = /* LUT   22 13  3 */ n2416;
assign n4351 = /* LUT   21 27  7 */ n2986;
assign n4352 = /* LUT   27  6  4 */ (n3330 ? (\rco[0]  ? (n3455 ? \rco[74]  : 1'b0) : 1'b0) : 1'b0);
assign n4353 = /* LUT   13 15  5 */ n1474;
assign n4354 = /* LUT   30 12  5 */ n3898;
assign n4355 = /* LUT    9 24  5 */ n1078;
assign n4356 = /* LUT   13 26  2 */ n1545;
assign n4357 = /* LUT   18 19  7 */ n2135;
assign n4358 = /* LUT    3 18  0 */ n326;
assign n4359 = /* LUT    6  8  1 */ n580;
assign n4360 = /* LUT   18 28  6 */ n2405;
assign n4361 = /* LUT   20 21  0 */ n2773;
assign n4362 = /* LUT    1 19  6 */ n109;
assign n4363 = /* LUT   28 17  3 */ n3768;
assign n4364 = /* LUT   16 15  0 */ n1948;
assign n4365 = /* LUT   19  7  1 */ n2452;
assign n4366 = /* LUT   23 13  4 */ n3211;
assign n4367 = /* LUT   10 25  7 */ n797;
assign n4368 = /* LUT   24 14  4 */ n3372;
assign n4369 = /* LUT   10 18  6 */ n1040;
assign n4370 = /* LUT    9 10  4 */ n837;
assign n4371 = /* LUT   13 12  1 */ n1449;
assign n4372 = /* LUT   31 25  1 */ (n336 ? \rco[127]  : 1'b0);
assign n4373 = /* LUT   18  5  2 */ n2227;
assign n4374 = /* LUT   20 27  3 */ n2816;
assign n4375 = /* LUT   14 21  6 */ (\rco[99]  ? (\rco[0]  ? (n335 ? n1671 : 1'b0) : 1'b0) : 1'b0);
assign n4376 = /* LUT   12 20  0 */ (n335 ? (\rco[0]  ? (n1337 ? \rco[99]  : 1'b0) : 1'b0) : 1'b0);
assign n4377 = /* LUT   14 14  7 */ n1790;
assign n4378 = /* LUT   17 11  3 */ n2070;
assign n4379 = /* LUT    1 16  0 */ n92;
assign n4380 = /* LUT   19 21  2 */ n2577;
assign n4381 = /* LUT   19  8  5 */ n2465;
assign n4382 = /* LUT   23 14  6 */ n3221;
assign n4383 = /* LUT   24 17  2 */ n3395;
assign n4384 = /* LUT   28  7  3 */ n3721;
assign n4385 = /* LUT    3 14  2 */ (n278 ? (n289 ? (n87 ? !n287 : 1'b1) : 1'b1) : 1'b1);
assign n4386 = /* LUT   21 10  3 */ (n2457 ? (n2671 ? (\rco[48]  ? \rco[0]  : 1'b0) : 1'b0) : 1'b0);
assign n1056 = /* LUT    9 20  0 */ (n114 ? (\rco[0]  ? (n696 ? !n1043 : 1'b1) : 1'b1) : 1'b1);
assign n4388 = /* LUT    7 19  2 */ n760;
assign n4389 = /* LUT   26 19  0 */ (\rco[35]  ? \rco[0]  : 1'b0);
assign n4390 = /* LUT   27  9  2 */ n3611;
assign n1873 = /* LUT   14 24  0 */ (n658 ? (n1709 ? (n563 ? n671 : 1'b0) : 1'b0) : 1'b0);
assign n4392 = /* LUT   17  5  4 */ (n2044 ? \rco[172]  : 1'b0);
assign n4393 = /* LUT   17  8  7 */ (\rco[93]  ? (n2057 ? \rco[0]  : 1'b0) : 1'b0);
assign n4394 = /* LUT    2  7  4 */ n250;
assign n4395 = /* LUT   11 18  2 */ n1180;
assign n4396 = /* LUT    4 12  5 */ n397;
assign n4397 = /* LUT   22 12  0 */ n2857;
assign n1213 = /* LUT   10 22  3 */ (n551 ? (n669 ? (n550 ? n769 : 1'b0) : 1'b0) : 1'b0);
assign n4399 = /* LUT   21 28  6 */ n2984;
assign n4400 = /* LUT   13 16  4 */ n1480;
assign n4401 = /* LUT   27  7  7 */ n3472;
assign n4402 = /* LUT    9 25  6 */ n940;
assign n4403 = /* LUT   27 10  4 */ (n1491 ? (n3525 ? (\rco[0]  ? \rco[59]  : 1'b0) : 1'b0) : 1'b0);
assign n4404 = /* LUT   13 27  5 */ n1555;
assign n4405 = /* LUT   18 18  0 */ n2337;
assign n4406 = /* LUT    3 19  3 */ n331;
assign n4407 = /* LUT    6 11  0 */ n604;
assign n4408 = /* LUT   23 18  0 */ n3247;
assign n4409 = /* LUT   14 10  4 */ n1607;
assign n4410 = /* LUT   19 17  7 */ n2547;
assign n4411 = /* LUT    5 17  1 */ n524;
assign n4412 = /* LUT    4 15  1 */ n412;
assign n4413 = /* LUT   10 24  4 */ n1075;
assign n4414 = /* LUT   28 11  6 */ (n3752 ? 1'b0 : n3848);
assign n4415 = /* LUT   24 13  5 */ n3365;
assign n4416 = /* LUT   10 21  7 */ n921;
assign n4417 = /* LUT   13 13  2 */ n1456;
assign n4418 = /* LUT   18  4  1 */ n2213;
assign n4419 = /* LUT   20 26  0 */ n2810;
assign n4420 = /* LUT   14 20  5 */ n1680;
assign n1559 = /* LUT   12 27  1 */ (n1543 ? (n1244 ? n1272 : 1'b0) : 1'b0);
assign n4422 = /* LUT   17 20  2 */ n2137;
assign n4423 = /* LUT   19 18  3 */ n2556;
assign n4424 = /* LUT   23 15  5 */ n3226;
assign n4425 = /* LUT   28  6  0 */ n3716;
assign n4426 = /* LUT    3 15  1 */ n293;
assign n4427 = /* LUT   21 16  5 */ n2891;
assign n4428 = /* LUT    7 16  3 */ n743;
assign n4429 = /* LUT    9 21  3 */ n916;
assign n4430 = /* LUT   21 11  4 */ n2862;
assign n4431 = /* LUT   26 18  7 */ (\rco[23]  ? (n2534 ? (n2537 ? n3555 : 1'b0) : 1'b0) : 1'b0);
assign n4432 = /* LUT   18 22  5 */ (n817 ? (n2574 ? (n2369 ? !n2589 : 1'b1) : 1'b1) : 1'b1);
assign n4433 = /* LUT   14 27  1 */ n1720;
assign n4434 = /* LUT   17  6  5 */ n2053;
assign n4435 = /* LUT   17  9  4 */ (\rco[23]  ? (\rco[0]  ? (n2270 ? n1933 : 1'b0) : 1'b0) : 1'b0);
assign n3876 = /* LUT   28 20  1 */ (n3259 ? n3093 : 1'b0);
assign n4436 = /* LUT   22 26  6 */ n3138;
assign n4437 = /* LUT   22 15  1 */ n3058;
assign n4438 = /* LUT    7  6  6 */ n579;
assign n4439 = /* LUT    9  7  0 */ (\rco[0]  ? en_in : 1'b0);
assign n4440 = /* LUT   13 17  7 */ n1469;
assign n4441 = /* LUT   13 28  4 */ n1564;
assign n4442 = /* LUT   18 21  1 */ n2349;
assign n4443 = /* LUT    3 16  2 */ n304;
assign n4444 = /* LUT   23 19  3 */ n3252;
assign n4445 = /* LUT   14  5  5 */ n1575;
assign n4446 = /* LUT   19 14  6 */ n2518;
assign n4447 = /* LUT   17 27  0 */ n2269;
assign n4448 = /* LUT   28 23  5 */ n3807;
assign n4449 = /* LUT    5 18  0 */ n536;
assign n513  = /* LUT    4 14  2 */ (n278 ? (n287 ? (n261 ? !n87 : 1'b1) : 1'b1) : 1'b1);
assign n4451 = /* LUT   19  5  7 */ n2225;
assign n4452 = /* LUT   10 27  5 */ n1097;
assign n4453 = /* LUT   22 25  0 */ n3130;
assign n4454 = /* LUT   24 12  2 */ n3354;
assign n4455 = /* LUT   28 10  5 */ n3745;
assign n4456 = /* LUT   10 20  4 */ n1051;
assign n4457 = /* LUT   13 14  3 */ n1464;
assign n4458 = /* LUT   18  7  0 */ n2243;
assign n4459 = /* LUT   20 25  1 */ n2798;
assign n4460 = /* LUT   15  5  6 */ n1731;
assign n4461 = /* LUT   14 23  4 */ n936;
assign n4462 = /* LUT   12 26  2 */ n1386;
assign n4463 = /* LUT   14  8  5 */ n1597;
assign n4464 = /* LUT    2 10  0 */ n167;
assign n4465 = /* LUT    1 18  2 */ n214;
assign n4466 = /* LUT   19 19  0 */ (n2759 ? (\rco[162]  ? (n807 ? n1409 : 1'b0) : 1'b0) : 1'b0);
assign n4467 = /* LUT   17 21  1 */ n2144;
assign n4468 = /* LUT   23 12  4 */ n3203;
assign n4469 = /* LUT   28  5  1 */ n3705;
assign n4470 = /* LUT    3 12  0 */ (n278 ? (\rco[0]  ? (n261 ? \rco[11]  : 1'b0) : 1'b0) : 1'b0);
assign n4471 = /* LUT   21 17  6 */ n2899;
assign n4472 = /* LUT    7 17  4 */ n754;
assign n4473 = /* LUT   21 12  5 */ n2871;
assign n4474 = /* LUT   12  8  7 */ n1280;
assign n4475 = /* LUT   26 21  6 */ n3568;
assign n4476 = /* LUT   15  6  0 */ n1739;
assign n4477 = /* LUT   17  7  2 */ n2047;
assign n4478 = /* LUT   18 25  4 */ n2380;
assign n4479 = /* LUT   17 10  5 */ n2063;
assign n4480 = /* LUT   11 16  0 */ n738;
assign n4481 = /* LUT   10  8  2 */ (n758 ? (n1130 ? (n823 ? \rco[145]  : 1'b0) : 1'b0) : 1'b0);
assign n4482 = /* LUT    1 12  2 */ n47;
assign n4483 = /* LUT   22 14  6 */ n3057;
assign n4484 = /* LUT    7  7  5 */ n715;
assign n4485 = /* LUT   13 18  6 */ n1497;
assign n4486 = /* LUT   27  5  1 */ n3585;
assign n4487 = /* LUT   27  8  6 */ n3609;
assign n3393 = /* LUT   23 16  2 */ (\rco[37]  ? n1047 : 1'b0);
assign n4488 = /* LUT   11 14  3 */ n1150;
assign n4489 = /* LUT    2 14  5 */ n191;
assign n4490 = /* LUT   16  7  4 */ n1910;
assign n4491 = /* LUT   19 15  5 */ n2529;
assign n4492 = /* LUT   28 22  6 */ n3801;
assign n4493 = /* LUT   16 12  5 */ n1939;
assign n4494 = /* LUT    5 19  7 */ n430;
assign n4495 = /* LUT    4 13  3 */ (\rco[0]  ? (n103 ? (\rco[17]  ? n291 : 1'b0) : 1'b0) : 1'b0);
assign n4496 = /* LUT   22 24  3 */ n3118;
assign n4497 = /* LUT   24 11  3 */ (\rco[48]  ? (n3465 ? (\rco[0]  ? n2725 : 1'b0) : 1'b0) : 1'b0);
assign n4498 = /* LUT   10 26  2 */ (\rco[99]  ? (n1087 ? (n1090 ? n1221 : 1'b0) : 1'b0) : 1'b0);
assign n4499 = /* LUT   28  9  4 */ n3737;
assign n4500 = /* LUT   10 23  5 */ n1067;
assign n4501 = /* LUT    7 21  1 */ n770;
assign n4502 = /* LUT    6  7  1 */ n571;
assign n4503 = /* LUT   20 24  6 */ n2793;
assign n4504 = /* LUT   26  9  5 */ n3502;
assign n4505 = /* LUT   29 17  4 */ n3860;
assign n4506 = /* LUT   14 22  3 */ n1689;
assign n4507 = /* LUT   12 25  3 */ n1378;
assign n4508 = /* LUT   14 11  4 */ n1615;
assign n4509 = /* LUT   17 22  0 */ n2361;
assign n4510 = /* LUT   19 16  1 */ (n2538 ? 1'b0 : (n2731 ? (n2535 ? 1'b0 : !n2536) : 1'b0));
assign n4511 = /* LUT   23  6  2 */ n3160;
assign n4512 = /* LUT   16 26  1 */ n2012;
assign n4513 = /* LUT    4 19  3 */ (n326 ? (\rco[0]  ? (n327 ? n336 : 1'b0) : 1'b0) : 1'b0);
assign n4514 = /* LUT    3 13  7 */ (n56 ? 1'b0 : (n290 ? 1'b0 : (n285 ? n403 : 1'b0)));
assign n4515 = /* LUT   21 18  7 */ n2903;
assign n4516 = /* LUT   22 10  3 */ n3024;
assign n4517 = /* LUT    7 22  5 */ n787;
assign n4518 = /* LUT    9 23  5 */ n929;
assign n4519 = /* LUT   21 13  6 */ n2885;
assign n4520 = /* LUT   12 15  6 */ n1301;
assign n3685 = /* LUT   26 20  5 */ (n2942 ? (n3684 ? (n3417 ? n2934 : 1'b0) : 1'b0) : 1'b0);
assign n1914 = /* LUT   15  7  3 */ (n1601 ? (n1460 ? (n1752 ? !n1602 : 1'b0) : 1'b0) : 1'b0);
assign n4521 = /* LUT   19 30  0 */ n2639;
assign n4522 = /* LUT   10 11  3 */ n992;
assign n4523 = /* LUT   16  8  2 */ n1916;
assign n4524 = /* LUT    1 13  1 */ n61;
assign n4525 = /* LUT   22  4  4 */ (n2278 ? \rco[44]  : 1'b0);
assign n4526 = /* LUT   13 19  1 */ (\rco[138]  ? (n667 ? n777 : 1'b0) : 1'b0);
assign n4527 = /* LUT   15 21  0 */ n667;
assign n4528 = /* LUT   20 28  3 */ n2825;
assign n4529 = /* LUT   18 23  3 */ n2364;
assign n4530 = /* LUT   23 17  5 */ n3238;
assign n4531 = /* LUT   11 15  0 */ (n817 ? (\rco[0]  ? (n732 ? \rco[145]  : 1'b0) : 1'b0) : 1'b0);
assign n4532 = /* LUT   26  6  1 */ n3473;
assign n4533 = /* LUT   14  7  7 */ n1745;
assign n4534 = /* LUT   16  6  7 */ n1903;
assign n4535 = /* LUT   19 12  4 */ n2500;
assign n4536 = /* LUT   28 21  7 */ n3797;
assign n4537 = /* LUT   19  3  5 */ n2431;
assign n4538 = /* LUT   22 27  2 */ n3144;
assign n4539 = /* LUT   10 29  3 */ n1108;
assign n4540 = /* LUT   24 10  0 */ n3337;
assign n4541 = /* LUT   28  8  3 */ n3728;
assign n4542 = /* LUT    3  9  4 */ n255;
assign n4543 = /* LUT    7 26  0 */ n800;
assign n4544 = /* LUT    9 19  2 */ n902;
assign n4545 = /* LUT   12 19  5 */ n1332;
assign n4546 = /* LUT   26  8  6 */ n3495;
assign n4547 = /* LUT   29 18  5 */ n3776;
assign n4548 = /* LUT   14 17  2 */ n1655;
assign n4549 = /* LUT   12 24  4 */ n1370;
assign n4550 = /* LUT   17 12  6 */ n2082;
assign n4551 = /* LUT    2 12  2 */ n177;
assign n4552 = /* LUT   23  7  1 */ n3166;
assign n4553 = /* LUT   22 21  1 */ n3096;
assign n4554 = /* LUT   24 24  1 */ n3439;
assign n4555 = /* LUT   16 25  0 */ (\rco[99]  ? (n1337 ? !n1521 : 1'b0) : 1'b0);
assign n4556 = /* LUT    4 18  0 */ n244;
assign n4557 = /* LUT    3 10  6 */ n269;
assign n4558 = /* LUT   21 19  0 */ n2917;
assign n4559 = /* LUT   13 23  6 */ n1529;
assign n4560 = /* LUT   27 14  7 */ n3646;
assign n4561 = /* LUT    7 23  6 */ n776;
assign n4562 = /* LUT    9 16  4 */ n874;
assign n4563 = /* LUT   12 14  5 */ n1148;
assign n4564 = /* LUT   26 23  4 */ n3579;
assign n4565 = /* LUT   18 27  6 */ n2399;
assign n4566 = /* LUT    5  8  0 */ n474;
assign n4567 = /* LUT   19 31  3 */ n2643;
assign n4568 = /* LUT   23 21  2 */ n3272;
assign n4569 = /* LUT   10 10  4 */ n986;
assign n4570 = /* LUT   16 23  3 */ n1993;
assign n4571 = /* LUT    1 14  0 */ n74;
assign n4572 = /* LUT   22  7  5 */ n2996;
assign n1178 = /* LUT   10 17  6 */ (n1031 ? n1177 : 1'b0);
assign n4573 = /* LUT   24  6  5 */ n3325;
assign n4574 = /* LUT   22  8  4 */ n3011;
assign n4575 = /* LUT   13 20  0 */ n137;
assign n4576 = /* LUT   15 10  1 */ n1756;
assign n4577 = /* LUT    2 16  0 */ n205;
assign n4578 = /* LUT   20 19  2 */ n2750;
assign n4579 = /* LUT   12 28  1 */ n1558;
assign n4580 = /* LUT   23 22  4 */ n3282;
assign n4581 = /* LUT   14  6  0 */ (n1584 ? (n1578 ? (\rco[0]  ? \rco[83]  : 1'b0) : 1'b0) : 1'b0);
assign n4582 = /* LUT   16  5  6 */ n1893;
assign n4583 = /* LUT   17 19  4 */ n2131;
assign n4584 = /* LUT   19 13  3 */ n2509;
assign n4585 = /* LUT   16 10  7 */ n1924;
assign n4586 = /* LUT    5 21  5 */ (n244 ? (n338 ? (n123 ? n361 : 1'b0) : 1'b0) : 1'b0);
assign n4587 = /* LUT   10 28  0 */ n148;
assign n4588 = /* LUT   24  9  1 */ n3332;
assign n4589 = /* LUT   27 17  0 */ n3655;
assign n4590 = /* LUT   15 24  0 */ n1868;
assign n4591 = /* LUT   21 23  5 */ n2947;
assign n4592 = /* LUT   12 18  6 */ n1325;
assign n4593 = /* LUT   26 11  7 */ n3514;
assign n4594 = /* LUT   29 19  2 */ n3862;
assign n4595 = /* LUT   14 16  1 */ n1646;
assign n4596 = /* LUT   17 13  5 */ n2090;
assign n2325 = /* LUT   17 16  6 */ (n813 ? (n2324 ? (n1960 ? n2119 : 1'b0) : 1'b0) : 1'b0);
assign n4597 = /* LUT    2 15  3 */ n196;
assign n4598 = /* LUT   22 20  2 */ n3089;
assign n4599 = /* LUT   10 14  1 */ n1007;
assign n4600 = /* LUT   24 23  0 */ n3437;
assign n4601 = /* LUT    4 17  1 */ n426;
assign n4602 = /* LUT    3 11  5 */ n274;
assign n4603 = /* LUT    7  9  0 */ (n87 ? (n154 ? n719 : 1'b0) : 1'b0);
assign n4604 = /* LUT   21 20  1 */ n2923;
assign n4605 = /* LUT   13 24  7 */ (n1337 ? (n338 ? !n335 : 1'b1) : 1'b1);
assign n4606 = /* LUT    9 17  7 */ n888;
assign n4607 = /* LUT   19 22  0 */ n2360;
assign n4608 = /* LUT   18 26  1 */ n2385;
assign n4609 = /* LUT   17  2  1 */ (n614 ? (n1583 ? \rco[83]  : 1'b0) : 1'b0);
assign n4610 = /* LUT   20 12  0 */ n2691;
assign n4611 = /* LUT    5  9  3 */ n473;
assign n4612 = /* LUT   28 19  4 */ n3780;
assign n4613 = /* LUT   10 13  5 */ n1005;
assign n4614 = /* LUT   16 22  0 */ (\rco[118]  ? (n129 ? \rco[0]  : 1'b0) : 1'b0);
assign n4615 = /* LUT   22  6  2 */ n2991;
assign n4616 = /* LUT   10 16  5 */ n1027;
assign n4617 = /* LUT   24  5  4 */ n3157;
assign n4618 = /* LUT   22 11  5 */ (n1491 ? (\rco[0]  ? (\rco[48]  ? n2725 : 1'b0) : 1'b0) : 1'b0);
assign n4619 = /* LUT   13 21  3 */ n1515;
assign n4620 = /* LUT   15 11  2 */ n1769;
assign n339  = /* LUT    2 19  1 */ (n326 ? n336 : 1'b0);
assign n4621 = /* LUT    6 13  2 */ n616;
assign n4622 = /* LUT   20 18  1 */ n2741;
assign n4623 = /* LUT   23 23  7 */ n3435;
assign n4624 = /* LUT   11 13  6 */ n1145;
assign n4625 = /* LUT   19 10  2 */ n2480;
assign n4626 = /* LUT    5 22  4 */ n558;
assign n4627 = /* LUT   28 14  1 */ n3761;
assign n4628 = /* LUT   13  7  0 */ n1420;
assign n4629 = /* LUT   15 25  7 */ n1875;
assign n4630 = /* LUT    7 13  5 */ (\rco[153]  ? (n738 ? n736 : 1'b0) : 1'b0);
assign n4631 = /* LUT   12 17  7 */ n1318;
assign n4632 = /* LUT   26 10  0 */ n3506;
assign n4633 = /* LUT   18 30  6 */ n2423;
assign n1826 = /* LUT   14 19  0 */ (n1813 ? (n1667 ? (n667 ? !n1684 : 1'b1) : 1'b1) : 1'b1);
assign n4635 = /* LUT   17 14  4 */ n2097;
assign n4636 = /* LUT   26  7  7 */ n3497;
assign n4637 = /* LUT   29 20  3 */ n3870;
assign n4638 = /* LUT   17 17  5 */ n2121;
assign n4639 = /* LUT   22 23  3 */ (n2173 ? (\rco[172]  ? (n2229 ? \rco[0]  : 1'b0) : 1'b0) : 1'b0);
assign n4640 = /* LUT   24 22  3 */ n3427;
assign n4641 = /* LUT    1 11  4 */ n40;
assign n4642 = /* LUT    7 14  1 */ n734;
assign n4643 = /* LUT   21 21  2 */ n2927;
assign n4644 = /* LUT   13 25  4 */ n1537;
assign n4645 = /* LUT   27 12  5 */ n3633;
assign n4646 = /* LUT    9 18  6 */ n897;
assign n4647 = /* LUT   18 29  0 */ n1872;
assign n4648 = /* LUT    6 18  0 */ n123;
assign n4649 = /* LUT    5 10  2 */ n475;
assign n4650 = /* LUT   19 29  5 */ n2633;
assign n4651 = /* LUT   11  9  3 */ n1132;
assign n4652 = /* LUT   23 27  0 */ n3316;
assign n4653 = /* LUT   24 25  7 */ n3452;
assign n4654 = /* LUT   16 21  1 */ n1983;
assign n4655 = /* LUT    1  8  6 */ n18;
assign n4656 = /* LUT   10 19  4 */ n1044;
assign n4657 = /* LUT   13 22  2 */ (n669 ? (n696 ? (n114 ? !n550 : 1'b1) : 1'b1) : 1'b1);
assign n4658 = /* LUT   15  8  3 */ n1599;
assign n4659 = /* LUT    3 22  0 */ n359;
assign n4660 = /* LUT   21  7  2 */ (n2440 ? (n3007 ? (\rco[0]  ? n2278 : 1'b0) : 1'b0) : 1'b0);
assign n4661 = /* LUT    6 12  1 */ n606;
assign n4662 = /* LUT   20 17  0 */ n2738;
assign n4663 = /* LUT   26 14  5 */ n3540;
assign n4664 = /* LUT   23 20  6 */ n3270;
assign n4665 = /* LUT   19 11  1 */ n2486;
assign n4666 = /* LUT    4 20  3 */ n442;
assign n4667 = /* LUT    7 18  4 */ n441;
assign n4668 = /* LUT    9 27  6 */ n951;
assign n4669 = /* LUT   21  9  7 */ n3021;
assign n4670 = /* LUT   12 16  0 */ n1309;
assign n3640 = /* LUT   26 13  1 */ (n3619 ? n3639 : 1'b0);
assign n4671 = /* LUT   29 21  0 */ n3880;
assign n4672 = /* LUT   17 15  3 */ n2107;
assign n4673 = /* LUT   19 25  2 */ n2605;
assign n4674 = /* LUT   22 22  4 */ n3105;
assign n4675 = /* LUT   24 21  2 */ (n3432 ? (n3470 ? (n2942 ? n3417 : 1'b0) : 1'b0) : 1'b0);
assign n4676 = /* LUT   22 13  6 */ n3048;
assign n814  = /* LUT    7 15  2 */ (n301 ? n740 : 1'b0);
assign n4677 = /* LUT    9 24  0 */ n937;
assign n4678 = /* LUT   13 26  5 */ n1548;
assign n4679 = /* LUT   21 22  3 */ n2937;
assign n4680 = /* LUT   27 13  2 */ n3461;
assign n4681 = /* LUT    2 22  3 */ n237;
assign n4682 = /* LUT   18 28  3 */ n2402;
assign n4683 = /* LUT   19 26  4 */ (\rco[0]  ? (n2813 ? (n1998 ? n1876 : 1'b0) : 1'b0) : 1'b0);
assign n4684 = /* LUT   23 24  1 */ n3296;
assign n4685 = /* LUT   11 22  2 */ n1207;
assign n4686 = /* LUT   28 17  6 */ n3772;
assign n4687 = /* LUT   16 15  7 */ n1167;
assign n4688 = /* LUT   10 15  7 */ n1019;
assign n4689 = /* LUT   16 20  6 */ n1981;
assign n4690 = /* LUT   10 18  3 */ n1035;
assign n4691 = /* LUT   15 18  5 */ n1812;
assign n4692 = /* LUT   20 27  6 */ n2819;
assign n2523 = /* LUT   18 14  0 */ (n2304 ? n2239 : 1'b0);
assign n4693 = /* LUT    2 21  7 */ n233;
assign n4694 = /* LUT    6 15  0 */ (\rco[8]  ? \rco[0]  : 1'b0);
assign n4695 = /* LUT   20 16  7 */ (n2725 ? (n2728 ? (\rco[0]  ? \rco[48]  : 1'b0) : 1'b0) : 1'b0);
assign n4696 = /* LUT   12 20  5 */ (n114 ? (n1337 ? (n696 ? n335 : 1'b0) : 1'b0) : 1'b0);
assign n4697 = /* LUT   19  8  0 */ n2476;
assign n4698 = /* LUT    4 11  1 */ n387;
assign n4699 = /* LUT   22 18  1 */ n3080;
assign n4700 = /* LUT   13  9  2 */ n1284;
assign n4701 = /* LUT    7 19  7 */ n646;
assign n4702 = /* LUT    9 20  7 */ n957;
assign n3030 = /* LUT   21 10  6 */ (\rco[37]  ? (n2679 ? 1'b0 : (n2306 ? n2510 : 1'b0)) : 1'b0);
assign n4703 = /* LUT   27  9  7 */ n3616;
assign n4704 = /* LUT   21  5  7 */ n2840;
assign n4705 = /* LUT   12 23  1 */ n1358;
assign n4706 = /* LUT   26 12  2 */ n3518;
assign n2257 = /* LUT   17  8  2 */ (n1583 ? (n587 ? (n1603 ? !n614 : 1'b1) : 1'b1) : 1'b1);
assign n4708 = /* LUT    5 15  2 */ n515;
assign n4709 = /* LUT   19 22  3 */ n2586;
assign n4710 = /* LUT   11 25  0 */ (\rco[104]  ? n1221 : 1'b0);
assign n4711 = /* LUT   22 17  5 */ n3076;
assign n4712 = /* LUT   24 20  5 */ n3416;
assign n4713 = /* LUT   16 16  3 */ n1955;
assign n4714 = /* LUT   22 12  5 */ n3040;
assign n4715 = /* LUT    4 22  4 */ n426;
assign n4716 = /* LUT    9 25  3 */ (\rco[120]  ? (n137 ? n1043 : 1'b0) : 1'b0);
assign n4717 = /* LUT   27 10  3 */ (\rco[59]  ? (n3749 ? (\rco[0]  ? n1491 : 1'b0) : 1'b0) : 1'b0);
assign n4718 = /* LUT   13 27  2 */ (n1543 ? (n1558 ? n1390 : 1'b0) : 1'b0);
assign n4719 = /* LUT   15 13  1 */ n1777;
assign n4720 = /* LUT   20 20  4 */ n2764;
assign n4721 = /* LUT   23 18  7 */ n3257;
assign n4722 = /* LUT    5 12  4 */ n487;
assign n4723 = /* LUT   19 27  7 */ n2622;
assign n4724 = /* LUT   11 23  1 */ n1214;
assign n4725 = /* LUT   23 25  6 */ n3309;
assign n4726 = /* LUT    1 10  4 */ n17;
assign n4727 = /* LUT   10 21  2 */ n1059;
assign n4728 = /* LUT    9 11  0 */ n848;
assign n4729 = /* LUT   15 19  6 */ n1822;
assign n4730 = /* LUT   20 26  5 */ n2809;
assign n4731 = /* LUT   18 17  1 */ n1047;
assign n4732 = /* LUT    3 20  2 */ n343;
assign n4733 = /* LUT    2 20  4 */ n220;
assign n4734 = /* LUT   20 23  6 */ (n2003 ? (n2011 ? n2599 : 1'b0) : 1'b0);
assign n4735 = /* LUT   15 14  5 */ n1787;
assign n4736 = /* LUT   12 27  4 */ (n1272 ? (n1087 ? (n1244 ? !n1221 : 1'b1) : 1'b1) : 1'b1);
assign n4737 = /* LUT   11  8  5 */ n1127;
assign n4738 = /* LUT   29  5  5 */ n3822;
assign n4739 = /* LUT    4 10  2 */ n380;
assign n4740 = /* LUT   24 16  2 */ n3385;
assign n4741 = /* LUT   27 22  5 */ n3699;
assign n4742 = /* LUT   13 10  3 */ n1436;
assign n4743 = /* LUT    7 16  6 */ n748;
assign n4744 = /* LUT    9 21  4 */ n917;
assign n4745 = /* LUT   21 11  1 */ n2860;
assign n4746 = /* LUT   21  6  6 */ n2838;
assign n4747 = /* LUT   12 22  2 */ n1349;
assign n4748 = /* LUT   26 15  3 */ n3542;
assign n4749 = /* LUT   17  9  1 */ (n1934 ? (\rco[0]  ? (\rco[39]  ? n2269 : 1'b0) : 1'b0) : 1'b0);
assign n4750 = /* LUT   19 23  0 */ (n2173 ? (\rco[172]  ? (n2229 ? n2784 : 1'b0) : 1'b0) : 1'b0);
assign n4751 = /* LUT   10  9  4 */ n981;
assign n4752 = /* LUT   28 20  6 */ (\rco[153]  ? (\rco[0]  ? (n3240 ? n2574 : 1'b0) : 1'b0) : 1'b0);
assign n4753 = /* LUT   22 15  4 */ n3061;
assign n4754 = /* LUT    4 21  5 */ n451;
assign n4755 = /* LUT   13 28  3 */ n1563;
assign n4756 = /* LUT   27 11  0 */ (n3619 ? (n3525 ? (n3646 ? n3033 : 1'b0) : 1'b0) : 1'b0);
assign n4757 = /* LUT    6 10  4 */ n594;
assign n4758 = /* LUT   20 11  5 */ n2694;
assign n4759 = /* LUT   23 19  4 */ n3253;
assign n4760 = /* LUT    5 13  7 */ n498;
assign n4761 = /* LUT   19 24  6 */ n2601;
assign n4762 = /* LUT   11 20  0 */ n1194;
assign n4763 = /* LUT   29  9  6 */ n3830;
assign n4764 = /* LUT   17 27  5 */ n2192;
assign n4765 = /* LUT   28 23  0 */ n3810;
assign n4766 = /* LUT   10 20  1 */ n1048;
assign n4767 = /* LUT   15 16  7 */ n1799;
assign n4768 = /* LUT   21 15  6 */ (n1601 ? (n3069 ? (n1491 ? n1752 : 1'b0) : 1'b0) : 1'b0);
assign n4769 = /* LUT   20 25  4 */ n2801;
assign n1954 = /* LUT   15 15  6 */ (n1340 ? n1953 : 1'b0);
assign n461  = /* LUT    3 21  5 */ (n121 ? (n123 ? (\rco[0]  ? n244 : 1'b0) : 1'b0) : 1'b0);
assign n4771 = /* LUT   18 16  2 */ n2315;
assign n4772 = /* LUT    6  9  6 */ (n403 ? (n728 ? 1'b0 : (n277 ? n87 : 1'b0)) : 1'b0);
assign n4773 = /* LUT   20 22  5 */ n2780;
assign n4774 = /* LUT   12 26  7 */ n1254;
assign n4775 = /* LUT   17 24  1 */ n2166;
assign n4776 = /* LUT    4  9  3 */ n373;
assign n4777 = /* LUT   24 15  3 */ n3379;
assign n4778 = /* LUT   13 11  4 */ n1444;
assign n4779 = /* LUT    7 17  1 */ n751;
assign n4780 = /* LUT   21 12  0 */ n2872;
assign n4781 = /* LUT   14 26  3 */ n1713;
assign n4782 = /* LUT   12 21  3 */ n1343;
assign n4783 = /* LUT   17 10  0 */ n2278;
assign n4784 = /* LUT   20  4  1 */ (n2057 ? \rco[93]  : 1'b0);
assign n4785 = /* LUT   19 20  1 */ n2565;
assign n4786 = /* LUT   22 19  7 */ (n811 ? (n737 ? n2354 : 1'b0) : 1'b0);
assign n4787 = /* LUT   10  5  4 */ n969;
assign n4788 = /* LUT   24 18  7 */ n3413;
assign n4789 = /* LUT   22 14  3 */ n3053;
assign n4790 = /* LUT   27  8  1 */ (\rco[66]  ? (n3733 ? (\rco[0]  ? n1752 : 1'b0) : 1'b0) : 1'b0);
assign n4791 = /* LUT    3 17  2 */ n311;
assign n4792 = /* LUT   14 25  7 */ n795;
assign n4793 = /* LUT    6 21  5 */ (n338 ? (n781 ? (n779 ? n670 : 1'b0) : 1'b0) : 1'b0);
assign n4794 = /* LUT   17  4  3 */ n2034;
assign n4795 = /* LUT   23 16  5 */ (n1543 ? \rco[99]  : 1'b0);
assign n4796 = /* LUT   11 14  6 */ n1153;
assign n4797 = /* LUT   20  7  5 */ n2665;
assign n4798 = /* LUT    5 14  6 */ n505;
assign n4799 = /* LUT   20 10  6 */ n2858;
assign n4800 = /* LUT   11 21  7 */ n924;
assign n4801 = /* LUT   28 22  3 */ n3812;
assign n4802 = /* LUT   16 12  2 */ n1772;
assign n4803 = /* LUT   16 17  5 */ n1963;
assign n4804 = /* LUT   10 23  0 */ (\rco[99]  ? (n1091 ? 1'b0 : (n148 ? n1090 : 1'b0)) : 1'b0);
assign n4805 = /* LUT   13 15  1 */ n1470;
assign n3718 = /* LUT   27  6  0 */ (n3330 ? (n3455 ? n2676 : 1'b0) : 1'b0);
assign n4806 = /* LUT   30 12  1 */ n3894;
assign n4807 = /* LUT   15 17  0 */ n1806;
assign n4808 = /* LUT   18  6  4 */ n2234;
assign n4809 = /* LUT    7 21  6 */ n775;
assign n4810 = /* LUT    6  7  4 */ n586;
assign n4811 = /* LUT   18 19  3 */ n2341;
assign n4812 = /* LUT    3 18  4 */ n321;
assign n4813 = /* LUT   20 24  3 */ n2790;
assign n4814 = /* LUT   20 21  4 */ n2771;
assign n4815 = /* LUT   12 25  6 */ n1381;
assign n4816 = /* LUT    1 19  2 */ n105;
assign n4817 = /* LUT   17 25  2 */ n2177;
assign n4818 = /* LUT   23 13  0 */ n2729;
assign n4819 = /* LUT   10 25  3 */ n1082;
assign n4820 = /* LUT   24 14  0 */ n3374;
assign n4821 = /* LUT   27 20  7 */ n3681;
assign n4822 = /* LUT    4 19  6 */ (n438 ? (n121 ? \rco[123]  : 1'b0) : 1'b0);
assign n4823 = /* LUT   13 12  5 */ n1455;
assign n4824 = /* LUT   18  5  6 */ n2226;
assign n4825 = /* LUT    7 22  0 */ n550;
assign n4826 = /* LUT    9 23  2 */ n926;
assign n4827 = /* LUT   21 13  3 */ n2876;
assign n4828 = /* LUT   14 21  2 */ (\rco[110]  ? (n1845 ? (n1684 ? \rco[0]  : 1'b0) : 1'b0) : 1'b0);
assign n4829 = /* LUT   19 30  7 */ n2648;
assign n4830 = /* LUT    1 16  4 */ n94;
assign n4831 = /* LUT   19 21  6 */ n2583;
assign n4832 = /* LUT   11 17  4 */ n1171;
assign n4833 = /* LUT   10 11  6 */ n995;
assign n4834 = /* LUT   16  8  7 */ n1762;
assign n4835 = /* LUT   24 17  6 */ n3399;
assign n4836 = /* LUT   28  7  7 */ n3710;
assign n4837 = /* LUT   22  9  2 */ n2281;
assign n4838 = /* LUT   15 21  5 */ n1840;
assign n4839 = /* LUT   14 24  4 */ (n117 ? (n338 ? (n780 ? n121 : 1'b0) : 1'b0) : 1'b0);
assign n4840 = /* LUT   17  5  0 */ (n777 ? \rco[138]  : 1'b0);
assign n4841 = /* LUT    6 20  6 */ n665;
assign n4842 = /* LUT   23 17  2 */ n3235;
assign n4843 = /* LUT   11 15  5 */ n1157;
assign n4844 = /* LUT   26  6  6 */ n3478;
assign n4845 = /* LUT   11 18  6 */ n1184;
assign n4846 = /* LUT   29 11  0 */ n3847;
assign n4847 = /* LUT   28 21  2 */ n3792;
assign n4848 = /* LUT    4 12  1 */ n393;
assign n4849 = /* LUT   13 16  0 */ n1043;
assign n4850 = /* LUT   27  7  3 */ n3599;
assign n4851 = /* LUT   15 22  1 */ n1846;
assign n4852 = /* LUT   18  9  5 */ n2265;
assign n4853 = /* LUT    9 19  7 */ n792;
assign n4854 = /* LUT    3 19  7 */ n99;
assign n4855 = /* LUT    6 11  4 */ n613;
assign n4856 = /* LUT   12 24  1 */ n1367;
assign n4857 = /* LUT   26  5  0 */ n3480;
assign n4858 = /* LUT   14 10  0 */ n614;
assign n4859 = /* LUT   19 17  3 */ n2543;
assign n4860 = /* LUT   22 21  4 */ n3099;
assign n4861 = /* LUT   24 24  6 */ n3440;
assign n4862 = /* LUT    4 15  5 */ n416;
assign n4863 = /* LUT   10 24  0 */ n1231;
assign n4864 = /* LUT   24 13  1 */ n3361;
assign n4865 = /* LUT   27 21  0 */ n3240;
assign n4866 = /* LUT    4 18  5 */ n434;
assign n4867 = /* LUT   18  4  5 */ n2217;
assign n4868 = /* LUT   21 14  2 */ n2883;
assign n4869 = /* LUT    9 16  3 */ n877;
assign n4870 = /* LUT   14 20  1 */ n1676;
assign n4871 = /* LUT    5  8  7 */ n155;
assign n4872 = /* LUT   19 31  4 */ n2644;
assign n4873 = /* LUT    2 11  3 */ n170;
assign n4874 = /* LUT   23 21  7 */ n3277;
assign n4875 = /* LUT   19 18  7 */ n2560;
assign n4876 = /* LUT   10 10  1 */ n87;
assign n4877 = /* LUT   16 23  6 */ n1997;
assign n4878 = /* LUT   28  6  4 */ n3714;
assign n4879 = /* LUT   21 16  1 */ n2887;
assign n4880 = /* LUT   15 10  4 */ n1757;
assign n4881 = /* LUT   18 22  1 */ n2580;
assign n4882 = /* LUT   17  6  1 */ n2038;
assign n4883 = /* LUT    6 23  7 */ n693;
assign n4884 = /* LUT   20  8  0 */ (n2457 ? (n2671 ? (n2247 ? n2689 : 1'b0) : 1'b0) : 1'b0);
assign n4885 = /* LUT   12 28  6 */ n1399;
assign n4886 = /* LUT   23 22  3 */ n3281;
assign n1335 = /* LUT   11 19  5 */ (n465 ? (n913 ? (n365 ? n1038 : 1'b0) : 1'b0) : 1'b0);
assign n4887 = /* LUT   29 12  1 */ n3849;
assign n4888 = /* LUT   16 10  0 */ n1931;
assign n4889 = /* LUT   22 26  2 */ n3134;
assign n4890 = /* LUT   27 17  5 */ n3552;
assign n4891 = /* LUT    9  7  4 */ n826;
assign n4892 = /* LUT   13 17  3 */ n1486;
assign n4893 = /* LUT   15 23  2 */ n1853;
assign n4894 = /* LUT   18  8  6 */ n2267;
assign n4895 = /* LUT   18 21  5 */ n2353;
assign n4896 = /* LUT    3 16  6 */ n309;
assign n4897 = /* LUT   14  5  1 */ n1571;
assign n4898 = /* LUT   19 14  2 */ n2514;
assign n4899 = /* LUT   22 20  7 */ n2918;
assign n4900 = /* LUT   10 14  6 */ n1014;
assign n4901 = /* LUT    4 14  6 */ n103;
assign n4902 = /* LUT   22 25  4 */ n3128;
assign n4903 = /* LUT   10 27  1 */ n1093;
assign n4904 = /* LUT   24 12  6 */ n3358;
assign n4905 = /* LUT   16 24  4 */ (\rco[118]  ? (n2175 ? 1'b0 : (n365 ? n1038 : 1'b0)) : 1'b0);
assign n4906 = /* LUT   27 18  1 */ n3657;
assign n4907 = /* LUT   28 10  1 */ n3741;
assign n4908 = /* LUT    4 17  4 */ n429;
assign n4909 = /* LUT   13 14  7 */ n1468;
assign n4910 = /* LUT   18  7  4 */ n2244;
assign n4911 = /* LUT    9 17  0 */ n889;
assign n4912 = /* LUT   26 22  0 */ n3573;
assign n4913 = /* LUT   15  5  2 */ n1726;
assign n4914 = /* LUT   14 23  0 */ (\rco[99]  ? (\rco[0]  ? (n335 ? n780 : 1'b0) : 1'b0) : 1'b0);
assign n4915 = /* LUT   20 12  5 */ n2702;
assign n4916 = /* LUT   19 28  5 */ n2625;
assign n4917 = /* LUT   19 19  4 */ (n2044 ? (n1710 ? (\rco[0]  ? \rco[162]  : 1'b0) : 1'b0) : 1'b0);
assign n4918 = /* LUT   10 13  0 */ (n817 ? (n912 ? (\rco[0]  ? \rco[99]  : 1'b0) : 1'b0) : 1'b0);
assign n4919 = /* LUT   28  5  5 */ n3709;
assign n4920 = /* LUT   22 11  0 */ (n2494 ? (n2859 ? (\rco[53]  ? n2857 : 1'b0) : 1'b0) : 1'b0);
assign n4921 = /* LUT   21 17  2 */ (\rco[59]  ? n2728 : 1'b0);
assign n4922 = /* LUT   30 10  4 */ n3888;
assign n4923 = /* LUT   15 11  7 */ n1754;
assign n341  = /* LUT    2 19  4 */ (n328 ? (n340 ? (n246 ? n118 : 1'b0) : 1'b0) : 1'b0);
assign n4925 = /* LUT   18 25  0 */ n1551;
assign n4926 = /* LUT   15  6  4 */ n1736;
assign n4927 = /* LUT   17  7  6 */ n2051;
assign n4928 = /* LUT    6 22  0 */ n685;
assign n4929 = /* LUT   20 15  1 */ n2722;
assign n4930 = /* LUT   23 23  0 */ n2539;
assign n4931 = /* LUT   11 13  3 */ n1142;
assign n4932 = /* LUT   11 16  4 */ n1162;
assign n4933 = /* LUT   16  9  1 */ n1923;
assign n4934 = /* LUT   13  7  5 */ n1427;
assign n4935 = /* LUT   13 18  2 */ n1493;
assign n4936 = /* LUT   27  5  5 */ n3589;
assign n4937 = /* LUT   18 11  7 */ (n2306 ? (\rco[41]  ? \rco[0]  : 1'b0) : 1'b0);
assign n4938 = /* LUT   15 20  3 */ n1829;
assign n4939 = /* LUT   18 20  6 */ (n809 ? (n1151 ? (\rco[0]  ? \rco[153]  : 1'b0) : 1'b0) : 1'b0);
assign n4940 = /* LUT   26  7  2 */ n3482;
assign n4941 = /* LUT    2 14  1 */ n187;
assign n4942 = /* LUT   16  7  0 */ n587;
assign n4943 = /* LUT   19 15  1 */ n2718;
assign n4944 = /* LUT   23  5  4 */ n3153;
assign n4945 = /* LUT   22 23  6 */ (\rco[172]  ? (n982 ? (n2539 ? \rco[0]  : 1'b0) : 1'b0) : 1'b0);
assign n4946 = /* LUT   24 22  4 */ n3428;
assign n4947 = /* LUT    4 13  7 */ n401;
assign n4948 = /* LUT   22 24  7 */ n3120;
assign n4949 = /* LUT   10 26  6 */ (\rco[99]  ? (n1246 ? \rco[0]  : 1'b0) : 1'b0);
assign n4950 = /* LUT   24 11  7 */ (n3348 ? (n3468 ? (n1752 ? \rco[0]  : 1'b0) : 1'b0) : 1'b0);
assign n4951 = /* LUT   27 19  2 */ n3668;
assign n4952 = /* LUT   28  9  0 */ n3739;
assign n4953 = /* LUT    4 16  3 */ n422;
assign n4954 = /* LUT    9 18  1 */ n890;
assign n4955 = /* LUT   26  9  1 */ n3498;
assign n4956 = /* LUT   29 17  0 */ n3857;
assign n4957 = /* LUT   14 22  7 */ n1693;
assign n4958 = /* LUT   17  3  3 */ n2027;
assign n4959 = /* LUT    6 18  5 */ n653;
assign n4960 = /* LUT    5 10  5 */ n478;
assign n4961 = /* LUT   19 29  2 */ (\rco[183]  ? (n1541 ? n1816 : 1'b0) : 1'b0);
assign n4962 = /* LUT   23 27  5 */ n3317;
assign n4963 = /* LUT   19 16  5 */ (n812 ? (n2333 ? (n880 ? n2537 : 1'b0) : 1'b0) : 1'b0);
assign n4964 = /* LUT   23  6  6 */ n3164;
assign n4965 = /* LUT   11 28  7 */ n1273;
assign n4966 = /* LUT   10 12  3 */ n999;
assign n4967 = /* LUT   24 25  2 */ n3447;
assign n4968 = /* LUT   16 21  4 */ n1990;
assign n4969 = /* LUT   16 26  5 */ n2185;
assign n4970 = /* LUT   21 18  3 */ n2906;
assign n4971 = /* LUT    9 28  0 */ n958;
assign n4972 = /* LUT   15  8  6 */ n1747;
assign n4973 = /* LUT    3 22  7 */ n355;
assign n4974 = /* LUT    2 18  3 */ n211;
assign n4975 = /* LUT   21  7  7 */ (n3009 ? \rco[44]  : 1'b0);
assign n4976 = /* LUT   15  7  7 */ (\rco[83]  ? (\rco[0]  ? (n1583 ? n614 : 1'b0) : 1'b0) : 1'b0);
assign n4977 = /* LUT   18 24  3 */ n2372;
assign n4978 = /* LUT    6 17  1 */ n757;
assign n4979 = /* LUT   20 14  2 */ n2705;
assign n4980 = /* LUT   23 20  1 */ n3263;
assign n3458 = /* LUT   24  7  2 */ (n3456 ? (n3457 ? (n3326 ? \rco[0]  : 1'b0) : 1'b0) : 1'b0);
assign n4982 = /* LUT    9 14  7 */ n856;
assign n4983 = /* LUT   13 19  5 */ (\rco[99]  ? (n1674 ? 1'b0 : n1671) : 1'b0);
assign n4984 = /* LUT   18 10  0 */ n2279;
assign n4985 = /* LUT   18 23  7 */ n2159;
assign n4986 = /* LUT   12 29  2 */ n1406;
assign n4987 = /* LUT   19 25  7 */ n2610;
assign n4988 = /* LUT   14  7  3 */ n1587;
assign n4989 = /* LUT   16  6  3 */ n1899;
assign n4990 = /* LUT   19 12  0 */ n2503;
assign n4991 = /* LUT   23 10  5 */ n3189;
assign n4992 = /* LUT   22 22  1 */ n2949;
assign n4993 = /* LUT   24 21  5 */ n3423;
assign n4994 = /* LUT   22 27  6 */ n3148;
assign n4995 = /* LUT   24 10  4 */ n3343;
assign n4996 = /* LUT   28  8  7 */ n3618;
assign n4997 = /* LUT   13  5  2 */ n1414;
assign n4998 = /* LUT    3  9  0 */ n376;
assign n4999 = /* LUT   12 19  1 */ n1328;
assign n5000 = /* LUT   26  8  2 */ n3491;
assign n5001 = /* LUT   14 17  6 */ n1658;
assign n5002 = /* LUT   17 12  2 */ n2078;
assign n2813 = /* LUT   19 26  3 */ (\rco[145]  ? (n2574 ? (n817 ? n1710 : 1'b0) : 1'b0) : 1'b0);
assign n5003 = /* LUT   23 24  4 */ n3299;
assign n5004 = /* LUT    2 12  6 */ n183;
assign n5005 = /* LUT   23  7  5 */ n3170;
assign n5006 = /* LUT   10 15  2 */ n1021;
assign n5007 = /* LUT   16 20  3 */ n1976;
assign n5008 = /* LUT   16 25  4 */ n2006;
assign n5009 = /* LUT   21 24  5 */ n2957;
assign n5010 = /* LUT   21 19  4 */ n2908;
assign n5011 = /* LUT   13 23  2 */ n1525;
assign n5012 = /* LUT   27 14  3 */ n3643;
assign n5013 = /* LUT   18 14  5 */ n2305;
assign n5014 = /* LUT    2 21  2 */ n228;
assign n5015 = /* LUT   18 27  2 */ n2394;
assign n5016 = /* LUT    6 16  2 */ n639;
assign n5017 = /* LUT   20 13  3 */ (n2510 ? !n2881 : 1'b1);
assign n5018 = /* LUT    4 11  4 */ n390;
assign n5019 = /* LUT   22 18  6 */ n3086;
assign n5020 = /* LUT   22  7  1 */ n2998;
assign n1176 = /* LUT   10 17  2 */ (\rco[0]  ? (n1032 ? (n1031 ? !n989 : 1'b1) : 1'b1) : 1'b1);
assign n5022 = /* LUT    9 15  0 */ n880;
assign n5023 = /* LUT   24  6  1 */ n3321;
assign n5024 = /* LUT   28 12  4 */ n3756;
assign n5025 = /* LUT   13 20  4 */ n1506;
assign n5026 = /* LUT   18 13  1 */ n2295;
assign n5027 = /* LUT   14 13  5 */ n1459;
assign n5028 = /* LUT   14  6  4 */ n1580;
assign n5029 = /* LUT   16  5  2 */ n1889;
assign n5030 = /* LUT   17 19  0 */ n2344;
assign n5031 = /* LUT   23 11  6 */ n3195;
assign n5032 = /* LUT   11 25  5 */ n1235;
assign n5033 = /* LUT   22 17  0 */ n2552;
assign n5034 = /* LUT   24 20  2 */ n3407;
assign n5035 = /* LUT   10 28  4 */ n1104;
assign n5036 = /* LUT   24  9  5 */ n3336;
assign n5037 = /* LUT   13  6  3 */ n1417;
assign n564  = /* LUT    4 22  1 */ (n463 ? (n120 ? n226 : 1'b0) : 1'b0);
assign n5038 = /* LUT   21 23  1 */ n2943;
assign n5039 = /* LUT   15 13  6 */ n1629;
assign n5040 = /* LUT   12 18  2 */ n1321;
assign n5041 = /* LUT   26 11  3 */ n3528;
assign n5042 = /* LUT   29 19  6 */ n3867;
assign n5043 = /* LUT   14 16  5 */ n1650;
assign n5044 = /* LUT   17 13  1 */ n2086;
assign n5045 = /* LUT    5 12  3 */ n400;
assign n5046 = /* LUT   19 27  0 */ n1816;
assign n5047 = /* LUT   23 25  3 */ n3306;
assign n5048 = /* LUT   11 26  1 */ n1236;
assign n5049 = /* LUT    7  2  5 */ (\rco[162]  ? n807 : 1'b0);
assign n5050 = /* LUT    9 11  5 */ n846;
assign n5051 = /* LUT   21 25  6 */ n2969;
assign n5052 = /* LUT    7  9  4 */ n721;
assign n5053 = /* LUT   21 20  5 */ n2922;
assign n5054 = /* LUT   13 24  3 */ (n1337 ? (n335 ? \rco[99]  : 1'b0) : 1'b0);
assign n5055 = /* LUT   15 14  0 */ n1130;
assign n5056 = /* LUT    3 20  5 */ n346;
assign n5057 = /* LUT    2 20  1 */ n217;
assign n5058 = /* LUT   18 17  4 */ n2328;
assign n5059 = /* LUT   18 26  5 */ n2389;
assign n766  = /* LUT    6 19  3 */ (n326 ? (n244 ? (n327 ? n123 : 1'b0) : 1'b0) : 1'b0);
assign n5061 = /* LUT   11  8  0 */ n1128;
assign n5062 = /* LUT   28 19  0 */ n3241;
assign n5063 = /* LUT   19  9  4 */ n2474;
assign n5064 = /* LUT    4 10  7 */ n385;
assign n5065 = /* LUT   24 16  7 */ n3390;
assign n5066 = /* LUT   22  6  6 */ n2995;
assign n5067 = /* LUT   10 16  1 */ n1023;
assign n5068 = /* LUT   13 10  6 */ n1440;
assign n5069 = /* LUT   13 21  7 */ n1686;
assign n5070 = /* LUT   31 22  7 */ (\rco[183]  ? (n3124 ? n2796 : 1'b0) : 1'b0);
assign n5071 = /* LUT   18 12  2 */ n2287;
assign n5072 = /* LUT   21  6  1 */ n2833;
assign n5073 = /* LUT   11  6  3 */ n1120;
assign n5074 = /* LUT   14 12  6 */ (n614 ? (n1603 ? n1583 : 1'b0) : 1'b0);
assign n2787 = /* LUT   19 23  5 */ (n1340 ? (n1710 ? (n768 ? 1'b1 : !n1375) : 1'b1) : 1'b1);
assign n5076 = /* LUT   19 10  6 */ n2485;
assign n5077 = /* LUT    4 21  0 */ n452;
assign n5078 = /* LUT    7 13  1 */ (\rco[153]  ? n811 : 1'b0);
assign n5079 = /* LUT   21  8  0 */ n3010;
assign n5080 = /* LUT   26 17  5 */ n3550;
assign n5081 = /* LUT   12 17  3 */ n1314;
assign n5082 = /* LUT   26 10  4 */ n3510;
assign n5083 = /* LUT   18 30  2 */ n2418;
assign n5084 = /* LUT   14 19  4 */ n1667;
assign n5085 = /* LUT   17 14  0 */ (n1950 ? (n2030 ? n2095 : 1'b0) : 1'b0);
assign n5086 = /* LUT   29 20  7 */ n3874;
assign n5087 = /* LUT    5 13  0 */ n494;
assign n5088 = /* LUT   19 24  1 */ n2594;
assign n5089 = /* LUT   11 27  2 */ n1248;
assign n5090 = /* LUT   16 18  1 */ n1971;
assign n5091 = /* LUT    1 11  0 */ (\rco[0]  ? !n56 : 1'b0);
assign n5092 = /* LUT   21 26  7 */ (n3114 ? 1'b0 : (n3142 ? (n2784 ? n2627 : 1'b0) : 1'b0));
assign n5093 = /* LUT   21 21  6 */ n2931;
assign n5094 = /* LUT   13 25  0 */ (\rco[198]  ? n1706 : 1'b0);
assign n5095 = /* LUT   27 12  1 */ n3631;
assign n5096 = /* LUT   15 15  3 */ (\rco[99]  ? (n1952 ? 1'b0 : n912) : 1'b0);
assign n459  = /* LUT    3 21  2 */ (n129 ? (n457 ? n121 : 1'b0) : 1'b0);
assign n5098 = /* LUT   18 16  7 */ n2320;
assign n5099 = /* LUT   18 29  4 */ n2411;
assign n5100 = /* LUT   28 18  3 */ n3775;
assign n5101 = /* LUT   19  6  5 */ n2447;
assign n5102 = /* LUT    4  9  6 */ n378;
assign n5103 = /* LUT   22 28  4 */ (n1043 ? \rco[120]  : 1'b0);
assign n5104 = /* LUT   10  6  7 */ n973;
assign n5105 = /* LUT   24 15  6 */ n3382;
assign n1188 = /* LUT   10 19  0 */ (n114 ? (\rco[0]  ? (n696 ? !n117 : 1'b1) : 1'b1) : 1'b1);
assign n5107 = /* LUT    9  9  2 */ n828;
assign n5108 = /* LUT   13 11  1 */ n1441;
assign n5109 = /* LUT   13 22  6 */ n1523;
assign n5110 = /* LUT   18 15  3 */ n2310;
assign n5111 = /* LUT   26 14  1 */ n3648;
assign n5112 = /* LUT   14 15  7 */ n1653;
assign n5113 = /* LUT    2  9  4 */ n158;
assign n5114 = /* LUT   20  4  6 */ n2655;
assign n5115 = /* LUT   19 20  4 */ n2568;
assign n5116 = /* LUT   19 11  5 */ n2490;
assign n5117 = /* LUT   23  9  0 */ n1934;
assign n3261 = /* LUT   22 19  2 */ (n809 ? (n3260 ? 1'b0 : (n738 ? n1979 : 1'b0)) : 1'b0);
assign n5118 = /* LUT   10  5  3 */ n968;
assign n5119 = /* LUT   24 18  0 */ n3412;
assign n5120 = /* LUT   21  9  3 */ n2847;
assign n5121 = /* LUT    9 27  2 */ n1099;
assign n5122 = /* LUT   12 11  5 */ (\rco[23]  ? n813 : 1'b0);
assign n5123 = /* LUT   26 16  6 */ n3651;
assign n5124 = /* LUT    3 17  7 */ n425;
assign n5125 = /* LUT   12 16  4 */ n1307;
assign n5126 = /* LUT   14 25  2 */ n1702;
assign n5127 = /* LUT   26 13  5 */ n3531;
assign n5128 = /* LUT   17 15  7 */ n2104;
assign n5129 = /* LUT   29 21  4 */ n3877;
assign n5130 = /* LUT   20  7  0 */ n2457;
assign n5131 = /* LUT    5 14  1 */ n504;
assign n5132 = /* LUT   11 24  3 */ n1225;
assign n5133 = /* LUT   16 17  0 */ n1959;
assign n5134 = /* LUT   21 27  0 */ n2977;
assign n5135 = /* LUT   13 15  6 */ n1475;
assign n5136 = /* LUT   27  6  7 */ n3595;
assign n5137 = /* LUT    7 15  6 */ (\rco[0]  ? (n812 ? \rco[25]  : 1'b0) : 1'b0);
assign n5138 = /* LUT    9 24  4 */ n935;
assign n5139 = /* LUT   13 26  1 */ n1544;
assign n5140 = /* LUT   21 22  7 */ n2783;
assign n5141 = /* LUT   18 19  6 */ n2346;
assign n5142 = /* LUT    3 18  3 */ n320;
assign n5143 = /* LUT   18 28  7 */ n2406;
assign n5144 = /* LUT    1 19  7 */ n110;
assign n5145 = /* LUT   28 17  2 */ n3767;
assign n5146 = /* LUT   16 15  3 */ n1945;
assign n5147 = /* LUT    5 16  5 */ n520;
assign n5148 = /* LUT   19  7  6 */ n2459;
assign n5149 = /* LUT   23 13  5 */ n3212;
assign n5150 = /* LUT   10 25  6 */ n1086;
assign n5151 = /* LUT   24 14  5 */ n3373;
assign n5152 = /* LUT   10 18  7 */ n1034;
assign n5153 = /* LUT    9 10  3 */ n836;
assign n5154 = /* LUT   13 12  0 */ n1454;
assign n5155 = /* LUT   15 18  1 */ n1808;
assign n5156 = /* LUT   20 27  2 */ n2815;
assign n5157 = /* LUT   12 20  1 */ (n243 ? (n361 ? n780 : 1'b0) : 1'b0);
assign n5158 = /* LUT   14 14  0 */ n1637;
assign n5159 = /* LUT   17 11  4 */ n2071;
assign n5160 = /* LUT    1 16  3 */ n90;
assign n5161 = /* LUT   19 21  3 */ n2578;
assign n5162 = /* LUT   19  8  4 */ n2464;
assign n5163 = /* LUT   23 14  1 */ n3217;
assign n5164 = /* LUT   24 17  1 */ n3394;
assign n5165 = /* LUT   28  7  2 */ n3720;
assign n5166 = /* LUT    3 14  5 */ (n287 ? (n87 ? (n289 ? !n31 : 1'b1) : 1'b1) : 1'b1);
assign n5167 = /* LUT    7 19  3 */ n761;
assign n1057 = /* LUT    9 20  3 */ (n465 ? (n696 ? (\rco[0]  ? !n114 : 1'b1) : 1'b1) : 1'b1);
assign n5169 = /* LUT   21 10  2 */ (n1934 ? (n2269 ? (n2306 ? !n1933 : 1'b1) : 1'b1) : 1'b1);
assign n5170 = /* LUT   27  9  3 */ n3612;
assign n5171 = /* LUT   17  5  5 */ (\rco[172]  ? n982 : 1'b0);
assign n5172 = /* LUT   12 23  5 */ n1362;
assign n1874 = /* LUT   14 24  1 */ (n1710 ? (n1873 ? (n1697 ? n1698 : 1'b0) : 1'b0) : 1'b0);
assign n5174 = /* LUT   26 12  6 */ n3622;
assign n5175 = /* LUT   17  8  6 */ (n2260 ? (n2240 ? \rco[0]  : 1'b0) : 1'b0);
assign n5176 = /* LUT    2  7  3 */ n150;
assign n5177 = /* LUT    4 12  6 */ n398;
assign n5178 = /* LUT   22 12  1 */ n3036;
assign n5179 = /* LUT   10 22  4 */ (\rco[0]  ? (n1213 ? (n114 ? n696 : 1'b0) : 1'b0) : 1'b0);
assign n5180 = /* LUT   21 28  1 */ n2979;
assign n5181 = /* LUT   13 16  7 */ n1483;
assign n5182 = /* LUT   27  7  4 */ n3600;
assign n5183 = /* LUT    9 25  7 */ n941;
assign n5184 = /* LUT   27 10  7 */ (\rco[0]  ? (n3528 ? (\rco[59]  ? n1491 : 1'b0) : 1'b0) : 1'b0);
assign n5185 = /* LUT   13 27  6 */ n1556;
assign n5186 = /* LUT   18 18  1 */ n2334;
assign n5187 = /* LUT    3 19  0 */ (n327 ? (n114 ? (n244 ? n123 : 1'b0) : 1'b0) : 1'b0);
assign n5188 = /* LUT   20 20  0 */ n2766;
assign n5189 = /* LUT   23 18  3 */ n3244;
assign n5190 = /* LUT   14 10  5 */ n1608;
assign n5191 = /* LUT    1  7  7 */ (n154 ? \rco[21]  : 1'b0);
assign n5192 = /* LUT    5 17  6 */ n530;
assign n5193 = /* LUT    4 15  0 */ n298;
assign n5194 = /* LUT   10 24  5 */ n1076;
assign n5195 = /* LUT   24 13  4 */ n3364;
assign n5196 = /* LUT   10 21  6 */ n1064;
assign n5197 = /* LUT   13 13  3 */ n1457;
assign n5198 = /* LUT   15 19  2 */ n1818;
assign n5199 = /* LUT   20 26  1 */ n2805;
assign n5200 = /* LUT   12 27  0 */ (n1272 ? (n1543 ? (n1244 ? \rco[99]  : 1'b0) : 1'b0) : 1'b0);
assign n5201 = /* LUT   17 20  5 */ n2140;
assign n5202 = /* LUT    2 11  6 */ n173;
assign n5203 = /* LUT   19 18  2 */ n2555;
assign n5204 = /* LUT   23 15  2 */ n3223;
assign n5205 = /* LUT   28  6  1 */ n3711;
assign n5206 = /* LUT   27 22  1 */ n3695;
assign n5207 = /* LUT    3 15  6 */ n300;
assign n5208 = /* LUT   21 16  4 */ n2890;
assign n5209 = /* LUT    7 16  2 */ n742;
assign n5210 = /* LUT    9 21  0 */ n365;
assign n5211 = /* LUT   21 11  5 */ n2863;
assign n3664 = /* LUT   26 18  0 */ (n2124 ? (n3555 ? \rco[23]  : 1'b0) : 1'b0);
assign n5212 = /* LUT   18 22  6 */ n2357;
assign n5213 = /* LUT   17  6  4 */ n2043;
assign n5214 = /* LUT   12 22  6 */ n1354;
assign n2272 = /* LUT   17  9  5 */ (n2266 ? (n2057 ? (n2236 ? !\rco[0]  : 1'b1) : 1'b1) : 1'b1);
assign n5216 = /* LUT   10  9  0 */ n987;
assign n5217 = /* LUT   28 20  2 */ (\rco[153]  ? (n3876 ? (\rco[0]  ? n2574 : 1'b0) : 1'b0) : 1'b0);
assign n5218 = /* LUT   22 26  7 */ n3139;
assign n5219 = /* LUT   22 15  0 */ n3063;
assign n5220 = /* LUT    7  6  1 */ n706;
assign n5221 = /* LUT    9  7  1 */ n717;
assign n5222 = /* LUT   13 17  4 */ n1487;
assign n5223 = /* LUT    9 26  6 */ n955;
assign n5224 = /* LUT   13 28  7 */ n1407;
assign n5225 = /* LUT   27 11  4 */ n3626;
assign n5226 = /* LUT   18 21  0 */ n2355;
assign n5227 = /* LUT    3 16  1 */ n303;
assign n5228 = /* LUT    6 10  0 */ n596;
assign n2866 = /* LUT   20 11  1 */ (n2416 ? n2865 : 1'b0);
assign n5229 = /* LUT   23 19  0 */ n1409;
assign n5230 = /* LUT   14  5  4 */ n1574;
assign n5231 = /* LUT   29  9  2 */ (n3330 ? \rco[74]  : 1'b0);
assign n5232 = /* LUT   17 27  1 */ n2188;
assign n5233 = /* LUT   28 23  4 */ n2796;
assign n5234 = /* LUT   19  5  0 */ n2441;
assign n514  = /* LUT    4 14  3 */ (n386 ? (n513 ? 1'b0 : (n376 ? \rco[9]  : 1'b0)) : 1'b0);
assign n5235 = /* LUT   22 25  3 */ n3127;
assign n5236 = /* LUT   10 27  4 */ n1096;
assign n5237 = /* LUT   24 12  3 */ n3355;
assign n5238 = /* LUT   10 20  5 */ n1052;
assign n5239 = /* LUT   13 14  2 */ n1463;
assign n5240 = /* LUT   15 16  3 */ n1795;
assign n3067 = /* LUT   21 15  2 */ (n2602 ? 1'b1 : (n982 ? (n2539 ? !n3066 : 1'b1) : 1'b1));
assign n5242 = /* LUT   20 25  0 */ n2803;
assign n5243 = /* LUT   26 22  5 */ n3574;
assign n5244 = /* LUT   15  5  7 */ n1895;
assign n5245 = /* LUT   12 26  3 */ n1387;
assign n5246 = /* LUT   14  8  2 */ n1594;
assign n5247 = /* LUT    2 10  1 */ n165;
assign n5248 = /* LUT    1 18  1 */ n98;
assign n5249 = /* LUT   19 19  1 */ (n1151 ? (n2758 ? (n2344 ? n809 : 1'b0) : 1'b0) : 1'b0);
assign n5250 = /* LUT   17 21  6 */ n2149;
assign n5251 = /* LUT   17 24  5 */ n2170;
assign n5252 = /* LUT   23 12  3 */ n3202;
assign n5253 = /* LUT   28  5  0 */ n3596;
assign n3815 = /* LUT   27 23  2 */ (n2797 ? (n3814 ? 1'b0 : n2603) : 1'b0);
assign n5254 = /* LUT    3 12  7 */ n166;
assign n5255 = /* LUT   21 17  7 */ n2900;
assign n5256 = /* LUT    7 17  5 */ n755;
assign n5257 = /* LUT    9 22  1 */ n923;
assign n5258 = /* LUT   21 12  4 */ n2870;
assign n5259 = /* LUT   12  8  0 */ n1282;
assign n5260 = /* LUT   26 21  1 */ n3562;
assign n5261 = /* LUT   15  6  3 */ n1735;
assign n5262 = /* LUT   17  7  3 */ n2048;
assign n5263 = /* LUT   12 21  7 */ n1341;
assign n5264 = /* LUT   18 25  7 */ n2382;
assign n5265 = /* LUT   17 10  4 */ n2062;
assign n5266 = /* LUT    9 32  7 */ (n803 ? \rco[106]  : 1'b0);
assign n5267 = /* LUT    1 12  5 */ n50;
assign n5268 = /* LUT   22 14  7 */ n3215;
assign n5269 = /* LUT    7  7  2 */ n712;
assign n5270 = /* LUT   13 18  5 */ n1496;
assign n5271 = /* LUT   27  5  2 */ n3586;
assign n5272 = /* LUT   27  8  5 */ n3608;
assign n2575 = /* LUT   18 20  3 */ (n1340 ? (n768 ? 1'b0 : (\rco[23]  ? !n1621 : 1'b0)) : 1'b0);
assign n5273 = /* LUT    6 21  1 */ n686;
assign n5274 = /* LUT   20 10  2 */ n2684;
assign n5275 = /* LUT   23 16  1 */ n2321;
assign n5276 = /* LUT   11 14  2 */ n1147;
assign n5277 = /* LUT    2 14  6 */ n192;
assign n5278 = /* LUT   16  7  7 */ n1913;
assign n5279 = /* LUT   29 10  3 */ n3836;
assign n5280 = /* LUT   28 22  7 */ n3804;
assign n5281 = /* LUT   16 12  6 */ n1940;
assign n5282 = /* LUT    5 19  0 */ n544;
assign n5283 = /* LUT    4 13  2 */ (n291 ? (n502 ? (n500 ? n103 : 1'b0) : 1'b0) : 1'b0);
assign n5284 = /* LUT   22 24  0 */ n3122;
assign n1245 = /* LUT   10 26  3 */ (n1221 ? (n1087 ? n1090 : 1'b0) : 1'b0);
assign n3465 = /* LUT   24 11  2 */ (n3050 ? (n2728 ? (n2729 ? n2740 : 1'b0) : 1'b0) : 1'b0);
assign n5285 = /* LUT   10 23  4 */ (n148 ? !n803 : 1'b1);
assign n5286 = /* LUT   15 17  4 */ n1804;
assign n5287 = /* LUT   18  6  0 */ n2237;
assign n5288 = /* LUT    7 21  2 */ n771;
assign n5289 = /* LUT    6  7  0 */ n576;
assign n5290 = /* LUT   20 24  7 */ n2794;
assign n5291 = /* LUT   26  9  4 */ n3501;
assign n5292 = /* LUT   12 25  2 */ n1377;
assign n5293 = /* LUT   14 11  3 */ n1614;
assign n5294 = /* LUT    2 13  0 */ n186;
assign n5295 = /* LUT   17 22  7 */ n2158;
assign n2731 = /* LUT   19 16  0 */ (n2124 ? (n1950 ? (n2521 ? n2122 : 1'b0) : 1'b0) : 1'b0);
assign n5296 = /* LUT   17 25  6 */ n2181;
assign n5297 = /* LUT   27 20  3 */ n3783;
assign n5298 = /* LUT    4 19  2 */ (n336 ? (n327 ? (\rco[127]  ? n326 : 1'b0) : 1'b0) : 1'b0);
assign n5299 = /* LUT    3 13  0 */ (n386 ? (\rco[13]  ? (\rco[0]  ? n376 : 1'b0) : 1'b0) : 1'b0);
assign n5300 = /* LUT   21 18  6 */ n2904;
assign n5301 = /* LUT   22 10  4 */ n3025;
assign n5302 = /* LUT    7 22  4 */ n786;
assign n5303 = /* LUT    9 23  6 */ n930;
assign n5304 = /* LUT   21 13  7 */ n2878;
assign n5305 = /* LUT   12 15  1 */ n1296;
assign n5306 = /* LUT   26 20  2 */ n3679;
assign n5307 = /* LUT   15  7  0 */ (n587 ? (\rco[83]  ? (n1738 ? n1623 : 1'b0) : 1'b0) : 1'b0);
assign n5308 = /* LUT   18 24  4 */ n2373;
assign n5309 = /* LUT   19 30  3 */ n2636;
assign n5310 = /* LUT   11 17  0 */ n1173;
assign n5311 = /* LUT   10 11  2 */ (\rco[99]  ? (n1136 ? (n912 ? \rco[0]  : 1'b0) : 1'b0) : 1'b0);
assign n5312 = /* LUT   16  8  3 */ n1917;
assign n5313 = /* LUT    1 13  6 */ n66;
assign n5314 = /* LUT   22  9  6 */ n3019;
assign n1673 = /* LUT   13 19  2 */ (n777 ? (n667 ? (\rco[0]  ? !n668 : 1'b1) : 1'b1) : 1'b1);
assign n5316 = /* LUT   15 21  1 */ n1836;
assign n5317 = /* LUT   20 28  4 */ n2826;
assign n5318 = /* LUT   18 23  2 */ n2363;
assign n5319 = /* LUT    6 20  2 */ n661;
assign n2853 = /* LUT   20  9  3 */ (n2680 ? (n2269 ? (n2510 ? !n1934 : 1'b1) : 1'b1) : 1'b1);
assign n5321 = /* LUT   23 17  6 */ n3239;
assign n5322 = /* LUT   11 15  1 */ (\rco[145]  ? (\rco[0]  ? (n736 ? n817 : 1'b0) : 1'b0) : 1'b0);
assign n5323 = /* LUT   26  6  2 */ n3474;
assign n5324 = /* LUT   14  7  6 */ n1591;
assign n5325 = /* LUT   16  6  4 */ n1900;
assign n5326 = /* LUT   29 11  4 */ n3842;
assign n5327 = /* LUT   28 21  6 */ n3796;
assign n5328 = /* LUT   19  3  2 */ n2428;
assign n5329 = /* LUT   22 27  1 */ n3143;
assign n5330 = /* LUT   10 29  2 */ n1111;
assign n5331 = /* LUT   24 10  1 */ n3340;
assign n5332 = /* LUT    3  9  5 */ n256;
assign n5333 = /* LUT   15 22  5 */ n1850;
assign n5334 = /* LUT   18  9  1 */ n2261;
assign n5335 = /* LUT    7 26  3 */ n798;
assign n5336 = /* LUT    9 19  3 */ n903;
assign n5337 = /* LUT   12 19  4 */ n1331;
assign n5338 = /* LUT   26  8  7 */ n3496;
assign n5339 = /* LUT   12 24  5 */ n1371;
assign n5340 = /* LUT   17 23  0 */ n2162;
assign n5341 = /* LUT    2 12  3 */ n178;
assign n5342 = /* LUT   22 21  0 */ n3102;
assign n5343 = /* LUT   24 24  2 */ n3300;
assign n5344 = /* LUT   27 21  4 */ n3690;
assign n5345 = /* LUT    4 18  1 */ n437;
assign n5346 = /* LUT    3 10  1 */ n262;
assign n5347 = /* LUT   13 23  7 */ n1530;
assign n5348 = /* LUT   27 14  6 */ n3538;
assign n5349 = /* LUT    9 16  7 */ n879;
assign n5350 = /* LUT   12 14  2 */ n1289;
assign n5351 = /* LUT   26 23  3 */ n3578;
assign n5352 = /* LUT   18 27  5 */ n2397;
assign n5353 = /* LUT   19 31  0 */ n2627;
assign n5354 = /* LUT   23 21  3 */ n3273;
assign n5355 = /* LUT   16 23  2 */ n1992;
assign n5356 = /* LUT    1 14  7 */ n91;
assign n5357 = /* LUT   22  7  4 */ n3001;
assign n5358 = /* LUT   22  8  5 */ n3012;
assign n5359 = /* LUT   13 20  3 */ n1505;
assign n5360 = /* LUT   15 10  0 */ n1768;
assign n5361 = /* LUT   20 19  5 */ n2753;
assign n5362 = /* LUT    6 23  3 */ n689;
assign n5363 = /* LUT   20  8  4 */ n2673;
assign n5364 = /* LUT   12 28  2 */ n1395;
assign n5365 = /* LUT   23 22  7 */ n3285;
assign n5366 = /* LUT   14  6  1 */ n1579;
assign n5367 = /* LUT   16  5  5 */ n1892;
assign n5368 = /* LUT   17 19  5 */ n2132;
assign n5369 = /* LUT   29 12  5 */ n3853;
assign n5370 = /* LUT   16 10  4 */ n1929;
assign n5371 = /* LUT    5 21  2 */ (\rco[110]  ? (n676 ? (n553 ? n554 : 1'b0) : 1'b0) : 1'b0);
assign n5372 = /* LUT   10 28  1 */ n1101;
assign n5373 = /* LUT    9 12  1 */ n1001;
assign n5374 = /* LUT   24  9  0 */ n3338;
assign n5375 = /* LUT   27 17  1 */ n3654;
assign n5376 = /* LUT   15 24  7 */ n1859;
assign n5377 = /* LUT   21 23  6 */ n2950;
assign n5378 = /* LUT   15 23  6 */ n1857;
assign n5379 = /* LUT   18  8  2 */ n2250;
assign n5380 = /* LUT   12 18  7 */ n1326;
assign n5381 = /* LUT   26 11  6 */ n3513;
assign n5382 = /* LUT   29 19  3 */ n3863;
assign n2322 = /* LUT   17 16  1 */ (n2109 ? \rco[23]  : 1'b0);
assign n5383 = /* LUT    2 15  2 */ (\rco[0]  ? n302 : 1'b0);
assign n5384 = /* LUT   22 20  3 */ n3090;
assign n5385 = /* LUT   10 14  2 */ n1010;
assign n5386 = /* LUT   24 23  3 */ n3293;
assign n5387 = /* LUT   16 24  0 */ (\rco[118]  ? (n117 ? (n121 ? n338 : 1'b0) : 1'b0) : 1'b0);
assign n5388 = /* LUT   27 18  5 */ n3669;
assign n5389 = /* LUT    4 17  0 */ (n327 ? (n225 ? (n120 ? \rco[0]  : 1'b0) : 1'b0) : 1'b0);
assign n5390 = /* LUT    3 11  2 */ n271;
assign n5391 = /* LUT    7  9  1 */ n595;
assign n5392 = /* LUT   21 20  0 */ n3093;
assign n5393 = /* LUT   13 24  6 */ (n669 ? \rco[110]  : 1'b0);
assign n5394 = /* LUT   27 15  5 */ n3649;
assign n5395 = /* LUT    9 17  4 */ n886;
assign n5396 = /* LUT   18 26  2 */ n2386;
assign n5397 = /* LUT   20 12  1 */ n2698;
assign n5398 = /* LUT   19 28  1 */ n2624;
assign n5399 = /* LUT   28 19  7 */ n3677;
assign n5400 = /* LUT   10 13  4 */ n1004;
assign n5401 = /* LUT   28 24  6 */ (n1684 ? \rco[138]  : 1'b0);
assign n5402 = /* LUT   16 22  1 */ (n129 ? \rco[118]  : 1'b0);
assign n202  = /* LUT    1 15  0 */ (n31 ? (n181 ? (n73 ? !n56 : 1'b0) : 1'b0) : 1'b0);
assign n5403 = /* LUT   22  6  3 */ n2992;
assign n5404 = /* LUT   22 11  4 */ (\rco[53]  ? n2859 : 1'b0);
assign n5405 = /* LUT   13 21  0 */ n1518;
assign n5406 = /* LUT   30 10  0 */ n3890;
assign n5407 = /* LUT   15 11  3 */ n1765;
assign n5408 = /* LUT    2 19  0 */ (\rco[123]  ? (n116 ? (n121 ? \rco[0]  : 1'b0) : 1'b0) : 1'b0);
assign n5409 = /* LUT    6 13  5 */ n619;
assign n5410 = /* LUT   20 18  6 */ n2747;
assign n5411 = /* LUT    6 22  4 */ n681;
assign n5412 = /* LUT   20 15  5 */ n2721;
assign n5413 = /* LUT   23 23  4 */ n3290;
assign n5414 = /* LUT   11 13  7 */ n735;
assign n5415 = /* LUT   16  4  2 */ n2033;
assign n5416 = /* LUT    5 22  3 */ n557;
assign n5417 = /* LUT    9 13  2 */ n1006;
assign n5418 = /* LUT   13  7  1 */ n1423;
assign n5419 = /* LUT   15 25  0 */ (n2011 ? (\rco[183]  ? n2003 : 1'b0) : 1'b0);
assign n5420 = /* LUT    7 13  6 */ n811;
assign n5421 = /* LUT   18 11  3 */ (\rco[9]  ? n2495 : 1'b0);
assign n5422 = /* LUT   15 20  7 */ n1833;
assign n5423 = /* LUT   12 17  6 */ n1317;
assign n5424 = /* LUT   26 10  1 */ n3507;
assign n5425 = /* LUT   18 30  7 */ n2409;
assign n5426 = /* LUT   29 20  2 */ n3869;
assign n5427 = /* LUT   26  7  6 */ n3487;
assign n5428 = /* LUT   17 17  2 */ n2115;
assign n5429 = /* LUT   22 23  2 */ (\rco[162]  ? (n982 ? (n1710 ? \rco[0]  : 1'b0) : 1'b0) : 1'b0);
assign n5430 = /* LUT   24 22  0 */ n3430;
assign n5431 = /* LUT    1 11  5 */ n41;
assign n5432 = /* LUT   27 19  6 */ n3674;
assign n5433 = /* LUT    7 14  0 */ n731;
assign n5434 = /* LUT   21 21  3 */ n2928;
assign n5435 = /* LUT   13 25  5 */ n1538;
assign n5436 = /* LUT   27 12  4 */ n3632;
assign n5437 = /* LUT    9 18  5 */ n896;
assign n5438 = /* LUT   18 29  3 */ n2410;
assign n5439 = /* LUT    6 18  1 */ n649;
assign n5440 = /* LUT    5 10  1 */ n287;
assign n5441 = /* LUT   19 29  6 */ n2626;
assign n5442 = /* LUT   11  9  4 */ n1133;
assign n5443 = /* LUT   23 27  1 */ n3312;
assign n5444 = /* LUT   11 28  3 */ n1257;
assign n5445 = /* LUT   10 12  7 */ n853;
assign n5446 = /* LUT   24 25  6 */ n3451;
assign n5447 = /* LUT   16 21  0 */ n1986;
assign n5448 = /* LUT    1  8  1 */ n14;
assign n5449 = /* LUT   13 22  1 */ n1522;
assign n5450 = /* LUT   31 23  1 */ (\rco[183]  ? n3124 : 1'b0);
assign n5451 = /* LUT   15  8  2 */ n1598;
assign n5452 = /* LUT    3 22  3 */ n354;
assign n3008 = /* LUT   21  7  3 */ (n2470 ? (\rco[0]  ? (n2270 ? !n2510 : 1'b1) : 1'b1) : 1'b1);
assign n5454 = /* LUT    6 12  6 */ n600;
assign n5455 = /* LUT   20 17  7 */ n2548;
assign n5456 = /* LUT   26 14  6 */ n3537;
assign n5457 = /* LUT   23 20  5 */ n3267;
assign n5458 = /* LUT    9 14  3 */ n861;
assign n5459 = /* LUT    4 20  4 */ n443;
assign n5460 = /* LUT   21  9  4 */ n2848;
assign n5461 = /* LUT    9 27  7 */ n952;
assign n5462 = /* LUT   18 10  4 */ n2276;
assign n5463 = /* LUT   12 16  1 */ n1299;
assign n3639 = /* LUT   26 13  0 */ (n3528 ? n3516 : 1'b0);
assign n5464 = /* LUT   14 18  0 */ n1664;
assign n5465 = /* LUT   12 29  6 */ n1382;
assign n5466 = /* LUT    1 20  3 */ n221;
assign n5467 = /* LUT   19 25  3 */ n2606;
assign n5468 = /* LUT   23 10  1 */ n3186;
assign n5469 = /* LUT   22 22  5 */ n3110;
assign n3470 = /* LUT   24 21  1 */ (\rco[145]  ? (\rco[0]  ? (n817 ? n2574 : 1'b0) : 1'b0) : 1'b0);
assign n5470 = /* LUT   13  5  6 */ n1413;
assign n815  = /* LUT    7 15  3 */ (n59 ? (n814 ? (n56 ? 1'b0 : n289) : 1'b0) : 1'b0);
assign n5471 = /* LUT    9 24  3 */ n934;
assign n5472 = /* LUT   13 26  4 */ n1547;
assign n5473 = /* LUT   21 22  2 */ n2936;
assign n5474 = /* LUT    2 22  4 */ n238;
assign n2628 = /* LUT   18 28  0 */ (\rco[183]  ? n1699 : 1'b0);
assign n5475 = /* LUT   19 26  7 */ (\rco[172]  ? (\rco[0]  ? (n2044 ? n2563 : 1'b0) : 1'b0) : 1'b0);
assign n5476 = /* LUT    5 11  6 */ n480;
assign n5477 = /* LUT   11 22  5 */ n1212;
assign n5478 = /* LUT   23 24  0 */ n2173;
assign n5479 = /* LUT   28 17  5 */ n3770;
assign n5480 = /* LUT   16 15  6 */ n1949;
assign n5481 = /* LUT   11 29  4 */ n1265;
assign n5482 = /* LUT   10 15  6 */ n1020;
assign n5483 = /* LUT   16 20  7 */ n1977;
assign n5484 = /* LUT   21 24  1 */ n2960;
assign n5485 = /* LUT   15 18  4 */ n1811;
assign n5486 = /* LUT   18 14  1 */ (n2521 ? (n2523 ? (n2122 ? !n2124 : 1'b1) : 1'b1) : 1'b1);
assign n5487 = /* LUT    2 21  6 */ n232;
assign n5488 = /* LUT    6 15  7 */ n636;
assign n5489 = /* LUT   12 20  6 */ (\rco[118]  ? (\rco[0]  ? (n117 ? n338 : 1'b0) : 1'b0) : 1'b0);
assign n5490 = /* LUT    6 16  6 */ n523;
assign n5491 = /* LUT   20 13  7 */ n2506;
assign n5492 = /* LUT   14  3  2 */ (n1623 ? (n587 ? \rco[83]  : 1'b0) : 1'b0);
assign n5493 = /* LUT    4 11  0 */ (n287 ? (n103 ? (n386 ? n376 : 1'b0) : 1'b0) : 1'b0);
assign n5494 = /* LUT   22 18  2 */ n3081;
assign n5495 = /* LUT    9 15  4 */ n870;
assign n5496 = /* LUT   28 12  0 */ n3758;
assign n5497 = /* LUT   21 10  5 */ (\rco[48]  ? (n2725 ? \rco[0]  : 1'b0) : 1'b0);
assign n5498 = /* LUT    7 19  4 */ n762;
assign n5499 = /* LUT    9 20  6 */ n911;
assign n5500 = /* LUT   18 13  5 */ n2299;
assign n5501 = /* LUT   12 23  0 */ n551;
assign n5502 = /* LUT   26 12  3 */ n3524;
assign n5503 = /* LUT    5 15  3 */ n516;
assign n5504 = /* LUT   19 22  2 */ n2585;
assign n5505 = /* LUT   23 11  2 */ n3191;
assign n5506 = /* LUT   11 25  1 */ n1221;
assign n5507 = /* LUT   22 17  4 */ n3075;
assign n5508 = /* LUT   24 20  6 */ n3419;
assign n5509 = /* LUT   16 16  4 */ n1962;
assign n5510 = /* LUT   13  6  7 */ n1430;
assign n5511 = /* LUT    9 25  0 */ (n658 ? (n117 ? (n121 ? \rco[120]  : 1'b0) : 1'b0) : 1'b0);
assign n5512 = /* LUT   13 27  3 */ (n1272 ? (n1558 ? (n1390 ? !n1543 : 1'b1) : 1'b1) : 1'b1);
assign n3749 = /* LUT   27 10  2 */ (n3646 ? (n3525 ? (n3619 ? n3622 : 1'b0) : 1'b0) : 1'b0);
assign n5513 = /* LUT   15 13  2 */ n1778;
assign n5514 = /* LUT   20 20  5 */ n2765;
assign n5515 = /* LUT   23 18  6 */ n3248;
assign n5516 = /* LUT    5 12  7 */ n486;
assign n5517 = /* LUT   19 27  4 */ n2619;
assign n5518 = /* LUT   11 23  6 */ n1220;
assign n5519 = /* LUT   23 25  7 */ n3453;
assign n5520 = /* LUT   11 26  5 */ n1240;
assign n5521 = /* LUT   16 19  6 */ n1879;
assign n5522 = /* LUT    1 10  3 */ n32;
assign n5523 = /* LUT   21 25  2 */ n2963;
assign n5524 = /* LUT    9 11  1 */ n842;
assign n5525 = /* LUT   15 19  7 */ n1823;
assign n5526 = /* LUT   18 17  0 */ (\rco[37]  ? \rco[0]  : 1'b0);
assign n5527 = /* LUT    3 20  1 */ n342;
assign n5528 = /* LUT   15 14  4 */ n1786;
assign n5529 = /* LUT    6 14  0 */ n627;
assign n5530 = /* LUT   20 23  1 */ n2772;
assign n5531 = /* LUT   12 27  7 */ (\rco[99]  ? !n1560 : 1'b0);
assign n5532 = /* LUT   11  8  4 */ n1126;
assign n5533 = /* LUT   29  5  2 */ n3819;
assign n5534 = /* LUT   19  9  0 */ n2477;
assign n5535 = /* LUT    4 10  3 */ n381;
assign n5536 = /* LUT   24 16  3 */ n3386;
assign n5537 = /* LUT   27 22  4 */ n3698;
assign n5538 = /* LUT   13 10  2 */ n1435;
assign n5539 = /* LUT   18  3  7 */ n2030;
assign n5540 = /* LUT    7 16  5 */ n747;
assign n5541 = /* LUT    9 21  5 */ n918;
assign n5542 = /* LUT   18 12  6 */ n2291;
assign n5543 = /* LUT   21 11  2 */ (n2691 ? n2416 : 1'b0);
assign n5544 = /* LUT   21  6  5 */ n2837;
assign n5545 = /* LUT   12 22  3 */ n1350;
assign n5546 = /* LUT   26 15  2 */ n3541;
assign n5547 = /* LUT   14 12  2 */ (n1666 ? (n1774 ? (n1375 ? !n817 : 1'b1) : 1'b1) : 1'b1);
assign n5548 = /* LUT   19 23  1 */ (\rco[172]  ? (n2229 ? n2173 : 1'b0) : 1'b0);
assign n5549 = /* LUT   10  9  7 */ n979;
assign n5550 = /* LUT   28 20  7 */ (\rco[162]  ? n3240 : 1'b0);
assign n5551 = /* LUT   31  9  1 */ (n3636 ? (\rco[66]  ? (n3034 ? n3463 : 1'b0) : 1'b0) : 1'b0);
assign n5552 = /* LUT    4 21  4 */ n450;
assign n5553 = /* LUT   13 28  2 */ n1562;
assign n5554 = /* LUT   26 17  1 */ n2333;
assign n5555 = /* LUT   27 11  1 */ n3623;
assign n5556 = /* LUT    6 10  5 */ n597;
assign n5557 = /* LUT   20 11  4 */ n2693;
assign n5558 = /* LUT   23 19  5 */ n3254;
assign n5559 = /* LUT    5 13  4 */ n492;
assign n5560 = /* LUT   19 24  5 */ n2598;
assign n5561 = /* LUT   11 20  7 */ n1204;
assign n5562 = /* LUT   29  9  7 */ n3831;
assign n5563 = /* LUT   17 27  6 */ n2193;
assign n5564 = /* LUT   28 23  3 */ n3806;
assign n5565 = /* LUT   11 27  6 */ n1252;
assign n5566 = /* LUT   21 26  3 */ (\rco[153]  ? (n3141 ? !n2602 : 1'b0) : 1'b0);
assign n5567 = /* LUT   15 16  6 */ n1798;
assign n5568 = /* LUT   21 15  7 */ (n3050 ? n2895 : 1'b0);
assign n5569 = /* LUT   15 15  7 */ (\rco[0]  ? (n1954 ? (n823 ? n758 : 1'b0) : 1'b0) : 1'b0);
assign n5570 = /* LUT    3 21  6 */ (\rco[123]  ? (n461 ? (n440 ? n455 : 1'b0) : 1'b0) : 1'b0);
assign n5571 = /* LUT   18 16  3 */ n2316;
assign n726  = /* LUT    6  9  1 */ (n56 ? 1'b0 : (n87 ? n403 : 1'b0));
assign n5573 = /* LUT   20 22  2 */ n2777;
assign n5574 = /* LUT   12 26  4 */ n1388;
assign n5575 = /* LUT   17 24  0 */ n913;
assign n5576 = /* LUT   19  6  1 */ n2443;
assign n5577 = /* LUT    4  9  2 */ n372;
assign n5578 = /* LUT   10  6  3 */ n972;
assign n5579 = /* LUT   24 15  2 */ n3378;
assign n5580 = /* LUT    9  9  6 */ n833;
assign n5581 = /* LUT   13 11  5 */ n1445;
assign n5582 = /* LUT   18  2  0 */ n2218;
assign n5583 = /* LUT    7 17  2 */ n752;
assign n5584 = /* LUT    9 22  4 */ n931;
assign n5585 = /* LUT   18 15  7 */ n1311;
assign n5586 = /* LUT   21 12  3 */ n2869;
assign n5587 = /* LUT   14 26  4 */ n1714;
assign n5588 = /* LUT   12 21  2 */ n1342;
assign n5589 = /* LUT   14 15  3 */ n1641;
assign n5590 = /* LUT    2  9  0 */ n261;
assign n5591 = /* LUT   20  4  2 */ (\rco[93]  ? n2240 : 1'b0);
assign n5592 = /* LUT   19 20  0 */ n2002;
assign n5593 = /* LUT    9 32  2 */ (n1115 ? n1113 : 1'b0);
assign n5594 = /* LUT   23  9  4 */ n3179;
assign n5595 = /* LUT   22 19  6 */ (\rco[99]  ? (n3262 ? 1'b0 : (n912 ? n809 : 1'b0)) : 1'b0);
assign n5596 = /* LUT   16 30  6 */ (n225 ? \rco[132]  : 1'b0);
assign n3733 = /* LUT   27  8  0 */ (n3348 ? n3337 : 1'b0);
assign n5597 = /* LUT    3 17  3 */ n312;
assign n5598 = /* LUT   14 25  6 */ n1708;
assign n781  = /* LUT    6 21  4 */ (n361 ? (n669 ? (n550 ? n243 : 1'b0) : 1'b0) : 1'b0);
assign n5600 = /* LUT   20 10  7 */ n2494;
assign n5601 = /* LUT   23 16  4 */ n3230;
assign n5602 = /* LUT   20  7  4 */ n2664;
assign n5603 = /* LUT    5 14  5 */ n508;
assign n5604 = /* LUT   11 21  0 */ (n769 ? (n361 ? (n551 ? n243 : 1'b0) : 1'b0) : 1'b0);
assign n5605 = /* LUT   29 10  6 */ n3832;
assign n5606 = /* LUT   28 22  0 */ n3800;
assign n5607 = /* LUT   16 12  3 */ n1937;
assign n5608 = /* LUT   11 24  7 */ n1229;
assign n5609 = /* LUT   16 17  4 */ n1966;
assign n5610 = /* LUT   21 27  4 */ n2975;
assign n5611 = /* LUT   13 15  2 */ n1471;
assign n5612 = /* LUT   30 12  6 */ n3899;
assign n5613 = /* LUT   15 17  1 */ n1801;
assign n5614 = /* LUT   18  6  5 */ n2235;
assign n5615 = /* LUT    7 21  7 */ n566;
assign n5616 = /* LUT   18 19  2 */ n2340;
assign n5617 = /* LUT    3 18  7 */ n324;
assign n5618 = /* LUT    6  8  2 */ n574;
assign n5619 = /* LUT   20 21  3 */ n2770;
assign n5620 = /* LUT   12 25  5 */ n1380;
assign n5621 = /* LUT    1 19  3 */ n106;
assign n5622 = /* LUT   17 25  3 */ n2178;
assign n5623 = /* LUT    5 16  1 */ n522;
assign n5624 = /* LUT   19  7  2 */ n2453;
assign n5625 = /* LUT   23 13  1 */ n3208;
assign n5626 = /* LUT   10 25  2 */ n1081;
assign n5627 = /* LUT   24 14  1 */ n3369;
assign n5628 = /* LUT   27 20  6 */ n3782;
assign n5629 = /* LUT    9 10  7 */ n840;
assign n5630 = /* LUT   13 12  4 */ n1452;
assign n5631 = /* LUT   18  5  1 */ n2221;
assign n5632 = /* LUT    7 22  3 */ n785;
assign n5633 = /* LUT    9 23  3 */ n927;
assign n5634 = /* LUT   21 13  0 */ n2879;
assign n5635 = /* LUT   14 21  5 */ (n1592 ? (\rco[0]  ? (n1671 ? \rco[110]  : 1'b0) : 1'b0) : 1'b0);
assign n5636 = /* LUT   19 30  6 */ n2640;
assign n5637 = /* LUT   17 11  0 */ (n962 ? (n2067 ? (n1491 ? !\rco[37]  : 1'b1) : 1'b1) : 1'b1);
assign n5638 = /* LUT    2  8  3 */ n156;
assign n5639 = /* LUT    1 16  7 */ n93;
assign n5640 = /* LUT   14 14  4 */ n1635;
assign n5641 = /* LUT   19 21  7 */ n2588;
assign n5642 = /* LUT   11 17  5 */ n1174;
assign n5643 = /* LUT   10 11  5 */ n994;
assign n5644 = /* LUT   23 14  5 */ n3220;
assign n5645 = /* LUT   24 17  5 */ n3398;
assign n5646 = /* LUT   28  7  6 */ n3725;
assign n5647 = /* LUT    3 14  1 */ (\rco[0]  ? n410 : 1'b0);
assign n5648 = /* LUT   15 21  6 */ n1841;
assign n5649 = /* LUT   12 10  2 */ n206;
assign n5650 = /* LUT   26 19  3 */ n3557;
assign n5651 = /* LUT   17  5  1 */ (n1592 ? \rco[138]  : 1'b0);
assign n5652 = /* LUT   14 24  5 */ (n1541 ? (n1816 ? n1872 : 1'b0) : 1'b0);
assign n5653 = /* LUT    6 20  7 */ n666;
assign n5654 = /* LUT   20  9  6 */ (n2854 ? n2669 : 1'b0);
assign n5655 = /* LUT   23 17  3 */ n3236;
assign n5656 = /* LUT    2  7  7 */ n151;
assign n5657 = /* LUT   26  6  7 */ n3479;
assign n5658 = /* LUT   11 18  1 */ n1037;
assign n5659 = /* LUT   29 11  1 */ n3839;
assign n5660 = /* LUT   28 21  1 */ n3791;
assign n5661 = /* LUT    4 12  2 */ n394;
assign n5662 = /* LUT   10 22  0 */ (\rco[0]  ? (n669 ? (\rco[110]  ? n550 : 1'b0) : 1'b0) : 1'b0);
assign n5663 = /* LUT   21 28  5 */ n2983;
assign n5664 = /* LUT   13 16  3 */ n1479;
assign n5665 = /* LUT   27  7  0 */ (n3455 ? (n3456 ? (n2676 ? !n3174 : 1'b1) : 1'b1) : 1'b1);
assign n5666 = /* LUT   15 22  0 */ n1851;
assign n5667 = /* LUT   18  9  4 */ n2264;
assign n5668 = /* LUT   18 18  5 */ n2126;
assign n5669 = /* LUT    3 19  4 */ n332;
assign n5670 = /* LUT    6 11  3 */ n601;
assign n5671 = /* LUT   12 24  2 */ n1368;
assign n5672 = /* LUT   14 10  1 */ n1604;
assign n5673 = /* LUT   19 17  4 */ n2544;
assign n5674 = /* LUT   22 21  7 */ n2933;
assign n5675 = /* LUT   24 24  7 */ n3302;
assign n5676 = /* LUT    5 17  2 */ n525;
assign n5677 = /* LUT    4 15  4 */ n415;
assign n5678 = /* LUT   10 24  1 */ n1072;
assign n5679 = /* LUT   24 13  0 */ n3366;
assign n3848 = /* LUT   28 11  5 */ (n3847 ? (n3528 ? (n3516 ? n3463 : 1'b0) : 1'b0) : 1'b0);
assign n5681 = /* LUT   27 21  1 */ n3687;
assign n5682 = /* LUT   18  4  2 */ n2214;
assign n5683 = /* LUT    7 23  0 */ n793;
assign n5684 = /* LUT    9 16  2 */ n876;
assign n5685 = /* LUT   21 14  1 */ n2882;
assign n5686 = /* LUT   14 20  6 */ n1682;
assign n5687 = /* LUT    5  8  6 */ n470;
assign n5688 = /* LUT   17 20  1 */ n2136;
assign n5689 = /* LUT    2 11  2 */ n169;
assign n5690 = /* LUT   19 31  5 */ n2645;
assign n5691 = /* LUT   19 18  6 */ n2559;
assign n5692 = /* LUT   10 10  2 */ n984;
assign n5693 = /* LUT   23 15  6 */ n3227;
assign n5694 = /* LUT   28  6  5 */ n3715;
assign n5695 = /* LUT    3 15  2 */ n294;
assign n5696 = /* LUT   21 16  0 */ n2740;
assign n5697 = /* LUT   26 18  4 */ (n2124 ? (n3666 ? (n2521 ? \rco[23]  : 1'b0) : 1'b0) : 1'b0);
assign n5698 = /* LUT   12  9  3 */ n1287;
assign n2590 = /* LUT   18 22  2 */ (n2037 ? n2357 : 1'b0);
assign n5699 = /* LUT   17  6  0 */ n2042;
assign n5700 = /* LUT    6 23  6 */ n692;
assign n5701 = /* LUT   20  8  1 */ n2672;
assign n5702 = /* LUT   12 28  7 */ n1400;
assign n5703 = /* LUT   23 22  2 */ n3280;
assign n5704 = /* LUT   29 12  0 */ n3854;
assign n5705 = /* LUT   16 10  1 */ n1926;
assign n5706 = /* LUT   22 26  3 */ n3135;
assign n5707 = /* LUT   27 17  6 */ n3656;
assign n5708 = /* LUT   13 17  0 */ n1489;
assign n5709 = /* LUT   15 23  3 */ n1854;
assign n5710 = /* LUT   18  8  7 */ n2255;
assign n5711 = /* LUT   18 21  4 */ n2352;
assign n5712 = /* LUT    3 16  5 */ n308;
assign n5713 = /* LUT   14  5  0 */ n1578;
assign n5714 = /* LUT   19 14  5 */ n2517;
assign n5715 = /* LUT   22 20  4 */ n3091;
assign n5716 = /* LUT   10 14  7 */ n1017;
assign n5717 = /* LUT    5 18  3 */ n533;
assign n5718 = /* LUT    4 14  7 */ n408;
assign n5719 = /* LUT   19  5  4 */ n2438;
assign n5720 = /* LUT   10 27  0 */ n1098;
assign n5721 = /* LUT   22 25  7 */ n3310;
assign n5722 = /* LUT   27 18  0 */ n2521;
assign n5723 = /* LUT   24 12  7 */ n3359;
assign n5724 = /* LUT   28 10  6 */ n3746;
assign n5725 = /* LUT   13 14  6 */ n1467;
assign n5726 = /* LUT   18  7  3 */ (n2057 ? (n2266 ? \rco[93]  : 1'b0) : 1'b0);
assign n5727 = /* LUT    9 17  1 */ n883;
assign n5728 = /* LUT   26 22  1 */ n3569;
assign n5729 = /* LUT   15  5  3 */ n1727;
assign n5730 = /* LUT   14 23  7 */ (n674 ? (n1863 ? (n1196 ? !n1383 : 1'b0) : 1'b0) : 1'b0);
assign n5731 = /* LUT   20 12  6 */ n2703;
assign n5732 = /* LUT   14  8  6 */ n1600;
assign n5733 = /* LUT   17 21  2 */ n2145;
assign n5734 = /* LUT   19 19  5 */ (\rco[162]  ? (\rco[0]  ? (n1710 ? n1998 : 1'b0) : 1'b0) : 1'b0);
assign n5735 = /* LUT   10 13  3 */ n1031;
assign n5736 = /* LUT   24 26  0 */ n3140;
assign n5737 = /* LUT   23 12  7 */ n3197;
assign n5738 = /* LUT   28  5  4 */ n3708;
assign n5739 = /* LUT   16 27  1 */ n2018;
assign n5740 = /* LUT    3 12  3 */ n281;
assign n5741 = /* LUT    7 10  0 */ n725;
assign n5742 = /* LUT   21 17  3 */ (n2910 ? \rco[59]  : 1'b0);
assign n5743 = /* LUT   30 10  5 */ n3889;
assign n5744 = /* LUT   15 11  4 */ n1766;
assign n5745 = /* LUT   12  8  4 */ n1281;
assign n5746 = /* LUT   26 21  5 */ n3566;
assign n5747 = /* LUT   15  6  7 */ n1904;
assign n5748 = /* LUT   17  7  7 */ n2052;
assign n5749 = /* LUT   18 25  3 */ n2379;
assign n5750 = /* LUT    6 22  1 */ n226;
assign n5751 = /* LUT   20 15  0 */ n2724;
assign n5752 = /* LUT   23 23  1 */ n3287;
assign n5753 = /* LUT   11 16  3 */ n1161;
assign n5754 = /* LUT   16  9  0 */ n1925;
assign n5755 = /* LUT    1 12  1 */ n46;
assign n5756 = /* LUT   13  7  6 */ n1428;
assign n5757 = /* LUT    7  7  6 */ n716;
assign n5758 = /* LUT   13 18  1 */ n1492;
assign n5759 = /* LUT   27  5  6 */ n3590;
assign n5760 = /* LUT   18 11  6 */ (n2278 ? (n2496 ? (\rco[0]  ? n2306 : 1'b0) : 1'b0) : 1'b0);
assign n5761 = /* LUT   15 20  2 */ n1828;
assign n5762 = /* LUT   18 20  7 */ (\rco[153]  ? (\rco[0]  ? (n811 ? n737 : 1'b0) : 1'b0) : 1'b0);
assign n5763 = /* LUT   12 30  0 */ n1401;
assign n5764 = /* LUT   26  7  1 */ n3481;
assign n5765 = /* LUT    2 14  2 */ n188;
assign n5766 = /* LUT   16  7  3 */ n1909;
assign n5767 = /* LUT   19 15  6 */ n2532;
assign n5768 = /* LUT   23  5  5 */ n3154;
assign n5769 = /* LUT   22 23  5 */ n3115;
assign n5770 = /* LUT   24 22  5 */ n3429;
assign n5771 = /* LUT    5 19  4 */ n542;
assign n5772 = /* LUT    4 13  6 */ (n291 ? (n503 ? (n500 ? n298 : 1'b0) : 1'b0) : 1'b0);
assign n5773 = /* LUT   22 24  4 */ n2959;
assign n5774 = /* LUT   10 26  7 */ (n1221 ? (\rco[0]  ? (n1087 ? !n803 : 1'b1) : 1'b1) : 1'b1);
assign n3468 = /* LUT   24 11  6 */ (\rco[37]  ? n3467 : 1'b0);
assign n5775 = /* LUT   28  9  7 */ n3617;
assign n5776 = /* LUT   27 19  3 */ n3661;
assign n5777 = /* LUT    9 18  0 */ n899;
assign n5778 = /* LUT   26  9  0 */ n3619;
assign n5779 = /* LUT   29 17  1 */ n3859;
assign n5780 = /* LUT   14 22  0 */ n1684;
assign n5781 = /* LUT   17  3  4 */ n2028;
assign n5782 = /* LUT    6 18  6 */ n654;
assign n5783 = /* LUT    5 10  4 */ n477;
assign n5784 = /* LUT   14 11  7 */ n1611;
assign n5785 = /* LUT   17 22  3 */ n2154;
assign n5786 = /* LUT   19 29  3 */ n2631;
assign n5787 = /* LUT   19 16  4 */ n2549;
assign n5788 = /* LUT   23  6  1 */ n3159;
assign n5789 = /* LUT   11 28  6 */ n1262;
assign n5790 = /* LUT   10 12  0 */ n989;
assign n5791 = /* LUT   24 25  1 */ n3446;
assign n407  = /* LUT    3 13  4 */ (n398 ? (n406 ? (n386 ? n376 : 1'b0) : 1'b0) : 1'b0);
assign n5792 = /* LUT   22 10  0 */ n2689;
assign n5793 = /* LUT    9 28  3 */ n945;
assign n5794 = /* LUT   21 18  2 */ n2915;
assign n5795 = /* LUT   15  8  5 */ n1751;
assign n5796 = /* LUT    3 22  6 */ n240;
assign n5797 = /* LUT   12 15  5 */ n1305;
assign n3686 = /* LUT   26 20  6 */ (n3093 ? (n3685 ? n3420 : 1'b0) : 1'b0);
assign n5798 = /* LUT   15  7  4 */ (n614 ? (n1914 ? \rco[0]  : 1'b0) : 1'b0);
assign n5799 = /* LUT   18 24  0 */ n2375;
assign n5800 = /* LUT    6 17  0 */ n647;
assign n5801 = /* LUT   23 20  0 */ n3269;
assign n5802 = /* LUT    1 13  2 */ n62;
assign n5803 = /* LUT   24  7  5 */ (\rco[74]  ? (n3175 ? (\rco[0]  ? n3456 : 1'b0) : 1'b0) : 1'b0);
assign n5804 = /* LUT    9 14  6 */ n866;
assign n1675 = /* LUT   13 19  6 */ (n1340 ? (n1620 ? (n1666 ? \rco[23]  : 1'b0) : 1'b0) : 1'b0);
assign n5805 = /* LUT   18 10  1 */ n2273;
assign n5806 = /* LUT   20 28  0 */ (\rco[183]  ? (n1877 ? (n2823 ? \rco[0]  : 1'b0) : 1'b0) : 1'b0);
assign n5807 = /* LUT   18 23  6 */ n2368;
assign n5808 = /* LUT   12 29  1 */ n1405;
assign n5809 = /* LUT   14  7  2 */ n1586;
assign n5810 = /* LUT   16  6  0 */ n1738;
assign n5811 = /* LUT   19 12  7 */ n2293;
assign n5812 = /* LUT   23 10  4 */ n3185;
assign n5813 = /* LUT   22 22  2 */ n3106;
assign n5814 = /* LUT   24 21  4 */ n3417;
assign n5815 = /* LUT   19  3  6 */ n2432;
assign n5816 = /* LUT   22 27  5 */ n3147;
assign n5817 = /* LUT   24 10  5 */ n3344;
assign n5818 = /* LUT   28  8  0 */ n3731;
assign n5819 = /* LUT    3  9  1 */ n252;
assign n5820 = /* LUT   12 19  0 */ n1333;
assign n5821 = /* LUT   26  8  3 */ n3492;
assign n5822 = /* LUT   14 17  1 */ n1654;
assign n5823 = /* LUT   17 12  5 */ n2081;
assign n5824 = /* LUT   19 26  2 */ (n2002 ? (\rco[172]  ? (n1998 ? \rco[0]  : 1'b0) : 1'b0) : 1'b0);
assign n5825 = /* LUT   17 23  4 */ n1531;
assign n5826 = /* LUT    2 12  7 */ n53;
assign n5827 = /* LUT   23  7  2 */ n3167;
assign n5828 = /* LUT   11 29  1 */ (\rco[100]  ? n1272 : 1'b0);
assign n5829 = /* LUT   10 15  1 */ n1022;
assign n5830 = /* LUT   16 25  3 */ n2005;
assign n5831 = /* LUT   21 24  4 */ n2956;
assign n5832 = /* LUT    3 10  5 */ n266;
assign n5833 = /* LUT   21 19  5 */ n2911;
assign n5834 = /* LUT   13 23  3 */ n1526;
assign n5835 = /* LUT   27 14  2 */ n3642;
assign n5836 = /* LUT   18 14  6 */ (n2124 ? (n2521 ? (\rco[31]  ? n2122 : 1'b0) : 1'b0) : 1'b0);
assign n5837 = /* LUT   12 14  6 */ n1293;
assign n5838 = /* LUT   26 23  7 */ n3702;
assign n5839 = /* LUT   18 27  1 */ n2393;
assign n5840 = /* LUT    6 16  3 */ n640;
assign n2881 = /* LUT   20 13  2 */ (n1772 ? (n1759 ? n2502 : 1'b0) : 1'b0);
assign n5841 = /* LUT    4 11  7 */ n482;
assign n5842 = /* LUT   22 18  7 */ n3079;
assign n5843 = /* LUT    1 14  3 */ n70;
assign n5844 = /* LUT   22  7  0 */ n3004;
assign n1177 = /* LUT   10 17  5 */ (n989 ? (n847 ? (n888 ? n1032 : 1'b0) : 1'b0) : 1'b0);
assign n5846 = /* LUT    9 15  1 */ n867;
assign n5847 = /* LUT   13  9  4 */ n1432;
assign n5848 = /* LUT   24  6  6 */ n3328;
assign n5849 = /* LUT   28 12  5 */ n3759;
assign n5850 = /* LUT   13 20  7 */ n1509;
assign n5851 = /* LUT   18 13  0 */ n2510;
assign n5852 = /* LUT   20 19  1 */ n2767;
assign n5853 = /* LUT   14  6  5 */ n1581;
assign n5854 = /* LUT   16  5  1 */ n1888;
assign n5855 = /* LUT   17 19  1 */ n2128;
assign n5856 = /* LUT   23 11  7 */ n3196;
assign n5857 = /* LUT   22 17  3 */ n3074;
assign n5858 = /* LUT   24 20  3 */ n3406;
assign n5859 = /* LUT   10 28  5 */ n1105;
assign n5860 = /* LUT   24  9  4 */ n3335;
assign n5861 = /* LUT   13  6  2 */ n1416;
assign n5862 = /* LUT   28 15  1 */ n3760;
assign n5863 = /* LUT   15 24  3 */ n1866;
assign n5864 = /* LUT   21 23  2 */ n2944;
assign n5865 = /* LUT   26 11  2 */ (\rco[66]  ? n3526 : 1'b0);
assign n5866 = /* LUT   12 18  3 */ n1322;
assign n5867 = /* LUT   29 19  7 */ n3875;
assign n5868 = /* LUT   14 16  2 */ n1647;
assign n5869 = /* LUT   17 13  6 */ n2093;
assign n5870 = /* LUT    5 12  2 */ n484;
assign n2324 = /* LUT   17 16  5 */ (n812 ? (n206 ? n880 : 1'b0) : 1'b0);
assign n5871 = /* LUT    2 15  6 */ n200;
assign n5872 = /* LUT   19 27  1 */ n2616;
assign n5873 = /* LUT   11 26  0 */ n1241;
assign n5874 = /* LUT   21 25  7 */ n3132;
assign n5875 = /* LUT    9 11  6 */ n849;
assign n5876 = /* LUT    3 11  6 */ n276;
assign n5877 = /* LUT    7  9  5 */ n722;
assign n5878 = /* LUT   21 20  4 */ n2921;
assign n5879 = /* LUT   13 24  2 */ (\rco[99]  ? (n1700 ? (n769 ? \rco[0]  : 1'b0) : 1'b0) : 1'b0);
assign n5880 = /* LUT   31 21  4 */ (\rco[183]  ? (n2369 ? (n2589 ? n2002 : 1'b0) : 1'b0) : 1'b0);
assign n5881 = /* LUT   27 15  1 */ n3545;
assign n5882 = /* LUT   15 14  3 */ n1785;
assign n5883 = /* LUT    3 20  4 */ n345;
assign n5884 = /* LUT   18 17  7 */ n2331;
assign n5885 = /* LUT   18 26  6 */ n2390;
assign n5886 = /* LUT    6 19  2 */ (\rco[123]  ? (n765 ? 1'b0 : (\rco[0]  ? n326 : 1'b0)) : 1'b0);
assign n5887 = /* LUT   28 19  3 */ n3779;
assign n5888 = /* LUT   19  9  5 */ n2475;
assign n5889 = /* LUT    4 10  4 */ n382;
assign n5890 = /* LUT    1 15  4 */ n73;
assign n5891 = /* LUT   22  6  7 */ n3002;
assign n5892 = /* LUT   10 16  6 */ n1029;
assign n5893 = /* LUT   13 10  5 */ n1438;
assign n5894 = /* LUT   13 21  4 */ n1516;
assign n5895 = /* LUT   18 12  3 */ n2288;
assign n5896 = /* LUT   21  6  0 */ n2669;
assign n5897 = /* LUT    6 13  1 */ n615;
assign n5898 = /* LUT   20 18  2 */ n2742;
assign n5899 = /* LUT   11  6  2 */ n1119;
assign n5900 = /* LUT   14 12  7 */ n1453;
assign n5901 = /* LUT   29  2  3 */ (\rco[48]  ? n2671 : 1'b0);
assign n5902 = /* LUT   19 10  1 */ n2479;
assign n5903 = /* LUT   22 16  0 */ n2894;
assign n5904 = /* LUT    5 22  7 */ n560;
assign n5905 = /* LUT   28 14  2 */ n3762;
assign n5906 = /* LUT   15 25  4 */ (n1877 ? \rco[183]  : 1'b0);
assign n5907 = /* LUT    7 13  2 */ (n809 ? \rco[153]  : 1'b0);
assign n5908 = /* LUT   21  8  3 */ n2842;
assign n5909 = /* LUT   26 17  4 */ n3549;
assign n5910 = /* LUT   12 17  2 */ n1313;
assign n5911 = /* LUT   26 10  5 */ n3515;
assign n5912 = /* LUT   18 30  3 */ n2419;
assign n5913 = /* LUT   14 19  3 */ (n1813 ? (n1684 ? n1667 : 1'b0) : 1'b0);
assign n5914 = /* LUT   17 14  7 */ n2100;
assign n5915 = /* LUT   29 20  6 */ n3873;
assign n5916 = /* LUT    5 13  1 */ n495;
assign n5917 = /* LUT   17 17  6 */ n2119;
assign n5918 = /* LUT   19 24  0 */ n2600;
assign n5919 = /* LUT   11 27  3 */ n1249;
assign n175  = /* LUT    1 11  1 */ (n31 ? !n56 : 1'b0);
assign n3142 = /* LUT   21 26  6 */ (n2044 ? (n2967 ? (n2563 ? n2400 : 1'b0) : 1'b0) : 1'b0);
assign n5920 = /* LUT   21 21  7 */ n2932;
assign n5921 = /* LUT   13 25  1 */ n1706;
assign n5922 = /* LUT   27 12  0 */ n3517;
assign n5923 = /* LUT   18 16  4 */ n2317;
assign n460  = /* LUT    3 21  3 */ (n117 ? (n459 ? (n120 ? n226 : 1'b0) : 1'b0) : 1'b0);
assign n5925 = /* LUT   18 29  7 */ n2408;
assign n5926 = /* LUT   11  9  0 */ (\rco[145]  ? (\rco[0]  ? (n989 ? n1031 : 1'b0) : 1'b0) : 1'b0);
assign n5927 = /* LUT   28 18  0 */ (\rco[31]  ? \rco[0]  : 1'b0);
assign n5928 = /* LUT   19  6  4 */ n2446;
assign n5929 = /* LUT    4  9  5 */ n375;
assign n5930 = /* LUT    9  9  3 */ n829;
assign n5931 = /* LUT   16 32  6 */ (n962 ? \rco[53]  : 1'b0);
assign n5932 = /* LUT   13 11  2 */ n1442;
assign n5933 = /* LUT   13 22  5 */ (n696 ? (\rco[0]  ? (n335 ? !n114 : 1'b1) : 1'b1) : 1'b1);
assign n5934 = /* LUT   18 15  2 */ n2311;
assign n5935 = /* LUT    6 12  2 */ n607;
assign n5936 = /* LUT   20 17  3 */ n2734;
assign n5937 = /* LUT   26 14  2 */ n3534;
assign n5938 = /* LUT   14 15  6 */ n1645;
assign n5939 = /* LUT    2  9  7 */ n163;
assign n5940 = /* LUT   20  4  7 */ n2656;
assign n5941 = /* LUT   17 29  3 */ (n2416 ? \rco[53]  : 1'b0);
assign n5942 = /* LUT   16  3  7 */ (\rco[83]  ? n1620 : 1'b0);
assign n5943 = /* LUT   19 11  2 */ n2487;
assign n5944 = /* LUT   23  9  1 */ n3176;
assign n3260 = /* LUT   22 19  1 */ (n1151 ? (n749 ? (n2344 ? !n2758 : 1'b1) : 1'b1) : 1'b1);
assign n5946 = /* LUT   10  5  2 */ n967;
assign n5947 = /* LUT   24 18  1 */ n3402;
assign n5948 = /* LUT    4 20  0 */ (n225 ? (n326 ? (n327 ? n336 : 1'b0) : 1'b0) : 1'b0);
assign n5949 = /* LUT   21  9  0 */ n2850;
assign n5950 = /* LUT    9 27  3 */ n948;
assign n5951 = /* LUT   12 16  5 */ n1308;
assign n5952 = /* LUT   26 13  4 */ n3530;
assign n5953 = /* LUT   29 21  5 */ n3879;
assign n5954 = /* LUT   17 15  0 */ n2108;
assign n5955 = /* LUT   20  7  3 */ n2663;
assign n5956 = /* LUT    5 14  0 */ n507;
assign n5957 = /* LUT   11 24  2 */ n1224;
assign n5958 = /* LUT   22 13  5 */ n3047;
assign n5959 = /* LUT   21 27  1 */ n2972;
assign n5960 = /* LUT   13 15  7 */ n1476;
assign n5961 = /* LUT   27  6  6 */ n2676;
assign n5962 = /* LUT    7 15  7 */ n745;
assign n5963 = /* LUT   21 22  6 */ n2941;
assign n5964 = /* LUT   13 26  0 */ n1718;
assign n5965 = /* LUT   18 19  5 */ n2343;
assign n5966 = /* LUT    3 18  2 */ n319;
assign n5967 = /* LUT    2 22  0 */ n242;
assign n5968 = /* LUT   18 28  4 */ n2403;
assign n5969 = /* LUT   11 22  1 */ n1206;
assign n5970 = /* LUT   28 17  1 */ n3766;
assign n5971 = /* LUT   16 15  2 */ n1944;
assign n5972 = /* LUT    5 16  4 */ n519;
assign n5973 = /* LUT   19  7  7 */ n2666;
assign n5974 = /* LUT   23 13  6 */ n3213;
assign n5975 = /* LUT   10 18  0 */ n1039;
assign n5976 = /* LUT    9 10  2 */ n835;
assign n5977 = /* LUT   13 12  3 */ n1451;
assign n5978 = /* LUT   15 18  0 */ n1814;
assign n5979 = /* LUT   20 27  5 */ n2818;
assign n5980 = /* LUT    6 15  3 */ n632;
assign n5981 = /* LUT   20 16  4 */ (n2886 ? (n2897 ? (n2740 ? n2729 : 1'b0) : 1'b0) : 1'b0);
assign n1511 = /* LUT   12 20  2 */ (n335 ? (n361 ? (n780 ? !n243 : 1'b1) : 1'b1) : 1'b1);
assign n5983 = /* LUT   14 14  1 */ n1632;
assign n5984 = /* LUT   17 11  5 */ n2072;
assign n5985 = /* LUT    1 16  2 */ n89;
assign n5986 = /* LUT   19  8  3 */ n2463;
assign n5987 = /* LUT   23 14  0 */ (n2740 ? (n2728 ? (\rco[0]  ? \rco[59]  : 1'b0) : 1'b0) : 1'b0);
assign n5988 = /* LUT   24 17  0 */ n2512;
assign n5989 = /* LUT    3 14  4 */ n292;
assign n5990 = /* LUT    7 19  0 */ (n326 ? (n336 ? (n244 ? n123 : 1'b0) : 1'b0) : 1'b0);
assign n5991 = /* LUT    9 20  2 */ n909;
assign n5992 = /* LUT   21 10  1 */ (n2457 ? (\rco[48]  ? n2671 : 1'b0) : 1'b0);
assign n5993 = /* LUT   26 19  6 */ n3560;
assign n5994 = /* LUT   27  9  4 */ n3613;
assign n5995 = /* LUT   12 23  4 */ n1361;
assign n5996 = /* LUT   26 12  7 */ n3522;
assign n5997 = /* LUT   17  8  1 */ (\rco[93]  ? (\rco[0]  ? n2239 : 1'b0) : 1'b0);
assign n5998 = /* LUT   20  6  0 */ n2660;
assign n5999 = /* LUT    4 12  7 */ n485;
assign n6000 = /* LUT   16 16  0 */ n1961;
assign n6001 = /* LUT   22 12  6 */ n3041;
assign n6002 = /* LUT   10 22  5 */ (n551 ? (n669 ? (n696 ? n769 : 1'b0) : 1'b0) : 1'b0);
assign n6003 = /* LUT   21 28  0 */ n2376;
assign n6004 = /* LUT   13 16  6 */ n1482;
assign n6005 = /* LUT   27  7  5 */ n3601;
assign n6006 = /* LUT    9 25  4 */ n225;
assign n6007 = /* LUT   27 10  6 */ (n1491 ? (n3750 ? (n1752 ? \rco[0]  : 1'b0) : 1'b0) : 1'b0);
assign n6008 = /* LUT   13 27  7 */ n1403;
assign n6009 = /* LUT   18 18  2 */ n2335;
assign n6010 = /* LUT    3 19  1 */ n330;
assign n6011 = /* LUT   20 20  1 */ n2761;
assign n6012 = /* LUT   23 18  2 */ n3243;
assign n6013 = /* LUT   14 10  6 */ n1609;
assign n6014 = /* LUT   11 23  2 */ n1215;
assign n6015 = /* LUT    5 17  7 */ n528;
assign n6016 = /* LUT    4 15  3 */ n414;
assign n6017 = /* LUT    1 10  7 */ n33;
assign n6018 = /* LUT   10 21  1 */ n1058;
assign n6019 = /* LUT   13 13  0 */ (\rco[23]  ? \rco[0]  : 1'b0);
assign n6020 = /* LUT   15 19  3 */ n1819;
assign n6021 = /* LUT   20 26  6 */ n2811;
assign n6022 = /* LUT   20 23  5 */ (\rco[0]  ? (n2953 ? (n2011 ? \rco[183]  : 1'b0) : 1'b0) : 1'b0);
assign n6023 = /* LUT    6 14  4 */ n626;
assign n6024 = /* LUT   12 27  3 */ n1259;
assign n6025 = /* LUT   17 20  4 */ n2139;
assign n6026 = /* LUT    2 11  5 */ n172;
assign n6027 = /* LUT   29  5  6 */ n3823;
assign n6028 = /* LUT   23 15  3 */ n3224;
assign n6029 = /* LUT   27 22  0 */ n2951;
assign n6030 = /* LUT    3 15  7 */ n419;
assign n6031 = /* LUT   21 16  7 */ n2893;
assign n6032 = /* LUT    7 16  1 */ n741;
assign n6033 = /* LUT    9 21  1 */ n914;
assign n6034 = /* LUT   21 11  6 */ n2864;
assign n6035 = /* LUT   26 18  1 */ (\rco[0]  ? n3664 : 1'b0);
assign n6036 = /* LUT   12  9  6 */ n1283;
assign n6037 = /* LUT   18 22  7 */ n2359;
assign n6038 = /* LUT   12 22  7 */ n1365;
assign n2271 = /* LUT   17  9  2 */ (\rco[23]  ? (n2270 ? n1933 : 1'b0) : 1'b0);
assign n6039 = /* LUT    6 24  0 */ (\rco[112]  ? n769 : 1'b0);
assign n6040 = /* LUT   20  5  1 */ n2659;
assign n6041 = /* LUT   10  9  3 */ n978;
assign n6042 = /* LUT   28 20  3 */ (n3259 ? \rco[162]  : 1'b0);
assign n6043 = /* LUT   22 15  7 */ n3229;
assign n6044 = /* LUT    7  6  0 */ n708;
assign n6045 = /* LUT    9  7  2 */ n824;
assign n6046 = /* LUT   13 17  5 */ n1488;
assign n6047 = /* LUT    9 26  5 */ n944;
assign n6048 = /* LUT   13 28  6 */ n1567;
assign n6049 = /* LUT   27 11  5 */ n3627;
assign n6050 = /* LUT   18 21  3 */ n2351;
assign n6051 = /* LUT    3 16  0 */ n307;
assign n6052 = /* LUT    6 10  1 */ n591;
assign n2865 = /* LUT   20 11  0 */ (n2494 ? (n2691 ? (n2706 ? n2857 : 1'b0) : 1'b0) : 1'b0);
assign n6054 = /* LUT   23 19  1 */ n3250;
assign n6055 = /* LUT   11 20  3 */ n1191;
assign n6056 = /* LUT   29  9  3 */ (n3175 ? \rco[74]  : 1'b0);
assign n6057 = /* LUT   17 27  2 */ n2189;
assign n6058 = /* LUT   28 23  7 */ n3811;
assign n6059 = /* LUT    5 18  6 */ n656;
assign n512  = /* LUT    4 14  0 */ (n398 ? (\rco[15]  ? (n194 ? n103 : 1'b0) : 1'b0) : 1'b0);
assign n6060 = /* LUT   19  5  1 */ n2223;
assign n6061 = /* LUT   22 25  2 */ n3126;
assign n6062 = /* LUT   10 20  2 */ n1049;
assign n6063 = /* LUT   13 14  1 */ n1462;
assign n6064 = /* LUT   15 16  2 */ n1794;
assign n6065 = /* LUT   21 15  3 */ (n1340 ? (n3067 ? 1'b0 : (n912 ? !n2593 : 1'b0)) : 1'b0);
assign n6066 = /* LUT   20 25  7 */ n2611;
assign n6067 = /* LUT   26 22  6 */ n3575;
assign n728  = /* LUT    6  9  5 */ (n717 ? (n590 ? !en_in : 1'b1) : 1'b1);
assign n6068 = /* LUT   20 22  6 */ n2781;
assign n6069 = /* LUT   12 26  0 */ n1391;
assign n6070 = /* LUT   14  8  3 */ n1595;
assign n6071 = /* LUT    2 10  2 */ n174;
assign n6072 = /* LUT    1 18  0 */ n101;
assign n6073 = /* LUT   17 21  7 */ n2150;
assign n6074 = /* LUT   17 24  4 */ n2169;
assign n6075 = /* LUT   23 12  2 */ n3201;
assign n6076 = /* LUT   27 23  3 */ (\rco[183]  ? (n3815 ? (n2796 ? \rco[0]  : 1'b0) : 1'b0) : 1'b0);
assign n6077 = /* LUT    3 12  6 */ n284;
assign n6078 = /* LUT   21 17  4 */ n2550;
assign n6079 = /* LUT   18  2  4 */ n2202;
assign n6080 = /* LUT    7 17  6 */ n756;
assign n6081 = /* LUT    9 22  0 */ n925;
assign n6082 = /* LUT   21 12  7 */ n3043;
assign n6083 = /* LUT   12  8  1 */ n1278;
assign n6084 = /* LUT   26 21  0 */ n3567;
assign n6085 = /* LUT   15  6  2 */ n1734;
assign n6086 = /* LUT   14 26  0 */ n1244;
assign n6087 = /* LUT   12 21  6 */ n1346;
assign n6088 = /* LUT   17 10  3 */ n2061;
assign n6089 = /* LUT    1 12  4 */ n49;
assign n6090 = /* LUT   22 14  0 */ n3056;
assign n6091 = /* LUT    7  7  3 */ n713;
assign n6092 = /* LUT   13 18  4 */ n1495;
assign n6093 = /* LUT   27  5  3 */ n3587;
assign n6094 = /* LUT   27  8  4 */ n3607;
assign n6095 = /* LUT   18 20  0 */ (n809 ? (\rco[153]  ? (n1151 ? n2344 : 1'b0) : 1'b0) : 1'b0);
assign n6096 = /* LUT    6 21  0 */ (\rco[110]  ? (n780 ? (\rco[0]  ? n243 : 1'b0) : 1'b0) : 1'b0);
assign n6097 = /* LUT   20 10  3 */ n2685;
assign n6098 = /* LUT   23 16  0 */ (\rco[29]  ? \rco[0]  : 1'b0);
assign n6099 = /* LUT   11 14  5 */ n1294;
assign n6100 = /* LUT   16  7  6 */ n1912;
assign n6101 = /* LUT   11 21  4 */ n1201;
assign n6102 = /* LUT   29 10  2 */ n3835;
assign n6103 = /* LUT   28 22  4 */ n3802;
assign n6104 = /* LUT    5 19  1 */ n539;
assign n502  = /* LUT    4 13  1 */ (n376 ? (n501 ? (n194 ? n398 : 1'b0) : 1'b0) : 1'b0);
assign n6105 = /* LUT   22 24  1 */ n3116;
assign n6106 = /* LUT   10 23  3 */ (\rco[99]  ? (n1222 ? 1'b0 : (n1090 ? !n1065 : 1'b0)) : 1'b0);
assign n6107 = /* LUT   30 12  2 */ n3895;
assign n6108 = /* LUT   15 17  5 */ n1805;
assign n6109 = /* LUT   18  6  1 */ n2231;
assign n6110 = /* LUT    7 21  3 */ n772;
assign n6111 = /* LUT    6  7  7 */ n581;
assign n6112 = /* LUT   20 24  0 */ n2599;
assign n6113 = /* LUT    6  8  6 */ n583;
assign n6114 = /* LUT   12 25  1 */ n1376;
assign n6115 = /* LUT   14 11  2 */ n1613;
assign n6116 = /* LUT   17 22  6 */ n2157;
assign n6117 = /* LUT   17 25  7 */ n2182;
assign n6118 = /* LUT   27 20  2 */ n3675;
assign n6119 = /* LUT    4 19  5 */ (n121 ? (n547 ? (n329 ? n350 : 1'b0) : 1'b0) : 1'b0);
assign n404  = /* LUT    3 13  1 */ (n181 ? (n73 ? n60 : 1'b0) : 1'b0);
assign n6120 = /* LUT   21 18  5 */ n2902;
assign n6121 = /* LUT   22 10  5 */ n3026;
assign n6122 = /* LUT   18  5  5 */ n2435;
assign n6123 = /* LUT    7 22  7 */ n789;
assign n6124 = /* LUT   21 13  4 */ n2877;
assign n6125 = /* LUT   12 15  0 */ n737;
assign n3683 = /* LUT   26 20  3 */ (n3241 ? (n3268 ? (n1409 ? n2759 : 1'b0) : 1'b0) : 1'b0);
assign n6127 = /* LUT   18 24  5 */ n2374;
assign n1845 = /* LUT   14 21  1 */ (n456 ? (n1844 ? (n658 ? n121 : 1'b0) : 1'b0) : 1'b0);
assign n6128 = /* LUT   19 30  2 */ n2635;
assign n6129 = /* LUT   11 17  1 */ n1168;
assign n1136 = /* LUT   10 11  1 */ (n989 ? (n1031 ? (n888 ? n1032 : 1'b0) : 1'b0) : 1'b0);
assign n6130 = /* LUT   16  8  4 */ n1918;
assign n6131 = /* LUT    1 13  7 */ n185;
assign n6132 = /* LUT   13 19  3 */ (\rco[99]  ? (n1673 ? 1'b0 : (n335 ? n1671 : 1'b0)) : 1'b0);
assign n6133 = /* LUT   15 21  2 */ n1837;
assign n6134 = /* LUT   20 28  5 */ n2827;
assign n6135 = /* LUT   18 23  1 */ n2362;
assign n6136 = /* LUT    6 20  3 */ n662;
assign n6137 = /* LUT   20  9  2 */ (n2470 ? (n2852 ? (n1934 ? !n2269 : 1'b1) : 1'b1) : 1'b1);
assign n6138 = /* LUT   23 17  7 */ n3232;
assign n6139 = /* LUT   11 15  6 */ n1158;
assign n6140 = /* LUT   26  6  3 */ n3475;
assign n6141 = /* LUT   14  7  5 */ n1589;
assign n6142 = /* LUT   16  6  5 */ n1901;
assign n6143 = /* LUT   11 18  5 */ n1183;
assign n6144 = /* LUT   29 11  5 */ n3843;
assign n6145 = /* LUT   28 21  5 */ n3795;
assign n6146 = /* LUT   19  3  3 */ n2429;
assign n6147 = /* LUT   22 27  0 */ n2967;
assign n6148 = /* LUT    3  9  6 */ n257;
assign n6149 = /* LUT   15 22  4 */ n1849;
assign n6150 = /* LUT   18  9  0 */ n2263;
assign n6151 = /* LUT    7 26  2 */ n799;
assign n6152 = /* LUT    9 19  4 */ n904;
assign n6153 = /* LUT   12 19  7 */ n1327;
assign n6154 = /* LUT   26  8  4 */ n3493;
assign n6155 = /* LUT    6 11  7 */ n602;
assign n6156 = /* LUT   12 24  6 */ n1372;
assign n6157 = /* LUT   17 23  1 */ n2160;
assign n6158 = /* LUT    2 12  0 */ n182;
assign n6159 = /* LUT   19 17  0 */ n2737;
assign n6160 = /* LUT   17 26  6 */ n2013;
assign n6161 = /* LUT   22 21  3 */ n3098;
assign n6162 = /* LUT   24 24  3 */ n3444;
assign n6163 = /* LUT   27 21  5 */ n3691;
assign n6164 = /* LUT    4 18  6 */ n435;
assign n6165 = /* LUT    3 10  0 */ n268;
assign n6166 = /* LUT   21 19  2 */ n2758;
assign n6167 = /* LUT   18  4  6 */ n2425;
assign n6168 = /* LUT   21 14  5 */ n2884;
assign n6169 = /* LUT    9 16  6 */ n878;
assign n6170 = /* LUT   12 14  3 */ n1290;
assign n6171 = /* LUT   26 23  2 */ n3577;
assign n6172 = /* LUT   18 27  4 */ n2396;
assign n6173 = /* LUT   14 20  2 */ n1677;
assign n6174 = /* LUT    5  8  2 */ n469;
assign n6175 = /* LUT   19 31  1 */ n2641;
assign n6176 = /* LUT   23 21  4 */ n3274;
assign n6177 = /* LUT   11 30  0 */ n1269;
assign n6178 = /* LUT   16 23  5 */ n1995;
assign n6179 = /* LUT    1 14  6 */ n75;
assign n6180 = /* LUT   22  8  2 */ n3020;
assign n6181 = /* LUT   13 20  2 */ n1504;
assign n6182 = /* LUT   15 10  3 */ n1753;
assign n6183 = /* LUT   20 19  4 */ n2752;
assign n6184 = /* LUT    6 23  2 */ n688;
assign n6185 = /* LUT   20  8  5 */ n2674;
assign n6186 = /* LUT   12 28  3 */ n1396;
assign n6187 = /* LUT   23 22  6 */ n3284;
assign n6188 = /* LUT   17 19  6 */ n2133;
assign n6189 = /* LUT   16  5  4 */ n1891;
assign n1336 = /* LUT   11 19  6 */ (n659 ? 1'b1 : (n1335 ? (n777 ? !n674 : 1'b1) : 1'b1));
assign n6191 = /* LUT   29 12  4 */ n3852;
assign n6192 = /* LUT   16 10  5 */ n1930;
assign n677  = /* LUT    5 21  3 */ (n669 ? (n550 ? (n551 ? n243 : 1'b0) : 1'b0) : 1'b0);
assign n6194 = /* LUT   27 17  2 */ n3773;
assign n6195 = /* LUT   15 24  6 */ n1870;
assign n6196 = /* LUT   21 23  7 */ n3111;
assign n6197 = /* LUT   15 23  7 */ n1858;
assign n6198 = /* LUT   18  8  3 */ n2251;
assign n6199 = /* LUT   12 18  4 */ n1323;
assign n6200 = /* LUT   26 11  5 */ n3512;
assign n6201 = /* LUT   17 16  0 */ (n813 ? (n880 ? (n206 ? n812 : 1'b0) : 1'b0) : 1'b0);
assign n302  = /* LUT    2 15  1 */ (n59 ? !n56 : 1'b0);
assign n6202 = /* LUT   19 14  1 */ n2513;
assign n6203 = /* LUT   22 20  0 */ n3094;
assign n6204 = /* LUT   10 14  3 */ n1012;
assign n6205 = /* LUT   24 23  2 */ n3434;
assign n6206 = /* LUT   28 10  2 */ n3742;
assign n6207 = /* LUT   27 18  4 */ n3660;
assign n6208 = /* LUT    3 11  3 */ n272;
assign n6209 = /* LUT    7  9  2 */ n719;
assign n6210 = /* LUT   21 20  3 */ n2920;
assign n6211 = /* LUT   18  7  7 */ n1896;
assign n6212 = /* LUT    7 20  5 */ (n777 ? (n660 ? 1'b1 : (n121 ? !n456 : 1'b1)) : 1'b1);
assign n6213 = /* LUT    9 17  5 */ n887;
assign n6214 = /* LUT   18 26  3 */ n2387;
assign n6215 = /* LUT   14 23  3 */ (n780 ? (n1861 ? \rco[99]  : 1'b0) : 1'b0);
assign n6216 = /* LUT   20 12  2 */ n2699;
assign n6217 = /* LUT    5  9  1 */ n471;
assign n6218 = /* LUT   19 28  0 */ n2623;
assign n6219 = /* LUT    1 15  1 */ (\rco[0]  ? n202 : 1'b0);
assign n6220 = /* LUT   22 11  3 */ (n2857 ? (n3198 ? (n2859 ? n2494 : 1'b0) : 1'b0) : 1'b0);
assign n6221 = /* LUT   13 21  1 */ n1513;
assign n6222 = /* LUT   30 10  1 */ n3885;
assign n6223 = /* LUT   15 11  0 */ n1759;
assign n6224 = /* LUT    6 13  4 */ n618;
assign n6225 = /* LUT   20 18  7 */ n2561;
assign n6226 = /* LUT    6 22  5 */ n679;
assign n6227 = /* LUT   20 15  4 */ n2720;
assign n6228 = /* LUT   23 23  5 */ n3291;
assign n6229 = /* LUT   11 13  0 */ n1140;
assign n6230 = /* LUT   11 16  7 */ n1165;
assign n6231 = /* LUT    5 22  2 */ n556;
assign n6232 = /* LUT   13  7  2 */ n1424;
assign n6233 = /* LUT   15 25  1 */ (n2003 ? \rco[183]  : 1'b0);
assign n6234 = /* LUT    7 13  7 */ n730;
assign n2495 = /* LUT   18 11  2 */ (n76 ? (n54 ? (n2270 ? n718 : 1'b0) : 1'b0) : 1'b0);
assign n6236 = /* LUT   15 20  6 */ n1832;
assign n6237 = /* LUT    7 24  0 */ n698;
assign n6238 = /* LUT   12 17  5 */ n1316;
assign n6239 = /* LUT   26 10  2 */ n3508;
assign n6240 = /* LUT   26  7  5 */ n3485;
assign n6241 = /* LUT   17 17  3 */ n2116;
assign n6242 = /* LUT   19 15  2 */ n2526;
assign n6243 = /* LUT   23  5  1 */ n3162;
assign n6244 = /* LUT   22 23  1 */ (\rco[162]  ? (n3295 ? (\rco[0]  ? n1710 : 1'b0) : 1'b0) : 1'b0);
assign n6245 = /* LUT   24 22  1 */ n3425;
assign n6246 = /* LUT   28  9  3 */ n3736;
assign n6247 = /* LUT   27 19  7 */ n3672;
assign n6248 = /* LUT    4 16  0 */ n409;
assign n6249 = /* LUT   21 21  0 */ n3101;
assign n6250 = /* LUT    9 18  4 */ n895;
assign n6251 = /* LUT   18 29  2 */ n2415;
assign n6252 = /* LUT   14 22  4 */ n1690;
assign n6253 = /* LUT   17  3  0 */ n2031;
assign n6254 = /* LUT    6 18  2 */ n650;
assign n6255 = /* LUT    5 10  0 */ (\rco[10]  ? \rco[0]  : 1'b0);
assign n6256 = /* LUT   23 27  6 */ n2183;
assign n6257 = /* LUT   23  6  5 */ n3151;
assign n6258 = /* LUT   11 28  2 */ n1256;
assign n6259 = /* LUT   10 12  4 */ n1000;
assign n6260 = /* LUT   24 25  5 */ n3450;
assign n6261 = /* LUT   16 21  7 */ n1985;
assign n6262 = /* LUT    1  8  0 */ n19;
assign n6263 = /* LUT   16 26  6 */ n2008;
assign n6264 = /* LUT   13 22  0 */ (\rco[0]  ? (n669 ? (\rco[99]  ? n335 : 1'b0) : 1'b0) : 1'b0);
assign n6265 = /* LUT   15  8  1 */ n1748;
assign n6266 = /* LUT    3 22  2 */ n358;
assign n6267 = /* LUT   21  7  4 */ (n3008 ? 1'b0 : (n2855 ? 1'b0 : \rco[23] ));
assign n6268 = /* LUT    2 18  0 */ n327;
assign n6269 = /* LUT    6 12  7 */ n612;
assign n6270 = /* LUT   20 17  6 */ n2739;
assign n6271 = /* LUT   26 14  7 */ n3539;
assign n6272 = /* LUT   23 20  4 */ n3266;
assign n3457 = /* LUT   24  7  1 */ (n3330 ? (n3174 ? (n3455 ? n2676 : 1'b0) : 1'b0) : 1'b0);
assign n6273 = /* LUT    9 14  2 */ n860;
assign n6274 = /* LUT    4 20  5 */ n444;
assign n6275 = /* LUT   21  9  5 */ n2849;
assign n6276 = /* LUT   18 10  5 */ n2277;
assign n6277 = /* LUT   12 16  2 */ n1310;
assign n6278 = /* LUT   26 13  3 */ n3529;
assign n6279 = /* LUT   14 18  1 */ n1661;
assign n6280 = /* LUT   19 25  4 */ n2607;
assign n6281 = /* LUT   17 18  2 */ n2336;
assign n6282 = /* LUT   19 12  3 */ n2499;
assign n6283 = /* LUT   23 10  0 */ n2285;
assign n6284 = /* LUT   22 22  6 */ n3108;
assign n6285 = /* LUT   24 21  0 */ (n3421 ? (n807 ? (n1409 ? n2759 : 1'b0) : 1'b0) : 1'b0);
assign n6286 = /* LUT   28  8  4 */ n3729;
assign n6287 = /* LUT    7 15  0 */ (\rco[23]  ? (n206 ? (n812 ? n813 : 1'b0) : 1'b0) : 1'b0);
assign n6288 = /* LUT    9 24  2 */ n933;
assign n6289 = /* LUT   21 22  1 */ n2935;
assign n6290 = /* LUT    2 22  5 */ n239;
assign n6291 = /* LUT   18 28  1 */ (n2628 ? n1709 : 1'b0);
assign n6292 = /* LUT   14 17  5 */ n1660;
assign n6293 = /* LUT   17 12  1 */ n2077;
assign n6294 = /* LUT   19 26  6 */ (n1541 ? (\rco[172]  ? (n1998 ? \rco[0]  : 1'b0) : 1'b0) : 1'b0);
assign n6295 = /* LUT   23 24  7 */ n3441;
assign n6296 = /* LUT   11 22  4 */ n1209;
assign n6297 = /* LUT   28 17  4 */ n3769;
assign n6298 = /* LUT   23  7  6 */ n3171;
assign n6299 = /* LUT   11 29  5 */ n1266;
assign n6300 = /* LUT   10 15  5 */ n1009;
assign n6301 = /* LUT   16 20  0 */ n1980;
assign n6302 = /* LUT   21 24  0 */ n3121;
assign n6303 = /* LUT   15 18  7 */ n1824;
assign n6304 = /* LUT   18 14  2 */ (n2248 ? (n2236 ? (n2091 ? n2266 : 1'b0) : 1'b0) : 1'b0);
assign n6305 = /* LUT    2 21  1 */ n227;
assign n6306 = /* LUT    6 15  6 */ n635;
assign n2896 = /* LUT   20 16  1 */ (n2550 ? n2722 : 1'b0);
assign n6307 = /* LUT   12 20  7 */ (\rco[0]  ? (n1043 ? (n338 ? \rco[118]  : 1'b0) : 1'b0) : 1'b0);
assign n6308 = /* LUT   20 13  6 */ n2711;
assign n6309 = /* LUT    4 11  3 */ n389;
assign n6310 = /* LUT   22 18  3 */ n3082;
assign n6311 = /* LUT   10 17  1 */ (n989 ? (\rco[145]  ? n1031 : 1'b0) : 1'b0);
assign n6312 = /* LUT    9 15  5 */ n871;
assign n6313 = /* LUT   24  6  2 */ n3322;
assign n6314 = /* LUT   28 12  1 */ n3753;
assign n6315 = /* LUT    7 19  5 */ n763;
assign n6316 = /* LUT   21 10  4 */ (n2680 ? (\rco[0]  ? (n2859 ? \rco[48]  : 1'b0) : 1'b0) : 1'b0);
assign n6317 = /* LUT   18 13  4 */ n2298;
assign n6318 = /* LUT    3 24  5 */ (\rco[123]  ? n465 : 1'b0);
assign n6319 = /* LUT   12 23  3 */ n1360;
assign n6320 = /* LUT   26 12  0 */ n3520;
assign n6321 = /* LUT   14 13  0 */ n1630;
assign n6322 = /* LUT    5 15  4 */ n517;
assign n6323 = /* LUT   23 11  3 */ n3192;
assign n6324 = /* LUT   11 25  2 */ n1232;
assign n6325 = /* LUT   22 17  7 */ n3078;
assign n6326 = /* LUT   24 20  7 */ n3405;
assign n6327 = /* LUT   16 16  5 */ n1967;
assign n6328 = /* LUT   13  6  6 */ n1422;
assign n6329 = /* LUT    4 22  2 */ (n113 ? (n564 ? (n122 ? n247 : 1'b0) : 1'b0) : 1'b0);
assign n6330 = /* LUT   15 13  3 */ n1779;
assign n6331 = /* LUT   20 20  6 */ n2749;
assign n6332 = /* LUT   14 16  6 */ n1651;
assign n6333 = /* LUT   17 13  2 */ n2087;
assign n6334 = /* LUT    5 12  6 */ n489;
assign n6335 = /* LUT   23 25  0 */ (\rco[183]  ? (\rco[0]  ? (n1876 ? n2797 : 1'b0) : 1'b0) : 1'b0);
assign n6336 = /* LUT   11 23  7 */ n1230;
assign n6337 = /* LUT   19 27  5 */ n2620;
assign n6338 = /* LUT   11 26  4 */ n1239;
assign n6339 = /* LUT   16 19  1 */ (n1684 ? n1813 : 1'b0);
assign n6340 = /* LUT    1 10  2 */ n29;
assign n6341 = /* LUT   21 25  3 */ n2964;
assign n6342 = /* LUT    9 11  2 */ n843;
assign n6343 = /* LUT   15 19  4 */ n1820;
assign n6344 = /* LUT   15 14  7 */ n1789;
assign n6345 = /* LUT    3 20  0 */ n347;
assign n6346 = /* LUT    2 20  2 */ n218;
assign n6347 = /* LUT   20 23  0 */ (\rco[183]  ? (\rco[0]  ? (n2002 ? n2369 : 1'b0) : 1'b0) : 1'b0);
assign n6348 = /* LUT    6 14  1 */ n623;
assign n1560 = /* LUT   12 27  6 */ (\rco[0]  ? (n1272 ? (n1244 ? !n1543 : 1'b1) : 1'b1) : 1'b1);
assign n6350 = /* LUT   18 17  3 */ n2327;
assign n6351 = /* LUT    6 19  6 */ (n446 ? (n668 ? (n658 ? !n667 : 1'b1) : 1'b1) : 1'b1);
assign n6352 = /* LUT   11  8  3 */ n1125;
assign n6353 = /* LUT   29  5  3 */ n3820;
assign n6354 = /* LUT   19  9  1 */ n2471;
assign n6355 = /* LUT    4 10  0 */ n386;
assign n6356 = /* LUT   24 16  4 */ n3387;
assign n6357 = /* LUT   27 22  7 */ n3701;
assign n6358 = /* LUT   10 16  2 */ n1024;
assign n6359 = /* LUT   13 10  1 */ n1434;
assign n6360 = /* LUT   18  3  6 */ (\rco[83]  ? n2054 : 1'b0);
assign n6361 = /* LUT   15 28  2 */ n1721;
assign n6362 = /* LUT    7 16  4 */ n744;
assign n6363 = /* LUT   21 11  3 */ n2861;
assign n6364 = /* LUT   18 12  7 */ n2292;
assign n6365 = /* LUT   21  6  4 */ n2836;
assign n6366 = /* LUT   12 22  0 */ n1353;
assign n6367 = /* LUT   26 15  1 */ n2122;
assign n1775 = /* LUT   14 12  3 */ (n1601 ? (n1752 ? n1460 : 1'b0) : 1'b0);
assign n6369 = /* LUT   19 23  6 */ (n2593 ? 1'b0 : (n2787 ? 1'b0 : (n1998 ? n2574 : 1'b0)));
assign n6370 = /* LUT   19 10  5 */ n2483;
assign n6371 = /* LUT    4 21  3 */ n449;
assign n6372 = /* LUT    9 26  0 */ n943;
assign n6373 = /* LUT   26 17  0 */ (\rco[36]  ? \rco[0]  : 1'b0);
assign n6374 = /* LUT   12  4  1 */ (\rco[145]  ? n990 : 1'b0);
assign n6375 = /* LUT    6 10  6 */ n598;
assign n6376 = /* LUT   20 11  7 */ n2712;
assign n6377 = /* LUT   17 14  3 */ n2096;
assign n6378 = /* LUT    5 13  5 */ n496;
assign n6379 = /* LUT   19 24  4 */ n2597;
assign n6380 = /* LUT   11 20  6 */ n1195;
assign n6381 = /* LUT   29  9  4 */ n3348;
assign n6382 = /* LUT   28 23  2 */ n3805;
assign n6383 = /* LUT   11 27  7 */ n1253;
assign n3141 = /* LUT   21 26  2 */ (n2044 ? (n2563 ? n2400 : 1'b0) : 1'b0);
assign n6385 = /* LUT   15 16  5 */ n1797;
assign n6386 = /* LUT   15 15  4 */ (n912 ? (n823 ? (\rco[0]  ? \rco[99]  : 1'b0) : 1'b0) : 1'b0);
assign n6387 = /* LUT   18 16  0 */ (\rco[23]  ? (n2533 ? n2113 : 1'b0) : 1'b0);
assign n6388 = /* LUT    6  9  0 */ (\rco[21]  ? \rco[0]  : 1'b0);
assign n6389 = /* LUT   20 22  3 */ n2778;
assign n6390 = /* LUT   12 26  5 */ n1389;
assign n6391 = /* LUT   17 24  3 */ n2168;
assign n6392 = /* LUT   19  6  0 */ n2236;
assign n6393 = /* LUT    4  9  1 */ n371;
assign n6394 = /* LUT   10  6  4 */ n976;
assign n6395 = /* LUT   24 15  5 */ n3381;
assign n6396 = /* LUT   10 19  3 */ n905;
assign n6397 = /* LUT    9  9  7 */ n980;
assign n6398 = /* LUT   13 11  6 */ n1446;
assign n6399 = /* LUT   18  2  1 */ n2199;
assign n6400 = /* LUT    7 17  3 */ n753;
assign n6401 = /* LUT   21 12  2 */ n2868;
assign n6402 = /* LUT   18 15  6 */ n2314;
assign n6403 = /* LUT   14 26  5 */ n1715;
assign n6404 = /* LUT   14 15  2 */ n1640;
assign n6405 = /* LUT    2  9  3 */ n159;
assign n6406 = /* LUT   20  4  3 */ n2239;
assign n6407 = /* LUT   19 20  7 */ n2571;
assign n6408 = /* LUT   19 11  6 */ n2491;
assign n6409 = /* LUT   23  9  5 */ n3180;
assign n3262 = /* LUT   22 19  5 */ (n817 ? (n1151 ? (\rco[0]  ? !n2344 : 1'b1) : 1'b1) : 1'b1);
assign n6411 = /* LUT   24 18  5 */ n3410;
assign n6412 = /* LUT    3 17  4 */ n313;
assign n6413 = /* LUT   14 25  1 */ n1701;
assign n6414 = /* LUT    6 21  7 */ (n672 ? (n782 ? (n325 ? \rco[110]  : 1'b0) : 1'b0) : 1'b0);
assign n6415 = /* LUT   17  4  5 */ n2220;
assign n6416 = /* LUT   17 15  4 */ n2103;
assign n6417 = /* LUT   20 10  4 */ n2686;
assign n6418 = /* LUT   20  7  7 */ n2667;
assign n6419 = /* LUT    5 14  4 */ n506;
assign n6420 = /* LUT   11 21  1 */ n1198;
assign n6421 = /* LUT   29 10  5 */ n3838;
assign n6422 = /* LUT   28 22  1 */ n3808;
assign n6423 = /* LUT   11 24  6 */ n1228;
assign n6424 = /* LUT   16 17  3 */ n1964;
assign n6425 = /* LUT   21 27  5 */ n2976;
assign n6426 = /* LUT   27  6  2 */ (n1752 ? (n3175 ? (\rco[66]  ? \rco[0]  : 1'b0) : 1'b0) : 1'b0);
assign n6427 = /* LUT   13 15  3 */ n1472;
assign n6428 = /* LUT   30 12  7 */ n3900;
assign n6429 = /* LUT   15 17  2 */ n1802;
assign n6430 = /* LUT   18  6  6 */ n2238;
assign n6431 = /* LUT   18 19  1 */ n2339;
assign n6432 = /* LUT    3 18  6 */ n323;
assign n6433 = /* LUT    6  8  3 */ n584;
assign n6434 = /* LUT   20 21  2 */ n2769;
assign n6435 = /* LUT   12 25  4 */ n1379;
assign n6436 = /* LUT    1 19  4 */ n107;
assign n6437 = /* LUT   17 25  0 */ n2044;
assign n6438 = /* LUT    5 16  0 */ n521;
assign n6439 = /* LUT   19  7  3 */ n2454;
assign n6440 = /* LUT   23 13  2 */ n3209;
assign n6441 = /* LUT   10 25  5 */ n1084;
assign n6442 = /* LUT   24 14  6 */ n3375;
assign n6443 = /* LUT   27 20  5 */ n3676;
assign n6444 = /* LUT   10 18  4 */ n1038;
assign n6445 = /* LUT    9 10  6 */ n839;
assign n6446 = /* LUT   18  5  0 */ n2440;
assign n6447 = /* LUT    7 22  2 */ n784;
assign n6448 = /* LUT   20 27  1 */ n2814;
assign n6449 = /* LUT   21 13  1 */ n2874;
assign n6450 = /* LUT   14 21  4 */ (\rco[110]  ? (\rco[0]  ? (n777 ? n1671 : 1'b0) : 1'b0) : 1'b0);
assign n6451 = /* LUT   14 14  5 */ n1636;
assign n6452 = /* LUT    2  8  0 */ n152;
assign n6453 = /* LUT    1 16  6 */ n86;
assign n6454 = /* LUT    6 26  3 */ n803;
assign n6455 = /* LUT   17 11  1 */ n2068;
assign n6456 = /* LUT   11 17  6 */ n1319;
assign n6457 = /* LUT   10 11  4 */ n993;
assign n6458 = /* LUT   19  8  7 */ n2467;
assign n6459 = /* LUT   19 21  0 */ n2581;
assign n6460 = /* LUT   23 14  4 */ n3219;
assign n6461 = /* LUT   24 17  4 */ n3397;
assign n6462 = /* LUT   28  7  1 */ n3719;
assign n410  = /* LUT    3 14  0 */ (n288 ? 1'b0 : (n59 ? (n56 ? 1'b0 : n403) : 1'b0));
assign n6463 = /* LUT   15 21  7 */ n1842;
assign n6464 = /* LUT   27  9  0 */ n3516;
assign n6465 = /* LUT   12 10  3 */ n1285;
assign n6466 = /* LUT   26 19  2 */ n3556;
assign n6467 = /* LUT   14 24  2 */ (\rco[99]  ? (n1874 ? (n1699 ? n1871 : 1'b0) : 1'b0) : 1'b0);
assign n6468 = /* LUT   17  5  6 */ (n2229 ? \rco[172]  : 1'b0);
assign n6469 = /* LUT    6 20  4 */ n663;
assign n2854 = /* LUT   20  9  5 */ (n2476 ? (n2689 ? (n2457 ? n2281 : 1'b0) : 1'b0) : 1'b0);
assign n2260 = /* LUT   17  8  5 */ (n1340 ? (n2259 ? (\rco[37]  ? n1933 : 1'b0) : 1'b0) : 1'b0);
assign n6471 = /* LUT    2  7  6 */ n149;
assign n6472 = /* LUT   23 28  3 */ (\rco[172]  ? (n3066 ? (n2539 ? n982 : 1'b0) : 1'b0) : 1'b0);
assign n6473 = /* LUT   11 18  0 */ n1036;
assign n6474 = /* LUT   29 11  2 */ n3840;
assign n6475 = /* LUT   28 21  0 */ n2942;
assign n6476 = /* LUT    4 12  3 */ n395;
assign n6477 = /* LUT   22 12  2 */ n3037;
assign n6478 = /* LUT   10 22  1 */ n1210;
assign n6479 = /* LUT   21 28  4 */ n2982;
assign n6480 = /* LUT   13 16  2 */ n1478;
assign n6481 = /* LUT   27  7  1 */ n3597;
assign n6482 = /* LUT   15 22  3 */ n1848;
assign n6483 = /* LUT   18  9  7 */ n2262;
assign n6484 = /* LUT   18 18  6 */ n2338;
assign n6485 = /* LUT    3 19  5 */ n333;
assign n6486 = /* LUT    6 11  2 */ n611;
assign n6487 = /* LUT   12 24  3 */ n1369;
assign n6488 = /* LUT   14 10  2 */ n1605;
assign n6489 = /* LUT   19 17  5 */ n2545;
assign n6490 = /* LUT   17 26  1 */ n2186;
assign n6491 = /* LUT   22 21  6 */ n3103;
assign n6492 = /* LUT    5 17  3 */ n526;
assign n6493 = /* LUT    4 15  7 */ n418;
assign n6494 = /* LUT   10 24  6 */ n1079;
assign n6495 = /* LUT   24 13  7 */ n3360;
assign n6496 = /* LUT   28 11  4 */ n3757;
assign n6497 = /* LUT   27 21  2 */ n3688;
assign n6498 = /* LUT   10 21  5 */ n1062;
assign n6499 = /* LUT   13 13  4 */ n1458;
assign n6500 = /* LUT   18  4  3 */ n2215;
assign n6501 = /* LUT    7 23  1 */ n790;
assign n6502 = /* LUT   20 26  2 */ n2806;
assign n6503 = /* LUT   21 14  0 */ n2901;
assign n6504 = /* LUT   14 20  7 */ n1834;
assign n6505 = /* LUT   17 20  0 */ n1979;
assign n6506 = /* LUT    2 11  1 */ n278;
assign n6507 = /* LUT   19 18  1 */ n2554;
assign n6508 = /* LUT   10 10  3 */ n985;
assign n6509 = /* LUT   23 15  7 */ n3228;
assign n6510 = /* LUT   28  6  2 */ n3712;
assign n6511 = /* LUT    3 15  3 */ n295;
assign n6512 = /* LUT   21 16  3 */ n2889;
assign n6513 = /* LUT   15 10  6 */ n1764;
assign n6514 = /* LUT   26 18  5 */ (\rco[23]  ? n3555 : 1'b0);
assign n2591 = /* LUT   18 22  3 */ (n1710 ? (n2590 ? (\rco[0]  ? !n2002 : 1'b1) : 1'b1) : 1'b1);
assign n6516 = /* LUT   14 27  3 */ n1694;
assign n6517 = /* LUT    6 23  5 */ n691;
assign n2844 = /* LUT   20  8  2 */ (n2281 ? n2669 : 1'b0);
assign n6518 = /* LUT   17  9  6 */ (n2054 ? (n2272 ? 1'b0 : (\rco[39]  ? n1340 : 1'b0)) : 1'b0);
assign n6519 = /* LUT   11 19  3 */ (\rco[0]  ? (n365 ? (n465 ? \rco[123]  : 1'b0) : 1'b0) : 1'b0);
assign n6520 = /* LUT   29 12  3 */ n3851;
assign n6521 = /* LUT   22 26  4 */ n3136;
assign n6522 = /* LUT    9 12  7 */ n852;
assign n6523 = /* LUT   27 17  7 */ n3652;
assign n6524 = /* LUT   22 15  3 */ n3060;
assign n6525 = /* LUT    7  6  4 */ n710;
assign n6526 = /* LUT   13 17  1 */ n1484;
assign n6527 = /* LUT   15 23  0 */ (\rco[114]  ? n243 : 1'b0);
assign n6528 = /* LUT   18  8  4 */ n2252;
assign n6529 = /* LUT   18 21  7 */ n2151;
assign n6530 = /* LUT    3 16  4 */ n306;
assign n6531 = /* LUT   14  5  3 */ n1573;
assign n6532 = /* LUT   19 14  4 */ n2516;
assign n6533 = /* LUT   22 20  5 */ n3092;
assign n6534 = /* LUT    5 18  2 */ n532;
assign n6535 = /* LUT    4 14  4 */ (n398 ? (n514 ? (n194 ? \rco[0]  : 1'b0) : 1'b0) : 1'b0);
assign n6536 = /* LUT   19  5  5 */ n2439;
assign n6537 = /* LUT   10 27  7 */ n946;
assign n6538 = /* LUT   24 12  0 */ n2895;
assign n6539 = /* LUT   16 24  6 */ n2001;
assign n6540 = /* LUT   22 25  6 */ n3131;
assign n6541 = /* LUT   10 20  6 */ n1054;
assign n6542 = /* LUT   27 18  3 */ n3659;
assign n6543 = /* LUT   13 14  5 */ n1466;
assign n6544 = /* LUT   28 10  7 */ n3747;
assign n6545 = /* LUT   18  7  2 */ (n2266 ? (n2460 ? (\rco[93]  ? \rco[0]  : 1'b0) : 1'b0) : 1'b0);
assign n6546 = /* LUT    7 20  0 */ (n769 ? (\rco[0]  ? (n114 ? n696 : 1'b0) : 1'b0) : 1'b0);
assign n6547 = /* LUT   20 25  3 */ n2800;
assign n6548 = /* LUT   26 22  2 */ n3570;
assign n6549 = /* LUT   15  5  4 */ n1728;
assign n1863 = /* LUT   14 23  6 */ (n1862 ? n1542 : 1'b0);
assign n6551 = /* LUT   20 12  7 */ n2704;
assign n6552 = /* LUT   14  8  7 */ n1746;
assign n6553 = /* LUT   17 21  3 */ n2146;
assign n6554 = /* LUT    1 18  4 */ n100;
assign n6555 = /* LUT   10 13  2 */ (n1031 ? (n912 ? (\rco[0]  ? \rco[99]  : 1'b0) : 1'b0) : 1'b0);
assign n6556 = /* LUT   24 26  1 */ n3454;
assign n6557 = /* LUT   23 12  6 */ n3206;
assign n6558 = /* LUT   28  5  3 */ n3707;
assign n6559 = /* LUT    3 12  2 */ n280;
assign n6560 = /* LUT   21 17  0 */ (\rco[59]  ? n2550 : 1'b0);
assign n6561 = /* LUT   26 24  7 */ n3561;
assign n6562 = /* LUT   30 10  6 */ n3891;
assign n6563 = /* LUT   15 11  5 */ n1767;
assign n6564 = /* LUT   26 21  4 */ n3565;
assign n6565 = /* LUT   15  6  6 */ n1740;
assign n6566 = /* LUT   17  7  0 */ n2248;
assign n6567 = /* LUT   18 25  2 */ n2378;
assign n6568 = /* LUT    6 22  2 */ n683;
assign n6569 = /* LUT   20 15  3 */ n2719;
assign n6570 = /* LUT   17 10  7 */ n2065;
assign n6571 = /* LUT   11 16  2 */ n1160;
assign n6572 = /* LUT    1 12  0 */ n181;
assign n6573 = /* LUT   24  8  5 */ (n3348 ? (n3337 ? n2681 : 1'b0) : 1'b0);
assign n6574 = /* LUT   13  7  7 */ n1429;
assign n6575 = /* LUT   22 14  4 */ n3054;
assign n6576 = /* LUT    7  7  7 */ n707;
assign n6577 = /* LUT   13 18  0 */ n114;
assign n6578 = /* LUT   27  5  7 */ n3591;
assign n6579 = /* LUT   30  9  0 */ (n3636 ? (\rco[66]  ? n3034 : 1'b0) : 1'b0);
assign n6580 = /* LUT   15 20  1 */ n1827;
assign n2496 = /* LUT   18 11  5 */ (n1934 ? (n2269 ? (\rco[37]  ? n1933 : 1'b0) : 1'b0) : 1'b0);
assign n6581 = /* LUT   18 20  4 */ (n736 ? (n2575 ? (\rco[0]  ? n738 : 1'b0) : 1'b0) : 1'b0);
assign n6582 = /* LUT   26  7  0 */ n3486;
assign n6583 = /* LUT   11 14  1 */ n1146;
assign n6584 = /* LUT    2 14  3 */ n189;
assign n6585 = /* LUT   16  7  2 */ n1908;
assign n6586 = /* LUT   19 15  7 */ n2525;
assign n6587 = /* LUT   23  5  6 */ n3319;
assign n6588 = /* LUT   22 23  4 */ (n2539 ? (n2173 ? (n3066 ? !n3101 : 1'b1) : 1'b1) : 1'b1);
assign n6589 = /* LUT    5 19  5 */ n543;
assign n503  = /* LUT    4 13  5 */ (n278 ? (n194 ? (n261 ? n398 : 1'b0) : 1'b0) : 1'b0);
assign n6591 = /* LUT   19  2  4 */ n2205;
assign n6592 = /* LUT   10 26  0 */ (\rco[99]  ? (\rco[0]  ? (n1090 ? n1221 : 1'b0) : 1'b0) : 1'b0);
assign n6593 = /* LUT   24 11  1 */ (n2740 ? (n2728 ? \rco[59]  : 1'b0) : 1'b0);
assign n6594 = /* LUT   13  4  3 */ (n1409 ? (n807 ? \rco[162]  : 1'b0) : 1'b0);
assign n6595 = /* LUT   22 24  5 */ n3119;
assign n6596 = /* LUT   10 23  7 */ n1070;
assign n6597 = /* LUT   27 19  0 */ n3673;
assign n6598 = /* LUT   28  9  6 */ n3740;
assign n6599 = /* LUT    6  7  3 */ n573;
assign n6600 = /* LUT   20 24  4 */ n2791;
assign n6601 = /* LUT   26  9  3 */ n3500;
assign n6602 = /* LUT   29 17  6 */ n3858;
assign n6603 = /* LUT   14 22  1 */ n1687;
assign n6604 = /* LUT   17  3  5 */ n2029;
assign n6605 = /* LUT    6 18  7 */ n655;
assign n6606 = /* LUT   14 11  6 */ n1618;
assign n6607 = /* LUT   17 22  2 */ n2153;
assign n6608 = /* LUT   19 16  3 */ (n2537 ? !n2333 : 1'b1);
assign n6609 = /* LUT   23  6  0 */ n3155;
assign n6610 = /* LUT   11 28  5 */ n1261;
assign n6611 = /* LUT   10 12  1 */ n997;
assign n6612 = /* LUT   24 25  0 */ n2603;
assign n6613 = /* LUT   16 26  3 */ n2187;
assign n6614 = /* LUT    4 19  1 */ (n546 ? \rco[127]  : 1'b0);
assign n6615 = /* LUT    3 13  5 */ (n103 ? (n407 ? (n194 ? \rco[0]  : 1'b0) : 1'b0) : 1'b0);
assign n6616 = /* LUT   21 18  1 */ n2907;
assign n6617 = /* LUT    9 28  2 */ n959;
assign n6618 = /* LUT   22 10  1 */ n3022;
assign n6619 = /* LUT   15  8  4 */ n1749;
assign n6620 = /* LUT   26 20  7 */ (n2574 ? (n3686 ? !\rco[0]  : 1'b1) : 1'b1);
assign n6621 = /* LUT   12 15  4 */ n1303;
assign n6622 = /* LUT   15  7  5 */ (\rco[83]  ? (n1623 ? \rco[0]  : 1'b0) : 1'b0);
assign n6623 = /* LUT   18 24  1 */ n2370;
assign n6624 = /* LUT   20 14  0 */ n2713;
assign n6625 = /* LUT   16  8  0 */ n1920;
assign n6626 = /* LUT    1 13  3 */ n63;
assign n6627 = /* LUT    5 23  2 */ (n114 ? n696 : 1'b0);
assign n6628 = /* LUT    9 14  5 */ n865;
assign n6629 = /* LUT   22  9  5 */ n3018;
assign n6630 = /* LUT   13 19  7 */ (n335 ? n1675 : 1'b0);
assign n6631 = /* LUT   18 10  2 */ n2274;
assign n6632 = /* LUT    2 17  1 */ n208;
assign n6633 = /* LUT   20 28  1 */ n2824;
assign n6634 = /* LUT   18 23  5 */ n2366;
assign n6635 = /* LUT   14 18  6 */ n1657;
assign n6636 = /* LUT   12 29  0 */ n1404;
assign n6637 = /* LUT   11 15  2 */ (n817 ? (\rco[0]  ? (n809 ? \rco[145]  : 1'b0) : 1'b0) : 1'b0);
assign n6638 = /* LUT   14  7  1 */ n1585;
assign n6639 = /* LUT   16  6  1 */ n1897;
assign n6640 = /* LUT   19 12  6 */ n2504;
assign n6641 = /* LUT   23 10  7 */ n3184;
assign n6642 = /* LUT   22 22  3 */ n3107;
assign n6643 = /* LUT   19  3  7 */ n2433;
assign n6644 = /* LUT   22 27  4 */ n3146;
assign n6645 = /* LUT   10 29  1 */ n1109;
assign n6646 = /* LUT   24 10  2 */ n3341;
assign n6647 = /* LUT   13  5  0 */ n1411;
assign n6648 = /* LUT   28  8  1 */ n3726;
assign n6649 = /* LUT    3  9  2 */ n253;
assign n6650 = /* LUT    9 19  0 */ n906;
assign n6651 = /* LUT   12 19  3 */ n1330;
assign n6652 = /* LUT   26  8  0 */ n3455;
assign n6653 = /* LUT   14 17  0 */ n1659;
assign n6654 = /* LUT   17 12  4 */ n2080;
assign n6655 = /* LUT    2 12  4 */ n179;
assign n6656 = /* LUT   23  7  3 */ n3168;
assign n6657 = /* LUT   11 29  2 */ n1272;
assign n6658 = /* LUT   10 15  0 */ n1016;
assign n6659 = /* LUT   16 25  2 */ n2004;
assign n6660 = /* LUT   21 24  7 */ n2784;
assign n6661 = /* LUT    4 18  2 */ n538;
assign n6662 = /* LUT    3 10  4 */ n265;
assign n6663 = /* LUT   21 19  6 */ n2914;
assign n6664 = /* LUT   13 23  4 */ n1527;
assign n6665 = /* LUT   27 14  5 */ n3645;
assign n6666 = /* LUT   15  9  3 */ n1755;
assign n6667 = /* LUT   18 14  7 */ n2041;
assign n6668 = /* LUT   12 14  7 */ n1149;
assign n6669 = /* LUT   26 23  6 */ n3582;
assign n6670 = /* LUT   18 27  0 */ n2398;
assign n6671 = /* LUT    6 16  0 */ n643;
assign n6672 = /* LUT   20 13  1 */ (n2270 ? (n2725 ? (n2510 ? !n2470 : 1'b1) : 1'b1) : 1'b1);
assign n6673 = /* LUT   23 21  0 */ n3268;
assign n6674 = /* LUT    4 11  6 */ n392;
assign n6675 = /* LUT   16 23  1 */ n1991;
assign n6676 = /* LUT    1 14  2 */ n69;
assign n6677 = /* LUT   22  7  7 */ n3003;
assign n6678 = /* LUT   10 17  4 */ n863;
assign n6679 = /* LUT    9 15  2 */ n868;
assign n6680 = /* LUT   24  6  7 */ n3173;
assign n6681 = /* LUT   22  8  6 */ n3015;
assign n6682 = /* LUT   28 12  6 */ n3748;
assign n6683 = /* LUT   13 20  6 */ n1508;
assign n6684 = /* LUT   31 17  0 */ n3408;
assign n6685 = /* LUT   18 13  3 */ n2297;
assign n6686 = /* LUT   20 19  0 */ n2756;
assign n6687 = /* LUT   14 13  7 */ n1627;
assign n6688 = /* LUT   14  6  6 */ n1582;
assign n6689 = /* LUT   16  5  0 */ n1583;
assign n6690 = /* LUT   17 19  2 */ n2129;
assign n6691 = /* LUT   19 13  1 */ n2302;
assign n6692 = /* LUT   23 11  4 */ n3193;
assign n6693 = /* LUT   22 17  2 */ n3073;
assign n6694 = /* LUT   10 28  2 */ n1102;
assign n6695 = /* LUT   24  9  3 */ n3334;
assign n6696 = /* LUT   13  6  1 */ n1415;
assign n6697 = /* LUT   15 24  2 */ n1865;
assign n6698 = /* LUT   21 23  3 */ n2945;
assign n6699 = /* LUT   12 18  0 */ n446;
assign n6700 = /* LUT   26 11  1 */ (n3525 ? \rco[66]  : 1'b0);
assign n6701 = /* LUT   30 21  2 */ n3572;
assign n6702 = /* LUT   14 16  3 */ n1648;
assign n6703 = /* LUT   17 13  7 */ n2084;
assign n6704 = /* LUT   29 19  0 */ n3866;
assign n6705 = /* LUT   17 16  4 */ (\rco[0]  ? n2323 : 1'b0);
assign n6706 = /* LUT    2 15  5 */ n199;
assign n6707 = /* LUT   11 26  3 */ n1238;
assign n6708 = /* LUT   21 25  4 */ n2965;
assign n6709 = /* LUT    9 11  7 */ n841;
assign n6710 = /* LUT    4 17  3 */ n428;
assign n6711 = /* LUT    3 11  7 */ n164;
assign n6712 = /* LUT    7  9  6 */ n723;
assign n6713 = /* LUT   21 20  7 */ n2919;
assign n6714 = /* LUT   13 24  5 */ (\rco[110]  ? (\rco[0]  ? (n114 ? n1337 : 1'b0) : 1'b0) : 1'b0);
assign n6715 = /* LUT   15 14  2 */ n1784;
assign n6716 = /* LUT   18 17  6 */ n2330;
assign n6717 = /* LUT   18 26  7 */ n2391;
assign n765  = /* LUT    6 19  1 */ (n327 ? (n121 ? (n244 ? !n336 : 1'b1) : 1'b1) : 1'b1);
assign n6719 = /* LUT   23 26  1 */ n3311;
assign n6720 = /* LUT   28 19  2 */ n3778;
assign n6721 = /* LUT   19  9  6 */ n2478;
assign n6722 = /* LUT    4 10  5 */ n264;
assign n6723 = /* LUT   16 22  2 */ n457;
assign n6724 = /* LUT   22  6  0 */ n2997;
assign n6725 = /* LUT   10 16  7 */ n1166;
assign n6726 = /* LUT   13 10  4 */ n1437;
assign n6727 = /* LUT   22 11  7 */ (n2470 ? (n3199 ? 1'b0 : (\rco[44]  ? n2859 : 1'b0)) : 1'b0);
assign n6728 = /* LUT   13 21  5 */ n1517;
assign n6729 = /* LUT   18 12  0 */ n2502;
assign n340  = /* LUT    2 19  3 */ (n120 ? (n225 ? (n226 ? \rco[0]  : 1'b0) : 1'b0) : 1'b0);
assign n6731 = /* LUT    6 13  0 */ n194;
assign n6732 = /* LUT   20 18  3 */ n2743;
assign n6733 = /* LUT   11  6  5 */ n1122;
assign n1776 = /* LUT   14 12  4 */ (n1602 ? 1'b0 : (n1775 ? \rco[0]  : 1'b0));
assign n6734 = /* LUT   11 13  4 */ n1143;
assign n6735 = /* LUT   19 10  0 */ n2484;
assign n6736 = /* LUT   22 16  1 */ n3070;
assign n6737 = /* LUT    5 22  6 */ n678;
assign n6738 = /* LUT   28 14  3 */ n3763;
assign n6739 = /* LUT   15 25  5 */ (\rco[183]  ? n1541 : 1'b0);
assign n6740 = /* LUT    7 13  3 */ (\rco[153]  ? n732 : 1'b0);
assign n6741 = /* LUT   12 17  1 */ n1312;
assign n6742 = /* LUT   18 30  4 */ n2420;
assign n6743 = /* LUT   14 19  2 */ n1665;
assign n6744 = /* LUT   17 14  6 */ n2099;
assign n6745 = /* LUT   29 20  1 */ n3868;
assign n6746 = /* LUT   17 17  7 */ n2117;
assign n6747 = /* LUT   11 27  0 */ n1390;
assign n6748 = /* LUT    1 11  2 */ (\rco[0]  ? n175 : 1'b0);
assign n6749 = /* LUT   21 26  5 */ (n2400 ? (n2563 ? (n2967 ? !n2044 : 1'b1) : 1'b1) : 1'b1);
assign n6750 = /* LUT    4 16  4 */ n423;
assign n6751 = /* LUT   21 21  4 */ n2929;
assign n6752 = /* LUT   13 25  6 */ n1539;
assign n6753 = /* LUT   27 12  7 */ n3630;
assign n6754 = /* LUT   18 16  5 */ n2318;
assign n6755 = /* LUT   18 29  6 */ n2413;
assign n6756 = /* LUT   23 27  2 */ n3313;
assign n6757 = /* LUT   28 18  1 */ n2124;
assign n6758 = /* LUT   19  6  7 */ n2449;
assign n6759 = /* LUT    4  9  4 */ n374;
assign n6760 = /* LUT    1  8  4 */ n30;
assign n6761 = /* LUT   10 19  6 */ n1046;
assign n6762 = /* LUT    9  9  0 */ n832;
assign n6763 = /* LUT   13 11  3 */ n1443;
assign n6764 = /* LUT   13 22  4 */ (\rco[0]  ? (\rco[99]  ? n335 : 1'b0) : 1'b0);
assign n6765 = /* LUT   18 15  1 */ n2310;
assign n6766 = /* LUT    2 18  4 */ n212;
assign n6767 = /* LUT    6 12  3 */ n608;
assign n6768 = /* LUT   20 17  2 */ n2733;
assign n6769 = /* LUT   26 14  3 */ n3535;
assign n6770 = /* LUT   14 15  5 */ n1643;
assign n6771 = /* LUT    2  9  6 */ n162;
assign n6772 = /* LUT   19 11  3 */ n2488;
assign n6773 = /* LUT   23  9  2 */ n3177;
assign n6774 = /* LUT   22 19  0 */ (\rco[153]  ? (n807 ? (n2574 ? \rco[0]  : 1'b0) : 1'b0) : 1'b0);
assign n6775 = /* LUT   21  9  1 */ n2845;
assign n6776 = /* LUT    9 27  4 */ n953;
assign n6777 = /* LUT   12 16  6 */ n1298;
assign n6778 = /* LUT   26 13  7 */ n3505;
assign n6779 = /* LUT   17 15  1 */ n2118;
assign n6780 = /* LUT   20  7  2 */ n2662;
assign n6781 = /* LUT   19 25  0 */ n2369;
assign n6782 = /* LUT   11 24  1 */ n1223;
assign n6783 = /* LUT   22 13  4 */ n3046;
assign n6784 = /* LUT   21 27  2 */ n2973;
assign n6785 = /* LUT    4 23  5 */ (\rco[132]  ? n462 : 1'b0);
assign n816  = /* LUT    7 15  4 */ (n76 ? (n815 ? (n718 ? n54 : 1'b0) : 1'b0) : 1'b0);
assign n6786 = /* LUT    9 24  6 */ n1077;
assign n6787 = /* LUT   13 26  7 */ n1549;
assign n6788 = /* LUT   21 22  5 */ n2939;
assign n6789 = /* LUT   27 13  0 */ n3638;
assign n6790 = /* LUT   15 12  0 */ n1631;
assign n6791 = /* LUT   18 19  4 */ n2342;
assign n6792 = /* LUT    2 22  1 */ n241;
assign n6793 = /* LUT   18 28  5 */ n2404;
assign n6794 = /* LUT   23 24  3 */ n3298;
assign n6795 = /* LUT   11 22  0 */ n1211;
assign n6796 = /* LUT   28 17  0 */ n3771;
assign n6797 = /* LUT   16 15  5 */ n1947;
assign n6798 = /* LUT   19  7  4 */ n2455;
assign n6799 = /* LUT   23 13  7 */ n3214;
assign n6800 = /* LUT   16 20  4 */ n2143;
assign n6801 = /* LUT   10 18  1 */ n1185;
assign n6802 = /* LUT    9 10  1 */ n834;
assign n6803 = /* LUT   13 12  2 */ n1450;
assign n6804 = /* LUT   15 18  3 */ n1810;
assign n6805 = /* LUT   20 27  4 */ n2817;
assign n6806 = /* LUT    2 21  5 */ n231;
assign n6807 = /* LUT    6 15  2 */ n631;
assign n1512 = /* LUT   12 20  3 */ (\rco[99]  ? (n1511 ? 1'b0 : (n114 ? n696 : 1'b0)) : 1'b0);
assign n6808 = /* LUT   14 14  2 */ n1633;
assign n6809 = /* LUT   17 11  6 */ n2073;
assign n6810 = /* LUT   17 30  1 */ n2197;
assign n6811 = /* LUT   19  8  2 */ n2462;
assign n6812 = /* LUT   23 14  3 */ n3218;
assign n6813 = /* LUT    3 14  7 */ (n301 ? n411 : 1'b0);
assign n6814 = /* LUT    7 19  1 */ n759;
assign n6815 = /* LUT    9 20  5 */ n910;
assign n6816 = /* LUT   21 10  0 */ (n2689 ? (\rco[48]  ? (n2671 ? n2457 : 1'b0) : 1'b0) : 1'b0);
assign n6817 = /* LUT   12 10  4 */ n1286;
assign n6818 = /* LUT   26 19  5 */ n3559;
assign n6819 = /* LUT   27  9  5 */ n3614;
assign n6820 = /* LUT   12 23  7 */ n1364;
assign n6821 = /* LUT   26 12  4 */ n3635;
assign n6822 = /* LUT   29 22  3 */ n3878;
assign n6823 = /* LUT   17  8  0 */ n810;
assign n6824 = /* LUT   20  6  1 */ n2839;
assign n6825 = /* LUT    5 15  0 */ (\rco[0]  ? \rco[7]  : 1'b0);
assign n6826 = /* LUT   19 22  1 */ n2584;
assign n6827 = /* LUT   16 16  1 */ n1960;
assign n6828 = /* LUT   22 12  7 */ n3042;
assign n6829 = /* LUT   21 28  3 */ n2981;
assign n6830 = /* LUT    4 22  6 */ (n225 ? (n226 ? (n122 ? n120 : 1'b0) : 1'b0) : 1'b0);
assign n6831 = /* LUT    9 25  5 */ n939;
assign n6832 = /* LUT   13 27  0 */ (\rco[99]  ? (\rco[0]  ? (n1543 ? n1272 : 1'b0) : 1'b0) : 1'b0);
assign n6833 = /* LUT   20 20  2 */ n2762;
assign n6834 = /* LUT   23 18  5 */ n3246;
assign n6835 = /* LUT   14 10  7 */ n1610;
assign n6836 = /* LUT   23 25  4 */ n3307;
assign n6837 = /* LUT   11 23  3 */ n1216;
assign n6838 = /* LUT    5 17  4 */ n527;
assign n6839 = /* LUT    4 15  2 */ n413;
assign n6840 = /* LUT   19  4  5 */ (\rco[145]  ? n1031 : 1'b0);
assign n6841 = /* LUT   16 19  5 */ n1973;
assign n6842 = /* LUT   10 21  0 */ n1063;
assign n6843 = /* LUT   13 13  1 */ n813;
assign n6844 = /* LUT   15 19  0 */ n1813;
assign n6845 = /* LUT   20 26  7 */ n2392;
assign n6846 = /* LUT    2 20  6 */ n223;
assign n6847 = /* LUT    6 14  5 */ n628;
assign n2953 = /* LUT   20 23  4 */ (n1876 ? (n2952 ? 1'b0 : (n2823 ? n2376 : 1'b0)) : 1'b0);
assign n6848 = /* LUT   12 27  2 */ (n1558 ? (n1559 ? (\rco[0]  ? \rco[99]  : 1'b0) : 1'b0) : 1'b0);
assign n6849 = /* LUT   17 20  7 */ n2142;
assign n6850 = /* LUT    2 11  4 */ n171;
assign n6851 = /* LUT   11  8  7 */ n1279;
assign n6852 = /* LUT   29  5  7 */ n3824;
assign n6853 = /* LUT   23 15  0 */ n3050;
assign n6854 = /* LUT   24 16  0 */ n1950;
assign n6855 = /* LUT   27 22  3 */ n3697;
assign n6856 = /* LUT    3 15  4 */ n296;
assign n6857 = /* LUT   21 16  6 */ n2892;
assign n6858 = /* LUT   18  3  2 */ (n1584 ? \rco[83]  : 1'b0);
assign n6859 = /* LUT    7 16  0 */ n746;
assign n6860 = /* LUT    9 21  6 */ n919;
assign n6861 = /* LUT   21 11  7 */ n3035;
assign n3665 = /* LUT   26 18  2 */ (n813 ? (n1960 ? n2119 : 1'b0) : 1'b0);
assign n6863 = /* LUT   12 22  4 */ n1351;
assign n6864 = /* LUT   26 15  5 */ n3544;
assign n6865 = /* LUT   17  9  3 */ (n1340 ? (n2271 ? (n2054 ? \rco[0]  : 1'b0) : 1'b0) : 1'b0);
assign n6866 = /* LUT   20  5  0 */ n2658;
assign n2786 = /* LUT   19 23  2 */ (n2602 ? 1'b1 : (n2784 ? (n2173 ? !n2229 : 1'b1) : 1'b1));
assign n6868 = /* LUT   28 20  4 */ (\rco[153]  ? (n3432 ? (\rco[0]  ? n2574 : 1'b0) : 1'b0) : 1'b0);
assign n6869 = /* LUT    4 24  0 */ (\rco[123]  ? (n465 ? n365 : 1'b0) : 1'b0);
assign n6870 = /* LUT   22 15  6 */ n3064;
assign n6871 = /* LUT    7  6  3 */ n709;
assign n6872 = /* LUT    9  7  3 */ n825;
assign n6873 = /* LUT    4 21  7 */ n362;
assign n6874 = /* LUT   13 28  1 */ n1561;
assign n6875 = /* LUT   27 11  2 */ n3624;
assign n6876 = /* LUT   18 21  2 */ n2350;
assign n6877 = /* LUT    6 10  2 */ n592;
assign n6878 = /* LUT   20 11  3 */ n2692;
assign n6879 = /* LUT   23 19  6 */ n3255;
assign n6880 = /* LUT   11 20  2 */ n1190;
assign n6881 = /* LUT   29  9  0 */ (n3348 ? \rco[74]  : 1'b0);
assign n6882 = /* LUT   17 27  3 */ n2190;
assign n6883 = /* LUT   28 23  6 */ n3813;
assign n6884 = /* LUT    5 18  5 */ n537;
assign n6885 = /* LUT    4 14  1 */ (n291 ? (n512 ? (n500 ? \rco[0]  : 1'b0) : 1'b0) : 1'b0);
assign n6886 = /* LUT   19  5  2 */ n2436;
assign n6887 = /* LUT   10 20  3 */ n1050;
assign n6888 = /* LUT   13 14  0 */ n668;
assign n6889 = /* LUT   15 16  1 */ n1793;
assign n3068 = /* LUT   21 15  4 */ (n2680 ? (n962 ? (n2510 ? !n2067 : 1'b1) : 1'b1) : 1'b1);
assign n6891 = /* LUT   20 25  6 */ n2804;
assign n6892 = /* LUT   26 22  7 */ n3583;
assign n6893 = /* LUT    6  9  4 */ n582;
assign n6894 = /* LUT   20 22  7 */ n2782;
assign n6895 = /* LUT   12 26  1 */ n1385;
assign n6896 = /* LUT   14  8  0 */ n1603;
assign n6897 = /* LUT   17 21  4 */ n2147;
assign n6898 = /* LUT   17 24  7 */ n2172;
assign n6899 = /* LUT   23 12  1 */ n3200;
assign n6900 = /* LUT   24 15  1 */ n3377;
assign n6901 = /* LUT    3 12  5 */ n283;
assign n6902 = /* LUT   21 17  5 */ n2898;
assign n6903 = /* LUT   18  2  5 */ n2203;
assign n6904 = /* LUT   21 12  6 */ n2873;
assign n6905 = /* LUT   26 21  3 */ n3564;
assign n6906 = /* LUT   14 26  1 */ n1711;
assign n6907 = /* LUT   12 21  5 */ n1345;
assign n6908 = /* LUT   17 10  2 */ n2060;
assign n6909 = /* LUT   19 20  3 */ n2567;
assign n1115 = /* LUT    9 32  1 */ (\rco[106]  ? (n803 ? n148 : 1'b0) : 1'b0);
assign n6910 = /* LUT    1 12  7 */ n52;
assign n6911 = /* LUT   22 14  1 */ n3051;
assign n6912 = /* LUT    7  7  0 */ (n717 ? (\rco[0]  ? en_in : 1'b0) : 1'b0);
assign n6913 = /* LUT   27  8  3 */ n3606;
assign n6914 = /* LUT   18 20  1 */ (\rco[153]  ? (n809 ? n1151 : 1'b0) : 1'b0);
assign n6915 = /* LUT    3 17  0 */ n315;
assign n6916 = /* LUT   14 25  5 */ n1705;
assign n6917 = /* LUT    6 21  3 */ (n243 ? (\rco[0]  ? (n674 ? n361 : 1'b0) : 1'b0) : 1'b0);
assign n6918 = /* LUT   17  4  1 */ n1886;
assign n6919 = /* LUT   23 16  7 */ (n3241 ? n3240 : 1'b0);
assign n6920 = /* LUT   11 14  4 */ n1292;
assign n6921 = /* LUT   20 10  0 */ n2688;
assign n6922 = /* LUT   14  4  5 */ (\rco[83]  ? n1623 : 1'b0);
assign n6923 = /* LUT   11 21  5 */ n1202;
assign n6924 = /* LUT   29 10  1 */ n3834;
assign n6925 = /* LUT   28 22  5 */ n3799;
assign n6926 = /* LUT   16 12  0 */ (n1759 ? (\rco[41]  ? n1772 : 1'b0) : 1'b0);
assign n6927 = /* LUT    5 19  2 */ n540;
assign n501  = /* LUT    4 13  0 */ (n386 ? (n261 ? (\rco[11]  ? n278 : 1'b0) : 1'b0) : 1'b0);
assign n6928 = /* LUT   16 17  7 */ n1969;
assign n1222 = /* LUT   10 23  2 */ (n1113 ? (\rco[0]  ? (n1087 ? !n1221 : 1'b1) : 1'b1) : 1'b1);
assign n6930 = /* LUT   30 12  3 */ n3896;
assign n6931 = /* LUT   15 17  6 */ n1807;
assign n6932 = /* LUT   18  6  2 */ n2232;
assign n6933 = /* LUT    7 21  4 */ n773;
assign n6934 = /* LUT    6  7  6 */ n578;
assign n6935 = /* LUT   20 24  1 */ n2788;
assign n6936 = /* LUT   26  9  6 */ n3503;
assign n6937 = /* LUT    6  8  7 */ n585;
assign n6938 = /* LUT   20 21  6 */ n2572;
assign n6939 = /* LUT   12 25  0 */ n1543;
assign n6940 = /* LUT   14 11  1 */ n1612;
assign n6941 = /* LUT   17 22  5 */ n2156;
assign n6942 = /* LUT    1 19  0 */ n122;
assign n6943 = /* LUT   17 25  4 */ n2179;
assign n6944 = /* LUT   10 25  1 */ n1080;
assign n6945 = /* LUT   24 14  2 */ n3370;
assign n6946 = /* LUT   27 20  1 */ n3682;
assign n547  = /* LUT    4 19  4 */ (\rco[99]  ? (n338 ? (n117 ? n545 : 1'b0) : 1'b0) : 1'b0);
assign n405  = /* LUT    3 13  2 */ (n289 ? (n404 ? n31 : 1'b0) : 1'b0);
assign n6947 = /* LUT   21 18  4 */ n2916;
assign n6948 = /* LUT   22 10  6 */ n3027;
assign n6949 = /* LUT   18  5  4 */ n2224;
assign n6950 = /* LUT    7 22  6 */ n788;
assign n6951 = /* LUT   21 13  5 */ n2880;
assign n6952 = /* LUT   26 20  0 */ (n3417 ? (\rco[162]  ? (n3432 ? n2942 : 1'b0) : 1'b0) : 1'b0);
assign n6953 = /* LUT   12 15  3 */ n1300;
assign n1844 = /* LUT   14 21  0 */ (n1683 ? n117 : 1'b0);
assign n6954 = /* LUT   19 30  5 */ n2638;
assign n6955 = /* LUT   19 21  4 */ n2579;
assign n6956 = /* LUT   11 17  2 */ n1169;
assign n6957 = /* LUT   10 11  0 */ n991;
assign n6958 = /* LUT   16  8  5 */ n1921;
assign n6959 = /* LUT    1 13  4 */ n64;
assign n6960 = /* LUT   28  7  5 */ n3723;
assign n6961 = /* LUT   16 29  2 */ (n114 ? \rco[116]  : 1'b0);
assign n6962 = /* LUT   22  9  0 */ (n2669 ? (\rco[48]  ? \rco[0]  : 1'b0) : 1'b0);
assign n6963 = /* LUT   15 21  3 */ n1838;
assign n6964 = /* LUT   20 28  6 */ n2828;
assign n6965 = /* LUT   18 23  0 */ n2367;
assign n2852 = /* LUT   20  9  1 */ (n1047 ? n2512 : 1'b0);
assign n6966 = /* LUT   23 17  0 */ (n2533 ? (\rco[29]  ? \rco[0]  : 1'b0) : 1'b0);
assign n6967 = /* LUT   11 15  7 */ n1139;
assign n6968 = /* LUT   26  6  4 */ n3476;
assign n6969 = /* LUT   14  7  4 */ n1588;
assign n6970 = /* LUT   11 18  4 */ n1182;
assign n6971 = /* LUT   29 11  6 */ n3844;
assign n6972 = /* LUT   28 21  4 */ n3794;
assign n6973 = /* LUT    5 20  3 */ n120;
assign n6974 = /* LUT   19  3  0 */ n2211;
assign n6975 = /* LUT    3  9  7 */ n258;
assign n6976 = /* LUT   15 22  7 */ n1984;
assign n6977 = /* LUT   18  9  3 */ n2249;
assign n6978 = /* LUT    9 19  5 */ n907;
assign n6979 = /* LUT   12 19  6 */ n1334;
assign n6980 = /* LUT   26  8  5 */ n3494;
assign n6981 = /* LUT    6 11  6 */ n605;
assign n6982 = /* LUT   12 24  7 */ n1373;
assign n6983 = /* LUT   17 23  2 */ n2161;
assign n6984 = /* LUT    2 12  1 */ n176;
assign n6985 = /* LUT   19 17  1 */ n2541;
assign n6986 = /* LUT   22 21  2 */ n3097;
assign n6987 = /* LUT   24 24  4 */ n3442;
assign n6988 = /* LUT   10 24  2 */ n1073;
assign n6989 = /* LUT   24 13  3 */ n3363;
assign n6990 = /* LUT   27 21  6 */ n3692;
assign n6991 = /* LUT    4 18  7 */ n436;
assign n6992 = /* LUT    3 10  3 */ n383;
assign n6993 = /* LUT    7  8  4 */ n711;
assign n6994 = /* LUT   21 19  3 */ n2912;
assign n6995 = /* LUT    9 16  1 */ n875;
assign n6996 = /* LUT   12 14  0 */ n1151;
assign n6997 = /* LUT   26 23  1 */ n3576;
assign n6998 = /* LUT   14 20  3 */ n1678;
assign n6999 = /* LUT   19 31  6 */ n2646;
assign n7000 = /* LUT   23 21  5 */ n3275;
assign n7001 = /* LUT   19 18  5 */ n2558;
assign n7002 = /* LUT   16 23  4 */ n1994;
assign n7003 = /* LUT    1 14  5 */ n72;
assign n7004 = /* LUT   28  6  6 */ n3717;
assign n7005 = /* LUT   15 10  2 */ n1760;
assign n7006 = /* LUT   20 19  7 */ n2755;
assign n7007 = /* LUT   17  6  3 */ n2040;
assign n7008 = /* LUT    6 23  1 */ n687;
assign n7009 = /* LUT   20  8  6 */ n2675;
assign n7010 = /* LUT   12 28  4 */ n1397;
assign n7011 = /* LUT   23 22  1 */ n3279;
assign n7012 = /* LUT   14  6  3 */ (\rco[83]  ? (\rco[0]  ? n1584 : 1'b0) : 1'b0);
assign n7013 = /* LUT   17 19  7 */ n2134;
assign n7014 = /* LUT   11 19  7 */ (n1196 ? (n1336 ? 1'b0 : (n335 ? n456 : 1'b0)) : 1'b0);
assign n7015 = /* LUT   29 12  7 */ n3846;
assign n7016 = /* LUT   16 10  2 */ n1927;
assign n675  = /* LUT    5 21  0 */ (n327 ? n225 : 1'b0);
assign n7018 = /* LUT   22 26  0 */ n2797;
assign n7019 = /* LUT    9 12  3 */ n851;
assign n7020 = /* LUT   27 17  3 */ n3653;
assign n7021 = /* LUT   15 24  5 */ n1869;
assign n7022 = /* LUT   15 23  4 */ n1855;
assign n7023 = /* LUT   18  8  0 */ n2256;
assign n7024 = /* LUT   12 18  5 */ n1324;
assign n7025 = /* LUT   26 11  4 */ n3511;
assign n2323 = /* LUT   17 16  3 */ (n1960 ? (n2109 ? \rco[23]  : 1'b0) : 1'b0);
assign n7026 = /* LUT    2 15  0 */ n289;
assign n7027 = /* LUT   19 14  0 */ (n813 ? (n2512 ? (n206 ? !n1047 : 1'b1) : 1'b1) : 1'b1);
assign n7028 = /* LUT   22 20  1 */ n3088;
assign n7029 = /* LUT   10 14  4 */ n1018;
assign n7030 = /* LUT   24 23  5 */ n3436;
assign n7031 = /* LUT   10 27  3 */ n1095;
assign n7032 = /* LUT   24 12  4 */ n3356;
assign n2174 = /* LUT   16 24  2 */ (n129 ? n457 : 1'b0);
assign n7033 = /* LUT   27 18  7 */ n3663;
assign n7034 = /* LUT   28 10  3 */ n3743;
assign n7035 = /* LUT    3 11  0 */ n275;
assign n7036 = /* LUT    7  9  3 */ n720;
assign n7037 = /* LUT   21 20  2 */ n3095;
assign n7038 = /* LUT   18  7  6 */ n2246;
assign n7039 = /* LUT    9 17  2 */ n884;
assign n7040 = /* LUT   15  5  0 */ n1730;
assign n1861 = /* LUT   14 23  2 */ (n1383 ? 1'b0 : (n1860 ? (n1542 ? n803 : 1'b0) : 1'b0));
assign n7041 = /* LUT   20 12  3 */ n2700;
assign n2760 = /* LUT   19 19  6 */ (\rco[99]  ? (n2574 ? (n912 ? n817 : 1'b0) : 1'b0) : 1'b0);
assign n203  = /* LUT    1 15  2 */ (n31 ? (n181 ? !n56 : 1'b0) : 1'b0);
assign n7042 = /* LUT   16 27  4 */ n2019;
assign n3198 = /* LUT   22 11  2 */ (n2680 ? (\rco[0]  ? \rco[48]  : 1'b0) : 1'b0);
assign n7043 = /* LUT   30 10  2 */ n3886;
assign n7044 = /* LUT   15 11  1 */ n1770;
assign n7045 = /* LUT    6 13  7 */ n621;
assign n7046 = /* LUT   20 18  4 */ n2744;
assign n7047 = /* LUT   17  7  4 */ n2049;
assign n7048 = /* LUT    6 22  6 */ n555;
assign n7049 = /* LUT   20 15  7 */ n2531;
assign n7050 = /* LUT   23 23  2 */ n3288;
assign n7051 = /* LUT   11 13  1 */ n1138;
assign n7052 = /* LUT   11 16  6 */ n1164;
assign n7053 = /* LUT    5 22  1 */ n561;
assign n7054 = /* LUT    9 13  0 */ n858;
assign n7055 = /* LUT   13  7  3 */ n1425;
assign n7056 = /* LUT   15 25  2 */ (n2002 ? \rco[183]  : 1'b0);
assign n7057 = /* LUT   18 11  1 */ (n1772 ? (\rco[41]  ? \rco[0]  : 1'b0) : 1'b0);
assign n7058 = /* LUT   15 20  5 */ n1831;
assign n7059 = /* LUT   12 17  4 */ n1315;
assign n7060 = /* LUT   26 10  3 */ n3509;
assign n7061 = /* LUT   26  7  4 */ n3484;
assign n7062 = /* LUT   17 17  0 */ n2101;
assign n7063 = /* LUT    5 24  0 */ n694;
assign n7064 = /* LUT   19 15  3 */ n2527;
assign n3295 = /* LUT   22 23  0 */ (n2539 ? (n2971 ? 1'b0 : (n3066 ? n3101 : 1'b0)) : 1'b0);
assign n7065 = /* LUT   23  5  2 */ n3156;
assign n7066 = /* LUT   24 22  6 */ n3431;
assign n7067 = /* LUT   10 26  4 */ (\rco[99]  ? (n1245 ? (n803 ? \rco[0]  : 1'b0) : 1'b0) : 1'b0);
assign n3467 = /* LUT   24 11  5 */ (n1491 ? (n3466 ? (n2679 ? 1'b0 : !n2307) : 1'b0) : 1'b0);
assign n7069 = /* LUT   27 19  4 */ n3670;
assign n7070 = /* LUT   28  9  2 */ n3735;
assign n7071 = /* LUT    4 16  1 */ n420;
assign n7072 = /* LUT   21 21  1 */ n2926;
assign n7073 = /* LUT    9 18  3 */ n894;
assign n7074 = /* LUT   14 22  5 */ n1691;
assign n7075 = /* LUT   17  3  1 */ n2025;
assign n7076 = /* LUT    6 18  3 */ n651;
assign n7077 = /* LUT   19 29  0 */ (\rco[183]  ? (n1816 ? (n1541 ? \rco[0]  : 1'b0) : 1'b0) : 1'b0);
assign n7078 = /* LUT   19 16  7 */ (n2533 ? (n2119 ? (n2552 ? n1960 : 1'b0) : 1'b0) : 1'b0);
assign n7079 = /* LUT   23  6  4 */ n3165;
assign n7080 = /* LUT   11 28  1 */ n1255;
assign n7081 = /* LUT   10 12  5 */ n1003;
assign n7082 = /* LUT   24 25  4 */ n3449;
assign n7083 = /* LUT    1  8  3 */ n16;
assign n7084 = /* LUT   27  1  0 */ (n3593 ? \rco[74]  : 1'b0);
assign n7085 = /* LUT   15  8  0 */ n1750;
assign n7086 = /* LUT    3 22  5 */ n357;
assign n7087 = /* LUT    2 18  1 */ n209;
assign n7088 = /* LUT    6 12  4 */ n609;
assign n7089 = /* LUT   20 17  5 */ n2736;
assign n7090 = /* LUT   23 20  3 */ n3265;
assign n7091 = /* LUT   24  7  0 */ (n3326 ? (n3456 ? (n3175 ? \rco[74]  : 1'b0) : 1'b0) : 1'b0);
assign n7092 = /* LUT    9 14  1 */ n859;
assign n7093 = /* LUT    4 20  6 */ n445;
assign n7094 = /* LUT   18 10  6 */ n2280;
assign n7095 = /* LUT   26 13  2 */ (n1491 ? (n3640 ? (\rco[0]  ? \rco[59]  : 1'b0) : 1'b0) : 1'b0);
assign n7096 = /* LUT   12 16  3 */ n1306;
assign n7097 = /* LUT   14 18  2 */ n1662;
assign n7098 = /* LUT   19 25  5 */ n2608;
assign n7099 = /* LUT   17 18  1 */ n2127;
assign n7100 = /* LUT   19 12  2 */ n2498;
assign n7101 = /* LUT   23 10  3 */ n3188;
assign n7102 = /* LUT   22 22  7 */ n3109;
assign n7103 = /* LUT   24 10  6 */ n3345;
assign n7104 = /* LUT   28  8  5 */ n3730;
assign n7105 = /* LUT    7 15  1 */ (\rco[25]  ? \rco[0]  : 1'b0);
assign n7106 = /* LUT   21 22  0 */ n2940;
assign n7107 = /* LUT   14 28  7 */ n1719;
assign n7108 = /* LUT    2 22  6 */ n247;
assign n7109 = /* LUT   14 17  4 */ n1663;
assign n7110 = /* LUT   17 12  0 */ n2091;
assign n7111 = /* LUT   19 26  1 */ (\rco[172]  ? (\rco[0]  ? (n1699 ? n1998 : 1'b0) : 1'b0) : 1'b0);
assign n7112 = /* LUT    5 11  0 */ n483;
assign n7113 = /* LUT   23 24  6 */ n3301;
assign n7114 = /* LUT   23  7  7 */ n3172;
assign n7115 = /* LUT   11 29  6 */ n1267;
assign n7116 = /* LUT   10 15  4 */ n1008;
assign n7117 = /* LUT   16 20  1 */ n1974;
assign n7118 = /* LUT   21 24  3 */ n2955;
assign n7119 = /* LUT   15 18  6 */ n1815;
assign n7120 = /* LUT   13 23  0 */ n669;
assign n7121 = /* LUT   27 14  1 */ n3641;
assign n2524 = /* LUT   18 14  3 */ (n2511 ? 1'b1 : !n2520);
assign n7123 = /* LUT   32  7  2 */ (n2669 ? \rco[48]  : 1'b0);
assign n7124 = /* LUT    2 21  0 */ n113;
assign n7125 = /* LUT   20 16  2 */ (\rco[48]  ? (n2896 ? (n2725 ? \rco[0]  : 1'b0) : 1'b0) : 1'b0);
assign n7126 = /* LUT    6 15  5 */ n634;
assign n7127 = /* LUT    6 16  4 */ n641;
assign n7128 = /* LUT   20 13  5 */ n2710;
assign n7129 = /* LUT    4 11  2 */ n388;
assign n7130 = /* LUT   22 18  4 */ n3083;
assign n7131 = /* LUT   22  7  3 */ n3000;
assign n7132 = /* LUT   10 17  0 */ (n1032 ? (\rco[145]  ? (n1031 ? n989 : 1'b0) : 1'b0) : 1'b0);
assign n7133 = /* LUT    9 15  6 */ n872;
assign n7134 = /* LUT   13  9  1 */ n1433;
assign n7135 = /* LUT   24  6  3 */ n3323;
assign n7136 = /* LUT   28 12  2 */ n3754;
assign n7137 = /* LUT   30 11  6 */ (n3636 ? (n3034 ? (\rco[66]  ? \rco[0]  : 1'b0) : 1'b0) : 1'b0);
assign n7138 = /* LUT   18 13  7 */ n2507;
assign n7139 = /* LUT   12 23  2 */ n1359;
assign n7140 = /* LUT   26 12  1 */ n3521;
assign n7141 = /* LUT   14 13  3 */ n1628;
assign n7142 = /* LUT    5 15  5 */ n518;
assign n7143 = /* LUT   19 22  4 */ n2587;
assign n7144 = /* LUT   19 13  5 */ n2301;
assign n7145 = /* LUT   23 11  0 */ n2706;
assign n7146 = /* LUT   11 25  3 */ n1233;
assign n7147 = /* LUT   22 17  6 */ n3077;
assign n7148 = /* LUT   24 20  0 */ n3418;
assign n7149 = /* LUT   16 16  6 */ n1965;
assign n7150 = /* LUT   10 28  6 */ n1106;
assign n7151 = /* LUT   24  9  7 */ n3347;
assign n7152 = /* LUT   13  6  5 */ n1419;
assign n7153 = /* LUT    4 22  3 */ (n462 ? (\rco[132]  ? n113 : 1'b0) : 1'b0);
assign n7154 = /* LUT   15 13  4 */ n1780;
assign n7155 = /* LUT   20 20  7 */ n2759;
assign n7156 = /* LUT   29 19  4 */ n3864;
assign n7157 = /* LUT   14 16  7 */ n1652;
assign n7158 = /* LUT   17 13  3 */ n2088;
assign n7159 = /* LUT    5 12  1 */ n399;
assign n7160 = /* LUT   19 27  2 */ n2617;
assign n7161 = /* LUT   11 23  4 */ n1217;
assign n7162 = /* LUT   23 25  1 */ n3305;
assign n7163 = /* LUT   11 26  7 */ n942;
assign n7164 = /* LUT   16 19  0 */ (n335 ? (n1671 ? \rco[99]  : 1'b0) : 1'b0);
assign n7165 = /* LUT    1 10  1 */ n28;
assign n7166 = /* LUT   21 25  0 */ n2968;
assign n7167 = /* LUT    9 11  3 */ n844;
assign n7168 = /* LUT   15 19  5 */ n1821;
assign n1700 = /* LUT   13 24  1 */ (n669 ? (n550 ? n335 : 1'b0) : 1'b0);
assign n7170 = /* LUT   15 14  6 */ n1788;
assign n7171 = /* LUT    3 20  7 */ n111;
assign n7172 = /* LUT    2 20  3 */ n219;
assign n7173 = /* LUT    6 14  2 */ n624;
assign n7174 = /* LUT   18 17  2 */ n2326;
assign n2952 = /* LUT   20 23  3 */ (n2797 ? (n2951 ? (n2603 ? !n2796 : 1'b1) : 1'b1) : 1'b1);
assign n7175 = /* LUT    6 19  5 */ (n667 ? (n767 ? (n668 ? !n446 : 1'b1) : 1'b1) : 1'b1);
assign n7176 = /* LUT   11  8  2 */ n1124;
assign n7177 = /* LUT   29  5  0 */ n2681;
assign n7178 = /* LUT   19  9  2 */ n2472;
assign n7179 = /* LUT    4 10  1 */ n379;
assign n7180 = /* LUT   24 16  5 */ n3388;
assign n7181 = /* LUT   27 22  6 */ n3700;
assign n7182 = /* LUT   22  6  4 */ n2993;
assign n7183 = /* LUT   10 16  3 */ n1025;
assign n7184 = /* LUT   13 10  0 */ n1439;
assign n7185 = /* LUT   18  3  5 */ (\rco[83]  ? (n2054 ? \rco[0]  : 1'b0) : 1'b0);
assign n7186 = /* LUT   31 22  5 */ (\rco[183]  ? (n2002 ? n2369 : 1'b0) : 1'b0);
assign n7187 = /* LUT   18 12  4 */ n2289;
assign n7188 = /* LUT   21  6  3 */ n2835;
assign n7189 = /* LUT   26 15  0 */ (\rco[33]  ? \rco[0]  : 1'b0);
assign n7190 = /* LUT   11  6  1 */ n974;
assign n7191 = /* LUT   12 22  1 */ n1348;
assign n1773 = /* LUT   14 12  0 */ (n1738 ? (n1578 ? (n1619 ? !n587 : 1'b1) : 1'b1) : 1'b1);
assign n7193 = /* LUT   19 23  7 */ (n1340 ? (n2602 ? 1'b0 : (n912 ? !n2593 : 1'b0)) : 1'b0);
assign n7194 = /* LUT   19 10  4 */ n2482;
assign n7195 = /* LUT    4 21  2 */ n448;
assign n7196 = /* LUT   26 17  3 */ n3548;
assign n7197 = /* LUT    6 10  7 */ n729;
assign n7198 = /* LUT   18 30  0 */ n2422;
assign n7199 = /* LUT   14 19  6 */ n1669;
assign n7200 = /* LUT   17 14  2 */ n2095;
assign n7201 = /* LUT   20 11  6 */ n2695;
assign n7202 = /* LUT    5 13  2 */ n493;
assign n7203 = /* LUT   19 24  3 */ n2596;
assign n7204 = /* LUT   11 20  5 */ n1193;
assign n7205 = /* LUT   29  9  5 */ n3829;
assign n7206 = /* LUT   29 20  5 */ n3872;
assign n7207 = /* LUT   11 27  4 */ n1250;
assign n7208 = /* LUT   21 26  1 */ (\rco[172]  ? (n2563 ? n2044 : 1'b0) : 1'b0);
assign n7209 = /* LUT   15 16  4 */ n1796;
assign n7210 = /* LUT   13 25  2 */ n1535;
assign n7211 = /* LUT   27 12  3 */ n3634;
assign n1953 = /* LUT   15 15  5 */ (n912 ? (n1620 ? (n1666 ? \rco[23]  : 1'b0) : 1'b0) : 1'b0);
assign n458  = /* LUT    3 21  0 */ (n244 ? n123 : 1'b0);
assign n7214 = /* LUT   18 16  1 */ n2533;
assign n7215 = /* LUT    6  9  3 */ (n154 ? (n727 ? \rco[0]  : 1'b0) : 1'b0);
assign n7216 = /* LUT   20 22  0 */ n2589;
assign n7217 = /* LUT   17 24  2 */ n2167;
assign n7218 = /* LUT   19  6  3 */ n2445;
assign n7219 = /* LUT    4  9  0 */ n377;
assign n7220 = /* LUT   10  6  5 */ n971;
assign n7221 = /* LUT   24 15  4 */ n3380;
assign n7222 = /* LUT   27 23  5 */ (\rco[172]  ? (n3124 ? (n1998 ? \rco[0]  : 1'b0) : 1'b0) : 1'b0);
assign n7223 = /* LUT   10 19  2 */ (n1043 ? (n137 ? n1044 : 1'b0) : 1'b0);
assign n7224 = /* LUT    9  9  4 */ n830;
assign n7225 = /* LUT   13 11  7 */ n1447;
assign n7226 = /* LUT   18  2  2 */ n2200;
assign n7227 = /* LUT   18 15  5 */ n2313;
assign n7228 = /* LUT   14 26  6 */ n1716;
assign n7229 = /* LUT   12 21  0 */ (\rco[99]  ? (n696 ? (n224 ? 1'b0 : n114) : 1'b0) : 1'b0);
assign n7230 = /* LUT   14 15  1 */ n1639;
assign n7231 = /* LUT    2  9  2 */ n161;
assign n7232 = /* LUT   20  4  4 */ n2653;
assign n7233 = /* LUT   19 20  6 */ n2570;
assign n7234 = /* LUT   19 11  7 */ n2492;
assign n7235 = /* LUT   23  9  6 */ n3181;
assign n7236 = /* LUT   22 19  4 */ n2909;
assign n7237 = /* LUT   10  5  1 */ n966;
assign n7238 = /* LUT   24 18  2 */ n3403;
assign n7239 = /* LUT    9 27  0 */ n1087;
assign n7240 = /* LUT   26 16  0 */ n3546;
assign n7241 = /* LUT    3 17  5 */ n314;
assign n7242 = /* LUT   14 25  0 */ n1707;
assign n782  = /* LUT    6 21  6 */ (n117 ? n121 : 1'b0);
assign n7244 = /* LUT   17  4  4 */ n2035;
assign n7245 = /* LUT   17 15  5 */ n2105;
assign n7246 = /* LUT   20 10  5 */ n2687;
assign n7247 = /* LUT   20  7  6 */ n2458;
assign n7248 = /* LUT    5 14  3 */ n510;
assign n7249 = /* LUT   29 21  6 */ n3883;
assign n7250 = /* LUT   11 21  2 */ n1199;
assign n7251 = /* LUT   29 10  4 */ n3837;
assign n7252 = /* LUT   11 24  5 */ n1227;
assign n7253 = /* LUT   16 17  2 */ n1970;
assign n7254 = /* LUT   22 13  0 */ (n2855 ? 1'b0 : (n2707 ? 1'b0 : \rco[23] ));
assign n7255 = /* LUT   21 27  6 */ n2978;
assign n7256 = /* LUT    9  5  1 */ (n758 ? (n823 ? \rco[145]  : 1'b0) : 1'b0);
assign n7257 = /* LUT   13 15  4 */ n1473;
assign n7258 = /* LUT   27  6  5 */ (\rco[74]  ? (n3330 ? n3455 : 1'b0) : 1'b0);
assign n7259 = /* LUT   30 12  4 */ n3897;
assign n7260 = /* LUT   15 17  3 */ n1803;
assign n7261 = /* LUT   13 26  3 */ n1546;
assign n7262 = /* LUT   18  6  7 */ n2450;
assign n7263 = /* LUT   27 13  4 */ n3637;
assign n7264 = /* LUT   18 19  0 */ n2345;
assign n7265 = /* LUT    3 18  1 */ n318;
assign n7266 = /* LUT    6  8  0 */ n590;
assign n7267 = /* LUT   20 21  1 */ n2768;
assign n7268 = /* LUT    1 19  5 */ n108;
assign n7269 = /* LUT   17 25  1 */ n2176;
assign n7270 = /* LUT   16 15  1 */ n1943;
assign n7271 = /* LUT   19  7  0 */ n2668;
assign n7272 = /* LUT   23 13  3 */ n3210;
assign n7273 = /* LUT   10 25  4 */ n1083;
assign n7274 = /* LUT   24 14  7 */ n3383;
assign n7275 = /* LUT   27 20  4 */ n3678;
assign n7276 = /* LUT   10 18  5 */ n1186;
assign n7277 = /* LUT    9 10  5 */ n838;
assign n7278 = /* LUT   13 12  6 */ n1448;
assign n7279 = /* LUT   18  5  3 */ n2228;
assign n7280 = /* LUT   20 27  0 */ n2823;
assign n7281 = /* LUT   14 21  7 */ (n1197 ? (n457 ? (n1520 ? 1'b0 : n129) : 1'b0) : 1'b0);
assign n7282 = /* LUT   14 14  6 */ n1638;
assign n7283 = /* LUT    2  8  1 */ n154;
assign n7284 = /* LUT    1 16  1 */ n88;
assign n7285 = /* LUT    6 26  4 */ n699;
assign n7286 = /* LUT   17 11  2 */ n2069;
assign n7287 = /* LUT   19 21  1 */ n2576;
assign n7288 = /* LUT   19  8  6 */ n2466;
assign n7289 = /* LUT   23 14  7 */ n3071;
assign n7290 = /* LUT   24 17  3 */ n3396;
assign n7291 = /* LUT   28  7  0 */ n3724;
assign n7292 = /* LUT    3 14  3 */ (n386 ? (\rco[12]  ? (\rco[0]  ? n261 : 1'b0) : 1'b0) : 1'b0);
assign n7293 = /* LUT    9 20  1 */ (\rco[99]  ? (n1056 ? 1'b0 : (n137 ? !n224 : 1'b0)) : 1'b0);
assign n7294 = /* LUT   27  9  1 */ n3610;
assign n7295 = /* LUT   12 10  0 */ (\rco[24]  ? \rco[0]  : 1'b0);
assign n7296 = /* LUT   26 19  1 */ n2537;
assign n7297 = /* LUT   14 24  3 */ (n335 ? (n456 ? n1592 : 1'b0) : 1'b0);
assign n7298 = /* LUT   17  5  7 */ (\rco[172]  ? n2037 : 1'b0);
assign n7299 = /* LUT    6 20  5 */ n664;
assign n7300 = /* LUT   20  9  4 */ (n2470 ? (n2853 ? 1'b0 : (n1933 ? n2306 : 1'b0)) : 1'b0);
assign n2259 = /* LUT   17  8  4 */ (n2030 ? (n2258 ? (n1578 ? n1420 : 1'b0) : 1'b0) : 1'b0);
assign n7301 = /* LUT   11 18  3 */ n1181;
assign n7302 = /* LUT   29 11  3 */ n3841;
assign n7303 = /* LUT    4 12  4 */ n396;
assign n7304 = /* LUT   22 12  3 */ n3038;
assign n7305 = /* LUT   10 22  2 */ (n669 ? (n550 ? (n769 ? n551 : 1'b0) : 1'b0) : 1'b0);
assign n7306 = /* LUT   21 28  7 */ n2985;
assign n7307 = /* LUT   13 16  5 */ n1481;
assign n7308 = /* LUT   27  7  6 */ n3602;
assign n7309 = /* LUT   15 22  2 */ n1847;
assign n3750 = /* LUT   27 10  5 */ (\rco[23]  ? (n2855 ? 1'b0 : !n2708) : 1'b0);
assign n7310 = /* LUT   13 27  4 */ n1554;
assign n7311 = /* LUT   18  9  6 */ n2268;
assign n7312 = /* LUT   18 18  7 */ n2125;
assign n7313 = /* LUT    3 19  2 */ (n327 ? \rco[0]  : 1'b0);
assign n7314 = /* LUT    6 11  1 */ n599;
assign n7315 = /* LUT   23 18  1 */ n3242;
assign n7316 = /* LUT   14 10  3 */ n1606;
assign n7317 = /* LUT   19 17  6 */ n2546;
assign n7318 = /* LUT    5 17  0 */ n648;
assign n7319 = /* LUT    4 15  6 */ n417;
assign n7320 = /* LUT   10 24  7 */ n938;
assign n7321 = /* LUT   24 13  6 */ n3367;
assign n7322 = /* LUT   28 11  7 */ (n3619 ? (n3636 ? (n3646 ? !n3622 : 1'b1) : 1'b1) : 1'b1);
assign n7323 = /* LUT   27 21  3 */ n3689;
assign n7324 = /* LUT   10 21  4 */ n1061;
assign n7325 = /* LUT   18  4  0 */ n2219;
assign n7326 = /* LUT   20 26  3 */ n2807;
assign n7327 = /* LUT   14 20  4 */ n1679;
assign n7328 = /* LUT   17 20  3 */ n2138;
assign n7329 = /* LUT    2 11  0 */ (\rco[0]  ? \rco[11]  : 1'b0);
assign n7330 = /* LUT   19 18  0 */ n2563;
assign n7331 = /* LUT   23 15  4 */ n3225;
assign n7332 = /* LUT   28  6  3 */ n3713;
assign n7333 = /* LUT    3 15  0 */ n299;
assign n7334 = /* LUT   21 16  2 */ n2888;
assign n7335 = /* LUT    9 21  2 */ n915;
assign n7336 = /* LUT   26 18  6 */ (n2534 ? (n3555 ? \rco[23]  : 1'b0) : 1'b0);
assign n7337 = /* LUT   18 22  4 */ (\rco[99]  ? (n2591 ? 1'b0 : (n912 ? !n2358 : 1'b0)) : 1'b0);
assign n7338 = /* LUT   20  8  3 */ (\rco[48]  ? (n2844 ? \rco[0]  : 1'b0) : 1'b0);
assign n7339 = /* LUT    6 23  4 */ n690;
assign n7340 = /* LUT   17  9  7 */ (n2236 ? (\rco[93]  ? (n2266 ? n2057 : 1'b0) : 1'b0) : 1'b0);
assign n7341 = /* LUT   11 19  0 */ (\rco[123]  ? (n365 ? (n1038 ? n465 : 1'b0) : 1'b0) : 1'b0);
assign n7342 = /* LUT   29 12  2 */ n3850;
assign n7343 = /* LUT   28 20  0 */ (n3785 ? \rco[162]  : 1'b0);
assign n7344 = /* LUT   22 26  5 */ n3137;
assign n7345 = /* LUT   22 15  2 */ n3059;
assign n7346 = /* LUT   13 17  6 */ n1490;
assign n7347 = /* LUT   15 23  1 */ n243;
assign n7348 = /* LUT   13 28  5 */ n1565;
assign n7349 = /* LUT   18  8  5 */ n2266;
assign n7350 = /* LUT   27 11  6 */ n3628;
assign n7351 = /* LUT   18 21  6 */ n2356;
assign n7352 = /* LUT    3 16  3 */ n305;
assign n7353 = /* LUT   23 19  2 */ n3251;
assign n7354 = /* LUT   14  5  2 */ n1572;
assign n7355 = /* LUT   19 14  7 */ n2716;
assign n7356 = /* LUT    5 18  1 */ n531;
assign n7357 = /* LUT    4 14  5 */ (n261 ? (n287 ? (n87 ? !n278 : 1'b1) : 1'b1) : 1'b1);
assign n7358 = /* LUT   19  5  6 */ n2442;
assign n7359 = /* LUT   10 27  6 */ n950;
assign n7360 = /* LUT   22 25  1 */ n3125;
assign n7361 = /* LUT   16 24  7 */ n2010;
assign n7362 = /* LUT   24 12  1 */ n3353;
assign n7363 = /* LUT   10 20  7 */ n1042;
assign n7364 = /* LUT   27 18  2 */ n3658;
assign n7365 = /* LUT   13 14  4 */ n1465;
assign n7366 = /* LUT   28 10  4 */ n3744;
assign n2460 = /* LUT   18  7  1 */ (n2248 ? n2239 : 1'b0);
assign n7367 = /* LUT   20 25  2 */ n2799;
assign n7368 = /* LUT   26 22  3 */ n3571;
assign n7369 = /* LUT   15  5  5 */ n1729;
assign n1862 = /* LUT   14 23  5 */ (n148 ? (n803 ? (n1113 ? n1231 : 1'b0) : 1'b0) : 1'b0);
assign n7371 = /* LUT   14  8  4 */ n1596;
assign n7372 = /* LUT   17 21  0 */ n2354;
assign n7373 = /* LUT   19 19  3 */ (\rco[162]  ? (n807 ? (n1409 ? \rco[0]  : 1'b0) : 1'b0) : 1'b0);
assign n7374 = /* LUT   23 12  5 */ n3204;
assign n7375 = /* LUT   28  5  2 */ n3706;
assign n7376 = /* LUT    3 12  1 */ n279;
assign n7377 = /* LUT   21 17  1 */ (n2726 ? \rco[59]  : 1'b0);
assign n7378 = /* LUT   30 10  7 */ n3893;
assign n7379 = /* LUT   12  8  6 */ n1134;
assign n7380 = /* LUT   26 21  7 */ n3694;
assign n7381 = /* LUT   15  6  1 */ n1733;
assign n7382 = /* LUT   17  7  1 */ n2046;
assign n7383 = /* LUT   18 25  5 */ n2381;
assign n7384 = /* LUT    6 22  3 */ n680;
assign n7385 = /* LUT   20 15  2 */ n2723;
assign n7386 = /* LUT   17 10  6 */ n2064;
assign n7387 = /* LUT   11 16  1 */ n1159;
assign n7388 = /* LUT    1 12  3 */ n48;
assign n7389 = /* LUT    9 13  5 */ n857;
assign n7390 = /* LUT   22 14  5 */ n3055;
assign n7391 = /* LUT    7  7  4 */ n714;
assign n7392 = /* LUT   13 18  7 */ n1498;
assign n7393 = /* LUT   27  5  0 */ n3456;
assign n7394 = /* LUT   18 11  4 */ (\rco[0]  ? (\rco[41]  ? (n1759 ? n1772 : 1'b0) : 1'b0) : 1'b0);
assign n7395 = /* LUT   15 20  0 */ n674;
assign n7396 = /* LUT   27  8  7 */ n3504;
assign n7397 = /* LUT   18 20  5 */ (n749 ? n732 : 1'b0);
assign n7398 = /* LUT   23 16  3 */ (\rco[0]  ? n3393 : 1'b0);
assign n7399 = /* LUT   11 14  0 */ n1152;
assign n7400 = /* LUT    2 14  4 */ n190;
assign n7401 = /* LUT   16  7  5 */ n1911;
assign n7402 = /* LUT   19 15  4 */ n2528;
assign n7403 = /* LUT   23  5  7 */ n3163;
assign n7404 = /* LUT   16 12  4 */ n1938;
assign n7405 = /* LUT    5 19  6 */ n431;
assign n7406 = /* LUT    4 13  4 */ (n398 ? (\rco[0]  ? (\rco[14]  ? n376 : 1'b0) : 1'b0) : 1'b0);
assign n7407 = /* LUT   22 24  2 */ n3117;
assign n7408 = /* LUT   10 26  1 */ (n1089 ? (\rco[0]  ? \rco[99]  : 1'b0) : 1'b0);
assign n7409 = /* LUT   24 11  0 */ (n2729 ? (n2740 ? (\rco[59]  ? n2728 : 1'b0) : 1'b0) : 1'b0);
assign n7410 = /* LUT   28  9  5 */ n3738;
assign n7411 = /* LUT   27 19  1 */ n3667;
assign n7412 = /* LUT   10 23  6 */ n1068;
assign n7413 = /* LUT    7 21  0 */ (n361 ? (n113 ? (n243 ? n550 : 1'b0) : 1'b0) : 1'b0);
assign n7414 = /* LUT    6  7  2 */ n572;
assign n7415 = /* LUT   20 24  5 */ n2792;
assign n7416 = /* LUT   26  9  2 */ n3499;
assign n7417 = /* LUT   14 22  2 */ n1688;
assign n7418 = /* LUT   17  3  6 */ n2212;
assign n7419 = /* LUT   14 11  5 */ n1616;
assign n7420 = /* LUT    2 13  6 */ n193;
assign n7421 = /* LUT   17 22  1 */ n2152;
assign n7422 = /* LUT   19 16  2 */ (n1960 ? (n2552 ? (n2119 ? !n2533 : 1'b1) : 1'b1) : 1'b1);
assign n7423 = /* LUT   23  6  3 */ n3161;
assign n7424 = /* LUT   11 28  4 */ n1258;
assign n7425 = /* LUT   16 26  0 */ n2014;
assign n546  = /* LUT    4 19  0 */ (n244 ? (n327 ? (n336 ? n326 : 1'b0) : 1'b0) : 1'b0);
assign n7427 = /* LUT    3 13  6 */ (n194 ? (n103 ? (n291 ? \rco[16]  : 1'b0) : 1'b0) : 1'b0);
assign n7428 = /* LUT   21 18  0 */ n2905;
assign n7429 = /* LUT   22 10  2 */ n3023;
assign n7430 = /* LUT    9 23  4 */ n928;
assign n7431 = /* LUT   12 15  7 */ n1304;
assign n3684 = /* LUT   26 20  4 */ (n3240 ? n3683 : 1'b0);
assign n7432 = /* LUT   18 24  6 */ n2383;
assign n7433 = /* LUT   20 14  1 */ n2714;
assign n7434 = /* LUT   19 30  1 */ n2634;
assign n7435 = /* LUT   16  8  1 */ n1915;
assign n7436 = /* LUT    1 13  0 */ (n31 ? (n60 ? (n181 ? n73 : 1'b0) : 1'b0) : 1'b0);
assign n7437 = /* LUT   24  7  7 */ (n3330 ? (n3155 ? (n3331 ? 1'b0 : n3326) : 1'b0) : 1'b0);
assign n7438 = /* LUT    9 14  4 */ n862;
assign n7439 = /* LUT   22  9  4 */ n3017;
assign n7440 = /* LUT   13 19  0 */ (n777 ? (n668 ? (n667 ? \rco[138]  : 1'b0) : 1'b0) : 1'b0);
assign n7441 = /* LUT   18 10  3 */ n2275;
assign n7442 = /* LUT    2 17  0 */ n317;
assign n7443 = /* LUT   20 28  2 */ (\rco[183]  ? (n2823 ? n1877 : 1'b0) : 1'b0);
assign n7444 = /* LUT   18 23  4 */ n2365;
assign n7445 = /* LUT   26  6  0 */ n3174;
assign n7446 = /* LUT   11 15  3 */ (\rco[145]  ? (\rco[0]  ? (n811 ? n817 : 1'b0) : 1'b0) : 1'b0);
assign n7447 = /* LUT   23 17  4 */ n3237;
assign n7448 = /* LUT   14  7  0 */ n1590;
assign n7449 = /* LUT   16  6  6 */ n1902;
assign n7450 = /* LUT   19 12  5 */ n2501;
assign n7451 = /* LUT   23 10  6 */ n3187;
assign n7452 = /* LUT   19  3  4 */ n2430;
assign n7453 = /* LUT   22 27  3 */ n3145;
assign n7454 = /* LUT   10 29  0 */ n1110;
assign n7455 = /* LUT   24 10  3 */ n3342;
assign n7456 = /* LUT   13  5  1 */ n1412;
assign n7457 = /* LUT   28  8  2 */ n3727;
assign n7458 = /* LUT    3  9  3 */ n254;
assign n7459 = /* LUT    7 26  1 */ n802;
assign n7460 = /* LUT    9 19  1 */ n901;
assign n7461 = /* LUT   12 19  2 */ n1329;
assign n7462 = /* LUT   26  8  1 */ n3490;
assign n7463 = /* LUT   14 17  3 */ n1656;
assign n7464 = /* LUT   17 12  7 */ n2083;
assign n7465 = /* LUT    2 12  5 */ n180;
assign n7466 = /* LUT   23  7  0 */ n3326;
assign n7467 = /* LUT   11 29  3 */ n1264;
assign n7468 = /* LUT   24 24  0 */ n3445;
assign n7469 = /* LUT   16 25  1 */ n129;
assign n7470 = /* LUT   21 24  6 */ n2958;
assign n7471 = /* LUT    4 18  3 */ n432;
assign n7472 = /* LUT    3 10  7 */ n267;
assign n7473 = /* LUT   21 19  7 */ n2913;
assign n7474 = /* LUT   13 23  5 */ n1528;
assign n7475 = /* LUT   27 14  4 */ n3644;
assign n7476 = /* LUT    9 16  5 */ n881;
assign n7477 = /* LUT   12 14  4 */ n1291;
assign n7478 = /* LUT   26 23  5 */ n3580;
assign n7479 = /* LUT   18 27  7 */ n2198;
assign n7480 = /* LUT    6 16  1 */ n638;
assign n7481 = /* LUT    5  8  1 */ n468;
assign n7482 = /* LUT   20 13  0 */ (n2680 ? (n2270 ? (n2470 ? !n2510 : 1'b1) : 1'b1) : 1'b1);
assign n7483 = /* LUT   19 31  2 */ n2642;
assign n7484 = /* LUT   23 21  1 */ n3271;
assign n7485 = /* LUT   16 23  0 */ n1996;
assign n7486 = /* LUT    1 14  1 */ n68;
assign n7487 = /* LUT   22  7  6 */ n3005;
assign n7488 = /* LUT   10 17  7 */ (n758 ? (n1178 ? (n1130 ? n1175 : 1'b0) : 1'b0) : 1'b0);
assign n7489 = /* LUT    9 15  3 */ n869;
assign n7490 = /* LUT   24  6  4 */ n3324;
assign n7491 = /* LUT   22  8  7 */ n3013;
assign n7492 = /* LUT   13 20  1 */ n1503;
assign n7493 = /* LUT   18 13  2 */ n2296;
assign n7494 = /* LUT   20 19  3 */ n2751;
assign n7495 = /* LUT   14 13  6 */ n1626;
assign n7496 = /* LUT   12 28  0 */ (\rco[102]  ? n1558 : 1'b0);
assign n7497 = /* LUT   23 22  5 */ n3283;
assign n7498 = /* LUT   14  6  7 */ n1410;
assign n7499 = /* LUT   16  5  7 */ n1894;
assign n7500 = /* LUT   17 19  3 */ n2130;
assign n7501 = /* LUT   19 13  2 */ n2508;
assign n7502 = /* LUT   23 11  5 */ n3194;
assign n7503 = /* LUT   16 10  6 */ n1932;
assign n7504 = /* LUT    5 21  4 */ (n117 ? (n677 ? n121 : 1'b0) : 1'b0);
assign n7505 = /* LUT   10 28  3 */ n1103;
assign n7506 = /* LUT   24  9  2 */ n3333;
assign n7507 = /* LUT   13  6  0 */ n1421;
assign n7508 = /* LUT   15 24  1 */ n1864;
assign n7509 = /* LUT   21 23  4 */ n2946;
assign n7510 = /* LUT   26 11  0 */ (\rco[66]  ? n3528 : 1'b0);
assign n7511 = /* LUT   12 18  1 */ n1320;
assign n7512 = /* LUT   29 19  1 */ n3861;
assign n7513 = /* LUT   14 16  0 */ n1175;
assign n7514 = /* LUT   17 13  4 */ n2089;
assign n7515 = /* LUT   17 16  7 */ (n2325 ? \rco[23]  : 1'b0);
assign n7516 = /* LUT    2 15  4 */ n198;
assign n7517 = /* LUT   11 26  2 */ n1237;
assign n7518 = /* LUT   10 14  0 */ n1013;
assign n7519 = /* LUT   24 23  1 */ n3433;
assign n7520 = /* LUT   21 25  5 */ n2966;
assign n7521 = /* LUT    4 17  2 */ n427;
assign n7522 = /* LUT    3 11  4 */ n273;
assign n7523 = /* LUT    7  9  7 */ n724;
assign n7524 = /* LUT   21 20  6 */ n2925;
assign n7525 = /* LUT    9 17  6 */ n892;
assign n7526 = /* LUT   18 26  0 */ n2400;
assign n7527 = /* LUT    6 19  0 */ n535;
assign n7528 = /* LUT   23 26  0 */ n2821;
assign n7529 = /* LUT   28 19  5 */ n3781;
assign n7530 = /* LUT   19  9  7 */ n2468;
assign n7531 = /* LUT   16 22  3 */ n1988;
assign n7532 = /* LUT   22  6  1 */ n2990;
assign n7533 = /* LUT   10 16  4 */ n1026;
assign n3199 = /* LUT   22 11  6 */ (\rco[0]  ? (n2494 ? (n2680 ? !n2510 : 1'b1) : 1'b1) : 1'b1);
assign n7535 = /* LUT   13 21  2 */ n1514;
assign n7536 = /* LUT   18 12  1 */ n2286;
assign n7537 = /* LUT    2 19  2 */ (n117 ? (n339 ? (n121 ? n338 : 1'b0) : 1'b0) : 1'b0);
assign n7538 = /* LUT    6 13  3 */ n617;
assign n7539 = /* LUT   20 18  0 */ n2746;
assign n7540 = /* LUT   11  6  4 */ n1121;
assign n7541 = /* LUT   14 12  5 */ (n1623 ? (n1776 ? (n587 ? n1738 : 1'b0) : 1'b0) : 1'b0);
assign n7542 = /* LUT   23 23  6 */ n3292;
assign n7543 = /* LUT   11 13  5 */ n1144;
assign n7544 = /* LUT   19 10  3 */ n2481;
assign n7545 = /* LUT   16  9  7 */ n1941;
assign n7546 = /* LUT    5 22  5 */ n559;
assign n7547 = /* LUT   28 14  0 */ n3044;
assign n7548 = /* LUT   15 25  6 */ n2011;
assign n7549 = /* LUT    3  7  1 */ n157;
assign n7550 = /* LUT    7 13  4 */ (n736 ? \rco[153]  : 1'b0);
assign n7551 = /* LUT   21  8  5 */ n2843;
assign n7552 = /* LUT   26 17  6 */ n3551;
assign n7553 = /* LUT   12 17  0 */ n465;
assign n7554 = /* LUT   18 30  5 */ n2421;
assign n7555 = /* LUT   14 19  1 */ (n668 ? (n1826 ? 1'b0 : n446) : 1'b0);
assign n7556 = /* LUT   17 14  5 */ n2098;
assign n7557 = /* LUT   29 20  0 */ n3420;
assign n7558 = /* LUT   17 17  4 */ n2120;
assign n7559 = /* LUT   11 27  1 */ n1247;
assign n7560 = /* LUT   24 22  2 */ n3426;
assign n7561 = /* LUT    1 11  3 */ n31;
assign n7562 = /* LUT   31 10  2 */ (\rco[66]  ? n3034 : 1'b0);
assign n7563 = /* LUT   21 26  4 */ n2822;
assign n7564 = /* LUT    4 16  5 */ n424;
assign n7565 = /* LUT   21 21  5 */ n2930;
assign n7566 = /* LUT   13 25  7 */ n1540;
assign n7567 = /* LUT   27 12  6 */ n3519;
assign n7568 = /* LUT    9 18  7 */ n898;
assign n7569 = /* LUT   18 29  1 */ n2414;
assign n7570 = /* LUT    5 10  3 */ n476;
assign n7571 = /* LUT   19 29  4 */ n2632;
assign n7572 = /* LUT   11  9  2 */ n1032;
assign n7573 = /* LUT   23 27  3 */ n3314;
assign n7574 = /* LUT   19  6  6 */ n2448;
assign n7575 = /* LUT   10 19  5 */ n1045;
assign n7576 = /* LUT    9  9  1 */ n827;
assign n7577 = /* LUT   13 22  3 */ (n550 ? (n669 ? (n335 ? \rco[99]  : 1'b0) : 1'b0) : 1'b0);
assign n7578 = /* LUT   18 15  0 */ (n2309 ? (n1934 ? n2218 : 1'b0) : 1'b0);
assign n7579 = /* LUT    3 22  1 */ n235;
assign n3007 = /* LUT   21  7  1 */ (n2270 ? (n2855 ? 1'b0 : \rco[23] ) : 1'b0);
assign n7580 = /* LUT    2 18  5 */ n213;
assign n7581 = /* LUT    6 12  0 */ n291;
assign n7582 = /* LUT   20 17  1 */ n2732;
assign n7583 = /* LUT   26 14  4 */ n3533;
assign n7584 = /* LUT   14 15  4 */ n1642;
assign n7585 = /* LUT   23 20  7 */ n3278;
assign n7586 = /* LUT   16  3  1 */ (\rco[83]  ? (n1584 ? n1578 : 1'b0) : 1'b0);
assign n7587 = /* LUT   19 11  0 */ n2067;
assign n7588 = /* LUT   23  9  3 */ n3178;
assign n7589 = /* LUT    4 20  2 */ (n327 ? (n326 ? (n113 ? n336 : 1'b0) : 1'b0) : 1'b0);
assign n7590 = /* LUT   21  9  6 */ n2851;
assign n7591 = /* LUT    9 27  5 */ n947;
assign n7592 = /* LUT    7 25  4 */ n801;
assign n7593 = /* LUT   21  4  5 */ (n2278 ? (\rco[44]  ? n2440 : 1'b0) : 1'b0);
assign n7594 = /* LUT   12 16  7 */ n1302;
assign n7595 = /* LUT   26 13  6 */ n3532;
assign n7596 = /* LUT   29 21  3 */ n3881;
assign n7597 = /* LUT   17 15  2 */ n2102;
assign n7598 = /* LUT   19 25  1 */ n2604;
assign n7599 = /* LUT   11 24  0 */ n1113;
assign n7600 = /* LUT   24 21  3 */ (\rco[162]  ? (n3432 ? (\rco[0]  ? n2942 : 1'b0) : 1'b0) : 1'b0);
assign n7601 = /* LUT   22 13  7 */ n3049;
assign n7602 = /* LUT   21 27  3 */ n2974;
assign n7603 = /* LUT    7 15  5 */ (n813 ? (n816 ? n206 : 1'b0) : 1'b0);
assign n7604 = /* LUT    9 24  1 */ n932;
assign n7605 = /* LUT   13 26  6 */ n1717;
assign n7606 = /* LUT   21 22  4 */ n2938;
assign n7607 = /* LUT   14 28  3 */ n1722;
assign n7608 = /* LUT    2 22  2 */ n236;
assign n7609 = /* LUT   18 28  2 */ n1709;
assign n7610 = /* LUT   19 26  5 */ (\rco[172]  ? (n1877 ? (\rco[0]  ? n1998 : 1'b0) : 1'b0) : 1'b0);
assign n7611 = /* LUT   23 24  2 */ n3297;
assign n7612 = /* LUT   11 22  3 */ n1208;
assign n7613 = /* LUT   28 17  7 */ n3856;
assign n7614 = /* LUT   16 15  4 */ n1946;
assign n7615 = /* LUT   19  7  5 */ n2456;
assign n7616 = /* LUT   16 20  5 */ n1978;
assign n7617 = /* LUT   10 18  2 */ n1033;
assign n7618 = /* LUT    9 10  0 */ n847;
assign n7619 = /* LUT   15 18  2 */ n1809;
assign n7620 = /* LUT   20 27  7 */ n2820;
assign n7621 = /* LUT    2 21  4 */ n230;
assign n7622 = /* LUT   20 16  6 */ (\rco[48]  ? (\rco[0]  ? (n2725 ? n2550 : 1'b0) : 1'b0) : 1'b0);
assign n7623 = /* LUT    6 15  1 */ n740;
assign n7624 = /* LUT   12 20  4 */ (n338 ? (n1512 ? \rco[0]  : 1'b0) : 1'b0);
assign n7625 = /* LUT   14 14  3 */ n1634;
assign n7626 = /* LUT   17 11  7 */ n1935;
assign n7627 = /* LUT   17 30  0 */ n2407;
assign n7628 = /* LUT   19  8  1 */ n2461;
assign n7629 = /* LUT   23 14  2 */ (n2519 ? (n2728 ? (n2740 ? n2729 : 1'b0) : 1'b0) : 1'b0);
assign n7630 = /* LUT   22 18  0 */ n3085;
assign n411  = /* LUT    3 14  6 */ (n31 ? (n285 ? (n56 ? 1'b0 : n289) : 1'b0) : 1'b0);
assign n7631 = /* LUT    7 19  6 */ n764;
assign n7632 = /* LUT    9 20  4 */ (n224 ? 1'b0 : (n1057 ? 1'b0 : (n117 ? \rco[99]  : 1'b0)));
assign n7633 = /* LUT   21 10  7 */ (n1491 ? (n3030 ? (n2725 ? n1752 : 1'b0) : 1'b0) : 1'b0);
assign n7634 = /* LUT   26 19  4 */ n3558;
assign n7635 = /* LUT   27  9  6 */ n3615;
assign n7636 = /* LUT   12 23  6 */ n1363;
assign n7637 = /* LUT   26 12  5 */ n3523;
assign n2258 = /* LUT   17  8  3 */ (n1738 ? (n2257 ? 1'b0 : n1619) : 1'b0);
assign n7638 = /* LUT    5 15  1 */ n301;
/* FF 24 20  4 */ always @(posedge clk) if (n3411) n3416 <= 1'b0 ? 1'b0 : n3911;
/* FF 16 16  2 */ always @(posedge clk) if (n2110) n1957 <= 1'b0 ? 1'b0 : n3912;
/* FF 22 12  4 */ always @(posedge clk) if (n3029) n3040 <= 1'b0 ? 1'b0 : n3913;
/* FF 10 22  7 */ assign n779 = n3914;
/* FF 21 28  2 */ always @(posedge clk) if (n2196) n2981 <= 1'b0 ? 1'b0 : n3915;
/* FF  4 22  7 */ assign \rco[134]  = n3916;
/* FF 13 27  1 */ always @(posedge clk) if (n1532) n1543 <= 1'b0 ? 1'b0 : n3917;
/* FF 27 10  0 */ assign \rco[70]  = n3918;
/* FF 15 13  0 */ always @(posedge clk) if (n1015) n1777 <= 1'b0 ? 1'b0 : n3919;
/* FF 20 20  3 */ always @(posedge clk) if (n2562) n2764 <= 1'b0 ? 1'b0 : n3920;
/* FF 23 18  4 */ always @(posedge clk) if (n2573) n3246 <= 1'b0 ? 1'b0 : n3921;
/* FF  5 12  5 */ always @(posedge clk) if (n77) n489 <= 1'b0 ? 1'b0 : n3922;
/* FF 19 27  6 */ always @(posedge clk) if (n2614) n2622 <= 1'b0 ? 1'b0 : n3923;
/* FF 11 23  0 */ always @(posedge clk) if (n796) n1214 <= 1'b0 ? 1'b0 : n3924;
/* FF 23 25  5 */ always @(posedge clk) if (n2613) n3307 <= 1'b0 ? 1'b0 : n3925;
/* FF 16 19  4 */ always @(posedge clk) if (n1402) n1684 <= 1'b0 ? 1'b0 : n3926;
/* FF  1 10  5 */ always @(posedge clk) if (n37) n33 <= 1'b0 ? 1'b0 : n3927;
/* FF 10 21  3 */ always @(posedge clk) if (n818) n1061 <= 1'b0 ? 1'b0 : n3928;
/* FF 15 19  1 */ always @(posedge clk) if (n1355) n1818 <= 1'b0 ? 1'b0 : n3929;
/* FF 20 26  4 */ always @(posedge clk) if (n2615) n2809 <= 1'b0 ? 1'b0 : n3930;
/* FF  3 20  3 */ always @(posedge clk) if (n119) n345 <= 1'b0 ? 1'b0 : n3931;
/* FF  2 20  7 */ always @(posedge clk) if (n126) n223 <= 1'b0 ? 1'b0 : n3932;
/* FF  6 14  6 */ always @(posedge clk) if (n78) n628 <= 1'b0 ? 1'b0 : n3933;
/* FF 20 23  7 */ assign n1877 = n3934;
/* FF 12 27  5 */ assign n1384 = n3935;
/* FF 17 20  6 */ always @(posedge clk) if (n1843) n2142 <= 1'b0 ? 1'b0 : n3936;
/* FF 11  8  6 */ always @(posedge clk) if (n1131) n1128 <= 1'b0 ? 1'b0 : n3937;
/* FF 29  5  4 */ always @(posedge clk) if (n3605) n3822 <= 1'b0 ? 1'b0 : n3938;
/* FF 23 15  1 */ always @(posedge clk) if (n3216) n3223 <= 1'b0 ? 1'b0 : n3939;
/* FF 24 16  1 */ always @(posedge clk) if (n3376) n3385 <= 1'b0 ? 1'b0 : n3940;
/* FF 27 22  2 */ always @(posedge clk) if (n3703) n3697 <= 1'b0 ? 1'b0 : n3941;
/* FF  3 15  5 */ always @(posedge clk) if (n207) n298 <= 1'b0 ? 1'b0 : n3942;
/* FF 18  3  1 */ assign \rco[84]  = n3943;
/* FF 21 11  0 */ assign n2682 = n3944;
/* FF  7 16  7 */ always @(posedge clk) if (n630) n748 <= 1'b0 ? 1'b0 : n3945;
/* FF  9 21  7 */ always @(posedge clk) if (n818) n921 <= 1'b0 ? 1'b0 : n3946;
/* FF 26 18  3 */ assign n3555 = n3666;
/* FF 12 22  5 */ always @(posedge clk) if (n1357) n551 <= 1'b0 ? 1'b0 : n3947;
/* FF 26 15  4 */ always @(posedge clk) if (n3233) n3544 <= 1'b0 ? 1'b0 : n3948;
/* FF 17  9  0 */ assign \rco[40]  = n3949;
/* FF 19 23  3 */ assign n2592 = n3950;
/* FF 28 20  5 */ assign \rco[167]  = n3951;
/* FF 22 15  5 */ always @(posedge clk) if (n3216) n3050 <= 1'b0 ? 1'b0 : n3952;
/* FF  4 21  6 */ always @(posedge clk) if (n552) n452 <= 1'b0 ? 1'b0 : n3953;
/* FF 13 28  0 */ always @(posedge clk) if (n1394) n1561 <= 1'b0 ? 1'b0 : n3954;
/* FF 27 11  3 */ always @(posedge clk) if (n3460) n3624 <= 1'b0 ? 1'b0 : n3955;
/* FF 20 11  2 */ assign n2076 = n3956;
/* FF  6 10  3 */ always @(posedge clk) if (n589) n594 <= 1'b0 ? 1'b0 : n3957;
/* FF 23 19  7 */ always @(posedge clk) if (n2573) n3257 <= 1'b0 ? 1'b0 : n3958;
/* FF  5 13  6 */ always @(posedge clk) if (n402) n498 <= 1'b0 ? 1'b0 : n3959;
/* FF 19 24  7 */ always @(posedge clk) if (n2775) n2601 <= 1'b0 ? 1'b0 : n3960;
/* FF 11 20  1 */ always @(posedge clk) if (n1339) n1190 <= 1'b0 ? 1'b0 : n3961;
/* FF 29  9  1 */ assign \rco[76]  = n3962;
/* FF 17 27  4 */ always @(posedge clk) if (n1) n2192 <= 1'b0 ? 1'b0 : n3963;
/* FF 28 23  1 */ always @(posedge clk) if (n3704) n3808 <= 1'b0 ? 1'b0 : n3964;
/* FF  5 18  4 */ always @(posedge clk) if (n657) n535 <= 1'b0 ? 1'b0 : n3965;
/* FF 19  5  3 */ always @(posedge clk) if (n2230) n2438 <= 1'b0 ? 1'b0 : n3966;
/* FF 10 20  0 */ always @(posedge clk) if (n922) n1048 <= 1'b0 ? 1'b0 : n3967;
/* FF 15 16  0 */ always @(posedge clk) if (n1500) n1793 <= 1'b0 ? 1'b0 : n3968;
/* FF 21 15  5 */ assign n3969 = n3069;
/* FF 20 25  5 */ always @(posedge clk) if (n2612) n2369 <= 1'b0 ? 1'b0 : n3970;
/* FF  3 21  4 */ assign n126 = n3971;
/* FF  6  9  7 */ assign \rco[2]  = n3972;
/* FF 20 22  4 */ always @(posedge clk) if (n2384) n2780 <= 1'b0 ? 1'b0 : n3973;
/* FF 12 26  6 */ always @(posedge clk) if (n1393) n1391 <= 1'b0 ? 1'b0 : n3974;
/* FF 14  8  1 */ always @(posedge clk) if (n1741) n1594 <= 1'b0 ? 1'b0 : n3975;
/* FF 17 21  5 */ always @(posedge clk) if (n2347) n2149 <= 1'b0 ? 1'b0 : n3976;
/* FF 17 24  6 */ always @(posedge clk) if (n2000) n2172 <= 1'b0 ? 1'b0 : n3977;
/* FF 23 12  0 */ always @(posedge clk) if (n3031) n3200 <= 1'b0 ? 1'b0 : n3978;
/* FF 24 15  0 */ assign n3376 = n3979;
/* FF 10  6  1 */ always @(posedge clk) if (en_in) n972 <= 1'b0 ? 1'b0 : n3980;
/* FF 27 23  1 */ assign n3981 = n3814;
/* FF  3 12  4 */ always @(posedge clk) if (n168) n281 <= 1'b0 ? 1'b0 : n3982;
/* FF 31 24  3 */ assign \rco[129]  = n3983;
/* FF 18  2  6 */ always @(posedge clk) if (n2207) n2205 <= 1'b0 ? 1'b0 : n3984;
/* FF  7 17  0 */ always @(posedge clk) if (n549) n751 <= 1'b0 ? 1'b0 : n3985;
/* FF 21 12  1 */ always @(posedge clk) if (n3029) n2868 <= 1'b0 ? 1'b0 : n3986;
/* FF 26 21  2 */ always @(posedge clk) if (n3421) n3564 <= 1'b0 ? 1'b0 : n3987;
/* FF 14 26  2 */ always @(posedge clk) if (n1271) n1713 <= 1'b0 ? 1'b0 : n3988;
/* FF 12 21  4 */ always @(posedge clk) if (n1205) n1343 <= 1'b0 ? 1'b0 : n3989;
/* FF 17 10  1 */ always @(posedge clk) if (n2282) n2060 <= 1'b0 ? 1'b0 : n3990;
/* FF 20  4  0 */ assign \rco[94]  = n3991;
/* FF 19 20  2 */ always @(posedge clk) if (n2553) n2567 <= 1'b0 ? 1'b0 : n3992;
/* FF  1 12  6 */ always @(posedge clk) if (n39) n52 <= 1'b0 ? 1'b0 : n3993;
/* FF 10  5  5 */ always @(posedge clk) if (en_in) n971 <= 1'b0 ? 1'b0 : n3994;
/* FF 22 14  2 */ always @(posedge clk) if (n3045) n3053 <= 1'b0 ? 1'b0 : n3995;
/* FF 27  8  2 */ assign n3603 = n3996;
/* FF  3 17  1 */ always @(posedge clk) if (n79) n311 <= 1'b0 ? 1'b0 : n3997;
/* FF 14 25  4 */ always @(posedge clk) if (n697) n1705 <= 1'b0 ? 1'b0 : n3998;
/* FF  6 21  2 */ assign n670 = n3999;
/* FF 17  4  0 */ always @(posedge clk) if (n1761) n1896 <= 1'b0 ? 1'b0 : n4000;
/* FF 23 16  6 */ assign \rco[104]  = n4001;
/* FF 11 14  7 */ always @(posedge clk) if (n1154) n1153 <= 1'b0 ? 1'b0 : n4002;
/* FF 20 10  1 */ always @(posedge clk) if (n2697) n2684 <= 1'b0 ? 1'b0 : n4003;
/* FF  5 14  7 */ always @(posedge clk) if (n402) n510 <= 1'b0 ? 1'b0 : n4004;
/* FF 11 21  6 */ always @(posedge clk) if (n819) n1202 <= 1'b0 ? 1'b0 : n4005;
/* FF 29 10  0 */ always @(posedge clk) if (n3464) n3504 <= 1'b0 ? 1'b0 : n4006;
/* FF 28 22  2 */ always @(posedge clk) if (n3704) n3801 <= 1'b0 ? 1'b0 : n4007;
/* FF 16 12  1 */ assign \rco[42]  = n4008;
/* FF  5 19  3 */ always @(posedge clk) if (n349) n542 <= 1'b0 ? 1'b0 : n4009;
/* FF 19  2  2 */ always @(posedge clk) if (n2207) n2425 <= 1'b0 ? 1'b0 : n4010;
/* FF 16 17  6 */ always @(posedge clk) if (n2110) n1969 <= 1'b0 ? 1'b0 : n4011;
/* FF 10 23  1 */ always @(posedge clk) if (n821) n148 <= 1'b0 ? 1'b0 : n4012;
/* FF 27  6  1 */ assign n3459 = n4013;
/* FF 13 15  0 */ always @(posedge clk) if (n739) n1470 <= 1'b0 ? 1'b0 : n4014;
/* FF 30 12  0 */ always @(posedge clk) if (n3892) n3894 <= 1'b0 ? 1'b0 : n4015;
/* FF 15 17  7 */ always @(posedge clk) if (n1500) n1807 <= 1'b0 ? 1'b0 : n4016;
/* FF 18  6  3 */ always @(posedge clk) if (n2241) n2234 <= 1'b0 ? 1'b0 : n4017;
/* FF  7 21  5 */ always @(posedge clk) if (n360) n773 <= 1'b0 ? 1'b0 : n4018;
/* FF  6  7  5 */ always @(posedge clk) if (n570) n576 <= 1'b0 ? 1'b0 : n4019;
/* FF 20 24  2 */ always @(posedge clk) if (n2775) n2790 <= 1'b0 ? 1'b0 : n4020;
/* FF  3 18  5 */ always @(posedge clk) if (n215) n323 <= 1'b0 ? 1'b0 : n4021;
/* FF  6  8  4 */ always @(posedge clk) if (n570) n584 <= 1'b0 ? 1'b0 : n4022;
/* FF 20 21  5 */ always @(posedge clk) if (n2553) n2773 <= 1'b0 ? 1'b0 : n4023;
/* FF 14 11  0 */ always @(posedge clk) if (n1622) n1612 <= 1'b0 ? 1'b0 : n4024;
/* FF 17 22  4 */ always @(posedge clk) if (n1999) n2156 <= 1'b0 ? 1'b0 : n4025;
/* FF  1 19  1 */ always @(posedge clk) if (n119) n105 <= 1'b0 ? 1'b0 : n4026;
/* FF 17 25  5 */ always @(posedge clk) if (n2017) n2181 <= 1'b0 ? 1'b0 : n4027;
/* FF 10 25  0 */ always @(posedge clk) if (n567) n1080 <= 1'b0 ? 1'b0 : n4028;
/* FF 24 14  3 */ always @(posedge clk) if (n3376) n3372 <= 1'b0 ? 1'b0 : n4029;
/* FF 27 20  0 */ always @(posedge clk) if (n3424) n3675 <= 1'b0 ? 1'b0 : n4030;
/* FF  4 19  7 */ assign n215 = n4031;
/* FF  3 13  3 */ assign \rco[13]  = n406;
/* FF 22 10  7 */ always @(posedge clk) if (n2856) n3021 <= 1'b0 ? 1'b0 : n4032;
/* FF 18  5  7 */ always @(posedge clk) if (n2230) n2228 <= 1'b0 ? 1'b0 : n4033;
/* FF  7 22  1 */ always @(posedge clk) if (n695) n784 <= 1'b0 ? 1'b0 : n4034;
/* FF  9 23  1 */ always @(posedge clk) if (n819) n926 <= 1'b0 ? 1'b0 : n4035;
/* FF 21 13  2 */ always @(posedge clk) if (n2519) n2876 <= 1'b0 ? 1'b0 : n4036;
/* FF 26 20  1 */ assign \rco[168]  = n4037;
/* FF 12 15  2 */ always @(posedge clk) if (n1155) n1298 <= 1'b0 ? 1'b0 : n4038;
/* FF 14 21  3 */ assign n1672 = n4039;
/* FF 19 30  4 */ always @(posedge clk) if (n2592) n2638 <= 1'b0 ? 1'b0 : n4040;
/* FF 19 21  5 */ always @(posedge clk) if (n2164) n2581 <= 1'b0 ? 1'b0 : n4041;
/* FF 11 17  3 */ always @(posedge clk) if (n900) n1171 <= 1'b0 ? 1'b0 : n4042;
/* FF 10 11  7 */ always @(posedge clk) if (n996) n995 <= 1'b0 ? 1'b0 : n4043;
/* FF 16  8  6 */ always @(posedge clk) if (n1625) n1921 <= 1'b0 ? 1'b0 : n4044;
/* FF  1 13  5 */ always @(posedge clk) if (n83) n64 <= 1'b0 ? 1'b0 : n4045;
/* FF 24 17  7 */ always @(posedge clk) if (n2123) n3401 <= 1'b0 ? 1'b0 : n4046;
/* FF 28  7  4 */ always @(posedge clk) if (n3488) n3723 <= 1'b0 ? 1'b0 : n4047;
/* FF 22  9  3 */ always @(posedge clk) if (n2989) n3017 <= 1'b0 ? 1'b0 : n4048;
/* FF 15 21  4 */ always @(posedge clk) if (n1356) n1840 <= 1'b0 ? 1'b0 : n4049;
/* FF 20 28  7 */ always @(posedge clk) if (n2195) n2828 <= 1'b0 ? 1'b0 : n4050;
/* FF 17  5  3 */ assign \rco[150]  = n4051;
/* FF 20  9  0 */ assign n2678 = n4052;
/* FF  6 20  1 */ always @(posedge clk) if (n552) n661 <= 1'b0 ? 1'b0 : n4053;
/* FF 23 17  1 */ always @(posedge clk) if (n2540) n2533 <= 1'b0 ? 1'b0 : n4054;
/* FF 11 15  4 */ always @(posedge clk) if (n733) n811 <= 1'b0 ? 1'b0 : n4055;
/* FF 26  6  5 */ always @(posedge clk) if (n3459) n3478 <= 1'b0 ? 1'b0 : n4056;
/* FF 11 18  7 */ always @(posedge clk) if (n1187) n1186 <= 1'b0 ? 1'b0 : n4057;
/* FF 29 11  7 */ always @(posedge clk) if (n3751) n3846 <= 1'b0 ? 1'b0 : n4058;
/* FF 28 21  3 */ always @(posedge clk) if (n3788) n3794 <= 1'b0 ? 1'b0 : n4059;
/* FF 16 11  0 */ always @(posedge clk) if (n2076) n1935 <= 1'b0 ? 1'b0 : n4060;
/* FF 19  3  1 */ always @(posedge clk) if (n1887) n2428 <= 1'b0 ? 1'b0 : n4061;
/* FF  4 12  0 */ always @(posedge clk) if (n77) n393 <= 1'b0 ? 1'b0 : n4062;
/* FF 13 16  1 */ always @(posedge clk) if (n922) n1478 <= 1'b0 ? 1'b0 : n4063;
/* FF 27  7  2 */ always @(posedge clk) if (n3459) n3597 <= 1'b0 ? 1'b0 : n4064;
/* FF 15 22  6 */ always @(posedge clk) if (n1835) n1851 <= 1'b0 ? 1'b0 : n4065;
/* FF 18  9  2 */ always @(posedge clk) if (n2055) n2263 <= 1'b0 ? 1'b0 : n4066;
/* FF  7 26  4 */ always @(posedge clk) if (n567) n802 <= 1'b0 ? 1'b0 : n4067;
/* FF  9 19  6 */ always @(posedge clk) if (n454) n907 <= 1'b0 ? 1'b0 : n4068;
/* FF  3 19  6 */ always @(posedge clk) if (n115) n333 <= 1'b0 ? 1'b0 : n4069;
/* FF  6 11  5 */ always @(posedge clk) if (n286) n291 <= 1'b0 ? 1'b0 : n4070;
/* FF 12 24  0 */ always @(posedge clk) if (n961) n1367 <= 1'b0 ? 1'b0 : n4071;
/* FF 17 23  3 */ always @(posedge clk) if (n1069) n2162 <= 1'b0 ? 1'b0 : n4072;
/* FF 19 17  2 */ always @(posedge clk) if (n2727) n2543 <= 1'b0 ? 1'b0 : n4073;
/* FF 17 26  4 */ always @(posedge clk) if (n1557) n2186 <= 1'b0 ? 1'b0 : n4074;
/* FF 22 21  5 */ always @(posedge clk) if (n2564) n3101 <= 1'b0 ? 1'b0 : n4075;
/* FF 24 24  5 */ always @(posedge clk) if (n3112) n2173 <= 1'b0 ? 1'b0 : n4076;
/* FF 10 24  3 */ always @(posedge clk) if (n820) n1075 <= 1'b0 ? 1'b0 : n4077;
/* FF 28 11  3 */ assign n3751 = n4078;
/* FF 24 13  2 */ always @(posedge clk) if (n3351) n3363 <= 1'b0 ? 1'b0 : n4079;
/* FF 27 21  7 */ always @(posedge clk) if (n3421) n3694 <= 1'b0 ? 1'b0 : n4080;
/* FF  4 18  4 */ always @(posedge clk) if (n349) n434 <= 1'b0 ? 1'b0 : n4081;
/* FF  3 10  2 */ always @(posedge clk) if (n251) n264 <= 1'b0 ? 1'b0 : n4082;
/* FF 18  4  4 */ always @(posedge clk) if (n2207) n2217 <= 1'b0 ? 1'b0 : n4083;
/* FF  7 23  2 */ always @(posedge clk) if (n454) n792 <= 1'b0 ? 1'b0 : n4084;
/* FF  9 16  0 */ always @(posedge clk) if (n645) n875 <= 1'b0 ? 1'b0 : n4085;
/* FF 12 14  1 */ always @(posedge clk) if (n1154) n1289 <= 1'b0 ? 1'b0 : n4086;
/* FF 26 23  0 */ always @(posedge clk) if (n3703) n3576 <= 1'b0 ? 1'b0 : n4087;
/* FF 14 20  0 */ always @(posedge clk) if (n1347) n1676 <= 1'b0 ? 1'b0 : n4088;
/* FF  5  8  4 */ always @(posedge clk) if (n21) n471 <= 1'b0 ? 1'b0 : n4089;
/* FF 19 31  7 */ always @(posedge clk) if (n2592) n2648 <= 1'b0 ? 1'b0 : n4090;
/* FF 23 21  6 */ always @(posedge clk) if (n3258) n3277 <= 1'b0 ? 1'b0 : n4091;
/* FF 19 18  4 */ always @(posedge clk) if (n2348) n2558 <= 1'b0 ? 1'b0 : n4092;
/* FF 10 10  0 */ assign n983 = n4093;
/* FF 16 23  7 */ always @(posedge clk) if (n2000) n1997 <= 1'b0 ? 1'b0 : n4094;
/* FF  1 14  4 */ always @(posedge clk) if (n85) n72 <= 1'b0 ? 1'b0 : n4095;
/* FF 28  6  7 */ always @(posedge clk) if (n3594) n3717 <= 1'b0 ? 1'b0 : n4096;
/* FF 22  8  0 */ always @(posedge clk) if (n2989) n3010 <= 1'b0 ? 1'b0 : n4097;
/* FF 15 10  5 */ always @(posedge clk) if (n1624) n1759 <= 1'b0 ? 1'b0 : n4098;
/* FF  2 16  4 */ always @(posedge clk) if (n197) n205 <= 1'b0 ? 1'b0 : n4099;
/* FF 20 19  6 */ always @(posedge clk) if (n2562) n2755 <= 1'b0 ? 1'b0 : n4100;
/* FF 18 22  0 */ assign n1871 = n4101;
/* FF 17  6  2 */ always @(posedge clk) if (n2045) n2040 <= 1'b0 ? 1'b0 : n4102;
/* FF  6 23  0 */ always @(posedge clk) if (n360) n687 <= 1'b0 ? 1'b0 : n4103;
/* FF 20  8  7 */ always @(posedge clk) if (n2247) n2675 <= 1'b0 ? 1'b0 : n4104;
/* FF 12 28  5 */ always @(posedge clk) if (n1394) n1399 <= 1'b0 ? 1'b0 : n4105;
/* FF 23 22  0 */ always @(posedge clk) if (n3422) n3279 <= 1'b0 ? 1'b0 : n4106;
/* FF 11 19  4 */ always @(posedge clk) if (n900) n465 <= 1'b0 ? 1'b0 : n4107;
/* FF 29 12  6 */ always @(posedge clk) if (n3751) n3854 <= 1'b0 ? 1'b0 : n4108;
/* FF 16 10  3 */ always @(posedge clk) if (n1771) n1929 <= 1'b0 ? 1'b0 : n4109;
/* FF  5 21  1 */ assign n4110 = n676;
/* FF 22 26  1 */ always @(posedge clk) if (n2613) n3134 <= 1'b0 ? 1'b0 : n4111;
/* FF 15 24  4 */ always @(posedge clk) if (n778) n686 <= 1'b0 ? 1'b0 : n4112;
/* FF 13 17  2 */ always @(posedge clk) if (n1461) n1486 <= 1'b0 ? 1'b0 : n4113;
/* FF 27  4  3 */ assign \rco[81]  = n4114;
/* FF 15 23  5 */ always @(posedge clk) if (n778) n1857 <= 1'b0 ? 1'b0 : n4115;
/* FF 18  8  1 */ always @(posedge clk) if (n2055) n2250 <= 1'b0 ? 1'b0 : n4116;
/* FF  3 16  7 */ always @(posedge clk) if (n197) n309 <= 1'b0 ? 1'b0 : n4117;
/* FF 17 16  2 */ assign n2110 = n4118;
/* FF 19 14  3 */ always @(posedge clk) if (n2123) n2514 <= 1'b0 ? 1'b0 : n4119;
/* FF 22 20  6 */ always @(posedge clk) if (n3087) n3094 <= 1'b0 ? 1'b0 : n4120;
/* FF 10 14  5 */ always @(posedge clk) if (n750) n1012 <= 1'b0 ? 1'b0 : n4121;
/* FF 24 23  4 */ always @(posedge clk) if (n3104) n3437 <= 1'b0 ? 1'b0 : n4122;
/* FF 22 25  5 */ always @(posedge clk) if (n2812) n2603 <= 1'b0 ? 1'b0 : n4123;
/* FF 10 27  2 */ always @(posedge clk) if (n804) n1095 <= 1'b0 ? 1'b0 : n4124;
/* FF 24 12  5 */ always @(posedge clk) if (n3351) n3358 <= 1'b0 ? 1'b0 : n4125;
/* FF 16 24  3 */ assign n4126 = n2175;
/* FF 28 10  0 */ always @(posedge clk) if (n3462) n3741 <= 1'b0 ? 1'b0 : n4127;
/* FF 27 18  6 */ always @(posedge clk) if (n3553) n3663 <= 1'b0 ? 1'b0 : n4128;
/* FF  4 17  5 */ always @(posedge clk) if (n2) n429 <= 1'b0 ? 1'b0 : n4129;
/* FF  3 11  1 */ always @(posedge clk) if (n153) n271 <= 1'b0 ? 1'b0 : n4130;
/* FF 18  7  5 */ always @(posedge clk) if (n1761) n2244 <= 1'b0 ? 1'b0 : n4131;
/* FF  9 17  3 */ always @(posedge clk) if (n1030) n886 <= 1'b0 ? 1'b0 : n4132;
/* FF 15  5  1 */ always @(posedge clk) if (n1742) n1726 <= 1'b0 ? 1'b0 : n4133;
/* FF 14 23  1 */ assign n4134 = n1860;
/* FF 20 12  4 */ always @(posedge clk) if (n2682) n2702 <= 1'b0 ? 1'b0 : n4135;
/* FF 19 19  7 */ assign n2164 = n4136;
/* FF 10 13  1 */ assign n629 = n4137;
/* FF 16 22  4 */ always @(posedge clk) if (n1835) n1990 <= 1'b0 ? 1'b0 : n4138;
/* FF  1 15  3 */ assign n85 = n4139;
/* FF 16 27  7 */ always @(posedge clk) if (n1) n2019 <= 1'b0 ? 1'b0 : n4140;
/* FF 22 11  1 */ assign \rco[56]  = n4141;
/* FF 30 10  3 */ always @(posedge clk) if (n3892) n3888 <= 1'b0 ? 1'b0 : n4142;
/* FF 15 11  6 */ always @(posedge clk) if (n1624) n1769 <= 1'b0 ? 1'b0 : n4143;
/* FF  2 19  5 */ assign n119 = n4144;
/* FF  6 13  6 */ always @(posedge clk) if (n78) n621 <= 1'b0 ? 1'b0 : n4145;
/* FF 15  6  5 */ always @(posedge clk) if (n1744) n1738 <= 1'b0 ? 1'b0 : n4146;
/* FF 17  7  5 */ always @(posedge clk) if (n2045) n2051 <= 1'b0 ? 1'b0 : n4147;
/* FF 18 25  1 */ always @(posedge clk) if (n1878) n2378 <= 1'b0 ? 1'b0 : n4148;
/* FF  6 22  7 */ always @(posedge clk) if (n673) n685 <= 1'b0 ? 1'b0 : n4149;
/* FF 20 18  5 */ always @(posedge clk) if (n2348) n2563 <= 1'b0 ? 1'b0 : n4150;
/* FF 20 15  6 */ always @(posedge clk) if (n2715) n2723 <= 1'b0 ? 1'b0 : n4151;
/* FF 11 13  2 */ always @(posedge clk) if (n733) n1140 <= 1'b0 ? 1'b0 : n4152;
/* FF 23 23  3 */ always @(posedge clk) if (n3104) n3290 <= 1'b0 ? 1'b0 : n4153;
/* FF 11 16  5 */ always @(posedge clk) if (n891) n1164 <= 1'b0 ? 1'b0 : n4154;
/* FF  5 22  0 */ always @(posedge clk) if (n673) n555 <= 1'b0 ? 1'b0 : n4155;
/* FF  9 13  1 */ always @(posedge clk) if (n629) n856 <= 1'b0 ? 1'b0 : n4156;
/* FF 13  7  4 */ always @(posedge clk) if (n977) n1427 <= 1'b0 ? 1'b0 : n4157;
/* FF 15 25  3 */ assign \rco[187]  = n4158;
/* FF 13 18  3 */ always @(posedge clk) if (n1205) n1495 <= 1'b0 ? 1'b0 : n4159;
/* FF 27  5  4 */ always @(posedge clk) if (n3594) n3589 <= 1'b0 ? 1'b0 : n4160;
/* FF 18 11  0 */ assign n2283 = n4161;
/* FF 15 20  4 */ always @(posedge clk) if (n1347) n1831 <= 1'b0 ? 1'b0 : n4162;
/* FF 26  7  3 */ always @(posedge clk) if (n3603) n3484 <= 1'b0 ? 1'b0 : n4163;
/* FF 17 17  1 */ always @(posedge clk) if (n2111) n2115 <= 1'b0 ? 1'b0 : n4164;
/* FF  2 14  0 */ always @(posedge clk) if (n83) n187 <= 1'b0 ? 1'b0 : n4165;
/* FF 16  7  1 */ always @(posedge clk) if (n1743) n1908 <= 1'b0 ? 1'b0 : n4166;
/* FF 19 15  0 */ always @(posedge clk) if (n2715) n2525 <= 1'b0 ? 1'b0 : n4167;
/* FF 23  5  3 */ always @(posedge clk) if (n3158) n3153 <= 1'b0 ? 1'b0 : n4168;
/* FF 22 23  7 */ always @(posedge clk) if (n3104) n3115 <= 1'b0 ? 1'b0 : n4169;
/* FF 24 22  7 */ always @(posedge clk) if (n3422) n3431 <= 1'b0 ? 1'b0 : n4170;
/* FF 22 24  6 */ always @(posedge clk) if (n3113) n3122 <= 1'b0 ? 1'b0 : n4171;
/* FF 24 11  4 */ assign n2725 = n3466;
/* FF 10 26  5 */ assign n1090 = n1246;
/* FF 27 19  5 */ always @(posedge clk) if (n3553) n3672 <= 1'b0 ? 1'b0 : n4172;
/* FF 28  9  1 */ always @(posedge clk) if (n3621) n3735 <= 1'b0 ? 1'b0 : n4173;
/* FF  4 16  2 */ always @(posedge clk) if (n79) n422 <= 1'b0 ? 1'b0 : n4174;
/* FF  9 18  2 */ always @(posedge clk) if (n1030) n894 <= 1'b0 ? 1'b0 : n4175;
/* FF 14 22  6 */ always @(posedge clk) if (n1402) n1693 <= 1'b0 ? 1'b0 : n4176;
/* FF 17  3  2 */ always @(posedge clk) if (n1887) n2027 <= 1'b0 ? 1'b0 : n4177;
/* FF  6 18  4 */ always @(posedge clk) if (n657) n653 <= 1'b0 ? 1'b0 : n4178;
/* FF  5 10  6 */ always @(posedge clk) if (n184) n480 <= 1'b0 ? 1'b0 : n4179;
/* FF 19 29  1 */ always @(posedge clk) if (n2614) n1816 <= 1'b0 ? 1'b0 : n4180;
/* FF 23 27  4 */ always @(posedge clk) if (n2017) n2822 <= 1'b0 ? 1'b0 : n4181;
/* FF 19 16  6 */ assign n2538 = n4182;
/* FF 11 28  0 */ always @(posedge clk) if (n1384) n1255 <= 1'b0 ? 1'b0 : n4183;
/* FF 10 12  2 */ always @(posedge clk) if (n996) n999 <= 1'b0 ? 1'b0 : n4184;
/* FF 24 25  3 */ always @(posedge clk) if (n2812) n3449 <= 1'b0 ? 1'b0 : n4185;
/* FF 16 21  5 */ always @(posedge clk) if (n1835) n1986 <= 1'b0 ? 1'b0 : n4186;
/* FF  1  8  2 */ always @(posedge clk) if (n37) n16 <= 1'b0 ? 1'b0 : n4187;
/* FF 16 26  4 */ always @(posedge clk) if (n1557) n2014 <= 1'b0 ? 1'b0 : n4188;
/* FF  9 28  1 */ always @(posedge clk) if (n961) n957 <= 1'b0 ? 1'b0 : n4189;
/* FF  3 22  4 */ always @(posedge clk) if (n352) n357 <= 1'b0 ? 1'b0 : n4190;
/* FF  2 18  2 */ always @(posedge clk) if (n115) n211 <= 1'b0 ? 1'b0 : n4191;
/* FF  6 12  5 */ always @(posedge clk) if (n286) n611 <= 1'b0 ? 1'b0 : n4192;
/* FF 15  7  6 */ assign n1744 = n4193;
/* FF 21  7  6 */ assign n2470 = n3009;
/* FF 18 24  2 */ always @(posedge clk) if (n1878) n2372 <= 1'b0 ? 1'b0 : n4194;
/* FF 20 17  4 */ always @(posedge clk) if (n2727) n2736 <= 1'b0 ? 1'b0 : n4195;
/* FF 23 20  2 */ always @(posedge clk) if (n3258) n3265 <= 1'b0 ? 1'b0 : n4196;
/* FF 11 10  3 */ assign \rco[1]  = n4197;
/* FF 24  7  3 */ assign n3158 = n4198;
/* FF  9 14  0 */ always @(posedge clk) if (n629) n859 <= 1'b0 ? 1'b0 : n4199;
/* FF  4 20  7 */ always @(posedge clk) if (n215) n445 <= 1'b0 ? 1'b0 : n4200;
/* FF 13 19  4 */ assign n4201 = n1674;
/* FF 18 10  7 */ always @(posedge clk) if (n2282) n2280 <= 1'b0 ? 1'b0 : n4202;
/* FF 14 18  3 */ always @(posedge clk) if (n1672) n1664 <= 1'b0 ? 1'b0 : n4203;
/* FF 19 25  6 */ always @(posedge clk) if (n2612) n2610 <= 1'b0 ? 1'b0 : n4204;
/* FF 17 18  0 */ always @(posedge clk) if (n1825) n2125 <= 1'b0 ? 1'b0 : n4205;
/* FF 16  6  2 */ always @(posedge clk) if (n1744) n1899 <= 1'b0 ? 1'b0 : n4206;
/* FF 19 12  1 */ always @(posedge clk) if (n1936) n2498 <= 1'b0 ? 1'b0 : n4207;
/* FF 23 10  2 */ always @(posedge clk) if (n2697) n3185 <= 1'b0 ? 1'b0 : n4208;
/* FF 22 22  0 */ always @(posedge clk) if (n2961) n3105 <= 1'b0 ? 1'b0 : n4209;
/* FF 22 27  7 */ always @(posedge clk) if (n2970) n3132 <= 1'b0 ? 1'b0 : n4210;
/* FF 24 10  7 */ always @(posedge clk) if (n3352) n3347 <= 1'b0 ? 1'b0 : n4211;
/* FF 28  8  6 */ always @(posedge clk) if (n3605) n3731 <= 1'b0 ? 1'b0 : n4212;
/* FF 13  5  5 */ always @(posedge clk) if (n1577) n1413 <= 1'b0 ? 1'b0 : n4213;
/* FF  2 22  7 */ always @(posedge clk) if (n352) n242 <= 1'b0 ? 1'b0 : n4214;
/* FF 17 12  3 */ always @(posedge clk) if (n2056) n2080 <= 1'b0 ? 1'b0 : n4215;
/* FF 19 26  0 */ assign n1878 = n4216;
/* FF  5 11  1 */ always @(posedge clk) if (n184) n482 <= 1'b0 ? 1'b0 : n4217;
/* FF 11 22  6 */ always @(posedge clk) if (n695) n1212 <= 1'b0 ? 1'b0 : n4218;
/* FF 23 24  5 */ always @(posedge clk) if (n3112) n3301 <= 1'b0 ? 1'b0 : n4219;
/* FF 23  7  4 */ always @(posedge clk) if (n3006) n3170 <= 1'b0 ? 1'b0 : n4220;
/* FF 11 29  7 */ always @(posedge clk) if (n1384) n1269 <= 1'b0 ? 1'b0 : n4221;
/* FF 10 15  3 */ always @(posedge clk) if (n750) n1018 <= 1'b0 ? 1'b0 : n4222;
/* FF 16 20  2 */ always @(posedge clk) if (n1843) n1976 <= 1'b0 ? 1'b0 : n4223;
/* FF  1  9  1 */ always @(posedge clk) if (n153) n24 <= 1'b0 ? 1'b0 : n4224;
/* FF 16 25  5 */ always @(posedge clk) if (n1557) n2008 <= 1'b0 ? 1'b0 : n4225;
/* FF 21 24  2 */ always @(posedge clk) if (n3113) n2955 <= 1'b0 ? 1'b0 : n4226;
/* FF 13 23  1 */ always @(posedge clk) if (n1069) n1525 <= 1'b0 ? 1'b0 : n4227;
/* FF 27 14  0 */ always @(posedge clk) if (n3527) n3641 <= 1'b0 ? 1'b0 : n4228;
/* FF 18 14  4 */ assign n1666 = n4229;
/* FF  2 21  3 */ always @(posedge clk) if (n126) n230 <= 1'b0 ? 1'b0 : n4230;
/* FF  6 15  4 */ always @(posedge clk) if (n630) n634 <= 1'b0 ? 1'b0 : n4231;
/* FF 18 27  3 */ always @(posedge clk) if (n2020) n2396 <= 1'b0 ? 1'b0 : n4232;
/* FF 20 16  3 */ assign n2728 = n2897;
/* FF  6 16  5 */ always @(posedge clk) if (n511) n301 <= 1'b0 ? 1'b0 : n4233;
/* FF 20 13  4 */ always @(posedge clk) if (n2283) n2510 <= 1'b0 ? 1'b0 : n4234;
/* FF  4 11  5 */ always @(posedge clk) if (n184) n390 <= 1'b0 ? 1'b0 : n4235;
/* FF 22 18  5 */ always @(posedge clk) if (n3065) n2552 <= 1'b0 ? 1'b0 : n4236;
/* FF 22  7  2 */ always @(posedge clk) if (n2841) n3000 <= 1'b0 ? 1'b0 : n4237;
/* FF 10 17  3 */ assign n1030 = n4238;
/* FF  9 15  7 */ always @(posedge clk) if (n645) n874 <= 1'b0 ? 1'b0 : n4239;
/* FF 24  6  0 */ always @(posedge clk) if (n3006) n3321 <= 1'b0 ? 1'b0 : n4240;
/* FF 28 12  3 */ always @(posedge clk) if (n3462) n3756 <= 1'b0 ? 1'b0 : n4241;
/* FF 13 20  5 */ always @(posedge clk) if (n1339) n1508 <= 1'b0 ? 1'b0 : n4242;
/* FF 18 13  6 */ always @(posedge clk) if (n2283) n2301 <= 1'b0 ? 1'b0 : n4243;
/* FF 16  5  3 */ always @(posedge clk) if (n1742) n1891 <= 1'b0 ? 1'b0 : n4244;
/* FF 23 11  1 */ always @(posedge clk) if (n3031) n3191 <= 1'b0 ? 1'b0 : n4245;
/* FF 11 25  4 */ always @(posedge clk) if (n954) n1235 <= 1'b0 ? 1'b0 : n4246;
/* FF 22 17  1 */ always @(posedge clk) if (n3065) n3073 <= 1'b0 ? 1'b0 : n4247;
/* FF 24 20  1 */ always @(posedge clk) if (n3411) n3410 <= 1'b0 ? 1'b0 : n4248;
/* FF 16 16  7 */ always @(posedge clk) if (n2110) n1962 <= 1'b0 ? 1'b0 : n4249;
/* FF 10 28  7 */ always @(posedge clk) if (n821) n1108 <= 1'b0 ? 1'b0 : n4250;
/* FF 24  9  6 */ always @(posedge clk) if (n3352) n3338 <= 1'b0 ? 1'b0 : n4251;
/* FF 13  6  4 */ always @(posedge clk) if (n977) n1419 <= 1'b0 ? 1'b0 : n4252;
/* FF  4 22  0 */ assign \rco[137]  = n4253;
/* FF 21 23  0 */ always @(posedge clk) if (n2961) n2943 <= 1'b0 ? 1'b0 : n4254;
/* FF 15 13  5 */ always @(posedge clk) if (n1015) n813 <= 1'b0 ? 1'b0 : n4255;
/* FF 29 19  5 */ always @(posedge clk) if (n3786) n3420 <= 1'b0 ? 1'b0 : n4256;
/* FF 14 16  4 */ always @(posedge clk) if (n1792) n1650 <= 1'b0 ? 1'b0 : n4257;
/* FF 17 13  0 */ always @(posedge clk) if (n2056) n2086 <= 1'b0 ? 1'b0 : n4258;
/* FF  5 12  0 */ always @(posedge clk) if (n77) n484 <= 1'b0 ? 1'b0 : n4259;
/* FF 23 25  2 */ assign \rco[188]  = n4260;
/* FF 11 23  5 */ always @(posedge clk) if (n796) n1113 <= 1'b0 ? 1'b0 : n4261;
/* FF 19 27  3 */ always @(posedge clk) if (n2614) n2619 <= 1'b0 ? 1'b0 : n4262;
/* FF 11 26  6 */ always @(posedge clk) if (n954) n1241 <= 1'b0 ? 1'b0 : n4263;
/* FF  1 10  0 */ always @(posedge clk) if (n37) n28 <= 1'b0 ? 1'b0 : n4264;
/* FF 21 25  1 */ always @(posedge clk) if (n2970) n2963 <= 1'b0 ? 1'b0 : n4265;
/* FF  9 11  4 */ always @(posedge clk) if (n988) n846 <= 1'b0 ? 1'b0 : n4266;
/* FF 13 24  0 */ assign n1532 = n4267;
/* FF 15 14  1 */ always @(posedge clk) if (n1791) n1784 <= 1'b0 ? 1'b0 : n4268;
/* FF  3 20  6 */ always @(posedge clk) if (n119) n347 <= 1'b0 ? 1'b0 : n4269;
/* FF  2 20  0 */ always @(posedge clk) if (n126) n217 <= 1'b0 ? 1'b0 : n4270;
/* FF  6 14  3 */ always @(posedge clk) if (n78) n626 <= 1'b0 ? 1'b0 : n4271;
/* FF 20 23  2 */ assign n1876 = n4272;
/* FF 18 17  5 */ always @(posedge clk) if (n1825) n2330 <= 1'b0 ? 1'b0 : n4273;
/* FF 18 26  4 */ always @(posedge clk) if (n2615) n2389 <= 1'b0 ? 1'b0 : n4274;
/* FF  6 19  4 */ assign n658 = n767;
/* FF 11  8  1 */ always @(posedge clk) if (n1131) n1124 <= 1'b0 ? 1'b0 : n4275;
/* FF 29  5  1 */ always @(posedge clk) if (n3605) n3819 <= 1'b0 ? 1'b0 : n4276;
/* FF 28 19  1 */ always @(posedge clk) if (n3424) n3778 <= 1'b0 ? 1'b0 : n4277;
/* FF 19  9  3 */ always @(posedge clk) if (n2451) n2474 <= 1'b0 ? 1'b0 : n4278;
/* FF  4 10  6 */ always @(posedge clk) if (n251) n385 <= 1'b0 ? 1'b0 : n4279;
/* FF 22 29  4 */ assign \rco[177]  = n4280;
/* FF 24 16  6 */ always @(posedge clk) if (n3376) n3390 <= 1'b0 ? 1'b0 : n4281;
/* FF 22  6  5 */ always @(posedge clk) if (n2841) n2995 <= 1'b0 ? 1'b0 : n4282;
/* FF 10 16  0 */ always @(posedge clk) if (n891) n1023 <= 1'b0 ? 1'b0 : n4283;
/* FF 24  5  1 */ always @(posedge clk) if (n3158) n3319 <= 1'b0 ? 1'b0 : n4284;
/* FF 13 10  7 */ always @(posedge clk) if (n850) n1440 <= 1'b0 ? 1'b0 : n4285;
/* FF 31 27  7 */ assign \rco[140]  = n4286;
/* FF 18  3  4 */ assign n1887 = n4287;
/* FF 13 21  6 */ always @(posedge clk) if (n1356) n1518 <= 1'b0 ? 1'b0 : n4288;
/* FF 18 12  5 */ always @(posedge clk) if (n1936) n2291 <= 1'b0 ? 1'b0 : n4289;
/* FF 21  6  2 */ always @(posedge clk) if (n2247) n2835 <= 1'b0 ? 1'b0 : n4290;
/* FF 29 23  2 */ always @(posedge clk) if (n3788) n3883 <= 1'b0 ? 1'b0 : n4291;
/* FF 14 12  1 */ assign n1620 = n1774;
/* FF 19 23  4 */ assign n2593 = n4292;
/* FF 19 10  7 */ always @(posedge clk) if (n2678) n2485 <= 1'b0 ? 1'b0 : n4293;
/* FF 24 19  0 */ always @(posedge clk) if (n2123) n2716 <= 1'b0 ? 1'b0 : n4294;
/* FF 28 14  4 */ always @(posedge clk) if (n2085) n3035 <= 1'b0 ? 1'b0 : n4295;
/* FF  4 21  1 */ always @(posedge clk) if (n552) n448 <= 1'b0 ? 1'b0 : n4296;
/* FF  7 13  0 */ assign \rco[155]  = n4297;
/* FF 21  8  1 */ always @(posedge clk) if (n2989) n2281 <= 1'b0 ? 1'b0 : n4298;
/* FF 26 17  2 */ always @(posedge clk) if (n3249) n3548 <= 1'b0 ? 1'b0 : n4299;
/* FF 18 30  1 */ always @(posedge clk) if (n1881) n2418 <= 1'b0 ? 1'b0 : n4300;
/* FF 14 19  5 */ always @(posedge clk) if (n1672) n1669 <= 1'b0 ? 1'b0 : n4301;
/* FF 17 14  1 */ always @(posedge clk) if (n1625) n2095 <= 1'b0 ? 1'b0 : n4302;
/* FF 29 20  4 */ always @(posedge clk) if (n3786) n3872 <= 1'b0 ? 1'b0 : n4303;
/* FF  5 13  3 */ always @(posedge clk) if (n402) n495 <= 1'b0 ? 1'b0 : n4304;
/* FF 19 24  2 */ always @(posedge clk) if (n2775) n2596 <= 1'b0 ? 1'b0 : n4305;
/* FF 11 20  4 */ always @(posedge clk) if (n1339) n1193 <= 1'b0 ? 1'b0 : n4306;
/* FF 11 27  5 */ always @(posedge clk) if (n1393) n1252 <= 1'b0 ? 1'b0 : n4307;
/* FF 16 18  0 */ always @(posedge clk) if (n1205) n1971 <= 1'b0 ? 1'b0 : n4308;
/* FF 21 26  0 */ assign \rco[175]  = n4309;
/* FF 13 25  3 */ always @(posedge clk) if (n697) n1537 <= 1'b0 ? 1'b0 : n4310;
/* FF 27 12  2 */ always @(posedge clk) if (n3368) n3631 <= 1'b0 ? 1'b0 : n4311;
/* FF 15 15  2 */ assign n4312 = n1952;
/* FF  3 21  1 */ assign n351 = n4313;
/* FF 18 16  6 */ always @(posedge clk) if (n2540) n2320 <= 1'b0 ? 1'b0 : n4314;
/* FF  6  9  2 */ assign \rco[21]  = n727;
/* FF 18 29  5 */ always @(posedge clk) if (n1881) n2413 <= 1'b0 ? 1'b0 : n4315;
/* FF 20 22  1 */ always @(posedge clk) if (n2384) n2777 <= 1'b0 ? 1'b0 : n4316;
/* FF 28 18  2 */ always @(posedge clk) if (n3765) n3775 <= 1'b0 ? 1'b0 : n4317;
/* FF 19  6  2 */ always @(posedge clk) if (n2241) n2445 <= 1'b0 ? 1'b0 : n4318;
/* FF  4  9  7 */ always @(posedge clk) if (n260) n378 <= 1'b0 ? 1'b0 : n4319;
/* FF 24 15  7 */ always @(posedge clk) if (n3233) n3382 <= 1'b0 ? 1'b0 : n4320;
/* FF 10 19  1 */ assign n549 = n4321;
/* FF  9  9  5 */ always @(posedge clk) if (n983) n87 <= 1'b0 ? 1'b0 : n4322;
/* FF 13 11  0 */ always @(posedge clk) if (n1137) n1441 <= 1'b0 ? 1'b0 : n4323;
/* FF 18  2  3 */ always @(posedge clk) if (n2207) n2202 <= 1'b0 ? 1'b0 : n4324;
/* FF 13 22  7 */ always @(posedge clk) if (n1069) n1523 <= 1'b0 ? 1'b0 : n4325;
/* FF 18 15  4 */ always @(posedge clk) if (n1) n2311 <= 1'b0 ? 1'b0 : n4326;
/* FF 14 26  7 */ always @(posedge clk) if (n1271) n1718 <= 1'b0 ? 1'b0 : n4327;
/* FF 26 14  0 */ always @(posedge clk) if (n3527) n3533 <= 1'b0 ? 1'b0 : n4328;
/* FF 14 15  0 */ always @(posedge clk) if (n1792) n1639 <= 1'b0 ? 1'b0 : n4329;
/* FF  2  9  5 */ always @(posedge clk) if (n153) n162 <= 1'b0 ? 1'b0 : n4330;
/* FF 20  4  5 */ always @(posedge clk) if (n1761) n2655 <= 1'b0 ? 1'b0 : n4331;
/* FF 19 20  5 */ always @(posedge clk) if (n2553) n2570 <= 1'b0 ? 1'b0 : n4332;
/* FF 19 11  4 */ always @(posedge clk) if (n2076) n2490 <= 1'b0 ? 1'b0 : n4333;
/* FF 23  9  7 */ always @(posedge clk) if (n2678) n2690 <= 1'b0 ? 1'b0 : n4334;
/* FF 22 19  3 */ assign n3087 = n4335;
/* FF 10  5  0 */ always @(posedge clk) if (en_in) n966 <= 1'b0 ? 1'b0 : n4336;
/* FF 24 18  3 */ always @(posedge clk) if (n3411) n3405 <= 1'b0 ? 1'b0 : n4337;
/* FF 28 13  5 */ always @(posedge clk) if (n3233) n3760 <= 1'b0 ? 1'b0 : n4338;
/* FF 21  9  2 */ always @(posedge clk) if (n2856) n2847 <= 1'b0 ? 1'b0 : n4339;
/* FF  9 27  1 */ always @(posedge clk) if (n804) n947 <= 1'b0 ? 1'b0 : n4340;
/* FF  3 17  6 */ always @(posedge clk) if (n79) n315 <= 1'b0 ? 1'b0 : n4341;
/* FF 14 25  3 */ always @(posedge clk) if (n697) n1704 <= 1'b0 ? 1'b0 : n4342;
/* FF 29 21  7 */ always @(posedge clk) if (n3788) n3881 <= 1'b0 ? 1'b0 : n4343;
/* FF 17 15  6 */ always @(posedge clk) if (n2111) n2107 <= 1'b0 ? 1'b0 : n4344;
/* FF 20  7  1 */ always @(posedge clk) if (n2670) n2662 <= 1'b0 ? 1'b0 : n4345;
/* FF  5 14  2 */ always @(posedge clk) if (n402) n506 <= 1'b0 ? 1'b0 : n4346;
/* FF 11 21  3 */ always @(posedge clk) if (n819) n1199 <= 1'b0 ? 1'b0 : n4347;
/* FF 11 24  4 */ always @(posedge clk) if (n796) n1227 <= 1'b0 ? 1'b0 : n4348;
/* FF 16 17  1 */ always @(posedge clk) if (n2110) n1964 <= 1'b0 ? 1'b0 : n4349;
/* FF 22 13  3 */ always @(posedge clk) if (n2085) n3046 <= 1'b0 ? 1'b0 : n4350;
/* FF 21 27  7 */ always @(posedge clk) if (n2196) n2978 <= 1'b0 ? 1'b0 : n4351;
/* FF 27  6  4 */ assign n3488 = n4352;
/* FF 13 15  5 */ always @(posedge clk) if (n739) n1475 <= 1'b0 ? 1'b0 : n4353;
/* FF 30 12  5 */ always @(posedge clk) if (n3892) n3899 <= 1'b0 ? 1'b0 : n4354;
/* FF  9 24  5 */ always @(posedge clk) if (n820) n937 <= 1'b0 ? 1'b0 : n4355;
/* FF 13 26  2 */ always @(posedge clk) if (n1271) n1546 <= 1'b0 ? 1'b0 : n4356;
/* FF 18 19  7 */ always @(posedge clk) if (n1982) n2346 <= 1'b0 ? 1'b0 : n4357;
/* FF  3 18  0 */ always @(posedge clk) if (n215) n318 <= 1'b0 ? 1'b0 : n4358;
/* FF  6  8  1 */ always @(posedge clk) if (n570) n581 <= 1'b0 ? 1'b0 : n4359;
/* FF 18 28  6 */ always @(posedge clk) if (n2020) n2406 <= 1'b0 ? 1'b0 : n4360;
/* FF 20 21  0 */ always @(posedge clk) if (n2553) n2768 <= 1'b0 ? 1'b0 : n4361;
/* FF  1 19  6 */ always @(posedge clk) if (n119) n110 <= 1'b0 ? 1'b0 : n4362;
/* FF 28 17  3 */ always @(posedge clk) if (n3765) n3769 <= 1'b0 ? 1'b0 : n4363;
/* FF 16 15  0 */ always @(posedge clk) if (n739) n1943 <= 1'b0 ? 1'b0 : n4364;
/* FF 19  7  1 */ always @(posedge clk) if (n2670) n2453 <= 1'b0 ? 1'b0 : n4365;
/* FF 23 13  4 */ always @(posedge clk) if (n3045) n3212 <= 1'b0 ? 1'b0 : n4366;
/* FF 10 25  7 */ always @(posedge clk) if (n567) n1086 <= 1'b0 ? 1'b0 : n4367;
/* FF 24 14  4 */ always @(posedge clk) if (n3376) n3373 <= 1'b0 ? 1'b0 : n4368;
/* FF 10 18  6 */ always @(posedge clk) if (n1187) n1039 <= 1'b0 ? 1'b0 : n4369;
/* FF  9 10  4 */ always @(posedge clk) if (n988) n838 <= 1'b0 ? 1'b0 : n4370;
/* FF 13 12  1 */ always @(posedge clk) if (n1137) n1450 <= 1'b0 ? 1'b0 : n4371;
/* FF 31 25  1 */ assign \rco[128]  = n4372;
/* FF 18  5  2 */ always @(posedge clk) if (n2230) n2223 <= 1'b0 ? 1'b0 : n4373;
/* FF 20 27  3 */ always @(posedge clk) if (n2195) n2817 <= 1'b0 ? 1'b0 : n4374;
/* FF 14 21  6 */ assign n1402 = n4375;
/* FF 12 20  0 */ assign n1205 = n4376;
/* FF 14 14  7 */ always @(posedge clk) if (n1791) n1638 <= 1'b0 ? 1'b0 : n4377;
/* FF 17 11  3 */ always @(posedge clk) if (n2076) n2069 <= 1'b0 ? 1'b0 : n4378;
/* FF  1 16  0 */ always @(posedge clk) if (n85) n88 <= 1'b0 ? 1'b0 : n4379;
/* FF 19 21  2 */ always @(posedge clk) if (n2164) n2578 <= 1'b0 ? 1'b0 : n4380;
/* FF 19  8  5 */ always @(posedge clk) if (n2451) n2466 <= 1'b0 ? 1'b0 : n4381;
/* FF 23 14  6 */ always @(posedge clk) if (n2551) n3220 <= 1'b0 ? 1'b0 : n4382;
/* FF 24 17  2 */ always @(posedge clk) if (n2123) n3396 <= 1'b0 ? 1'b0 : n4383;
/* FF 28  7  3 */ always @(posedge clk) if (n3488) n3722 <= 1'b0 ? 1'b0 : n4384;
/* FF  3 14  2 */ assign n288 = n4385;
/* FF 21 10  3 */ assign n2856 = n4386;
/* FF  9 20  0 */ assign n4387 = n1056;
/* FF  7 19  2 */ always @(posedge clk) if (n549) n759 <= 1'b0 ? 1'b0 : n4388;
/* FF 26 19  0 */ assign n2730 = n4389;
/* FF 27  9  2 */ always @(posedge clk) if (n3621) n3612 <= 1'b0 ? 1'b0 : n4390;
/* FF 14 24  0 */ assign n4391 = n1873;
/* FF 17  5  4 */ assign \rco[173]  = n4392;
/* FF 17  8  7 */ assign n2055 = n4393;
/* FF  2  7  4 */ always @(posedge clk) if (n21) n150 <= 1'b0 ? 1'b0 : n4394;
/* FF 11 18  2 */ always @(posedge clk) if (n1187) n1181 <= 1'b0 ? 1'b0 : n4395;
/* FF  4 12  5 */ always @(posedge clk) if (n77) n398 <= 1'b0 ? 1'b0 : n4396;
/* FF 22 12  0 */ always @(posedge clk) if (n3029) n3036 <= 1'b0 ? 1'b0 : n4397;
/* FF 10 22  3 */ assign n4398 = n1213;
/* FF 21 28  6 */ always @(posedge clk) if (n2196) n2985 <= 1'b0 ? 1'b0 : n4399;
/* FF 13 16  4 */ always @(posedge clk) if (n922) n1481 <= 1'b0 ? 1'b0 : n4400;
/* FF 27  7  7 */ always @(posedge clk) if (n3459) n3602 <= 1'b0 ? 1'b0 : n4401;
/* FF  9 25  6 */ always @(posedge clk) if (n2) n941 <= 1'b0 ? 1'b0 : n4402;
/* FF 27 10  4 */ assign n3460 = n4403;
/* FF 13 27  5 */ always @(posedge clk) if (n1532) n1554 <= 1'b0 ? 1'b0 : n4404;
/* FF 18 18  0 */ always @(posedge clk) if (n1825) n2334 <= 1'b0 ? 1'b0 : n4405;
/* FF  3 19  3 */ always @(posedge clk) if (n115) n330 <= 1'b0 ? 1'b0 : n4406;
/* FF  6 11  0 */ always @(posedge clk) if (n286) n599 <= 1'b0 ? 1'b0 : n4407;
/* FF 23 18  0 */ always @(posedge clk) if (n2573) n3242 <= 1'b0 ? 1'b0 : n4408;
/* FF 14 10  4 */ always @(posedge clk) if (n1622) n1608 <= 1'b0 ? 1'b0 : n4409;
/* FF 19 17  7 */ always @(posedge clk) if (n2727) n2548 <= 1'b0 ? 1'b0 : n4410;
/* FF  5 17  1 */ always @(posedge clk) if (n2) n525 <= 1'b0 ? 1'b0 : n4411;
/* FF  4 15  1 */ always @(posedge clk) if (n207) n413 <= 1'b0 ? 1'b0 : n4412;
/* FF 10 24  4 */ always @(posedge clk) if (n820) n1076 <= 1'b0 ? 1'b0 : n4413;
/* FF 28 11  6 */ assign n1752 = n4414;
/* FF 24 13  5 */ always @(posedge clk) if (n3351) n2895 <= 1'b0 ? 1'b0 : n4415;
/* FF 10 21  7 */ always @(posedge clk) if (n818) n1064 <= 1'b0 ? 1'b0 : n4416;
/* FF 13 13  2 */ always @(posedge clk) if (n1015) n1457 <= 1'b0 ? 1'b0 : n4417;
/* FF 18  4  1 */ always @(posedge clk) if (n2207) n2214 <= 1'b0 ? 1'b0 : n4418;
/* FF 20 26  0 */ always @(posedge clk) if (n2615) n2805 <= 1'b0 ? 1'b0 : n4419;
/* FF 14 20  5 */ always @(posedge clk) if (n1347) n674 <= 1'b0 ? 1'b0 : n4420;
/* FF 12 27  1 */ assign n4421 = n1559;
/* FF 17 20  2 */ always @(posedge clk) if (n1843) n2138 <= 1'b0 ? 1'b0 : n4422;
/* FF 19 18  3 */ always @(posedge clk) if (n2348) n2557 <= 1'b0 ? 1'b0 : n4423;
/* FF 23 15  5 */ always @(posedge clk) if (n3216) n3227 <= 1'b0 ? 1'b0 : n4424;
/* FF 28  6  0 */ always @(posedge clk) if (n3594) n3711 <= 1'b0 ? 1'b0 : n4425;
/* FF  3 15  1 */ always @(posedge clk) if (n207) n294 <= 1'b0 ? 1'b0 : n4426;
/* FF 21 16  5 */ always @(posedge clk) if (n2551) n2892 <= 1'b0 ? 1'b0 : n4427;
/* FF  7 16  3 */ always @(posedge clk) if (n630) n744 <= 1'b0 ? 1'b0 : n4428;
/* FF  9 21  3 */ always @(posedge clk) if (n818) n917 <= 1'b0 ? 1'b0 : n4429;
/* FF 21 11  4 */ always @(posedge clk) if (n2085) n2861 <= 1'b0 ? 1'b0 : n4430;
/* FF 26 18  7 */ assign \rco[36]  = n4431;
/* FF 18 22  5 */ assign n2358 = n4432;
/* FF 14 27  1 */ always @(posedge clk) if (n1402) n1719 <= 1'b0 ? 1'b0 : n4433;
/* FF 17  6  5 */ always @(posedge clk) if (n2045) n2043 <= 1'b0 ? 1'b0 : n4434;
/* FF 17  9  4 */ assign n1 = n4435;
/* FF 28 20  1 */ assign n3785 = n3876;
/* FF 22 26  6 */ always @(posedge clk) if (n2613) n3139 <= 1'b0 ? 1'b0 : n4436;
/* FF 22 15  1 */ always @(posedge clk) if (n3216) n3059 <= 1'b0 ? 1'b0 : n4437;
/* FF  7  6  6 */ always @(posedge clk) if (n588) n710 <= 1'b0 ? 1'b0 : n4438;
/* FF  9  7  0 */ assign n588 = n4439;
/* FF 13 17  7 */ always @(posedge clk) if (n1461) n1490 <= 1'b0 ? 1'b0 : n4440;
/* FF 13 28  4 */ always @(posedge clk) if (n1394) n1565 <= 1'b0 ? 1'b0 : n4441;
/* FF 18 21  1 */ always @(posedge clk) if (n2347) n2350 <= 1'b0 ? 1'b0 : n4442;
/* FF  3 16  2 */ always @(posedge clk) if (n197) n305 <= 1'b0 ? 1'b0 : n4443;
/* FF 23 19  3 */ always @(posedge clk) if (n2573) n3253 <= 1'b0 ? 1'b0 : n4444;
/* FF 14  5  5 */ always @(posedge clk) if (n1577) n1576 <= 1'b0 ? 1'b0 : n4445;
/* FF 19 14  6 */ always @(posedge clk) if (n2123) n2517 <= 1'b0 ? 1'b0 : n4446;
/* FF 17 27  0 */ always @(posedge clk) if (n1) n2188 <= 1'b0 ? 1'b0 : n4447;
/* FF 28 23  5 */ always @(posedge clk) if (n3704) n2796 <= 1'b0 ? 1'b0 : n4448;
/* FF  5 18  0 */ always @(posedge clk) if (n657) n531 <= 1'b0 ? 1'b0 : n4449;
/* FF  4 14  2 */ assign n4450 = n513;
/* FF 19  5  7 */ always @(posedge clk) if (n2230) n2442 <= 1'b0 ? 1'b0 : n4451;
/* FF 10 27  5 */ always @(posedge clk) if (n804) n1087 <= 1'b0 ? 1'b0 : n4452;
/* FF 22 25  0 */ always @(posedge clk) if (n2812) n3125 <= 1'b0 ? 1'b0 : n4453;
/* FF 24 12  2 */ always @(posedge clk) if (n3351) n3355 <= 1'b0 ? 1'b0 : n4454;
/* FF 28 10  5 */ always @(posedge clk) if (n3462) n3746 <= 1'b0 ? 1'b0 : n4455;
/* FF 10 20  4 */ always @(posedge clk) if (n922) n1052 <= 1'b0 ? 1'b0 : n4456;
/* FF 13 14  3 */ always @(posedge clk) if (n1461) n1465 <= 1'b0 ? 1'b0 : n4457;
/* FF 18  7  0 */ always @(posedge clk) if (n1761) n2239 <= 1'b0 ? 1'b0 : n4458;
/* FF 20 25  1 */ always @(posedge clk) if (n2612) n2799 <= 1'b0 ? 1'b0 : n4459;
/* FF 15  5  6 */ always @(posedge clk) if (n1742) n1730 <= 1'b0 ? 1'b0 : n4460;
/* FF 14 23  4 */ always @(posedge clk) if (n820) n1231 <= 1'b0 ? 1'b0 : n4461;
/* FF 12 26  2 */ always @(posedge clk) if (n1393) n1387 <= 1'b0 ? 1'b0 : n4462;
/* FF 14  8  5 */ always @(posedge clk) if (n1741) n1598 <= 1'b0 ? 1'b0 : n4463;
/* FF  2 10  0 */ always @(posedge clk) if (n168) n165 <= 1'b0 ? 1'b0 : n4464;
/* FF  1 18  2 */ always @(posedge clk) if (n115) n100 <= 1'b0 ? 1'b0 : n4465;
/* FF 19 19  0 */ assign \rco[166]  = n4466;
/* FF 17 21  1 */ always @(posedge clk) if (n2347) n2145 <= 1'b0 ? 1'b0 : n4467;
/* FF 23 12  4 */ always @(posedge clk) if (n3031) n3204 <= 1'b0 ? 1'b0 : n4468;
/* FF 28  5  1 */ always @(posedge clk) if (n3488) n3706 <= 1'b0 ? 1'b0 : n4469;
/* FF  3 12  0 */ assign n251 = n4470;
/* FF 21 17  6 */ always @(posedge clk) if (n2519) n2900 <= 1'b0 ? 1'b0 : n4471;
/* FF  7 17  4 */ always @(posedge clk) if (n549) n755 <= 1'b0 ? 1'b0 : n4472;
/* FF 21 12  5 */ always @(posedge clk) if (n3029) n2857 <= 1'b0 ? 1'b0 : n4473;
/* FF 12  8  7 */ always @(posedge clk) if (n1131) n1282 <= 1'b0 ? 1'b0 : n4474;
/* FF 26 21  6 */ always @(posedge clk) if (n3421) n3567 <= 1'b0 ? 1'b0 : n4475;
/* FF 15  6  0 */ always @(posedge clk) if (n1744) n1733 <= 1'b0 ? 1'b0 : n4476;
/* FF 17  7  2 */ always @(posedge clk) if (n2045) n2048 <= 1'b0 ? 1'b0 : n4477;
/* FF 18 25  4 */ always @(posedge clk) if (n1878) n2381 <= 1'b0 ? 1'b0 : n4478;
/* FF 17 10  5 */ always @(posedge clk) if (n2282) n2064 <= 1'b0 ? 1'b0 : n4479;
/* FF 11 16  0 */ always @(posedge clk) if (n891) n1159 <= 1'b0 ? 1'b0 : n4480;
/* FF 10  8  2 */ assign \rco[152]  = n4481;
/* FF  1 12  2 */ always @(posedge clk) if (n39) n48 <= 1'b0 ? 1'b0 : n4482;
/* FF 22 14  6 */ always @(posedge clk) if (n3045) n3056 <= 1'b0 ? 1'b0 : n4483;
/* FF  7  7  5 */ always @(posedge clk) if (n588) n714 <= 1'b0 ? 1'b0 : n4484;
/* FF 13 18  6 */ always @(posedge clk) if (n1205) n1498 <= 1'b0 ? 1'b0 : n4485;
/* FF 27  5  1 */ always @(posedge clk) if (n3594) n3586 <= 1'b0 ? 1'b0 : n4486;
/* FF 27  8  6 */ always @(posedge clk) if (n3464) n3608 <= 1'b0 ? 1'b0 : n4487;
/* FF 23 16  2 */ assign \rco[38]  = n3393;
/* FF 11 14  3 */ always @(posedge clk) if (n1154) n1149 <= 1'b0 ? 1'b0 : n4488;
/* FF  2 14  5 */ always @(posedge clk) if (n83) n192 <= 1'b0 ? 1'b0 : n4489;
/* FF 16  7  4 */ always @(posedge clk) if (n1743) n1911 <= 1'b0 ? 1'b0 : n4490;
/* FF 19 15  5 */ always @(posedge clk) if (n2715) n2530 <= 1'b0 ? 1'b0 : n4491;
/* FF 28 22  6 */ always @(posedge clk) if (n3704) n3805 <= 1'b0 ? 1'b0 : n4492;
/* FF 16 12  5 */ always @(posedge clk) if (n1771) n1940 <= 1'b0 ? 1'b0 : n4493;
/* FF  5 19  7 */ always @(posedge clk) if (n349) n538 <= 1'b0 ? 1'b0 : n4494;
/* FF  4 13  3 */ assign n402 = n4495;
/* FF 22 24  3 */ always @(posedge clk) if (n3113) n3119 <= 1'b0 ? 1'b0 : n4496;
/* FF 24 11  3 */ assign n3351 = n4497;
/* FF 10 26  2 */ assign \rco[106]  = n4498;
/* FF 28  9  4 */ always @(posedge clk) if (n3621) n3738 <= 1'b0 ? 1'b0 : n4499;
/* FF 10 23  5 */ always @(posedge clk) if (n821) n1066 <= 1'b0 ? 1'b0 : n4500;
/* FF  7 21  1 */ always @(posedge clk) if (n360) n361 <= 1'b0 ? 1'b0 : n4501;
/* FF  6  7  1 */ always @(posedge clk) if (n570) n572 <= 1'b0 ? 1'b0 : n4502;
/* FF 20 24  6 */ always @(posedge clk) if (n2775) n2794 <= 1'b0 ? 1'b0 : n4503;
/* FF 26  9  5 */ always @(posedge clk) if (n3460) n3503 <= 1'b0 ? 1'b0 : n4504;
/* FF 29 17  4 */ always @(posedge clk) if (n3765) n3858 <= 1'b0 ? 1'b0 : n4505;
/* FF 14 22  3 */ always @(posedge clk) if (n1402) n1690 <= 1'b0 ? 1'b0 : n4506;
/* FF 12 25  3 */ always @(posedge clk) if (n1532) n1379 <= 1'b0 ? 1'b0 : n4507;
/* FF 14 11  4 */ always @(posedge clk) if (n1622) n1616 <= 1'b0 ? 1'b0 : n4508;
/* FF 17 22  0 */ always @(posedge clk) if (n1999) n2152 <= 1'b0 ? 1'b0 : n4509;
/* FF 19 16  1 */ assign n2270 = n4510;
/* FF 23  6  2 */ always @(posedge clk) if (n3158) n3161 <= 1'b0 ? 1'b0 : n4511;
/* FF 16 26  1 */ always @(posedge clk) if (n1557) n2013 <= 1'b0 ? 1'b0 : n4512;
/* FF  4 19  3 */ assign n438 = n4513;
/* FF  3 13  7 */ assign \rco[11]  = n4514;
/* FF 21 18  7 */ always @(posedge clk) if (n2757) n2909 <= 1'b0 ? 1'b0 : n4515;
/* FF 22 10  3 */ always @(posedge clk) if (n2856) n3025 <= 1'b0 ? 1'b0 : n4516;
/* FF  7 22  5 */ always @(posedge clk) if (n695) n788 <= 1'b0 ? 1'b0 : n4517;
/* FF  9 23  5 */ always @(posedge clk) if (n819) n930 <= 1'b0 ? 1'b0 : n4518;
/* FF 21 13  6 */ always @(posedge clk) if (n2519) n2880 <= 1'b0 ? 1'b0 : n4519;
/* FF 12 15  6 */ always @(posedge clk) if (n1155) n1302 <= 1'b0 ? 1'b0 : n4520;
/* FF 26 20  5 */ assign n3259 = n3685;
/* FF 15  7  3 */ assign \rco[83]  = n1914;
/* FF 19 30  0 */ always @(posedge clk) if (n2592) n2634 <= 1'b0 ? 1'b0 : n4521;
/* FF 10 11  3 */ always @(posedge clk) if (n996) n991 <= 1'b0 ? 1'b0 : n4522;
/* FF 16  8  2 */ always @(posedge clk) if (n1625) n1917 <= 1'b0 ? 1'b0 : n4523;
/* FF  1 13  1 */ always @(posedge clk) if (n83) n60 <= 1'b0 ? 1'b0 : n4524;
/* FF 22  4  4 */ assign \rco[45]  = n4525;
/* FF 13 19  1 */ assign \rco[142]  = n4526;
/* FF 15 21  0 */ always @(posedge clk) if (n1356) n1836 <= 1'b0 ? 1'b0 : n4527;
/* FF 20 28  3 */ always @(posedge clk) if (n2195) n2824 <= 1'b0 ? 1'b0 : n4528;
/* FF 18 23  3 */ always @(posedge clk) if (n1999) n2365 <= 1'b0 ? 1'b0 : n4529;
/* FF 23 17  5 */ always @(posedge clk) if (n2540) n3237 <= 1'b0 ? 1'b0 : n4530;
/* FF 11 15  0 */ assign n750 = n4531;
/* FF 26  6  1 */ always @(posedge clk) if (n3459) n3474 <= 1'b0 ? 1'b0 : n4532;
/* FF 14  7  7 */ always @(posedge clk) if (n1743) n1591 <= 1'b0 ? 1'b0 : n4533;
/* FF 16  6  7 */ always @(posedge clk) if (n1744) n1904 <= 1'b0 ? 1'b0 : n4534;
/* FF 19 12  4 */ always @(posedge clk) if (n1936) n2501 <= 1'b0 ? 1'b0 : n4535;
/* FF 28 21  7 */ always @(posedge clk) if (n3788) n3798 <= 1'b0 ? 1'b0 : n4536;
/* FF 19  3  5 */ always @(posedge clk) if (n1887) n2432 <= 1'b0 ? 1'b0 : n4537;
/* FF 22 27  2 */ always @(posedge clk) if (n2970) n3145 <= 1'b0 ? 1'b0 : n4538;
/* FF 10 29  3 */ always @(posedge clk) if (n821) n1111 <= 1'b0 ? 1'b0 : n4539;
/* FF 24 10  0 */ always @(posedge clk) if (n3352) n3340 <= 1'b0 ? 1'b0 : n4540;
/* FF 28  8  3 */ always @(posedge clk) if (n3605) n3729 <= 1'b0 ? 1'b0 : n4541;
/* FF  3  9  4 */ always @(posedge clk) if (n260) n256 <= 1'b0 ? 1'b0 : n4542;
/* FF  7 26  0 */ always @(posedge clk) if (n567) n798 <= 1'b0 ? 1'b0 : n4543;
/* FF  9 19  2 */ always @(posedge clk) if (n454) n903 <= 1'b0 ? 1'b0 : n4544;
/* FF 12 19  5 */ always @(posedge clk) if (n1501) n446 <= 1'b0 ? 1'b0 : n4545;
/* FF 26  8  6 */ always @(posedge clk) if (n3603) n3496 <= 1'b0 ? 1'b0 : n4546;
/* FF 29 18  5 */ always @(posedge clk) if (n3765) n3860 <= 1'b0 ? 1'b0 : n4547;
/* FF 14 17  2 */ always @(posedge clk) if (n1672) n1656 <= 1'b0 ? 1'b0 : n4548;
/* FF 12 24  4 */ always @(posedge clk) if (n961) n1371 <= 1'b0 ? 1'b0 : n4549;
/* FF 17 12  6 */ always @(posedge clk) if (n2056) n2083 <= 1'b0 ? 1'b0 : n4550;
/* FF  2 12  2 */ always @(posedge clk) if (n39) n178 <= 1'b0 ? 1'b0 : n4551;
/* FF 23  7  1 */ always @(posedge clk) if (n3006) n3167 <= 1'b0 ? 1'b0 : n4552;
/* FF 22 21  1 */ always @(posedge clk) if (n2564) n3097 <= 1'b0 ? 1'b0 : n4553;
/* FF 24 24  1 */ always @(posedge clk) if (n3112) n3440 <= 1'b0 ? 1'b0 : n4554;
/* FF 16 25  0 */ assign n1557 = n4555;
/* FF  4 18  0 */ always @(posedge clk) if (n349) n430 <= 1'b0 ? 1'b0 : n4556;
/* FF  3 10  6 */ always @(posedge clk) if (n251) n268 <= 1'b0 ? 1'b0 : n4557;
/* FF 21 19  0 */ always @(posedge clk) if (n2757) n2911 <= 1'b0 ? 1'b0 : n4558;
/* FF 13 23  6 */ always @(posedge clk) if (n1069) n1530 <= 1'b0 ? 1'b0 : n4559;
/* FF 27 14  7 */ always @(posedge clk) if (n3527) n3648 <= 1'b0 ? 1'b0 : n4560;
/* FF  7 23  6 */ always @(posedge clk) if (n454) n793 <= 1'b0 ? 1'b0 : n4561;
/* FF  9 16  4 */ always @(posedge clk) if (n645) n879 <= 1'b0 ? 1'b0 : n4562;
/* FF 12 14  5 */ always @(posedge clk) if (n1154) n1293 <= 1'b0 ? 1'b0 : n4563;
/* FF 26 23  4 */ always @(posedge clk) if (n3703) n3580 <= 1'b0 ? 1'b0 : n4564;
/* FF 18 27  6 */ always @(posedge clk) if (n2020) n2398 <= 1'b0 ? 1'b0 : n4565;
/* FF  5  8  0 */ always @(posedge clk) if (n21) n468 <= 1'b0 ? 1'b0 : n4566;
/* FF 19 31  3 */ always @(posedge clk) if (n2592) n2644 <= 1'b0 ? 1'b0 : n4567;
/* FF 23 21  2 */ always @(posedge clk) if (n3258) n3273 <= 1'b0 ? 1'b0 : n4568;
/* FF 10 10  4 */ always @(posedge clk) if (n983) n987 <= 1'b0 ? 1'b0 : n4569;
/* FF 16 23  3 */ always @(posedge clk) if (n2000) n1994 <= 1'b0 ? 1'b0 : n4570;
/* FF  1 14  0 */ always @(posedge clk) if (n85) n68 <= 1'b0 ? 1'b0 : n4571;
/* FF 22  7  5 */ always @(posedge clk) if (n2841) n3003 <= 1'b0 ? 1'b0 : n4572;
/* FF 10 17  6 */ assign n823 = n1178;
/* FF 24  6  5 */ always @(posedge clk) if (n3006) n3326 <= 1'b0 ? 1'b0 : n4573;
/* FF 22  8  4 */ always @(posedge clk) if (n2989) n3012 <= 1'b0 ? 1'b0 : n4574;
/* FF 13 20  0 */ always @(posedge clk) if (n1339) n1503 <= 1'b0 ? 1'b0 : n4575;
/* FF 15 10  1 */ always @(posedge clk) if (n1624) n1755 <= 1'b0 ? 1'b0 : n4576;
/* FF  2 16  0 */ always @(posedge clk) if (n197) n204 <= 1'b0 ? 1'b0 : n4577;
/* FF 20 19  2 */ always @(posedge clk) if (n2562) n2751 <= 1'b0 ? 1'b0 : n4578;
/* FF 12 28  1 */ always @(posedge clk) if (n1394) n1395 <= 1'b0 ? 1'b0 : n4579;
/* FF 23 22  4 */ always @(posedge clk) if (n3422) n3283 <= 1'b0 ? 1'b0 : n4580;
/* FF 14  6  0 */ assign n977 = n4581;
/* FF 16  5  6 */ always @(posedge clk) if (n1742) n1894 <= 1'b0 ? 1'b0 : n4582;
/* FF 17 19  4 */ always @(posedge clk) if (n1982) n2132 <= 1'b0 ? 1'b0 : n4583;
/* FF 19 13  3 */ always @(posedge clk) if (n2283) n2508 <= 1'b0 ? 1'b0 : n4584;
/* FF 16 10  7 */ always @(posedge clk) if (n1771) n1932 <= 1'b0 ? 1'b0 : n4585;
/* FF  5 21  5 */ assign n554 = n4586;
/* FF 10 28  0 */ always @(posedge clk) if (n821) n1101 <= 1'b0 ? 1'b0 : n4587;
/* FF 24  9  1 */ always @(posedge clk) if (n3352) n3333 <= 1'b0 ? 1'b0 : n4588;
/* FF 27 17  0 */ always @(posedge clk) if (n3249) n3408 <= 1'b0 ? 1'b0 : n4589;
/* FF 15 24  0 */ always @(posedge clk) if (n778) n1864 <= 1'b0 ? 1'b0 : n4590;
/* FF 21 23  5 */ always @(posedge clk) if (n2961) n2948 <= 1'b0 ? 1'b0 : n4591;
/* FF 12 18  6 */ always @(posedge clk) if (n1501) n1326 <= 1'b0 ? 1'b0 : n4592;
/* FF 26 11  7 */ always @(posedge clk) if (n3033) n3515 <= 1'b0 ? 1'b0 : n4593;
/* FF 29 19  2 */ always @(posedge clk) if (n3786) n3863 <= 1'b0 ? 1'b0 : n4594;
/* FF 14 16  1 */ always @(posedge clk) if (n1792) n1647 <= 1'b0 ? 1'b0 : n4595;
/* FF 17 13  5 */ always @(posedge clk) if (n2056) n2091 <= 1'b0 ? 1'b0 : n4596;
/* FF 17 16  6 */ assign n2113 = n2325;
/* FF  2 15  3 */ always @(posedge clk) if (n197) n198 <= 1'b0 ? 1'b0 : n4597;
/* FF 22 20  2 */ always @(posedge clk) if (n3087) n3090 <= 1'b0 ? 1'b0 : n4598;
/* FF 10 14  1 */ always @(posedge clk) if (n750) n1008 <= 1'b0 ? 1'b0 : n4599;
/* FF 24 23  0 */ always @(posedge clk) if (n3104) n3433 <= 1'b0 ? 1'b0 : n4600;
/* FF  4 17  1 */ always @(posedge clk) if (n2) n225 <= 1'b0 ? 1'b0 : n4601;
/* FF  3 11  5 */ always @(posedge clk) if (n153) n261 <= 1'b0 ? 1'b0 : n4602;
/* FF  7  9  0 */ assign n718 = n4603;
/* FF 21 20  1 */ always @(posedge clk) if (n3087) n2919 <= 1'b0 ? 1'b0 : n4604;
/* FF 13 24  7 */ assign n224 = n4605;
/* FF  9 17  7 */ always @(posedge clk) if (n1030) n890 <= 1'b0 ? 1'b0 : n4606;
/* FF 19 22  0 */ always @(posedge clk) if (n2164) n2584 <= 1'b0 ? 1'b0 : n4607;
/* FF 18 26  1 */ always @(posedge clk) if (n2615) n2386 <= 1'b0 ? 1'b0 : n4608;
/* FF 17  2  1 */ assign \rco[85]  = n4609;
/* FF 20 12  0 */ always @(posedge clk) if (n2682) n2698 <= 1'b0 ? 1'b0 : n4610;
/* FF  5  9  3 */ always @(posedge clk) if (n21) n474 <= 1'b0 ? 1'b0 : n4611;
/* FF 28 19  4 */ always @(posedge clk) if (n3424) n3781 <= 1'b0 ? 1'b0 : n4612;
/* FF 10 13  5 */ always @(posedge clk) if (n629) n1006 <= 1'b0 ? 1'b0 : n4613;
/* FF 16 22  0 */ assign n1835 = n4614;
/* FF 22  6  2 */ always @(posedge clk) if (n2841) n2992 <= 1'b0 ? 1'b0 : n4615;
/* FF 10 16  5 */ always @(posedge clk) if (n891) n738 <= 1'b0 ? 1'b0 : n4616;
/* FF 24  5  4 */ always @(posedge clk) if (n3158) n3320 <= 1'b0 ? 1'b0 : n4617;
/* FF 22 11  5 */ assign n3033 = n4618;
/* FF 13 21  3 */ always @(posedge clk) if (n1356) n1516 <= 1'b0 ? 1'b0 : n4619;
/* FF 15 11  2 */ always @(posedge clk) if (n1624) n1765 <= 1'b0 ? 1'b0 : n4620;
/* FF  2 19  1 */ assign n116 = n339;
/* FF  6 13  2 */ always @(posedge clk) if (n78) n617 <= 1'b0 ? 1'b0 : n4621;
/* FF 20 18  1 */ always @(posedge clk) if (n2348) n2742 <= 1'b0 ? 1'b0 : n4622;
/* FF 23 23  7 */ always @(posedge clk) if (n3104) n3294 <= 1'b0 ? 1'b0 : n4623;
/* FF 11 13  6 */ always @(posedge clk) if (n733) n1144 <= 1'b0 ? 1'b0 : n4624;
/* FF 19 10  2 */ always @(posedge clk) if (n2678) n2481 <= 1'b0 ? 1'b0 : n4625;
/* FF  5 22  4 */ always @(posedge clk) if (n673) n559 <= 1'b0 ? 1'b0 : n4626;
/* FF 28 14  1 */ always @(posedge clk) if (n2085) n3762 <= 1'b0 ? 1'b0 : n4627;
/* FF 13  7  0 */ always @(posedge clk) if (n977) n1423 <= 1'b0 ? 1'b0 : n4628;
/* FF 15 25  7 */ always @(posedge clk) if (n1878) n1551 <= 1'b0 ? 1'b0 : n4629;
/* FF  7 13  5 */ assign \rco[161]  = n4630;
/* FF 12 17  7 */ always @(posedge clk) if (n900) n1319 <= 1'b0 ? 1'b0 : n4631;
/* FF 26 10  0 */ always @(posedge clk) if (n3033) n3505 <= 1'b0 ? 1'b0 : n4632;
/* FF 18 30  6 */ always @(posedge clk) if (n1881) n2422 <= 1'b0 ? 1'b0 : n4633;
/* FF 14 19  0 */ assign n4634 = n1826;
/* FF 17 14  4 */ always @(posedge clk) if (n1625) n2098 <= 1'b0 ? 1'b0 : n4635;
/* FF 26  7  7 */ always @(posedge clk) if (n3603) n3487 <= 1'b0 ? 1'b0 : n4636;
/* FF 29 20  3 */ always @(posedge clk) if (n3786) n3871 <= 1'b0 ? 1'b0 : n4637;
/* FF 17 17  5 */ always @(posedge clk) if (n2111) n2119 <= 1'b0 ? 1'b0 : n4638;
/* FF 22 23  3 */ assign n3113 = n4639;
/* FF 24 22  3 */ always @(posedge clk) if (n3422) n3428 <= 1'b0 ? 1'b0 : n4640;
/* FF  1 11  4 */ always @(posedge clk) if (n37) n41 <= 1'b0 ? 1'b0 : n4641;
/* FF  7 14  1 */ always @(posedge clk) if (n733) n735 <= 1'b0 ? 1'b0 : n4642;
/* FF 21 21  2 */ always @(posedge clk) if (n2564) n2928 <= 1'b0 ? 1'b0 : n4643;
/* FF 13 25  4 */ always @(posedge clk) if (n697) n1538 <= 1'b0 ? 1'b0 : n4644;
/* FF 27 12  5 */ always @(posedge clk) if (n3368) n3622 <= 1'b0 ? 1'b0 : n4645;
/* FF  9 18  6 */ always @(posedge clk) if (n1030) n898 <= 1'b0 ? 1'b0 : n4646;
/* FF 18 29  0 */ always @(posedge clk) if (n1881) n2408 <= 1'b0 ? 1'b0 : n4647;
/* FF  6 18  0 */ always @(posedge clk) if (n657) n649 <= 1'b0 ? 1'b0 : n4648;
/* FF  5 10  2 */ always @(posedge clk) if (n184) n476 <= 1'b0 ? 1'b0 : n4649;
/* FF 19 29  5 */ always @(posedge clk) if (n2614) n2632 <= 1'b0 ? 1'b0 : n4650;
/* FF 11  9  3 */ always @(posedge clk) if (n1131) n1133 <= 1'b0 ? 1'b0 : n4651;
/* FF 23 27  0 */ always @(posedge clk) if (n2017) n3312 <= 1'b0 ? 1'b0 : n4652;
/* FF 24 25  7 */ always @(posedge clk) if (n2812) n3310 <= 1'b0 ? 1'b0 : n4653;
/* FF 16 21  1 */ always @(posedge clk) if (n1835) n1984 <= 1'b0 ? 1'b0 : n4654;
/* FF  1  8  6 */ always @(posedge clk) if (n37) n19 <= 1'b0 ? 1'b0 : n4655;
/* FF 10 19  4 */ always @(posedge clk) if (n454) n1045 <= 1'b0 ? 1'b0 : n4656;
/* FF 13 22  2 */ assign n1520 = n4657;
/* FF 15  8  3 */ always @(posedge clk) if (n1741) n1749 <= 1'b0 ? 1'b0 : n4658;
/* FF  3 22  0 */ always @(posedge clk) if (n352) n353 <= 1'b0 ? 1'b0 : n4659;
/* FF 21  7  2 */ assign n2841 = n4660;
/* FF  6 12  1 */ always @(posedge clk) if (n286) n607 <= 1'b0 ? 1'b0 : n4661;
/* FF 20 17  0 */ always @(posedge clk) if (n2727) n2732 <= 1'b0 ? 1'b0 : n4662;
/* FF 26 14  5 */ always @(posedge clk) if (n3527) n3538 <= 1'b0 ? 1'b0 : n4663;
/* FF 23 20  6 */ always @(posedge clk) if (n3258) n3269 <= 1'b0 ? 1'b0 : n4664;
/* FF 19 11  1 */ always @(posedge clk) if (n2076) n2487 <= 1'b0 ? 1'b0 : n4665;
/* FF  4 20  3 */ always @(posedge clk) if (n215) n441 <= 1'b0 ? 1'b0 : n4666;
/* FF  7 18  4 */ always @(posedge clk) if (n215) n326 <= 1'b0 ? 1'b0 : n4667;
/* FF  9 27  6 */ always @(posedge clk) if (n804) n952 <= 1'b0 ? 1'b0 : n4668;
/* FF 21  9  7 */ always @(posedge clk) if (n2856) n2851 <= 1'b0 ? 1'b0 : n4669;
/* FF 12 16  0 */ always @(posedge clk) if (n1155) n1304 <= 1'b0 ? 1'b0 : n4670;
/* FF 26 13  1 */ assign n3526 = n3640;
/* FF 29 21  0 */ always @(posedge clk) if (n3788) n3877 <= 1'b0 ? 1'b0 : n4671;
/* FF 17 15  3 */ always @(posedge clk) if (n2111) n2104 <= 1'b0 ? 1'b0 : n4672;
/* FF 19 25  2 */ always @(posedge clk) if (n2612) n2606 <= 1'b0 ? 1'b0 : n4673;
/* FF 22 22  4 */ always @(posedge clk) if (n2961) n3109 <= 1'b0 ? 1'b0 : n4674;
/* FF 24 21  2 */ assign n3422 = n4675;
/* FF 22 13  6 */ always @(posedge clk) if (n2085) n3049 <= 1'b0 ? 1'b0 : n4676;
/* FF  7 15  2 */ assign n403 = n814;
/* FF  9 24  0 */ always @(posedge clk) if (n820) n932 <= 1'b0 ? 1'b0 : n4677;
/* FF 13 26  5 */ always @(posedge clk) if (n1271) n1244 <= 1'b0 ? 1'b0 : n4678;
/* FF 21 22  3 */ always @(posedge clk) if (n2384) n2938 <= 1'b0 ? 1'b0 : n4679;
/* FF 27 13  2 */ always @(posedge clk) if (n3460) n3638 <= 1'b0 ? 1'b0 : n4680;
/* FF  2 22  3 */ always @(posedge clk) if (n352) n238 <= 1'b0 ? 1'b0 : n4681;
/* FF 18 28  3 */ always @(posedge clk) if (n2020) n2403 <= 1'b0 ? 1'b0 : n4682;
/* FF 19 26  4 */ assign n2613 = n4683;
/* FF 23 24  1 */ always @(posedge clk) if (n3112) n3297 <= 1'b0 ? 1'b0 : n4684;
/* FF 11 22  2 */ always @(posedge clk) if (n695) n1208 <= 1'b0 ? 1'b0 : n4685;
/* FF 28 17  6 */ always @(posedge clk) if (n3765) n3771 <= 1'b0 ? 1'b0 : n4686;
/* FF 16 15  7 */ always @(posedge clk) if (n739) n1949 <= 1'b0 ? 1'b0 : n4687;
/* FF 10 15  7 */ always @(posedge clk) if (n750) n1022 <= 1'b0 ? 1'b0 : n4688;
/* FF 16 20  6 */ always @(posedge clk) if (n1843) n1980 <= 1'b0 ? 1'b0 : n4689;
/* FF 10 18  3 */ always @(posedge clk) if (n1187) n1036 <= 1'b0 ? 1'b0 : n4690;
/* FF 15 18  5 */ always @(posedge clk) if (n1355) n1813 <= 1'b0 ? 1'b0 : n4691;
/* FF 20 27  6 */ always @(posedge clk) if (n2195) n2820 <= 1'b0 ? 1'b0 : n4692;
/* FF 18 14  0 */ assign n2240 = n2523;
/* FF  2 21  7 */ always @(posedge clk) if (n126) n234 <= 1'b0 ? 1'b0 : n4693;
/* FF  6 15  0 */ assign n630 = n4694;
/* FF 20 16  7 */ assign n2551 = n4695;
/* FF 12 20  5 */ assign n545 = n4696;
/* FF 19  8  0 */ always @(posedge clk) if (n2451) n2461 <= 1'b0 ? 1'b0 : n4697;
/* FF  4 11  1 */ always @(posedge clk) if (n184) n287 <= 1'b0 ? 1'b0 : n4698;
/* FF 22 18  1 */ always @(posedge clk) if (n3065) n3081 <= 1'b0 ? 1'b0 : n4699;
/* FF 13  9  2 */ always @(posedge clk) if (n850) n1432 <= 1'b0 ? 1'b0 : n4700;
/* FF  7 19  7 */ always @(posedge clk) if (n549) n764 <= 1'b0 ? 1'b0 : n4701;
/* FF  9 20  7 */ always @(posedge clk) if (n961) n911 <= 1'b0 ? 1'b0 : n4702;
/* FF 21 10  6 */ assign \rco[48]  = n3030;
/* FF 27  9  7 */ always @(posedge clk) if (n3621) n3617 <= 1'b0 ? 1'b0 : n4703;
/* FF 21  5  7 */ always @(posedge clk) if (n2989) n2832 <= 1'b0 ? 1'b0 : n4704;
/* FF 12 23  1 */ always @(posedge clk) if (n1357) n1359 <= 1'b0 ? 1'b0 : n4705;
/* FF 26 12  2 */ always @(posedge clk) if (n3368) n3519 <= 1'b0 ? 1'b0 : n4706;
/* FF 17  8  2 */ assign n4707 = n2257;
/* FF  5 15  2 */ always @(posedge clk) if (n511) n516 <= 1'b0 ? 1'b0 : n4708;
/* FF 19 22  3 */ always @(posedge clk) if (n2164) n2587 <= 1'b0 ? 1'b0 : n4709;
/* FF 11 25  0 */ assign \rco[105]  = n4710;
/* FF 22 17  5 */ always @(posedge clk) if (n3065) n3077 <= 1'b0 ? 1'b0 : n4711;
/* FF 24 20  5 */ always @(posedge clk) if (n3411) n3417 <= 1'b0 ? 1'b0 : n4712;
/* FF 16 16  3 */ always @(posedge clk) if (n2110) n1958 <= 1'b0 ? 1'b0 : n4713;
/* FF 22 12  5 */ always @(posedge clk) if (n3029) n3041 <= 1'b0 ? 1'b0 : n4714;
/* FF  4 22  4 */ always @(posedge clk) if (n2) n463 <= 1'b0 ? 1'b0 : n4715;
/* FF  9 25  3 */ assign \rco[122]  = n4716;
/* FF 27 10  3 */ assign n3462 = n4717;
/* FF 13 27  2 */ assign n1542 = n4718;
/* FF 15 13  1 */ always @(posedge clk) if (n1015) n1778 <= 1'b0 ? 1'b0 : n4719;
/* FF 20 20  4 */ always @(posedge clk) if (n2562) n2765 <= 1'b0 ? 1'b0 : n4720;
/* FF 23 18  7 */ always @(posedge clk) if (n2573) n3248 <= 1'b0 ? 1'b0 : n4721;
/* FF  5 12  4 */ always @(posedge clk) if (n77) n488 <= 1'b0 ? 1'b0 : n4722;
/* FF 19 27  7 */ always @(posedge clk) if (n2614) n2623 <= 1'b0 ? 1'b0 : n4723;
/* FF 11 23  1 */ always @(posedge clk) if (n796) n1215 <= 1'b0 ? 1'b0 : n4724;
/* FF 23 25  6 */ always @(posedge clk) if (n2613) n3308 <= 1'b0 ? 1'b0 : n4725;
/* FF  1 10  4 */ always @(posedge clk) if (n37) n32 <= 1'b0 ? 1'b0 : n4726;
/* FF 10 21  2 */ always @(posedge clk) if (n818) n1060 <= 1'b0 ? 1'b0 : n4727;
/* FF  9 11  0 */ always @(posedge clk) if (n988) n842 <= 1'b0 ? 1'b0 : n4728;
/* FF 15 19  6 */ always @(posedge clk) if (n1355) n1823 <= 1'b0 ? 1'b0 : n4729;
/* FF 20 26  5 */ always @(posedge clk) if (n2615) n2400 <= 1'b0 ? 1'b0 : n4730;
/* FF 18 17  1 */ always @(posedge clk) if (n1825) n2326 <= 1'b0 ? 1'b0 : n4731;
/* FF  3 20  2 */ always @(posedge clk) if (n119) n344 <= 1'b0 ? 1'b0 : n4732;
/* FF  2 20  4 */ always @(posedge clk) if (n126) n221 <= 1'b0 ? 1'b0 : n4733;
/* FF 20 23  6 */ assign n1541 = n4734;
/* FF 15 14  5 */ always @(posedge clk) if (n1791) n1788 <= 1'b0 ? 1'b0 : n4735;
/* FF 12 27  4 */ assign n1383 = n4736;
/* FF 11  8  5 */ always @(posedge clk) if (n1131) n1032 <= 1'b0 ? 1'b0 : n4737;
/* FF 29  5  5 */ always @(posedge clk) if (n3605) n3823 <= 1'b0 ? 1'b0 : n4738;
/* FF  4 10  2 */ always @(posedge clk) if (n251) n381 <= 1'b0 ? 1'b0 : n4739;
/* FF 24 16  2 */ always @(posedge clk) if (n3376) n3386 <= 1'b0 ? 1'b0 : n4740;
/* FF 27 22  5 */ always @(posedge clk) if (n3703) n3700 <= 1'b0 ? 1'b0 : n4741;
/* FF 13 10  3 */ always @(posedge clk) if (n850) n1437 <= 1'b0 ? 1'b0 : n4742;
/* FF  7 16  6 */ always @(posedge clk) if (n630) n747 <= 1'b0 ? 1'b0 : n4743;
/* FF  9 21  4 */ always @(posedge clk) if (n818) n918 <= 1'b0 ? 1'b0 : n4744;
/* FF 21 11  1 */ always @(posedge clk) if (n2085) n2416 <= 1'b0 ? 1'b0 : n4745;
/* FF 21  6  6 */ always @(posedge clk) if (n2247) n2839 <= 1'b0 ? 1'b0 : n4746;
/* FF 12 22  2 */ always @(posedge clk) if (n1357) n1350 <= 1'b0 ? 1'b0 : n4747;
/* FF 26 15  3 */ always @(posedge clk) if (n3233) n3543 <= 1'b0 ? 1'b0 : n4748;
/* FF 17  9  1 */ assign n1771 = n4749;
/* FF 19 23  0 */ assign \rco[181]  = n4750;
/* FF 10  9  4 */ always @(posedge clk) if (n983) n980 <= 1'b0 ? 1'b0 : n4751;
/* FF 28 20  6 */ assign n3424 = n4752;
/* FF 22 15  4 */ always @(posedge clk) if (n3216) n3062 <= 1'b0 ? 1'b0 : n4753;
/* FF  4 21  5 */ always @(posedge clk) if (n552) n120 <= 1'b0 ? 1'b0 : n4754;
/* FF 13 28  3 */ always @(posedge clk) if (n1394) n1564 <= 1'b0 ? 1'b0 : n4755;
/* FF 27 11  0 */ assign n3368 = n4756;
/* FF  6 10  4 */ always @(posedge clk) if (n589) n595 <= 1'b0 ? 1'b0 : n4757;
/* FF 20 11  5 */ always @(posedge clk) if (n2682) n2693 <= 1'b0 ? 1'b0 : n4758;
/* FF 23 19  4 */ always @(posedge clk) if (n2573) n3254 <= 1'b0 ? 1'b0 : n4759;
/* FF  5 13  7 */ always @(posedge clk) if (n402) n499 <= 1'b0 ? 1'b0 : n4760;
/* FF 19 24  6 */ always @(posedge clk) if (n2775) n2600 <= 1'b0 ? 1'b0 : n4761;
/* FF 11 20  0 */ always @(posedge clk) if (n1339) n1189 <= 1'b0 ? 1'b0 : n4762;
/* FF 29  9  6 */ always @(posedge clk) if (n3464) n3831 <= 1'b0 ? 1'b0 : n4763;
/* FF 17 27  5 */ always @(posedge clk) if (n1) n2193 <= 1'b0 ? 1'b0 : n4764;
/* FF 28 23  0 */ always @(posedge clk) if (n3704) n3807 <= 1'b0 ? 1'b0 : n4765;
/* FF 10 20  1 */ always @(posedge clk) if (n922) n1049 <= 1'b0 ? 1'b0 : n4766;
/* FF 15 16  7 */ always @(posedge clk) if (n1500) n1800 <= 1'b0 ? 1'b0 : n4767;
/* FF 21 15  6 */ assign n1340 = n4768;
/* FF 20 25  4 */ always @(posedge clk) if (n2612) n2802 <= 1'b0 ? 1'b0 : n4769;
/* FF 15 15  6 */ assign \rco[145]  = n1954;
/* FF  3 21  5 */ assign n4770 = n461;
/* FF 18 16  2 */ always @(posedge clk) if (n2540) n2316 <= 1'b0 ? 1'b0 : n4771;
/* FF  6  9  6 */ assign \rco[10]  = n4772;
/* FF 20 22  5 */ always @(posedge clk) if (n2384) n2781 <= 1'b0 ? 1'b0 : n4773;
/* FF 12 26  7 */ always @(posedge clk) if (n1393) n1392 <= 1'b0 ? 1'b0 : n4774;
/* FF 17 24  1 */ always @(posedge clk) if (n2000) n2167 <= 1'b0 ? 1'b0 : n4775;
/* FF  4  9  3 */ always @(posedge clk) if (n260) n374 <= 1'b0 ? 1'b0 : n4776;
/* FF 24 15  3 */ always @(posedge clk) if (n3233) n3378 <= 1'b0 ? 1'b0 : n4777;
/* FF 13 11  4 */ always @(posedge clk) if (n1137) n1445 <= 1'b0 ? 1'b0 : n4778;
/* FF  7 17  1 */ always @(posedge clk) if (n549) n752 <= 1'b0 ? 1'b0 : n4779;
/* FF 21 12  0 */ always @(posedge clk) if (n3029) n2867 <= 1'b0 ? 1'b0 : n4780;
/* FF 14 26  3 */ always @(posedge clk) if (n1271) n1714 <= 1'b0 ? 1'b0 : n4781;
/* FF 12 21  3 */ always @(posedge clk) if (n1205) n1342 <= 1'b0 ? 1'b0 : n4782;
/* FF 17 10  0 */ always @(posedge clk) if (n2282) n2059 <= 1'b0 ? 1'b0 : n4783;
/* FF 20  4  1 */ assign \rco[95]  = n4784;
/* FF 19 20  1 */ always @(posedge clk) if (n2553) n2566 <= 1'b0 ? 1'b0 : n4785;
/* FF 22 19  7 */ assign n809 = n4786;
/* FF 10  5  4 */ always @(posedge clk) if (en_in) n970 <= 1'b0 ? 1'b0 : n4787;
/* FF 24 18  7 */ always @(posedge clk) if (n3411) n3407 <= 1'b0 ? 1'b0 : n4788;
/* FF 22 14  3 */ always @(posedge clk) if (n3045) n3054 <= 1'b0 ? 1'b0 : n4789;
/* FF 27  8  1 */ assign n3605 = n4790;
/* FF  3 17  2 */ always @(posedge clk) if (n79) n312 <= 1'b0 ? 1'b0 : n4791;
/* FF 14 25  7 */ always @(posedge clk) if (n697) n1708 <= 1'b0 ? 1'b0 : n4792;
/* FF  6 21  5 */ assign n672 = n4793;
/* FF 17  4  3 */ always @(posedge clk) if (n1761) n2033 <= 1'b0 ? 1'b0 : n4794;
/* FF 23 16  5 */ assign \rco[100]  = n4795;
/* FF 11 14  6 */ always @(posedge clk) if (n1154) n1152 <= 1'b0 ? 1'b0 : n4796;
/* FF 20  7  5 */ always @(posedge clk) if (n2670) n2666 <= 1'b0 ? 1'b0 : n4797;
/* FF  5 14  6 */ always @(posedge clk) if (n402) n509 <= 1'b0 ? 1'b0 : n4798;
/* FF 20 10  6 */ always @(posedge clk) if (n2697) n2688 <= 1'b0 ? 1'b0 : n4799;
/* FF 11 21  7 */ always @(posedge clk) if (n819) n1203 <= 1'b0 ? 1'b0 : n4800;
/* FF 28 22  3 */ always @(posedge clk) if (n3704) n3802 <= 1'b0 ? 1'b0 : n4801;
/* FF 16 12  2 */ always @(posedge clk) if (n1771) n1937 <= 1'b0 ? 1'b0 : n4802;
/* FF 16 17  5 */ always @(posedge clk) if (n2110) n1968 <= 1'b0 ? 1'b0 : n4803;
/* FF 10 23  0 */ assign n796 = n4804;
/* FF 13 15  1 */ always @(posedge clk) if (n739) n1471 <= 1'b0 ? 1'b0 : n4805;
/* FF 27  6  0 */ assign n3593 = n3718;
/* FF 30 12  1 */ always @(posedge clk) if (n3892) n3895 <= 1'b0 ? 1'b0 : n4806;
/* FF 15 17  0 */ always @(posedge clk) if (n1500) n1801 <= 1'b0 ? 1'b0 : n4807;
/* FF 18  6  4 */ always @(posedge clk) if (n2241) n2235 <= 1'b0 ? 1'b0 : n4808;
/* FF  7 21  6 */ always @(posedge clk) if (n360) n774 <= 1'b0 ? 1'b0 : n4809;
/* FF  6  7  4 */ always @(posedge clk) if (n570) n575 <= 1'b0 ? 1'b0 : n4810;
/* FF 18 19  3 */ always @(posedge clk) if (n1982) n2342 <= 1'b0 ? 1'b0 : n4811;
/* FF  3 18  4 */ always @(posedge clk) if (n215) n322 <= 1'b0 ? 1'b0 : n4812;
/* FF 20 24  3 */ always @(posedge clk) if (n2775) n2791 <= 1'b0 ? 1'b0 : n4813;
/* FF 20 21  4 */ always @(posedge clk) if (n2553) n2772 <= 1'b0 ? 1'b0 : n4814;
/* FF 12 25  6 */ always @(posedge clk) if (n1532) n1382 <= 1'b0 ? 1'b0 : n4815;
/* FF  1 19  2 */ always @(posedge clk) if (n119) n106 <= 1'b0 ? 1'b0 : n4816;
/* FF 17 25  2 */ always @(posedge clk) if (n2017) n2178 <= 1'b0 ? 1'b0 : n4817;
/* FF 23 13  0 */ always @(posedge clk) if (n3045) n3208 <= 1'b0 ? 1'b0 : n4818;
/* FF 10 25  3 */ always @(posedge clk) if (n567) n1083 <= 1'b0 ? 1'b0 : n4819;
/* FF 24 14  0 */ always @(posedge clk) if (n3376) n3369 <= 1'b0 ? 1'b0 : n4820;
/* FF 27 20  7 */ always @(posedge clk) if (n3424) n3682 <= 1'b0 ? 1'b0 : n4821;
/* FF  4 19  6 */ assign n349 = n4822;
/* FF 13 12  5 */ always @(posedge clk) if (n1137) n1454 <= 1'b0 ? 1'b0 : n4823;
/* FF 18  5  6 */ always @(posedge clk) if (n2230) n2227 <= 1'b0 ? 1'b0 : n4824;
/* FF  7 22  0 */ always @(posedge clk) if (n695) n783 <= 1'b0 ? 1'b0 : n4825;
/* FF  9 23  2 */ always @(posedge clk) if (n819) n927 <= 1'b0 ? 1'b0 : n4826;
/* FF 21 13  3 */ always @(posedge clk) if (n2519) n2877 <= 1'b0 ? 1'b0 : n4827;
/* FF 14 21  2 */ assign n1355 = n4828;
/* FF 19 30  7 */ always @(posedge clk) if (n2592) n2640 <= 1'b0 ? 1'b0 : n4829;
/* FF  1 16  4 */ always @(posedge clk) if (n85) n92 <= 1'b0 ? 1'b0 : n4830;
/* FF 19 21  6 */ always @(posedge clk) if (n2164) n2582 <= 1'b0 ? 1'b0 : n4831;
/* FF 11 17  4 */ always @(posedge clk) if (n900) n1172 <= 1'b0 ? 1'b0 : n4832;
/* FF 10 11  6 */ always @(posedge clk) if (n996) n994 <= 1'b0 ? 1'b0 : n4833;
/* FF 16  8  7 */ always @(posedge clk) if (n1625) n1922 <= 1'b0 ? 1'b0 : n4834;
/* FF 24 17  6 */ always @(posedge clk) if (n2123) n3400 <= 1'b0 ? 1'b0 : n4835;
/* FF 28  7  7 */ always @(posedge clk) if (n3488) n3725 <= 1'b0 ? 1'b0 : n4836;
/* FF 22  9  2 */ always @(posedge clk) if (n2989) n3016 <= 1'b0 ? 1'b0 : n4837;
/* FF 15 21  5 */ always @(posedge clk) if (n1356) n1841 <= 1'b0 ? 1'b0 : n4838;
/* FF 14 24  4 */ assign n1698 = n4839;
/* FF 17  5  0 */ assign \rco[141]  = n4840;
/* FF  6 20  6 */ always @(posedge clk) if (n552) n666 <= 1'b0 ? 1'b0 : n4841;
/* FF 23 17  2 */ always @(posedge clk) if (n2540) n3234 <= 1'b0 ? 1'b0 : n4842;
/* FF 11 15  5 */ always @(posedge clk) if (n733) n1156 <= 1'b0 ? 1'b0 : n4843;
/* FF 26  6  6 */ always @(posedge clk) if (n3459) n3479 <= 1'b0 ? 1'b0 : n4844;
/* FF 11 18  6 */ always @(posedge clk) if (n1187) n1185 <= 1'b0 ? 1'b0 : n4845;
/* FF 29 11  0 */ always @(posedge clk) if (n3751) n3839 <= 1'b0 ? 1'b0 : n4846;
/* FF 28 21  2 */ always @(posedge clk) if (n3788) n3793 <= 1'b0 ? 1'b0 : n4847;
/* FF  4 12  1 */ always @(posedge clk) if (n77) n394 <= 1'b0 ? 1'b0 : n4848;
/* FF 13 16  0 */ always @(posedge clk) if (n922) n1477 <= 1'b0 ? 1'b0 : n4849;
/* FF 27  7  3 */ always @(posedge clk) if (n3459) n3598 <= 1'b0 ? 1'b0 : n4850;
/* FF 15 22  1 */ always @(posedge clk) if (n1835) n1847 <= 1'b0 ? 1'b0 : n4851;
/* FF 18  9  5 */ always @(posedge clk) if (n2055) n2266 <= 1'b0 ? 1'b0 : n4852;
/* FF  9 19  7 */ always @(posedge clk) if (n454) n908 <= 1'b0 ? 1'b0 : n4853;
/* FF  3 19  7 */ always @(posedge clk) if (n115) n334 <= 1'b0 ? 1'b0 : n4854;
/* FF  6 11  4 */ always @(posedge clk) if (n286) n603 <= 1'b0 ? 1'b0 : n4855;
/* FF 12 24  1 */ always @(posedge clk) if (n961) n1368 <= 1'b0 ? 1'b0 : n4856;
/* FF 26  5  0 */ always @(posedge clk) if (n3459) n3472 <= 1'b0 ? 1'b0 : n4857;
/* FF 14 10  0 */ always @(posedge clk) if (n1622) n1604 <= 1'b0 ? 1'b0 : n4858;
/* FF 19 17  3 */ always @(posedge clk) if (n2727) n2544 <= 1'b0 ? 1'b0 : n4859;
/* FF 22 21  4 */ always @(posedge clk) if (n2564) n3100 <= 1'b0 ? 1'b0 : n4860;
/* FF 24 24  6 */ always @(posedge clk) if (n3112) n3444 <= 1'b0 ? 1'b0 : n4861;
/* FF  4 15  5 */ always @(posedge clk) if (n207) n417 <= 1'b0 ? 1'b0 : n4862;
/* FF 10 24  0 */ always @(posedge clk) if (n820) n1072 <= 1'b0 ? 1'b0 : n4863;
/* FF 24 13  1 */ always @(posedge clk) if (n3351) n3362 <= 1'b0 ? 1'b0 : n4864;
/* FF 27 21  0 */ always @(posedge clk) if (n3421) n3687 <= 1'b0 ? 1'b0 : n4865;
/* FF  4 18  5 */ always @(posedge clk) if (n349) n435 <= 1'b0 ? 1'b0 : n4866;
/* FF 18  4  5 */ always @(posedge clk) if (n2207) n2218 <= 1'b0 ? 1'b0 : n4867;
/* FF 21 14  2 */ always @(posedge clk) if (n2519) n2884 <= 1'b0 ? 1'b0 : n4868;
/* FF  9 16  3 */ always @(posedge clk) if (n645) n878 <= 1'b0 ? 1'b0 : n4869;
/* FF 14 20  1 */ always @(posedge clk) if (n1347) n1677 <= 1'b0 ? 1'b0 : n4870;
/* FF  5  8  7 */ always @(posedge clk) if (n21) n473 <= 1'b0 ? 1'b0 : n4871;
/* FF 19 31  4 */ always @(posedge clk) if (n2592) n2645 <= 1'b0 ? 1'b0 : n4872;
/* FF  2 11  3 */ always @(posedge clk) if (n168) n171 <= 1'b0 ? 1'b0 : n4873;
/* FF 23 21  7 */ always @(posedge clk) if (n3258) n3278 <= 1'b0 ? 1'b0 : n4874;
/* FF 19 18  7 */ always @(posedge clk) if (n2348) n2561 <= 1'b0 ? 1'b0 : n4875;
/* FF 10 10  1 */ always @(posedge clk) if (n983) n984 <= 1'b0 ? 1'b0 : n4876;
/* FF 16 23  6 */ always @(posedge clk) if (n2000) n1996 <= 1'b0 ? 1'b0 : n4877;
/* FF 28  6  4 */ always @(posedge clk) if (n3594) n3715 <= 1'b0 ? 1'b0 : n4878;
/* FF 21 16  1 */ always @(posedge clk) if (n2551) n2888 <= 1'b0 ? 1'b0 : n4879;
/* FF 15 10  4 */ always @(posedge clk) if (n1624) n1758 <= 1'b0 ? 1'b0 : n4880;
/* FF 18 22  1 */ always @(posedge clk) if (n2164) n2357 <= 1'b0 ? 1'b0 : n4881;
/* FF 17  6  1 */ always @(posedge clk) if (n2045) n2039 <= 1'b0 ? 1'b0 : n4882;
/* FF  6 23  7 */ always @(posedge clk) if (n360) n694 <= 1'b0 ? 1'b0 : n4883;
/* FF 20  8  0 */ assign n2451 = n4884;
/* FF 12 28  6 */ always @(posedge clk) if (n1394) n1400 <= 1'b0 ? 1'b0 : n4885;
/* FF 23 22  3 */ always @(posedge clk) if (n3422) n3282 <= 1'b0 ? 1'b0 : n4886;
/* FF 11 19  5 */ assign n121 = n1335;
/* FF 29 12  1 */ always @(posedge clk) if (n3751) n3850 <= 1'b0 ? 1'b0 : n4887;
/* FF 16 10  0 */ always @(posedge clk) if (n1771) n1926 <= 1'b0 ? 1'b0 : n4888;
/* FF 22 26  2 */ always @(posedge clk) if (n2613) n3135 <= 1'b0 ? 1'b0 : n4889;
/* FF 27 17  5 */ always @(posedge clk) if (n3249) n3654 <= 1'b0 ? 1'b0 : n4890;
/* FF  9  7  4 */ always @(posedge clk) if (n588) n579 <= 1'b0 ? 1'b0 : n4891;
/* FF 13 17  3 */ always @(posedge clk) if (n1461) n1487 <= 1'b0 ? 1'b0 : n4892;
/* FF 15 23  2 */ always @(posedge clk) if (n778) n1854 <= 1'b0 ? 1'b0 : n4893;
/* FF 18  8  6 */ always @(posedge clk) if (n2055) n2255 <= 1'b0 ? 1'b0 : n4894;
/* FF 18 21  5 */ always @(posedge clk) if (n2347) n2354 <= 1'b0 ? 1'b0 : n4895;
/* FF  3 16  6 */ always @(posedge clk) if (n197) n308 <= 1'b0 ? 1'b0 : n4896;
/* FF 14  5  1 */ always @(posedge clk) if (n1577) n1572 <= 1'b0 ? 1'b0 : n4897;
/* FF 19 14  2 */ always @(posedge clk) if (n2123) n2513 <= 1'b0 ? 1'b0 : n4898;
/* FF 22 20  7 */ always @(posedge clk) if (n3087) n3095 <= 1'b0 ? 1'b0 : n4899;
/* FF 10 14  6 */ always @(posedge clk) if (n750) n1013 <= 1'b0 ? 1'b0 : n4900;
/* FF  4 14  6 */ always @(posedge clk) if (n79) n408 <= 1'b0 ? 1'b0 : n4901;
/* FF 22 25  4 */ always @(posedge clk) if (n2812) n3129 <= 1'b0 ? 1'b0 : n4902;
/* FF 10 27  1 */ always @(posedge clk) if (n804) n1094 <= 1'b0 ? 1'b0 : n4903;
/* FF 24 12  6 */ always @(posedge clk) if (n3351) n3359 <= 1'b0 ? 1'b0 : n4904;
/* FF 16 24  4 */ assign n2000 = n4905;
/* FF 27 18  1 */ always @(posedge clk) if (n3553) n3658 <= 1'b0 ? 1'b0 : n4906;
/* FF 28 10  1 */ always @(posedge clk) if (n3462) n3742 <= 1'b0 ? 1'b0 : n4907;
/* FF  4 17  4 */ always @(posedge clk) if (n2) n428 <= 1'b0 ? 1'b0 : n4908;
/* FF 13 14  7 */ always @(posedge clk) if (n1461) n1469 <= 1'b0 ? 1'b0 : n4909;
/* FF 18  7  4 */ always @(posedge clk) if (n1761) n2243 <= 1'b0 ? 1'b0 : n4910;
/* FF  9 17  0 */ always @(posedge clk) if (n1030) n883 <= 1'b0 ? 1'b0 : n4911;
/* FF 26 22  0 */ always @(posedge clk) if (n2730) n3569 <= 1'b0 ? 1'b0 : n4912;
/* FF 15  5  2 */ always @(posedge clk) if (n1742) n1727 <= 1'b0 ? 1'b0 : n4913;
/* FF 14 23  0 */ assign n778 = n4914;
/* FF 20 12  5 */ always @(posedge clk) if (n2682) n2703 <= 1'b0 ? 1'b0 : n4915;
/* FF 19 28  5 */ always @(posedge clk) if (n2614) n2626 <= 1'b0 ? 1'b0 : n4916;
/* FF 19 19  4 */ assign n2348 = n4917;
/* FF 10 13  0 */ assign n733 = n4918;
/* FF 28  5  5 */ always @(posedge clk) if (n3488) n3710 <= 1'b0 ? 1'b0 : n4919;
/* FF 22 11  0 */ assign \rco[57]  = n4920;
/* FF 21 17  2 */ assign \rco[62]  = n4921;
/* FF 30 10  4 */ always @(posedge clk) if (n3892) n3889 <= 1'b0 ? 1'b0 : n4922;
/* FF 15 11  7 */ always @(posedge clk) if (n1624) n1770 <= 1'b0 ? 1'b0 : n4923;
/* FF  2 19  4 */ assign n4924 = n341;
/* FF 18 25  0 */ always @(posedge clk) if (n1878) n2377 <= 1'b0 ? 1'b0 : n4925;
/* FF 15  6  4 */ always @(posedge clk) if (n1744) n1737 <= 1'b0 ? 1'b0 : n4926;
/* FF 17  7  6 */ always @(posedge clk) if (n2045) n2052 <= 1'b0 ? 1'b0 : n4927;
/* FF  6 22  0 */ always @(posedge clk) if (n673) n678 <= 1'b0 ? 1'b0 : n4928;
/* FF 20 15  1 */ always @(posedge clk) if (n2715) n2718 <= 1'b0 ? 1'b0 : n4929;
/* FF 23 23  0 */ always @(posedge clk) if (n3104) n3287 <= 1'b0 ? 1'b0 : n4930;
/* FF 11 13  3 */ always @(posedge clk) if (n733) n1141 <= 1'b0 ? 1'b0 : n4931;
/* FF 11 16  4 */ always @(posedge clk) if (n891) n1163 <= 1'b0 ? 1'b0 : n4932;
/* FF 16  9  1 */ always @(posedge clk) if (n1771) n1924 <= 1'b0 ? 1'b0 : n4933;
/* FF 13  7  5 */ always @(posedge clk) if (n977) n1428 <= 1'b0 ? 1'b0 : n4934;
/* FF 13 18  2 */ always @(posedge clk) if (n1205) n1494 <= 1'b0 ? 1'b0 : n4935;
/* FF 27  5  5 */ always @(posedge clk) if (n3594) n3590 <= 1'b0 ? 1'b0 : n4936;
/* FF 18 11  7 */ assign n2282 = n4937;
/* FF 15 20  3 */ always @(posedge clk) if (n1347) n1830 <= 1'b0 ? 1'b0 : n4938;
/* FF 18 20  6 */ assign n1982 = n4939;
/* FF 26  7  2 */ always @(posedge clk) if (n3603) n3483 <= 1'b0 ? 1'b0 : n4940;
/* FF  2 14  1 */ always @(posedge clk) if (n83) n188 <= 1'b0 ? 1'b0 : n4941;
/* FF 16  7  0 */ always @(posedge clk) if (n1743) n1907 <= 1'b0 ? 1'b0 : n4942;
/* FF 19 15  1 */ always @(posedge clk) if (n2715) n2526 <= 1'b0 ? 1'b0 : n4943;
/* FF 23  5  4 */ always @(posedge clk) if (n3158) n3154 <= 1'b0 ? 1'b0 : n4944;
/* FF 22 23  6 */ assign n2961 = n4945;
/* FF 24 22  4 */ always @(posedge clk) if (n3422) n3429 <= 1'b0 ? 1'b0 : n4946;
/* FF  4 13  7 */ always @(posedge clk) if (n78) n194 <= 1'b0 ? 1'b0 : n4947;
/* FF 22 24  7 */ always @(posedge clk) if (n3113) n3123 <= 1'b0 ? 1'b0 : n4948;
/* FF 10 26  6 */ assign n954 = n4949;
/* FF 24 11  7 */ assign n3352 = n4950;
/* FF 27 19  2 */ always @(posedge clk) if (n3553) n3669 <= 1'b0 ? 1'b0 : n4951;
/* FF 28  9  0 */ always @(posedge clk) if (n3621) n3734 <= 1'b0 ? 1'b0 : n4952;
/* FF  4 16  3 */ always @(posedge clk) if (n79) n423 <= 1'b0 ? 1'b0 : n4953;
/* FF  9 18  1 */ always @(posedge clk) if (n1030) n893 <= 1'b0 ? 1'b0 : n4954;
/* FF 26  9  1 */ always @(posedge clk) if (n3460) n3499 <= 1'b0 ? 1'b0 : n4955;
/* FF 29 17  0 */ always @(posedge clk) if (n3765) n3856 <= 1'b0 ? 1'b0 : n4956;
/* FF 14 22  7 */ always @(posedge clk) if (n1402) n1694 <= 1'b0 ? 1'b0 : n4957;
/* FF 17  3  3 */ always @(posedge clk) if (n1887) n2028 <= 1'b0 ? 1'b0 : n4958;
/* FF  6 18  5 */ always @(posedge clk) if (n657) n654 <= 1'b0 ? 1'b0 : n4959;
/* FF  5 10  5 */ always @(posedge clk) if (n184) n479 <= 1'b0 ? 1'b0 : n4960;
/* FF 19 29  2 */ assign \rco[196]  = n4961;
/* FF 23 27  5 */ always @(posedge clk) if (n2017) n3316 <= 1'b0 ? 1'b0 : n4962;
/* FF 19 16  5 */ assign n2520 = n4963;
/* FF 23  6  6 */ always @(posedge clk) if (n3158) n3165 <= 1'b0 ? 1'b0 : n4964;
/* FF 11 28  7 */ always @(posedge clk) if (n1384) n1262 <= 1'b0 ? 1'b0 : n4965;
/* FF 10 12  3 */ always @(posedge clk) if (n996) n1000 <= 1'b0 ? 1'b0 : n4966;
/* FF 24 25  2 */ always @(posedge clk) if (n2812) n3448 <= 1'b0 ? 1'b0 : n4967;
/* FF 16 21  4 */ always @(posedge clk) if (n1835) n1985 <= 1'b0 ? 1'b0 : n4968;
/* FF 16 26  5 */ always @(posedge clk) if (n1557) n2015 <= 1'b0 ? 1'b0 : n4969;
/* FF 21 18  3 */ always @(posedge clk) if (n2757) n2905 <= 1'b0 ? 1'b0 : n4970;
/* FF  9 28  0 */ always @(posedge clk) if (n961) n956 <= 1'b0 ? 1'b0 : n4971;
/* FF 15  8  6 */ always @(posedge clk) if (n1741) n1751 <= 1'b0 ? 1'b0 : n4972;
/* FF  3 22  7 */ always @(posedge clk) if (n352) n359 <= 1'b0 ? 1'b0 : n4973;
/* FF  2 18  3 */ always @(posedge clk) if (n115) n212 <= 1'b0 ? 1'b0 : n4974;
/* FF 21  7  7 */ assign \rco[47]  = n4975;
/* FF 15  7  7 */ assign n1741 = n4976;
/* FF 18 24  3 */ always @(posedge clk) if (n1878) n2373 <= 1'b0 ? 1'b0 : n4977;
/* FF  6 17  1 */ always @(posedge clk) if (n549) n647 <= 1'b0 ? 1'b0 : n4978;
/* FF 20 14  2 */ always @(posedge clk) if (n2682) n2714 <= 1'b0 ? 1'b0 : n4979;
/* FF 23 20  1 */ always @(posedge clk) if (n3258) n3264 <= 1'b0 ? 1'b0 : n4980;
/* FF 24  7  2 */ assign n4981 = n3458;
/* FF  9 14  7 */ always @(posedge clk) if (n629) n866 <= 1'b0 ? 1'b0 : n4982;
/* FF 13 19  5 */ assign n1461 = n4983;
/* FF 18 10  0 */ always @(posedge clk) if (n2282) n2273 <= 1'b0 ? 1'b0 : n4984;
/* FF 18 23  7 */ always @(posedge clk) if (n1999) n2368 <= 1'b0 ? 1'b0 : n4985;
/* FF 12 29  2 */ always @(posedge clk) if (n1532) n1405 <= 1'b0 ? 1'b0 : n4986;
/* FF 19 25  7 */ always @(posedge clk) if (n2612) n2611 <= 1'b0 ? 1'b0 : n4987;
/* FF 14  7  3 */ always @(posedge clk) if (n1743) n1588 <= 1'b0 ? 1'b0 : n4988;
/* FF 16  6  3 */ always @(posedge clk) if (n1744) n1900 <= 1'b0 ? 1'b0 : n4989;
/* FF 19 12  0 */ always @(posedge clk) if (n1936) n2497 <= 1'b0 ? 1'b0 : n4990;
/* FF 23 10  5 */ always @(posedge clk) if (n2697) n3188 <= 1'b0 ? 1'b0 : n4991;
/* FF 22 22  1 */ always @(posedge clk) if (n2961) n3106 <= 1'b0 ? 1'b0 : n4992;
/* FF 24 21  5 */ always @(posedge clk) if (n3411) n3413 <= 1'b0 ? 1'b0 : n4993;
/* FF 22 27  6 */ always @(posedge clk) if (n2970) n3149 <= 1'b0 ? 1'b0 : n4994;
/* FF 24 10  4 */ always @(posedge clk) if (n3352) n3344 <= 1'b0 ? 1'b0 : n4995;
/* FF 28  8  7 */ always @(posedge clk) if (n3605) n3732 <= 1'b0 ? 1'b0 : n4996;
/* FF 13  5  2 */ always @(posedge clk) if (n1577) n1412 <= 1'b0 ? 1'b0 : n4997;
/* FF  3  9  0 */ always @(posedge clk) if (n260) n252 <= 1'b0 ? 1'b0 : n4998;
/* FF 12 19  1 */ always @(posedge clk) if (n1501) n1329 <= 1'b0 ? 1'b0 : n4999;
/* FF 26  8  2 */ always @(posedge clk) if (n3603) n3492 <= 1'b0 ? 1'b0 : n5000;
/* FF 14 17  6 */ always @(posedge clk) if (n1672) n1660 <= 1'b0 ? 1'b0 : n5001;
/* FF 17 12  2 */ always @(posedge clk) if (n2056) n2079 <= 1'b0 ? 1'b0 : n5002;
/* FF 19 26  3 */ assign \rco[172]  = n2813;
/* FF 23 24  4 */ always @(posedge clk) if (n3112) n3300 <= 1'b0 ? 1'b0 : n5003;
/* FF  2 12  6 */ always @(posedge clk) if (n39) n182 <= 1'b0 ? 1'b0 : n5004;
/* FF 23  7  5 */ always @(posedge clk) if (n3006) n3171 <= 1'b0 ? 1'b0 : n5005;
/* FF 10 15  2 */ always @(posedge clk) if (n750) n1017 <= 1'b0 ? 1'b0 : n5006;
/* FF 16 20  3 */ always @(posedge clk) if (n1843) n1977 <= 1'b0 ? 1'b0 : n5007;
/* FF 16 25  4 */ always @(posedge clk) if (n1557) n2007 <= 1'b0 ? 1'b0 : n5008;
/* FF 21 24  5 */ always @(posedge clk) if (n3113) n2958 <= 1'b0 ? 1'b0 : n5009;
/* FF 21 19  4 */ always @(posedge clk) if (n2757) n2914 <= 1'b0 ? 1'b0 : n5010;
/* FF 13 23  2 */ always @(posedge clk) if (n1069) n1526 <= 1'b0 ? 1'b0 : n5011;
/* FF 27 14  3 */ always @(posedge clk) if (n3527) n3644 <= 1'b0 ? 1'b0 : n5012;
/* FF 18 14  5 */ always @(posedge clk) if (n2045) n2248 <= 1'b0 ? 1'b0 : n5013;
/* FF  2 21  2 */ always @(posedge clk) if (n126) n229 <= 1'b0 ? 1'b0 : n5014;
/* FF 18 27  2 */ always @(posedge clk) if (n2020) n2395 <= 1'b0 ? 1'b0 : n5015;
/* FF  6 16  2 */ always @(posedge clk) if (n511) n640 <= 1'b0 ? 1'b0 : n5016;
/* FF 20 13  3 */ assign n2307 = n5017;
/* FF  4 11  4 */ always @(posedge clk) if (n184) n389 <= 1'b0 ? 1'b0 : n5018;
/* FF 22 18  6 */ always @(posedge clk) if (n3065) n3085 <= 1'b0 ? 1'b0 : n5019;
/* FF 22  7  1 */ always @(posedge clk) if (n2841) n2999 <= 1'b0 ? 1'b0 : n5020;
/* FF 10 17  2 */ assign n5021 = n1176;
/* FF  9 15  0 */ always @(posedge clk) if (n645) n867 <= 1'b0 ? 1'b0 : n5022;
/* FF 24  6  1 */ always @(posedge clk) if (n3006) n3322 <= 1'b0 ? 1'b0 : n5023;
/* FF 28 12  4 */ always @(posedge clk) if (n3462) n3757 <= 1'b0 ? 1'b0 : n5024;
/* FF 13 20  4 */ always @(posedge clk) if (n1339) n1507 <= 1'b0 ? 1'b0 : n5025;
/* FF 18 13  1 */ always @(posedge clk) if (n2283) n2296 <= 1'b0 ? 1'b0 : n5026;
/* FF 14 13  5 */ always @(posedge clk) if (n1015) n1628 <= 1'b0 ? 1'b0 : n5027;
/* FF 14  6  4 */ always @(posedge clk) if (n1577) n1579 <= 1'b0 ? 1'b0 : n5028;
/* FF 16  5  2 */ always @(posedge clk) if (n1742) n1890 <= 1'b0 ? 1'b0 : n5029;
/* FF 17 19  0 */ always @(posedge clk) if (n1982) n2128 <= 1'b0 ? 1'b0 : n5030;
/* FF 23 11  6 */ always @(posedge clk) if (n3031) n3196 <= 1'b0 ? 1'b0 : n5031;
/* FF 11 25  5 */ always @(posedge clk) if (n954) n955 <= 1'b0 ? 1'b0 : n5032;
/* FF 22 17  0 */ always @(posedge clk) if (n3065) n3072 <= 1'b0 ? 1'b0 : n5033;
/* FF 24 20  2 */ always @(posedge clk) if (n3411) n3412 <= 1'b0 ? 1'b0 : n5034;
/* FF 10 28  4 */ always @(posedge clk) if (n821) n1105 <= 1'b0 ? 1'b0 : n5035;
/* FF 24  9  5 */ always @(posedge clk) if (n3352) n3337 <= 1'b0 ? 1'b0 : n5036;
/* FF 13  6  3 */ always @(posedge clk) if (n977) n1418 <= 1'b0 ? 1'b0 : n5037;
/* FF  4 22  1 */ assign n462 = n564;
/* FF 21 23  1 */ always @(posedge clk) if (n2961) n2944 <= 1'b0 ? 1'b0 : n5038;
/* FF 15 13  6 */ always @(posedge clk) if (n1015) n1782 <= 1'b0 ? 1'b0 : n5039;
/* FF 12 18  2 */ always @(posedge clk) if (n1501) n1322 <= 1'b0 ? 1'b0 : n5040;
/* FF 26 11  3 */ always @(posedge clk) if (n3033) n3511 <= 1'b0 ? 1'b0 : n5041;
/* FF 29 19  6 */ always @(posedge clk) if (n3786) n3866 <= 1'b0 ? 1'b0 : n5042;
/* FF 14 16  5 */ always @(posedge clk) if (n1792) n1651 <= 1'b0 ? 1'b0 : n5043;
/* FF 17 13  1 */ always @(posedge clk) if (n2056) n2087 <= 1'b0 ? 1'b0 : n5044;
/* FF  5 12  3 */ always @(posedge clk) if (n77) n487 <= 1'b0 ? 1'b0 : n5045;
/* FF 19 27  0 */ always @(posedge clk) if (n2614) n2616 <= 1'b0 ? 1'b0 : n5046;
/* FF 23 25  3 */ always @(posedge clk) if (n2613) n3305 <= 1'b0 ? 1'b0 : n5047;
/* FF 11 26  1 */ always @(posedge clk) if (n954) n1237 <= 1'b0 ? 1'b0 : n5048;
/* FF  7  2  5 */ assign \rco[164]  = n5049;
/* FF  9 11  5 */ always @(posedge clk) if (n988) n847 <= 1'b0 ? 1'b0 : n5050;
/* FF 21 25  6 */ always @(posedge clk) if (n2970) n2968 <= 1'b0 ? 1'b0 : n5051;
/* FF  7  9  4 */ always @(posedge clk) if (n589) n722 <= 1'b0 ? 1'b0 : n5052;
/* FF 21 20  5 */ always @(posedge clk) if (n3087) n2923 <= 1'b0 ? 1'b0 : n5053;
/* FF 13 24  3 */ assign \rco[116]  = n5054;
/* FF 15 14  0 */ always @(posedge clk) if (n1791) n1783 <= 1'b0 ? 1'b0 : n5055;
/* FF  3 20  5 */ always @(posedge clk) if (n119) n122 <= 1'b0 ? 1'b0 : n5056;
/* FF  2 20  1 */ always @(posedge clk) if (n126) n218 <= 1'b0 ? 1'b0 : n5057;
/* FF 18 17  4 */ always @(posedge clk) if (n1825) n2329 <= 1'b0 ? 1'b0 : n5058;
/* FF 18 26  5 */ always @(posedge clk) if (n2615) n2390 <= 1'b0 ? 1'b0 : n5059;
/* FF  6 19  3 */ assign n5060 = n766;
/* FF 11  8  0 */ always @(posedge clk) if (n1131) n1123 <= 1'b0 ? 1'b0 : n5061;
/* FF 28 19  0 */ always @(posedge clk) if (n3424) n3777 <= 1'b0 ? 1'b0 : n5062;
/* FF 19  9  4 */ always @(posedge clk) if (n2451) n2475 <= 1'b0 ? 1'b0 : n5063;
/* FF  4 10  7 */ always @(posedge clk) if (n251) n386 <= 1'b0 ? 1'b0 : n5064;
/* FF 24 16  7 */ always @(posedge clk) if (n3376) n3383 <= 1'b0 ? 1'b0 : n5065;
/* FF 22  6  6 */ always @(posedge clk) if (n2841) n2996 <= 1'b0 ? 1'b0 : n5066;
/* FF 10 16  1 */ always @(posedge clk) if (n891) n1024 <= 1'b0 ? 1'b0 : n5067;
/* FF 13 10  6 */ always @(posedge clk) if (n850) n1439 <= 1'b0 ? 1'b0 : n5068;
/* FF 13 21  7 */ always @(posedge clk) if (n1356) n1519 <= 1'b0 ? 1'b0 : n5069;
/* FF 31 22  7 */ assign \rco[190]  = n5070;
/* FF 18 12  2 */ always @(posedge clk) if (n1936) n2288 <= 1'b0 ? 1'b0 : n5071;
/* FF 21  6  1 */ always @(posedge clk) if (n2247) n2834 <= 1'b0 ? 1'b0 : n5072;
/* FF 11  6  3 */ always @(posedge clk) if (en_in) n1121 <= 1'b0 ? 1'b0 : n5073;
/* FF 14 12  6 */ assign n1623 = n5074;
/* FF 19 23  5 */ assign n5075 = n2787;
/* FF 19 10  6 */ always @(posedge clk) if (n2678) n2484 <= 1'b0 ? 1'b0 : n5076;
/* FF  4 21  0 */ always @(posedge clk) if (n552) n447 <= 1'b0 ? 1'b0 : n5077;
/* FF  7 13  1 */ assign \rco[154]  = n5078;
/* FF 21  8  0 */ always @(posedge clk) if (n2989) n2842 <= 1'b0 ? 1'b0 : n5079;
/* FF 26 17  5 */ always @(posedge clk) if (n3249) n3551 <= 1'b0 ? 1'b0 : n5080;
/* FF 12 17  3 */ always @(posedge clk) if (n900) n1315 <= 1'b0 ? 1'b0 : n5081;
/* FF 26 10  4 */ always @(posedge clk) if (n3033) n3509 <= 1'b0 ? 1'b0 : n5082;
/* FF 18 30  2 */ always @(posedge clk) if (n1881) n2419 <= 1'b0 ? 1'b0 : n5083;
/* FF 14 19  4 */ always @(posedge clk) if (n1672) n1668 <= 1'b0 ? 1'b0 : n5084;
/* FF 17 14  0 */ assign n2094 = n5085;
/* FF 29 20  7 */ always @(posedge clk) if (n3786) n3875 <= 1'b0 ? 1'b0 : n5086;
/* FF  5 13  0 */ always @(posedge clk) if (n402) n492 <= 1'b0 ? 1'b0 : n5087;
/* FF 19 24  1 */ always @(posedge clk) if (n2775) n2595 <= 1'b0 ? 1'b0 : n5088;
/* FF 11 27  2 */ always @(posedge clk) if (n1393) n1249 <= 1'b0 ? 1'b0 : n5089;
/* FF 16 18  1 */ always @(posedge clk) if (n1205) n1341 <= 1'b0 ? 1'b0 : n5090;
/* FF  1 11  0 */ assign n37 = n5091;
/* FF 21 26  7 */ assign n2037 = n5092;
/* FF 21 21  6 */ always @(posedge clk) if (n2564) n2932 <= 1'b0 ? 1'b0 : n5093;
/* FF 13 25  0 */ assign \rco[199]  = n5094;
/* FF 27 12  1 */ always @(posedge clk) if (n3368) n3630 <= 1'b0 ? 1'b0 : n5095;
/* FF 15 15  3 */ assign n1792 = n5096;
/* FF  3 21  2 */ assign n5097 = n459;
/* FF 18 16  7 */ always @(posedge clk) if (n2540) n2321 <= 1'b0 ? 1'b0 : n5098;
/* FF 18 29  4 */ always @(posedge clk) if (n1881) n2412 <= 1'b0 ? 1'b0 : n5099;
/* FF 28 18  3 */ always @(posedge clk) if (n3765) n3776 <= 1'b0 ? 1'b0 : n5100;
/* FF 19  6  5 */ always @(posedge clk) if (n2241) n2448 <= 1'b0 ? 1'b0 : n5101;
/* FF  4  9  6 */ always @(posedge clk) if (n260) n377 <= 1'b0 ? 1'b0 : n5102;
/* FF 22 28  4 */ assign \rco[121]  = n5103;
/* FF 10  6  7 */ always @(posedge clk) if (en_in) n976 <= 1'b0 ? 1'b0 : n5104;
/* FF 24 15  6 */ always @(posedge clk) if (n3233) n3381 <= 1'b0 ? 1'b0 : n5105;
/* FF 10 19  0 */ assign n5106 = n1188;
/* FF  9  9  2 */ always @(posedge clk) if (n983) n829 <= 1'b0 ? 1'b0 : n5107;
/* FF 13 11  1 */ always @(posedge clk) if (n1137) n1442 <= 1'b0 ? 1'b0 : n5108;
/* FF 13 22  6 */ always @(posedge clk) if (n1069) n1522 <= 1'b0 ? 1'b0 : n5109;
/* FF 18 15  3 */ always @(posedge clk) if (n1) n2269 <= 1'b0 ? 1'b0 : n5110;
/* FF 26 14  1 */ always @(posedge clk) if (n3527) n3534 <= 1'b0 ? 1'b0 : n5111;
/* FF 14 15  7 */ always @(posedge clk) if (n1792) n1645 <= 1'b0 ? 1'b0 : n5112;
/* FF  2  9  4 */ always @(posedge clk) if (n153) n161 <= 1'b0 ? 1'b0 : n5113;
/* FF 20  4  6 */ always @(posedge clk) if (n1761) n2656 <= 1'b0 ? 1'b0 : n5114;
/* FF 19 20  4 */ always @(posedge clk) if (n2553) n2569 <= 1'b0 ? 1'b0 : n5115;
/* FF 19 11  5 */ always @(posedge clk) if (n2076) n2491 <= 1'b0 ? 1'b0 : n5116;
/* FF 23  9  0 */ always @(posedge clk) if (n2678) n3176 <= 1'b0 ? 1'b0 : n5117;
/* FF 22 19  2 */ assign n2574 = n3261;
/* FF 10  5  3 */ always @(posedge clk) if (en_in) n969 <= 1'b0 ? 1'b0 : n5118;
/* FF 24 18  0 */ always @(posedge clk) if (n3411) n3402 <= 1'b0 ? 1'b0 : n5119;
/* FF 21  9  3 */ always @(posedge clk) if (n2856) n2848 <= 1'b0 ? 1'b0 : n5120;
/* FF  9 27  2 */ always @(posedge clk) if (n804) n948 <= 1'b0 ? 1'b0 : n5121;
/* FF 12 11  5 */ assign \rco[24]  = n5122;
/* FF 26 16  6 */ always @(posedge clk) if (n3249) n3546 <= 1'b0 ? 1'b0 : n5123;
/* FF  3 17  7 */ always @(posedge clk) if (n79) n316 <= 1'b0 ? 1'b0 : n5124;
/* FF 12 16  4 */ always @(posedge clk) if (n1155) n1308 <= 1'b0 ? 1'b0 : n5125;
/* FF 14 25  2 */ always @(posedge clk) if (n697) n1703 <= 1'b0 ? 1'b0 : n5126;
/* FF 26 13  5 */ always @(posedge clk) if (n3033) n3530 <= 1'b0 ? 1'b0 : n5127;
/* FF 17 15  7 */ always @(posedge clk) if (n2111) n2108 <= 1'b0 ? 1'b0 : n5128;
/* FF 29 21  4 */ always @(posedge clk) if (n3788) n3879 <= 1'b0 ? 1'b0 : n5129;
/* FF 20  7  0 */ always @(posedge clk) if (n2670) n2661 <= 1'b0 ? 1'b0 : n5130;
/* FF  5 14  1 */ always @(posedge clk) if (n402) n505 <= 1'b0 ? 1'b0 : n5131;
/* FF 11 24  3 */ always @(posedge clk) if (n796) n1226 <= 1'b0 ? 1'b0 : n5132;
/* FF 16 17  0 */ always @(posedge clk) if (n2110) n1963 <= 1'b0 ? 1'b0 : n5133;
/* FF 21 27  0 */ always @(posedge clk) if (n2196) n2972 <= 1'b0 ? 1'b0 : n5134;
/* FF 13 15  6 */ always @(posedge clk) if (n739) n1476 <= 1'b0 ? 1'b0 : n5135;
/* FF 27  6  7 */ always @(posedge clk) if (n3488) n3596 <= 1'b0 ? 1'b0 : n5136;
/* FF  7 15  6 */ assign n645 = n5137;
/* FF  9 24  4 */ always @(posedge clk) if (n820) n936 <= 1'b0 ? 1'b0 : n5138;
/* FF 13 26  1 */ always @(posedge clk) if (n1271) n1545 <= 1'b0 ? 1'b0 : n5139;
/* FF 21 22  7 */ always @(posedge clk) if (n2384) n2941 <= 1'b0 ? 1'b0 : n5140;
/* FF 18 19  6 */ always @(posedge clk) if (n1982) n2345 <= 1'b0 ? 1'b0 : n5141;
/* FF  3 18  3 */ always @(posedge clk) if (n215) n321 <= 1'b0 ? 1'b0 : n5142;
/* FF 18 28  7 */ always @(posedge clk) if (n2020) n2407 <= 1'b0 ? 1'b0 : n5143;
/* FF  1 19  7 */ always @(posedge clk) if (n119) n111 <= 1'b0 ? 1'b0 : n5144;
/* FF 28 17  2 */ always @(posedge clk) if (n3765) n3768 <= 1'b0 ? 1'b0 : n5145;
/* FF 16 15  3 */ always @(posedge clk) if (n739) n1946 <= 1'b0 ? 1'b0 : n5146;
/* FF  5 16  5 */ always @(posedge clk) if (n511) n523 <= 1'b0 ? 1'b0 : n5147;
/* FF 19  7  6 */ always @(posedge clk) if (n2670) n2458 <= 1'b0 ? 1'b0 : n5148;
/* FF 23 13  5 */ always @(posedge clk) if (n3045) n3213 <= 1'b0 ? 1'b0 : n5149;
/* FF 10 25  6 */ always @(posedge clk) if (n567) n1085 <= 1'b0 ? 1'b0 : n5150;
/* FF 24 14  5 */ always @(posedge clk) if (n3376) n1950 <= 1'b0 ? 1'b0 : n5151;
/* FF 10 18  7 */ always @(posedge clk) if (n1187) n1040 <= 1'b0 ? 1'b0 : n5152;
/* FF  9 10  3 */ always @(posedge clk) if (n988) n837 <= 1'b0 ? 1'b0 : n5153;
/* FF 13 12  0 */ always @(posedge clk) if (n1137) n1449 <= 1'b0 ? 1'b0 : n5154;
/* FF 15 18  1 */ always @(posedge clk) if (n1355) n1809 <= 1'b0 ? 1'b0 : n5155;
/* FF 20 27  2 */ always @(posedge clk) if (n2195) n2816 <= 1'b0 ? 1'b0 : n5156;
/* FF 12 20  1 */ assign n1337 = n5157;
/* FF 14 14  0 */ always @(posedge clk) if (n1791) n1632 <= 1'b0 ? 1'b0 : n5158;
/* FF 17 11  4 */ always @(posedge clk) if (n2076) n2070 <= 1'b0 ? 1'b0 : n5159;
/* FF  1 16  3 */ always @(posedge clk) if (n85) n91 <= 1'b0 ? 1'b0 : n5160;
/* FF 19 21  3 */ always @(posedge clk) if (n2164) n2579 <= 1'b0 ? 1'b0 : n5161;
/* FF 19  8  4 */ always @(posedge clk) if (n2451) n2465 <= 1'b0 ? 1'b0 : n5162;
/* FF 23 14  1 */ always @(posedge clk) if (n2551) n2740 <= 1'b0 ? 1'b0 : n5163;
/* FF 24 17  1 */ always @(posedge clk) if (n2123) n3395 <= 1'b0 ? 1'b0 : n5164;
/* FF 28  7  2 */ always @(posedge clk) if (n3488) n3721 <= 1'b0 ? 1'b0 : n5165;
/* FF  3 14  5 */ assign n290 = n5166;
/* FF  7 19  3 */ always @(posedge clk) if (n549) n760 <= 1'b0 ? 1'b0 : n5167;
/* FF  9 20  3 */ assign n5168 = n1057;
/* FF 21 10  2 */ assign n2855 = n5169;
/* FF 27  9  3 */ always @(posedge clk) if (n3621) n3613 <= 1'b0 ? 1'b0 : n5170;
/* FF 17  5  5 */ assign \rco[176]  = n5171;
/* FF 12 23  5 */ always @(posedge clk) if (n1357) n1363 <= 1'b0 ? 1'b0 : n5172;
/* FF 14 24  1 */ assign n5173 = n1874;
/* FF 26 12  6 */ always @(posedge clk) if (n3368) n3523 <= 1'b0 ? 1'b0 : n5174;
/* FF 17  8  6 */ assign n1625 = n5175;
/* FF  2  7  3 */ always @(posedge clk) if (n21) n149 <= 1'b0 ? 1'b0 : n5176;
/* FF  4 12  6 */ always @(posedge clk) if (n77) n399 <= 1'b0 ? 1'b0 : n5177;
/* FF 22 12  1 */ always @(posedge clk) if (n3029) n3037 <= 1'b0 ? 1'b0 : n5178;
/* FF 10 22  4 */ assign n363 = n5179;
/* FF 21 28  1 */ always @(posedge clk) if (n2196) n2980 <= 1'b0 ? 1'b0 : n5180;
/* FF 13 16  7 */ always @(posedge clk) if (n922) n1042 <= 1'b0 ? 1'b0 : n5181;
/* FF 27  7  4 */ always @(posedge clk) if (n3459) n3599 <= 1'b0 ? 1'b0 : n5182;
/* FF  9 25  7 */ always @(posedge clk) if (n2) n648 <= 1'b0 ? 1'b0 : n5183;
/* FF 27 10  7 */ assign n3621 = n5184;
/* FF 13 27  6 */ always @(posedge clk) if (n1532) n1555 <= 1'b0 ? 1'b0 : n5185;
/* FF 18 18  1 */ always @(posedge clk) if (n1825) n2335 <= 1'b0 ? 1'b0 : n5186;
/* FF  3 19  0 */ assign n328 = n5187;
/* FF 20 20  0 */ always @(posedge clk) if (n2562) n2761 <= 1'b0 ? 1'b0 : n5188;
/* FF 23 18  3 */ always @(posedge clk) if (n2573) n3245 <= 1'b0 ? 1'b0 : n5189;
/* FF 14 10  5 */ always @(posedge clk) if (n1622) n1609 <= 1'b0 ? 1'b0 : n5190;
/* FF  1  7  7 */ assign \rco[22]  = n5191;
/* FF  5 17  6 */ always @(posedge clk) if (n2) n529 <= 1'b0 ? 1'b0 : n5192;
/* FF  4 15  0 */ always @(posedge clk) if (n207) n412 <= 1'b0 ? 1'b0 : n5193;
/* FF 10 24  5 */ always @(posedge clk) if (n820) n1077 <= 1'b0 ? 1'b0 : n5194;
/* FF 24 13  4 */ always @(posedge clk) if (n3351) n3365 <= 1'b0 ? 1'b0 : n5195;
/* FF 10 21  6 */ always @(posedge clk) if (n818) n1063 <= 1'b0 ? 1'b0 : n5196;
/* FF 13 13  3 */ always @(posedge clk) if (n1015) n1458 <= 1'b0 ? 1'b0 : n5197;
/* FF 15 19  2 */ always @(posedge clk) if (n1355) n1819 <= 1'b0 ? 1'b0 : n5198;
/* FF 20 26  1 */ always @(posedge clk) if (n2615) n2806 <= 1'b0 ? 1'b0 : n5199;
/* FF 12 27  0 */ assign \rco[102]  = n5200;
/* FF 17 20  5 */ always @(posedge clk) if (n1843) n2141 <= 1'b0 ? 1'b0 : n5201;
/* FF  2 11  6 */ always @(posedge clk) if (n168) n174 <= 1'b0 ? 1'b0 : n5202;
/* FF 19 18  2 */ always @(posedge clk) if (n2348) n2556 <= 1'b0 ? 1'b0 : n5203;
/* FF 23 15  2 */ always @(posedge clk) if (n3216) n3224 <= 1'b0 ? 1'b0 : n5204;
/* FF 28  6  1 */ always @(posedge clk) if (n3594) n3712 <= 1'b0 ? 1'b0 : n5205;
/* FF 27 22  1 */ always @(posedge clk) if (n3703) n3696 <= 1'b0 ? 1'b0 : n5206;
/* FF  3 15  6 */ always @(posedge clk) if (n207) n299 <= 1'b0 ? 1'b0 : n5207;
/* FF 21 16  4 */ always @(posedge clk) if (n2551) n2891 <= 1'b0 ? 1'b0 : n5208;
/* FF  7 16  2 */ always @(posedge clk) if (n630) n743 <= 1'b0 ? 1'b0 : n5209;
/* FF  9 21  0 */ always @(posedge clk) if (n818) n914 <= 1'b0 ? 1'b0 : n5210;
/* FF 21 11  5 */ always @(posedge clk) if (n2085) n2862 <= 1'b0 ? 1'b0 : n5211;
/* FF 26 18  0 */ assign \rco[32]  = n3664;
/* FF 18 22  6 */ always @(posedge clk) if (n2164) n2359 <= 1'b0 ? 1'b0 : n5212;
/* FF 17  6  4 */ always @(posedge clk) if (n2045) n2042 <= 1'b0 ? 1'b0 : n5213;
/* FF 12 22  6 */ always @(posedge clk) if (n1357) n1353 <= 1'b0 ? 1'b0 : n5214;
/* FF 17  9  5 */ assign n5215 = n2272;
/* FF 10  9  0 */ always @(posedge clk) if (n983) n978 <= 1'b0 ? 1'b0 : n5216;
/* FF 28 20  2 */ assign n3786 = n5217;
/* FF 22 26  7 */ always @(posedge clk) if (n2613) n3140 <= 1'b0 ? 1'b0 : n5218;
/* FF 22 15  0 */ always @(posedge clk) if (n3216) n3058 <= 1'b0 ? 1'b0 : n5219;
/* FF  7  6  1 */ always @(posedge clk) if (n588) n707 <= 1'b0 ? 1'b0 : n5220;
/* FF  9  7  1 */ always @(posedge clk) if (n588) n824 <= 1'b0 ? 1'b0 : n5221;
/* FF 13 17  4 */ always @(posedge clk) if (n1461) n1488 <= 1'b0 ? 1'b0 : n5222;
/* FF  9 26  6 */ always @(posedge clk) if (n954) n944 <= 1'b0 ? 1'b0 : n5223;
/* FF 13 28  7 */ always @(posedge clk) if (n1394) n1567 <= 1'b0 ? 1'b0 : n5224;
/* FF 27 11  4 */ always @(posedge clk) if (n3460) n3625 <= 1'b0 ? 1'b0 : n5225;
/* FF 18 21  0 */ always @(posedge clk) if (n2347) n2349 <= 1'b0 ? 1'b0 : n5226;
/* FF  3 16  1 */ always @(posedge clk) if (n197) n304 <= 1'b0 ? 1'b0 : n5227;
/* FF  6 10  0 */ always @(posedge clk) if (n589) n591 <= 1'b0 ? 1'b0 : n5228;
/* FF 20 11  1 */ assign n962 = n2866;
/* FF 23 19  0 */ always @(posedge clk) if (n2573) n3250 <= 1'b0 ? 1'b0 : n5229;
/* FF 14  5  4 */ always @(posedge clk) if (n1577) n1575 <= 1'b0 ? 1'b0 : n5230;
/* FF 29  9  2 */ assign \rco[77]  = n5231;
/* FF 17 27  1 */ always @(posedge clk) if (n1) n2189 <= 1'b0 ? 1'b0 : n5232;
/* FF 28 23  4 */ always @(posedge clk) if (n3704) n3811 <= 1'b0 ? 1'b0 : n5233;
/* FF 19  5  0 */ always @(posedge clk) if (n2230) n2435 <= 1'b0 ? 1'b0 : n5234;
/* FF  4 14  3 */ assign \rco[15]  = n514;
/* FF 22 25  3 */ always @(posedge clk) if (n2812) n3128 <= 1'b0 ? 1'b0 : n5235;
/* FF 10 27  4 */ always @(posedge clk) if (n804) n1097 <= 1'b0 ? 1'b0 : n5236;
/* FF 24 12  3 */ always @(posedge clk) if (n3351) n3356 <= 1'b0 ? 1'b0 : n5237;
/* FF 10 20  5 */ always @(posedge clk) if (n922) n1043 <= 1'b0 ? 1'b0 : n5238;
/* FF 13 14  2 */ always @(posedge clk) if (n1461) n1464 <= 1'b0 ? 1'b0 : n5239;
/* FF 15 16  3 */ always @(posedge clk) if (n1500) n1796 <= 1'b0 ? 1'b0 : n5240;
/* FF 21 15  2 */ assign n5241 = n3067;
/* FF 20 25  0 */ always @(posedge clk) if (n2612) n2798 <= 1'b0 ? 1'b0 : n5242;
/* FF 26 22  5 */ always @(posedge clk) if (n2730) n3573 <= 1'b0 ? 1'b0 : n5243;
/* FF 15  5  7 */ always @(posedge clk) if (n1742) n1731 <= 1'b0 ? 1'b0 : n5244;
/* FF 12 26  3 */ always @(posedge clk) if (n1393) n1388 <= 1'b0 ? 1'b0 : n5245;
/* FF 14  8  2 */ always @(posedge clk) if (n1741) n1595 <= 1'b0 ? 1'b0 : n5246;
/* FF  2 10  1 */ always @(posedge clk) if (n168) n166 <= 1'b0 ? 1'b0 : n5247;
/* FF  1 18  1 */ always @(posedge clk) if (n115) n99 <= 1'b0 ? 1'b0 : n5248;
/* FF 19 19  1 */ assign n732 = n5249;
/* FF 17 21  6 */ always @(posedge clk) if (n2347) n2150 <= 1'b0 ? 1'b0 : n5250;
/* FF 17 24  5 */ always @(posedge clk) if (n2000) n2171 <= 1'b0 ? 1'b0 : n5251;
/* FF 23 12  3 */ always @(posedge clk) if (n3031) n3203 <= 1'b0 ? 1'b0 : n5252;
/* FF 28  5  0 */ always @(posedge clk) if (n3488) n3705 <= 1'b0 ? 1'b0 : n5253;
/* FF 27 23  2 */ assign n3124 = n3815;
/* FF  3 12  7 */ always @(posedge clk) if (n168) n284 <= 1'b0 ? 1'b0 : n5254;
/* FF 21 17  7 */ always @(posedge clk) if (n2519) n2901 <= 1'b0 ? 1'b0 : n5255;
/* FF  7 17  5 */ always @(posedge clk) if (n549) n756 <= 1'b0 ? 1'b0 : n5256;
/* FF  9 22  1 */ always @(posedge clk) if (n819) n924 <= 1'b0 ? 1'b0 : n5257;
/* FF 21 12  4 */ always @(posedge clk) if (n3029) n2871 <= 1'b0 ? 1'b0 : n5258;
/* FF 12  8  0 */ always @(posedge clk) if (n1131) n1278 <= 1'b0 ? 1'b0 : n5259;
/* FF 26 21  1 */ always @(posedge clk) if (n3421) n3563 <= 1'b0 ? 1'b0 : n5260;
/* FF 15  6  3 */ always @(posedge clk) if (n1744) n1736 <= 1'b0 ? 1'b0 : n5261;
/* FF 17  7  3 */ always @(posedge clk) if (n2045) n2049 <= 1'b0 ? 1'b0 : n5262;
/* FF 12 21  7 */ always @(posedge clk) if (n1205) n1346 <= 1'b0 ? 1'b0 : n5263;
/* FF 18 25  7 */ always @(posedge clk) if (n1878) n2383 <= 1'b0 ? 1'b0 : n5264;
/* FF 17 10  4 */ always @(posedge clk) if (n2282) n2063 <= 1'b0 ? 1'b0 : n5265;
/* FF  9 32  7 */ assign \rco[107]  = n5266;
/* FF  1 12  5 */ always @(posedge clk) if (n39) n51 <= 1'b0 ? 1'b0 : n5267;
/* FF 22 14  7 */ always @(posedge clk) if (n3045) n3057 <= 1'b0 ? 1'b0 : n5268;
/* FF  7  7  2 */ always @(posedge clk) if (n588) n711 <= 1'b0 ? 1'b0 : n5269;
/* FF 13 18  5 */ always @(posedge clk) if (n1205) n1497 <= 1'b0 ? 1'b0 : n5270;
/* FF 27  5  2 */ always @(posedge clk) if (n3594) n3587 <= 1'b0 ? 1'b0 : n5271;
/* FF 27  8  5 */ always @(posedge clk) if (n3464) n3607 <= 1'b0 ? 1'b0 : n5272;
/* FF 18 20  3 */ assign \rco[153]  = n2575;
/* FF  6 21  1 */ always @(posedge clk) if (n778) n243 <= 1'b0 ? 1'b0 : n5273;
/* FF 20 10  2 */ always @(posedge clk) if (n2697) n2685 <= 1'b0 ? 1'b0 : n5274;
/* FF 23 16  1 */ always @(posedge clk) if (n2540) n3230 <= 1'b0 ? 1'b0 : n5275;
/* FF 11 14  2 */ always @(posedge clk) if (n1154) n1148 <= 1'b0 ? 1'b0 : n5276;
/* FF  2 14  6 */ always @(posedge clk) if (n83) n193 <= 1'b0 ? 1'b0 : n5277;
/* FF 16  7  7 */ always @(posedge clk) if (n1743) n1745 <= 1'b0 ? 1'b0 : n5278;
/* FF 29 10  3 */ always @(posedge clk) if (n3464) n3835 <= 1'b0 ? 1'b0 : n5279;
/* FF 28 22  7 */ always @(posedge clk) if (n3704) n3806 <= 1'b0 ? 1'b0 : n5280;
/* FF 16 12  6 */ always @(posedge clk) if (n1771) n1941 <= 1'b0 ? 1'b0 : n5281;
/* FF  5 19  0 */ always @(posedge clk) if (n349) n539 <= 1'b0 ? 1'b0 : n5282;
/* FF  4 13  2 */ assign \rco[20]  = n5283;
/* FF 22 24  0 */ always @(posedge clk) if (n3113) n3116 <= 1'b0 ? 1'b0 : n5284;
/* FF 10 26  3 */ assign n1089 = n1245;
/* FF 24 11  2 */ assign n2910 = n3465;
/* FF 10 23  4 */ assign n1065 = n5285;
/* FF 15 17  4 */ always @(posedge clk) if (n1500) n1805 <= 1'b0 ? 1'b0 : n5286;
/* FF 18  6  0 */ always @(posedge clk) if (n2241) n2231 <= 1'b0 ? 1'b0 : n5287;
/* FF  7 21  2 */ always @(posedge clk) if (n360) n770 <= 1'b0 ? 1'b0 : n5288;
/* FF  6  7  0 */ always @(posedge clk) if (n570) n571 <= 1'b0 ? 1'b0 : n5289;
/* FF 20 24  7 */ always @(posedge clk) if (n2775) n2795 <= 1'b0 ? 1'b0 : n5290;
/* FF 26  9  4 */ always @(posedge clk) if (n3460) n3502 <= 1'b0 ? 1'b0 : n5291;
/* FF 12 25  2 */ always @(posedge clk) if (n1532) n1378 <= 1'b0 ? 1'b0 : n5292;
/* FF 14 11  3 */ always @(posedge clk) if (n1622) n1615 <= 1'b0 ? 1'b0 : n5293;
/* FF  2 13  0 */ always @(posedge clk) if (n83) n185 <= 1'b0 ? 1'b0 : n5294;
/* FF 17 22  7 */ always @(posedge clk) if (n1999) n2159 <= 1'b0 ? 1'b0 : n5295;
/* FF 19 16  0 */ assign n2534 = n2731;
/* FF 17 25  6 */ always @(posedge clk) if (n2017) n2182 <= 1'b0 ? 1'b0 : n5296;
/* FF 27 20  3 */ always @(posedge clk) if (n3424) n3678 <= 1'b0 ? 1'b0 : n5297;
/* FF  4 19  2 */ assign \rco[130]  = n5298;
/* FF  3 13  0 */ assign n77 = n5299;
/* FF 21 18  6 */ always @(posedge clk) if (n2757) n2908 <= 1'b0 ? 1'b0 : n5300;
/* FF 22 10  4 */ always @(posedge clk) if (n2856) n3026 <= 1'b0 ? 1'b0 : n5301;
/* FF  7 22  4 */ always @(posedge clk) if (n695) n787 <= 1'b0 ? 1'b0 : n5302;
/* FF  9 23  6 */ always @(posedge clk) if (n819) n931 <= 1'b0 ? 1'b0 : n5303;
/* FF 21 13  7 */ always @(posedge clk) if (n2519) n2550 <= 1'b0 ? 1'b0 : n5304;
/* FF 12 15  1 */ always @(posedge clk) if (n1155) n1297 <= 1'b0 ? 1'b0 : n5305;
/* FF 26 20  2 */ always @(posedge clk) if (n3424) n3241 <= 1'b0 ? 1'b0 : n5306;
/* FF 15  7  0 */ assign \rco[88]  = n5307;
/* FF 18 24  4 */ always @(posedge clk) if (n1878) n2374 <= 1'b0 ? 1'b0 : n5308;
/* FF 19 30  3 */ always @(posedge clk) if (n2592) n2637 <= 1'b0 ? 1'b0 : n5309;
/* FF 11 17  0 */ always @(posedge clk) if (n900) n1168 <= 1'b0 ? 1'b0 : n5310;
/* FF 10 11  2 */ assign n988 = n5311;
/* FF 16  8  3 */ always @(posedge clk) if (n1625) n1918 <= 1'b0 ? 1'b0 : n5312;
/* FF  1 13  6 */ always @(posedge clk) if (n83) n65 <= 1'b0 ? 1'b0 : n5313;
/* FF 22  9  6 */ always @(posedge clk) if (n2989) n3020 <= 1'b0 ? 1'b0 : n5314;
/* FF 13 19  2 */ assign n5315 = n1673;
/* FF 15 21  1 */ always @(posedge clk) if (n1356) n1837 <= 1'b0 ? 1'b0 : n5316;
/* FF 20 28  4 */ always @(posedge clk) if (n2195) n2825 <= 1'b0 ? 1'b0 : n5317;
/* FF 18 23  2 */ always @(posedge clk) if (n1999) n2364 <= 1'b0 ? 1'b0 : n5318;
/* FF  6 20  2 */ always @(posedge clk) if (n552) n662 <= 1'b0 ? 1'b0 : n5319;
/* FF 20  9  3 */ assign n5320 = n2853;
/* FF 23 17  6 */ always @(posedge clk) if (n2540) n3238 <= 1'b0 ? 1'b0 : n5321;
/* FF 11 15  1 */ assign n891 = n5322;
/* FF 26  6  2 */ always @(posedge clk) if (n3459) n3475 <= 1'b0 ? 1'b0 : n5323;
/* FF 14  7  6 */ always @(posedge clk) if (n1743) n1590 <= 1'b0 ? 1'b0 : n5324;
/* FF 16  6  4 */ always @(posedge clk) if (n1744) n1901 <= 1'b0 ? 1'b0 : n5325;
/* FF 29 11  4 */ always @(posedge clk) if (n3751) n3843 <= 1'b0 ? 1'b0 : n5326;
/* FF 28 21  6 */ always @(posedge clk) if (n3788) n3797 <= 1'b0 ? 1'b0 : n5327;
/* FF 19  3  2 */ always @(posedge clk) if (n1887) n2429 <= 1'b0 ? 1'b0 : n5328;
/* FF 22 27  1 */ always @(posedge clk) if (n2970) n3144 <= 1'b0 ? 1'b0 : n5329;
/* FF 10 29  2 */ always @(posedge clk) if (n821) n1110 <= 1'b0 ? 1'b0 : n5330;
/* FF 24 10  1 */ always @(posedge clk) if (n3352) n3341 <= 1'b0 ? 1'b0 : n5331;
/* FF  3  9  5 */ always @(posedge clk) if (n260) n257 <= 1'b0 ? 1'b0 : n5332;
/* FF 15 22  5 */ always @(posedge clk) if (n1835) n457 <= 1'b0 ? 1'b0 : n5333;
/* FF 18  9  1 */ always @(posedge clk) if (n2055) n2262 <= 1'b0 ? 1'b0 : n5334;
/* FF  7 26  3 */ always @(posedge clk) if (n567) n801 <= 1'b0 ? 1'b0 : n5335;
/* FF  9 19  3 */ always @(posedge clk) if (n454) n904 <= 1'b0 ? 1'b0 : n5336;
/* FF 12 19  4 */ always @(posedge clk) if (n1501) n1332 <= 1'b0 ? 1'b0 : n5337;
/* FF 26  8  7 */ always @(posedge clk) if (n3603) n3497 <= 1'b0 ? 1'b0 : n5338;
/* FF 12 24  5 */ always @(posedge clk) if (n961) n1372 <= 1'b0 ? 1'b0 : n5339;
/* FF 17 23  0 */ always @(posedge clk) if (n1069) n2160 <= 1'b0 ? 1'b0 : n5340;
/* FF  2 12  3 */ always @(posedge clk) if (n39) n179 <= 1'b0 ? 1'b0 : n5341;
/* FF 22 21  0 */ always @(posedge clk) if (n2564) n3096 <= 1'b0 ? 1'b0 : n5342;
/* FF 24 24  2 */ always @(posedge clk) if (n3112) n3441 <= 1'b0 ? 1'b0 : n5343;
/* FF 27 21  4 */ always @(posedge clk) if (n3421) n3691 <= 1'b0 ? 1'b0 : n5344;
/* FF  4 18  1 */ always @(posedge clk) if (n349) n431 <= 1'b0 ? 1'b0 : n5345;
/* FF  3 10  1 */ always @(posedge clk) if (n251) n263 <= 1'b0 ? 1'b0 : n5346;
/* FF 13 23  7 */ always @(posedge clk) if (n1069) n1531 <= 1'b0 ? 1'b0 : n5347;
/* FF 27 14  6 */ always @(posedge clk) if (n3527) n3647 <= 1'b0 ? 1'b0 : n5348;
/* FF  9 16  7 */ always @(posedge clk) if (n645) n882 <= 1'b0 ? 1'b0 : n5349;
/* FF 12 14  2 */ always @(posedge clk) if (n1154) n1290 <= 1'b0 ? 1'b0 : n5350;
/* FF 26 23  3 */ always @(posedge clk) if (n3703) n3579 <= 1'b0 ? 1'b0 : n5351;
/* FF 18 27  5 */ always @(posedge clk) if (n2020) n1709 <= 1'b0 ? 1'b0 : n5352;
/* FF 19 31  0 */ always @(posedge clk) if (n2592) n2641 <= 1'b0 ? 1'b0 : n5353;
/* FF 23 21  3 */ always @(posedge clk) if (n3258) n3274 <= 1'b0 ? 1'b0 : n5354;
/* FF 16 23  2 */ always @(posedge clk) if (n2000) n1993 <= 1'b0 ? 1'b0 : n5355;
/* FF  1 14  7 */ always @(posedge clk) if (n85) n75 <= 1'b0 ? 1'b0 : n5356;
/* FF 22  7  4 */ always @(posedge clk) if (n2841) n3002 <= 1'b0 ? 1'b0 : n5357;
/* FF 22  8  5 */ always @(posedge clk) if (n2989) n3013 <= 1'b0 ? 1'b0 : n5358;
/* FF 13 20  3 */ always @(posedge clk) if (n1339) n1506 <= 1'b0 ? 1'b0 : n5359;
/* FF 15 10  0 */ always @(posedge clk) if (n1624) n1754 <= 1'b0 ? 1'b0 : n5360;
/* FF 20 19  5 */ always @(posedge clk) if (n2562) n2754 <= 1'b0 ? 1'b0 : n5361;
/* FF  6 23  3 */ always @(posedge clk) if (n360) n690 <= 1'b0 ? 1'b0 : n5362;
/* FF 20  8  4 */ always @(posedge clk) if (n2247) n2672 <= 1'b0 ? 1'b0 : n5363;
/* FF 12 28  2 */ always @(posedge clk) if (n1394) n1396 <= 1'b0 ? 1'b0 : n5364;
/* FF 23 22  7 */ always @(posedge clk) if (n3422) n3286 <= 1'b0 ? 1'b0 : n5365;
/* FF 14  6  1 */ always @(posedge clk) if (n1577) n1578 <= 1'b0 ? 1'b0 : n5366;
/* FF 16  5  5 */ always @(posedge clk) if (n1742) n1893 <= 1'b0 ? 1'b0 : n5367;
/* FF 17 19  5 */ always @(posedge clk) if (n1982) n2133 <= 1'b0 ? 1'b0 : n5368;
/* FF 29 12  5 */ always @(posedge clk) if (n3751) n3847 <= 1'b0 ? 1'b0 : n5369;
/* FF 16 10  4 */ always @(posedge clk) if (n1771) n1930 <= 1'b0 ? 1'b0 : n5370;
/* FF  5 21  2 */ assign n552 = n5371;
/* FF 10 28  1 */ always @(posedge clk) if (n821) n1102 <= 1'b0 ? 1'b0 : n5372;
/* FF  9 12  1 */ always @(posedge clk) if (n996) n851 <= 1'b0 ? 1'b0 : n5373;
/* FF 24  9  0 */ always @(posedge clk) if (n3352) n3332 <= 1'b0 ? 1'b0 : n5374;
/* FF 27 17  1 */ always @(posedge clk) if (n3249) n3652 <= 1'b0 ? 1'b0 : n5375;
/* FF 15 24  7 */ always @(posedge clk) if (n778) n1870 <= 1'b0 ? 1'b0 : n5376;
/* FF 21 23  6 */ always @(posedge clk) if (n2961) n2949 <= 1'b0 ? 1'b0 : n5377;
/* FF 15 23  6 */ always @(posedge clk) if (n778) n1858 <= 1'b0 ? 1'b0 : n5378;
/* FF 18  8  2 */ always @(posedge clk) if (n2055) n2251 <= 1'b0 ? 1'b0 : n5379;
/* FF 12 18  7 */ always @(posedge clk) if (n1501) n1327 <= 1'b0 ? 1'b0 : n5380;
/* FF 26 11  6 */ always @(posedge clk) if (n3033) n3514 <= 1'b0 ? 1'b0 : n5381;
/* FF 29 19  3 */ always @(posedge clk) if (n3786) n3864 <= 1'b0 ? 1'b0 : n5382;
/* FF 17 16  1 */ assign \rco[27]  = n2322;
/* FF  2 15  2 */ assign n197 = n5383;
/* FF 22 20  3 */ always @(posedge clk) if (n3087) n3091 <= 1'b0 ? 1'b0 : n5384;
/* FF 10 14  2 */ always @(posedge clk) if (n750) n1009 <= 1'b0 ? 1'b0 : n5385;
/* FF 24 23  3 */ always @(posedge clk) if (n3104) n3436 <= 1'b0 ? 1'b0 : n5386;
/* FF 16 24  0 */ assign \rco[127]  = n5387;
/* FF 27 18  5 */ always @(posedge clk) if (n3553) n3662 <= 1'b0 ? 1'b0 : n5388;
/* FF  4 17  0 */ assign n325 = n5389;
/* FF  3 11  2 */ always @(posedge clk) if (n153) n272 <= 1'b0 ? 1'b0 : n5390;
/* FF  7  9  1 */ always @(posedge clk) if (n589) n719 <= 1'b0 ? 1'b0 : n5391;
/* FF 21 20  0 */ always @(posedge clk) if (n3087) n2918 <= 1'b0 ? 1'b0 : n5392;
/* FF 13 24  6 */ assign \rco[111]  = n5393;
/* FF 27 15  5 */ always @(posedge clk) if (n3233) n3650 <= 1'b0 ? 1'b0 : n5394;
/* FF  9 17  4 */ always @(posedge clk) if (n1030) n887 <= 1'b0 ? 1'b0 : n5395;
/* FF 18 26  2 */ always @(posedge clk) if (n2615) n2387 <= 1'b0 ? 1'b0 : n5396;
/* FF 20 12  1 */ always @(posedge clk) if (n2682) n2699 <= 1'b0 ? 1'b0 : n5397;
/* FF 19 28  1 */ always @(posedge clk) if (n2614) n2625 <= 1'b0 ? 1'b0 : n5398;
/* FF 28 19  7 */ always @(posedge clk) if (n3424) n3783 <= 1'b0 ? 1'b0 : n5399;
/* FF 10 13  4 */ always @(posedge clk) if (n629) n1005 <= 1'b0 ? 1'b0 : n5400;
/* FF 28 24  6 */ assign \rco[139]  = n5401;
/* FF 16 22  1 */ assign \rco[119]  = n5402;
/* FF  1 15  0 */ assign \rco[5]  = n202;
/* FF 22  6  3 */ always @(posedge clk) if (n2841) n2993 <= 1'b0 ? 1'b0 : n5403;
/* FF 22 11  4 */ assign \rco[55]  = n5404;
/* FF 13 21  0 */ always @(posedge clk) if (n1356) n1513 <= 1'b0 ? 1'b0 : n5405;
/* FF 30 10  0 */ always @(posedge clk) if (n3892) n3885 <= 1'b0 ? 1'b0 : n5406;
/* FF 15 11  3 */ always @(posedge clk) if (n1624) n1766 <= 1'b0 ? 1'b0 : n5407;
/* FF  2 19  0 */ assign n115 = n5408;
/* FF  6 13  5 */ always @(posedge clk) if (n78) n620 <= 1'b0 ? 1'b0 : n5409;
/* FF 20 18  6 */ always @(posedge clk) if (n2348) n2746 <= 1'b0 ? 1'b0 : n5410;
/* FF  6 22  4 */ always @(posedge clk) if (n673) n682 <= 1'b0 ? 1'b0 : n5411;
/* FF 20 15  5 */ always @(posedge clk) if (n2715) n2722 <= 1'b0 ? 1'b0 : n5412;
/* FF 23 23  4 */ always @(posedge clk) if (n3104) n3291 <= 1'b0 ? 1'b0 : n5413;
/* FF 11 13  7 */ always @(posedge clk) if (n733) n1145 <= 1'b0 ? 1'b0 : n5414;
/* FF 16  4  2 */ always @(posedge clk) if (n1761) n1886 <= 1'b0 ? 1'b0 : n5415;
/* FF  5 22  3 */ always @(posedge clk) if (n673) n558 <= 1'b0 ? 1'b0 : n5416;
/* FF  9 13  2 */ always @(posedge clk) if (n629) n857 <= 1'b0 ? 1'b0 : n5417;
/* FF 13  7  1 */ always @(posedge clk) if (n977) n1424 <= 1'b0 ? 1'b0 : n5418;
/* FF 15 25  0 */ assign \rco[194]  = n5419;
/* FF  7 13  6 */ always @(posedge clk) if (n733) n730 <= 1'b0 ? 1'b0 : n5420;
/* FF 18 11  3 */ assign \rco[37]  = n5421;
/* FF 15 20  7 */ always @(posedge clk) if (n1347) n1834 <= 1'b0 ? 1'b0 : n5422;
/* FF 12 17  6 */ always @(posedge clk) if (n900) n1318 <= 1'b0 ? 1'b0 : n5423;
/* FF 26 10  1 */ always @(posedge clk) if (n3033) n3506 <= 1'b0 ? 1'b0 : n5424;
/* FF 18 30  7 */ always @(posedge clk) if (n1881) n2423 <= 1'b0 ? 1'b0 : n5425;
/* FF 29 20  2 */ always @(posedge clk) if (n3786) n3870 <= 1'b0 ? 1'b0 : n5426;
/* FF 26  7  6 */ always @(posedge clk) if (n3603) n3486 <= 1'b0 ? 1'b0 : n5427;
/* FF 17 17  2 */ always @(posedge clk) if (n2111) n2116 <= 1'b0 ? 1'b0 : n5428;
/* FF 22 23  2 */ assign n3104 = n5429;
/* FF 24 22  0 */ always @(posedge clk) if (n3422) n3425 <= 1'b0 ? 1'b0 : n5430;
/* FF  1 11  5 */ always @(posedge clk) if (n37) n42 <= 1'b0 ? 1'b0 : n5431;
/* FF 27 19  6 */ always @(posedge clk) if (n3553) n3673 <= 1'b0 ? 1'b0 : n5432;
/* FF  7 14  0 */ always @(posedge clk) if (n733) n734 <= 1'b0 ? 1'b0 : n5433;
/* FF 21 21  3 */ always @(posedge clk) if (n2564) n2929 <= 1'b0 ? 1'b0 : n5434;
/* FF 13 25  5 */ always @(posedge clk) if (n697) n1539 <= 1'b0 ? 1'b0 : n5435;
/* FF 27 12  4 */ always @(posedge clk) if (n3368) n3633 <= 1'b0 ? 1'b0 : n5436;
/* FF  9 18  5 */ always @(posedge clk) if (n1030) n897 <= 1'b0 ? 1'b0 : n5437;
/* FF 18 29  3 */ always @(posedge clk) if (n1881) n2411 <= 1'b0 ? 1'b0 : n5438;
/* FF  6 18  1 */ always @(posedge clk) if (n657) n650 <= 1'b0 ? 1'b0 : n5439;
/* FF  5 10  1 */ always @(posedge clk) if (n184) n475 <= 1'b0 ? 1'b0 : n5440;
/* FF 19 29  6 */ always @(posedge clk) if (n2614) n2633 <= 1'b0 ? 1'b0 : n5441;
/* FF 11  9  4 */ always @(posedge clk) if (n1131) n1134 <= 1'b0 ? 1'b0 : n5442;
/* FF 23 27  1 */ always @(posedge clk) if (n2017) n3313 <= 1'b0 ? 1'b0 : n5443;
/* FF 11 28  3 */ always @(posedge clk) if (n1384) n1258 <= 1'b0 ? 1'b0 : n5444;
/* FF 10 12  7 */ always @(posedge clk) if (n996) n1003 <= 1'b0 ? 1'b0 : n5445;
/* FF 24 25  6 */ always @(posedge clk) if (n2812) n3452 <= 1'b0 ? 1'b0 : n5446;
/* FF 16 21  0 */ always @(posedge clk) if (n1835) n1983 <= 1'b0 ? 1'b0 : n5447;
/* FF  1  8  1 */ always @(posedge clk) if (n37) n15 <= 1'b0 ? 1'b0 : n5448;
/* FF 13 22  1 */ always @(posedge clk) if (n1069) n669 <= 1'b0 ? 1'b0 : n5449;
/* FF 31 23  1 */ assign \rco[189]  = n5450;
/* FF 15  8  2 */ always @(posedge clk) if (n1741) n1748 <= 1'b0 ? 1'b0 : n5451;
/* FF  3 22  3 */ always @(posedge clk) if (n352) n356 <= 1'b0 ? 1'b0 : n5452;
/* FF 21  7  3 */ assign n5453 = n3008;
/* FF  6 12  6 */ always @(posedge clk) if (n286) n612 <= 1'b0 ? 1'b0 : n5454;
/* FF 20 17  7 */ always @(posedge clk) if (n2727) n2739 <= 1'b0 ? 1'b0 : n5455;
/* FF 26 14  6 */ always @(posedge clk) if (n3527) n3539 <= 1'b0 ? 1'b0 : n5456;
/* FF 23 20  5 */ always @(posedge clk) if (n3258) n3268 <= 1'b0 ? 1'b0 : n5457;
/* FF  9 14  3 */ always @(posedge clk) if (n629) n862 <= 1'b0 ? 1'b0 : n5458;
/* FF  4 20  4 */ always @(posedge clk) if (n215) n442 <= 1'b0 ? 1'b0 : n5459;
/* FF 21  9  4 */ always @(posedge clk) if (n2856) n2849 <= 1'b0 ? 1'b0 : n5460;
/* FF  9 27  7 */ always @(posedge clk) if (n804) n953 <= 1'b0 ? 1'b0 : n5461;
/* FF 18 10  4 */ always @(posedge clk) if (n2282) n2277 <= 1'b0 ? 1'b0 : n5462;
/* FF 12 16  1 */ always @(posedge clk) if (n1155) n1305 <= 1'b0 ? 1'b0 : n5463;
/* FF 26 13  0 */ assign n3525 = n3639;
/* FF 14 18  0 */ always @(posedge clk) if (n1672) n1661 <= 1'b0 ? 1'b0 : n5464;
/* FF 12 29  6 */ always @(posedge clk) if (n1532) n1406 <= 1'b0 ? 1'b0 : n5465;
/* FF  1 20  3 */ always @(posedge clk) if (n126) n113 <= 1'b0 ? 1'b0 : n5466;
/* FF 19 25  3 */ always @(posedge clk) if (n2612) n2607 <= 1'b0 ? 1'b0 : n5467;
/* FF 23 10  1 */ always @(posedge clk) if (n2697) n3184 <= 1'b0 ? 1'b0 : n5468;
/* FF 22 22  5 */ always @(posedge clk) if (n2961) n3066 <= 1'b0 ? 1'b0 : n5469;
/* FF 24 21  1 */ assign n3421 = n3470;
/* FF 13  5  6 */ always @(posedge clk) if (n1577) n1414 <= 1'b0 ? 1'b0 : n5470;
/* FF  7 15  3 */ assign \rco[9]  = n815;
/* FF  9 24  3 */ always @(posedge clk) if (n820) n935 <= 1'b0 ? 1'b0 : n5471;
/* FF 13 26  4 */ always @(posedge clk) if (n1271) n1548 <= 1'b0 ? 1'b0 : n5472;
/* FF 21 22  2 */ always @(posedge clk) if (n2384) n2937 <= 1'b0 ? 1'b0 : n5473;
/* FF  2 22  4 */ always @(posedge clk) if (n352) n239 <= 1'b0 ? 1'b0 : n5474;
/* FF 18 28  0 */ assign \rco[197]  = n2628;
/* FF 19 26  7 */ assign n2615 = n5475;
/* FF  5 11  6 */ always @(posedge clk) if (n184) n483 <= 1'b0 ? 1'b0 : n5476;
/* FF 11 22  5 */ always @(posedge clk) if (n695) n1211 <= 1'b0 ? 1'b0 : n5477;
/* FF 23 24  0 */ always @(posedge clk) if (n3112) n3296 <= 1'b0 ? 1'b0 : n5478;
/* FF 28 17  5 */ always @(posedge clk) if (n3765) n2124 <= 1'b0 ? 1'b0 : n5479;
/* FF 16 15  6 */ always @(posedge clk) if (n739) n1948 <= 1'b0 ? 1'b0 : n5480;
/* FF 11 29  4 */ always @(posedge clk) if (n1384) n1266 <= 1'b0 ? 1'b0 : n5481;
/* FF 10 15  6 */ always @(posedge clk) if (n750) n1021 <= 1'b0 ? 1'b0 : n5482;
/* FF 16 20  7 */ always @(posedge clk) if (n1843) n1981 <= 1'b0 ? 1'b0 : n5483;
/* FF 21 24  1 */ always @(posedge clk) if (n3113) n2954 <= 1'b0 ? 1'b0 : n5484;
/* FF 15 18  4 */ always @(posedge clk) if (n1355) n1812 <= 1'b0 ? 1'b0 : n5485;
/* FF 18 14  1 */ assign n2303 = n5486;
/* FF  2 21  6 */ always @(posedge clk) if (n126) n233 <= 1'b0 ? 1'b0 : n5487;
/* FF  6 15  7 */ always @(posedge clk) if (n630) n637 <= 1'b0 ? 1'b0 : n5488;
/* FF 12 20  6 */ assign n900 = n5489;
/* FF  6 16  6 */ always @(posedge clk) if (n511) n643 <= 1'b0 ? 1'b0 : n5490;
/* FF 20 13  7 */ always @(posedge clk) if (n2283) n2711 <= 1'b0 ? 1'b0 : n5491;
/* FF 14  3  2 */ assign \rco[87]  = n5492;
/* FF  4 11  0 */ assign n54 = n5493;
/* FF 22 18  2 */ always @(posedge clk) if (n3065) n3082 <= 1'b0 ? 1'b0 : n5494;
/* FF  9 15  4 */ always @(posedge clk) if (n645) n871 <= 1'b0 ? 1'b0 : n5495;
/* FF 28 12  0 */ always @(posedge clk) if (n3462) n3753 <= 1'b0 ? 1'b0 : n5496;
/* FF 21 10  5 */ assign n2519 = n5497;
/* FF  7 19  4 */ always @(posedge clk) if (n549) n761 <= 1'b0 ? 1'b0 : n5498;
/* FF  9 20  6 */ always @(posedge clk) if (n961) n910 <= 1'b0 ? 1'b0 : n5499;
/* FF 18 13  5 */ always @(posedge clk) if (n2283) n2300 <= 1'b0 ? 1'b0 : n5500;
/* FF 12 23  0 */ always @(posedge clk) if (n1357) n1358 <= 1'b0 ? 1'b0 : n5501;
/* FF 26 12  3 */ always @(posedge clk) if (n3368) n3520 <= 1'b0 ? 1'b0 : n5502;
/* FF  5 15  3 */ always @(posedge clk) if (n511) n517 <= 1'b0 ? 1'b0 : n5503;
/* FF 19 22  2 */ always @(posedge clk) if (n2164) n2586 <= 1'b0 ? 1'b0 : n5504;
/* FF 23 11  2 */ always @(posedge clk) if (n3031) n3192 <= 1'b0 ? 1'b0 : n5505;
/* FF 11 25  1 */ always @(posedge clk) if (n954) n1232 <= 1'b0 ? 1'b0 : n5506;
/* FF 22 17  4 */ always @(posedge clk) if (n3065) n3076 <= 1'b0 ? 1'b0 : n5507;
/* FF 24 20  6 */ always @(posedge clk) if (n3411) n3418 <= 1'b0 ? 1'b0 : n5508;
/* FF 16 16  4 */ always @(posedge clk) if (n2110) n1959 <= 1'b0 ? 1'b0 : n5509;
/* FF 13  6  7 */ always @(posedge clk) if (n977) n1422 <= 1'b0 ? 1'b0 : n5510;
/* FF  9 25  0 */ assign \rco[132]  = n5511;
/* FF 13 27  3 */ assign n1243 = n5512;
/* FF 27 10  2 */ assign n3034 = n3749;
/* FF 15 13  2 */ always @(posedge clk) if (n1015) n1779 <= 1'b0 ? 1'b0 : n5513;
/* FF 20 20  5 */ always @(posedge clk) if (n2562) n2759 <= 1'b0 ? 1'b0 : n5514;
/* FF 23 18  6 */ always @(posedge clk) if (n2573) n3247 <= 1'b0 ? 1'b0 : n5515;
/* FF  5 12  7 */ always @(posedge clk) if (n77) n491 <= 1'b0 ? 1'b0 : n5516;
/* FF 19 27  4 */ always @(posedge clk) if (n2614) n2620 <= 1'b0 ? 1'b0 : n5517;
/* FF 11 23  6 */ always @(posedge clk) if (n796) n1219 <= 1'b0 ? 1'b0 : n5518;
/* FF 23 25  7 */ always @(posedge clk) if (n2613) n3309 <= 1'b0 ? 1'b0 : n5519;
/* FF 11 26  5 */ always @(posedge clk) if (n954) n1221 <= 1'b0 ? 1'b0 : n5520;
/* FF 16 19  6 */ always @(posedge clk) if (n1402) n1973 <= 1'b0 ? 1'b0 : n5521;
/* FF  1 10  3 */ always @(posedge clk) if (n37) n31 <= 1'b0 ? 1'b0 : n5522;
/* FF 21 25  2 */ always @(posedge clk) if (n2970) n2964 <= 1'b0 ? 1'b0 : n5523;
/* FF  9 11  1 */ always @(posedge clk) if (n988) n843 <= 1'b0 ? 1'b0 : n5524;
/* FF 15 19  7 */ always @(posedge clk) if (n1355) n1824 <= 1'b0 ? 1'b0 : n5525;
/* FF 18 17  0 */ assign n1825 = n5526;
/* FF  3 20  1 */ always @(posedge clk) if (n119) n343 <= 1'b0 ? 1'b0 : n5527;
/* FF 15 14  4 */ always @(posedge clk) if (n1791) n1787 <= 1'b0 ? 1'b0 : n5528;
/* FF  6 14  0 */ always @(posedge clk) if (n78) n623 <= 1'b0 ? 1'b0 : n5529;
/* FF 20 23  1 */ always @(posedge clk) if (n2553) n2002 <= 1'b0 ? 1'b0 : n5530;
/* FF 12 27  7 */ assign n1394 = n5531;
/* FF 11  8  4 */ always @(posedge clk) if (n1131) n1127 <= 1'b0 ? 1'b0 : n5532;
/* FF 29  5  2 */ always @(posedge clk) if (n3605) n3820 <= 1'b0 ? 1'b0 : n5533;
/* FF 19  9  0 */ always @(posedge clk) if (n2451) n2471 <= 1'b0 ? 1'b0 : n5534;
/* FF  4 10  3 */ always @(posedge clk) if (n251) n382 <= 1'b0 ? 1'b0 : n5535;
/* FF 24 16  3 */ always @(posedge clk) if (n3376) n3387 <= 1'b0 ? 1'b0 : n5536;
/* FF 27 22  4 */ always @(posedge clk) if (n3703) n3699 <= 1'b0 ? 1'b0 : n5537;
/* FF 13 10  2 */ always @(posedge clk) if (n850) n1436 <= 1'b0 ? 1'b0 : n5538;
/* FF 18  3  7 */ always @(posedge clk) if (n1887) n2211 <= 1'b0 ? 1'b0 : n5539;
/* FF  7 16  5 */ always @(posedge clk) if (n630) n746 <= 1'b0 ? 1'b0 : n5540;
/* FF  9 21  5 */ always @(posedge clk) if (n818) n919 <= 1'b0 ? 1'b0 : n5541;
/* FF 18 12  6 */ always @(posedge clk) if (n1936) n2292 <= 1'b0 ? 1'b0 : n5542;
/* FF 21 11  2 */ assign n2859 = n5543;
/* FF 21  6  5 */ always @(posedge clk) if (n2247) n2838 <= 1'b0 ? 1'b0 : n5544;
/* FF 12 22  3 */ always @(posedge clk) if (n1357) n1351 <= 1'b0 ? 1'b0 : n5545;
/* FF 26 15  2 */ always @(posedge clk) if (n3233) n3542 <= 1'b0 ? 1'b0 : n5546;
/* FF 14 12  2 */ assign n1621 = n5547;
/* FF 19 23  1 */ assign \rco[180]  = n5548;
/* FF 10  9  7 */ always @(posedge clk) if (n983) n981 <= 1'b0 ? 1'b0 : n5549;
/* FF 28 20  7 */ assign \rco[163]  = n5550;
/* FF 31  9  1 */ assign \rco[73]  = n5551;
/* FF  4 21  4 */ always @(posedge clk) if (n552) n451 <= 1'b0 ? 1'b0 : n5552;
/* FF 13 28  2 */ always @(posedge clk) if (n1394) n1563 <= 1'b0 ? 1'b0 : n5553;
/* FF 26 17  1 */ always @(posedge clk) if (n3249) n3547 <= 1'b0 ? 1'b0 : n5554;
/* FF 27 11  1 */ always @(posedge clk) if (n3460) n3619 <= 1'b0 ? 1'b0 : n5555;
/* FF  6 10  5 */ always @(posedge clk) if (n589) n596 <= 1'b0 ? 1'b0 : n5556;
/* FF 20 11  4 */ always @(posedge clk) if (n2682) n2692 <= 1'b0 ? 1'b0 : n5557;
/* FF 23 19  5 */ always @(posedge clk) if (n2573) n3255 <= 1'b0 ? 1'b0 : n5558;
/* FF  5 13  4 */ always @(posedge clk) if (n402) n496 <= 1'b0 ? 1'b0 : n5559;
/* FF 19 24  5 */ always @(posedge clk) if (n2775) n2599 <= 1'b0 ? 1'b0 : n5560;
/* FF 11 20  7 */ always @(posedge clk) if (n1339) n1195 <= 1'b0 ? 1'b0 : n5561;
/* FF 29  9  7 */ always @(posedge clk) if (n3464) n3832 <= 1'b0 ? 1'b0 : n5562;
/* FF 17 27  6 */ always @(posedge clk) if (n1) n2194 <= 1'b0 ? 1'b0 : n5563;
/* FF 28 23  3 */ always @(posedge clk) if (n3704) n3810 <= 1'b0 ? 1'b0 : n5564;
/* FF 11 27  6 */ always @(posedge clk) if (n1393) n1253 <= 1'b0 ? 1'b0 : n5565;
/* FF 21 26  3 */ assign n2970 = n5566;
/* FF 15 16  6 */ always @(posedge clk) if (n1500) n1799 <= 1'b0 ? 1'b0 : n5567;
/* FF 21 15  7 */ assign n2886 = n5568;
/* FF 15 15  7 */ assign n1791 = n5569;
/* FF  3 21  6 */ assign n352 = n5570;
/* FF 18 16  3 */ always @(posedge clk) if (n2540) n2317 <= 1'b0 ? 1'b0 : n5571;
/* FF  6  9  1 */ assign n5572 = n726;
/* FF 20 22  2 */ always @(posedge clk) if (n2384) n2778 <= 1'b0 ? 1'b0 : n5573;
/* FF 12 26  4 */ always @(posedge clk) if (n1393) n1389 <= 1'b0 ? 1'b0 : n5574;
/* FF 17 24  0 */ always @(posedge clk) if (n2000) n2166 <= 1'b0 ? 1'b0 : n5575;
/* FF 19  6  1 */ always @(posedge clk) if (n2241) n2444 <= 1'b0 ? 1'b0 : n5576;
/* FF  4  9  2 */ always @(posedge clk) if (n260) n373 <= 1'b0 ? 1'b0 : n5577;
/* FF 10  6  3 */ always @(posedge clk) if (en_in) n973 <= 1'b0 ? 1'b0 : n5578;
/* FF 24 15  2 */ always @(posedge clk) if (n3233) n3377 <= 1'b0 ? 1'b0 : n5579;
/* FF  9  9  6 */ always @(posedge clk) if (n983) n832 <= 1'b0 ? 1'b0 : n5580;
/* FF 13 11  5 */ always @(posedge clk) if (n1137) n1446 <= 1'b0 ? 1'b0 : n5581;
/* FF 18  2  0 */ always @(posedge clk) if (n2207) n2199 <= 1'b0 ? 1'b0 : n5582;
/* FF  7 17  2 */ always @(posedge clk) if (n549) n753 <= 1'b0 ? 1'b0 : n5583;
/* FF  9 22  4 */ always @(posedge clk) if (n819) n925 <= 1'b0 ? 1'b0 : n5584;
/* FF 18 15  7 */ always @(posedge clk) if (n1) n2314 <= 1'b0 ? 1'b0 : n5585;
/* FF 21 12  3 */ always @(posedge clk) if (n3029) n2870 <= 1'b0 ? 1'b0 : n5586;
/* FF 14 26  4 */ always @(posedge clk) if (n1271) n1715 <= 1'b0 ? 1'b0 : n5587;
/* FF 12 21  2 */ always @(posedge clk) if (n1205) n114 <= 1'b0 ? 1'b0 : n5588;
/* FF 14 15  3 */ always @(posedge clk) if (n1792) n1642 <= 1'b0 ? 1'b0 : n5589;
/* FF  2  9  0 */ always @(posedge clk) if (n153) n158 <= 1'b0 ? 1'b0 : n5590;
/* FF 20  4  2 */ assign \rco[98]  = n5591;
/* FF 19 20  0 */ always @(posedge clk) if (n2553) n2565 <= 1'b0 ? 1'b0 : n5592;
/* FF  9 32  2 */ assign \rco[109]  = n5593;
/* FF 23  9  4 */ always @(posedge clk) if (n2678) n3180 <= 1'b0 ? 1'b0 : n5594;
/* FF 22 19  6 */ assign n2757 = n5595;
/* FF 16 30  6 */ assign \rco[133]  = n5596;
/* FF 27  8  0 */ assign n3604 = n3733;
/* FF  3 17  3 */ always @(posedge clk) if (n79) n313 <= 1'b0 ? 1'b0 : n5597;
/* FF 14 25  6 */ always @(posedge clk) if (n697) n1707 <= 1'b0 ? 1'b0 : n5598;
/* FF  6 21  4 */ assign n5599 = n781;
/* FF 20 10  7 */ always @(posedge clk) if (n2697) n2285 <= 1'b0 ? 1'b0 : n5600;
/* FF 23 16  4 */ always @(posedge clk) if (n2540) n3232 <= 1'b0 ? 1'b0 : n5601;
/* FF 20  7  4 */ always @(posedge clk) if (n2670) n2665 <= 1'b0 ? 1'b0 : n5602;
/* FF  5 14  5 */ always @(posedge clk) if (n402) n500 <= 1'b0 ? 1'b0 : n5603;
/* FF 11 21  0 */ assign n1197 = n5604;
/* FF 29 10  6 */ always @(posedge clk) if (n3464) n3838 <= 1'b0 ? 1'b0 : n5605;
/* FF 28 22  0 */ always @(posedge clk) if (n3704) n3799 <= 1'b0 ? 1'b0 : n5606;
/* FF 16 12  3 */ always @(posedge clk) if (n1771) n1938 <= 1'b0 ? 1'b0 : n5607;
/* FF 11 24  7 */ always @(posedge clk) if (n796) n1230 <= 1'b0 ? 1'b0 : n5608;
/* FF 16 17  4 */ always @(posedge clk) if (n2110) n1967 <= 1'b0 ? 1'b0 : n5609;
/* FF 21 27  4 */ always @(posedge clk) if (n2196) n2976 <= 1'b0 ? 1'b0 : n5610;
/* FF 13 15  2 */ always @(posedge clk) if (n739) n1472 <= 1'b0 ? 1'b0 : n5611;
/* FF 30 12  6 */ always @(posedge clk) if (n3892) n3900 <= 1'b0 ? 1'b0 : n5612;
/* FF 15 17  1 */ always @(posedge clk) if (n1500) n1802 <= 1'b0 ? 1'b0 : n5613;
/* FF 18  6  5 */ always @(posedge clk) if (n2241) n2236 <= 1'b0 ? 1'b0 : n5614;
/* FF  7 21  7 */ always @(posedge clk) if (n360) n775 <= 1'b0 ? 1'b0 : n5615;
/* FF 18 19  2 */ always @(posedge clk) if (n1982) n2341 <= 1'b0 ? 1'b0 : n5616;
/* FF  3 18  7 */ always @(posedge clk) if (n215) n317 <= 1'b0 ? 1'b0 : n5617;
/* FF  6  8  2 */ always @(posedge clk) if (n570) n582 <= 1'b0 ? 1'b0 : n5618;
/* FF 20 21  3 */ always @(posedge clk) if (n2553) n2771 <= 1'b0 ? 1'b0 : n5619;
/* FF 12 25  5 */ always @(posedge clk) if (n1532) n1381 <= 1'b0 ? 1'b0 : n5620;
/* FF  1 19  3 */ always @(posedge clk) if (n119) n107 <= 1'b0 ? 1'b0 : n5621;
/* FF 17 25  3 */ always @(posedge clk) if (n2017) n2179 <= 1'b0 ? 1'b0 : n5622;
/* FF  5 16  1 */ always @(posedge clk) if (n511) n521 <= 1'b0 ? 1'b0 : n5623;
/* FF 19  7  2 */ always @(posedge clk) if (n2670) n2454 <= 1'b0 ? 1'b0 : n5624;
/* FF 23 13  1 */ always @(posedge clk) if (n3045) n3209 <= 1'b0 ? 1'b0 : n5625;
/* FF 10 25  2 */ always @(posedge clk) if (n567) n1082 <= 1'b0 ? 1'b0 : n5626;
/* FF 24 14  1 */ always @(posedge clk) if (n3376) n3370 <= 1'b0 ? 1'b0 : n5627;
/* FF 27 20  6 */ always @(posedge clk) if (n3424) n3681 <= 1'b0 ? 1'b0 : n5628;
/* FF  9 10  7 */ always @(posedge clk) if (n988) n841 <= 1'b0 ? 1'b0 : n5629;
/* FF 13 12  4 */ always @(posedge clk) if (n1137) n1453 <= 1'b0 ? 1'b0 : n5630;
/* FF 18  5  1 */ always @(posedge clk) if (n2230) n2222 <= 1'b0 ? 1'b0 : n5631;
/* FF  7 22  3 */ always @(posedge clk) if (n695) n786 <= 1'b0 ? 1'b0 : n5632;
/* FF  9 23  3 */ always @(posedge clk) if (n819) n928 <= 1'b0 ? 1'b0 : n5633;
/* FF 21 13  0 */ always @(posedge clk) if (n2519) n2874 <= 1'b0 ? 1'b0 : n5634;
/* FF 14 21  5 */ assign n1347 = n5635;
/* FF 19 30  6 */ always @(posedge clk) if (n2592) n2639 <= 1'b0 ? 1'b0 : n5636;
/* FF 17 11  0 */ assign n1602 = n5637;
/* FF  2  8  3 */ always @(posedge clk) if (n21) n157 <= 1'b0 ? 1'b0 : n5638;
/* FF  1 16  7 */ always @(posedge clk) if (n85) n94 <= 1'b0 ? 1'b0 : n5639;
/* FF 14 14  4 */ always @(posedge clk) if (n1791) n1636 <= 1'b0 ? 1'b0 : n5640;
/* FF 19 21  7 */ always @(posedge clk) if (n2164) n2583 <= 1'b0 ? 1'b0 : n5641;
/* FF 11 17  5 */ always @(posedge clk) if (n900) n1173 <= 1'b0 ? 1'b0 : n5642;
/* FF 10 11  5 */ always @(posedge clk) if (n996) n993 <= 1'b0 ? 1'b0 : n5643;
/* FF 23 14  5 */ always @(posedge clk) if (n2551) n3219 <= 1'b0 ? 1'b0 : n5644;
/* FF 24 17  5 */ always @(posedge clk) if (n2123) n3399 <= 1'b0 ? 1'b0 : n5645;
/* FF 28  7  6 */ always @(posedge clk) if (n3488) n3724 <= 1'b0 ? 1'b0 : n5646;
/* FF  3 14  1 */ assign n153 = n5647;
/* FF 15 21  6 */ always @(posedge clk) if (n1356) n1842 <= 1'b0 ? 1'b0 : n5648;
/* FF 12 10  2 */ always @(posedge clk) if (n850) n1285 <= 1'b0 ? 1'b0 : n5649;
/* FF 26 19  3 */ always @(posedge clk) if (n2730) n3558 <= 1'b0 ? 1'b0 : n5650;
/* FF 17  5  1 */ assign \rco[144]  = n5651;
/* FF 14 24  5 */ assign n1699 = n5652;
/* FF  6 20  7 */ always @(posedge clk) if (n552) n362 <= 1'b0 ? 1'b0 : n5653;
/* FF 20  9  6 */ assign n2680 = n5654;
/* FF 23 17  3 */ always @(posedge clk) if (n2540) n3235 <= 1'b0 ? 1'b0 : n5655;
/* FF  2  7  7 */ always @(posedge clk) if (n21) n152 <= 1'b0 ? 1'b0 : n5656;
/* FF 26  6  7 */ always @(posedge clk) if (n3459) n3480 <= 1'b0 ? 1'b0 : n5657;
/* FF 11 18  1 */ always @(posedge clk) if (n1187) n1180 <= 1'b0 ? 1'b0 : n5658;
/* FF 29 11  1 */ always @(posedge clk) if (n3751) n3840 <= 1'b0 ? 1'b0 : n5659;
/* FF 28 21  1 */ always @(posedge clk) if (n3788) n3792 <= 1'b0 ? 1'b0 : n5660;
/* FF  4 12  2 */ always @(posedge clk) if (n77) n395 <= 1'b0 ? 1'b0 : n5661;
/* FF 10 22  0 */ assign n819 = n5662;
/* FF 21 28  5 */ always @(posedge clk) if (n2196) n2984 <= 1'b0 ? 1'b0 : n5663;
/* FF 13 16  3 */ always @(posedge clk) if (n922) n1480 <= 1'b0 ? 1'b0 : n5664;
/* FF 27  7  0 */ assign n3331 = n5665;
/* FF 15 22  0 */ always @(posedge clk) if (n1835) n1846 <= 1'b0 ? 1'b0 : n5666;
/* FF 18  9  4 */ always @(posedge clk) if (n2055) n2265 <= 1'b0 ? 1'b0 : n5667;
/* FF 18 18  5 */ always @(posedge clk) if (n1825) n1047 <= 1'b0 ? 1'b0 : n5668;
/* FF  3 19  4 */ always @(posedge clk) if (n115) n331 <= 1'b0 ? 1'b0 : n5669;
/* FF  6 11  3 */ always @(posedge clk) if (n286) n602 <= 1'b0 ? 1'b0 : n5670;
/* FF 12 24  2 */ always @(posedge clk) if (n961) n1369 <= 1'b0 ? 1'b0 : n5671;
/* FF 14 10  1 */ always @(posedge clk) if (n1622) n1605 <= 1'b0 ? 1'b0 : n5672;
/* FF 19 17  4 */ always @(posedge clk) if (n2727) n2545 <= 1'b0 ? 1'b0 : n5673;
/* FF 22 21  7 */ always @(posedge clk) if (n2564) n3103 <= 1'b0 ? 1'b0 : n5674;
/* FF 24 24  7 */ always @(posedge clk) if (n3112) n3445 <= 1'b0 ? 1'b0 : n5675;
/* FF  5 17  2 */ always @(posedge clk) if (n2) n526 <= 1'b0 ? 1'b0 : n5676;
/* FF  4 15  4 */ always @(posedge clk) if (n207) n416 <= 1'b0 ? 1'b0 : n5677;
/* FF 10 24  1 */ always @(posedge clk) if (n820) n1073 <= 1'b0 ? 1'b0 : n5678;
/* FF 24 13  0 */ always @(posedge clk) if (n3351) n3361 <= 1'b0 ? 1'b0 : n5679;
/* FF 28 11  5 */ assign n5680 = n3848;
/* FF 27 21  1 */ always @(posedge clk) if (n3421) n3688 <= 1'b0 ? 1'b0 : n5681;
/* FF 18  4  2 */ always @(posedge clk) if (n2207) n2215 <= 1'b0 ? 1'b0 : n5682;
/* FF  7 23  0 */ always @(posedge clk) if (n454) n790 <= 1'b0 ? 1'b0 : n5683;
/* FF  9 16  2 */ always @(posedge clk) if (n645) n877 <= 1'b0 ? 1'b0 : n5684;
/* FF 21 14  1 */ always @(posedge clk) if (n2519) n2883 <= 1'b0 ? 1'b0 : n5685;
/* FF 14 20  6 */ always @(posedge clk) if (n1347) n1681 <= 1'b0 ? 1'b0 : n5686;
/* FF  5  8  6 */ always @(posedge clk) if (n21) n472 <= 1'b0 ? 1'b0 : n5687;
/* FF 17 20  1 */ always @(posedge clk) if (n1843) n2137 <= 1'b0 ? 1'b0 : n5688;
/* FF  2 11  2 */ always @(posedge clk) if (n168) n170 <= 1'b0 ? 1'b0 : n5689;
/* FF 19 31  5 */ always @(posedge clk) if (n2592) n2646 <= 1'b0 ? 1'b0 : n5690;
/* FF 19 18  6 */ always @(posedge clk) if (n2348) n2560 <= 1'b0 ? 1'b0 : n5691;
/* FF 10 10  2 */ always @(posedge clk) if (n983) n985 <= 1'b0 ? 1'b0 : n5692;
/* FF 23 15  6 */ always @(posedge clk) if (n3216) n3228 <= 1'b0 ? 1'b0 : n5693;
/* FF 28  6  5 */ always @(posedge clk) if (n3594) n3456 <= 1'b0 ? 1'b0 : n5694;
/* FF  3 15  2 */ always @(posedge clk) if (n207) n295 <= 1'b0 ? 1'b0 : n5695;
/* FF 21 16  0 */ always @(posedge clk) if (n2551) n2887 <= 1'b0 ? 1'b0 : n5696;
/* FF 26 18  4 */ assign \rco[33]  = n5697;
/* FF 12  9  3 */ always @(posedge clk) if (n850) n1283 <= 1'b0 ? 1'b0 : n5698;
/* FF 18 22  2 */ assign n1998 = n2590;
/* FF 17  6  0 */ always @(posedge clk) if (n2045) n2038 <= 1'b0 ? 1'b0 : n5699;
/* FF  6 23  6 */ always @(posedge clk) if (n360) n693 <= 1'b0 ? 1'b0 : n5700;
/* FF 20  8  1 */ always @(posedge clk) if (n2247) n2669 <= 1'b0 ? 1'b0 : n5701;
/* FF 12 28  7 */ always @(posedge clk) if (n1394) n1401 <= 1'b0 ? 1'b0 : n5702;
/* FF 23 22  2 */ always @(posedge clk) if (n3422) n3281 <= 1'b0 ? 1'b0 : n5703;
/* FF 29 12  0 */ always @(posedge clk) if (n3751) n3849 <= 1'b0 ? 1'b0 : n5704;
/* FF 16 10  1 */ always @(posedge clk) if (n1771) n1927 <= 1'b0 ? 1'b0 : n5705;
/* FF 22 26  3 */ always @(posedge clk) if (n2613) n3136 <= 1'b0 ? 1'b0 : n5706;
/* FF 27 17  6 */ always @(posedge clk) if (n3249) n3655 <= 1'b0 ? 1'b0 : n5707;
/* FF 13 17  0 */ always @(posedge clk) if (n1461) n1484 <= 1'b0 ? 1'b0 : n5708;
/* FF 15 23  3 */ always @(posedge clk) if (n778) n1855 <= 1'b0 ? 1'b0 : n5709;
/* FF 18  8  7 */ always @(posedge clk) if (n2055) n2256 <= 1'b0 ? 1'b0 : n5710;
/* FF 18 21  4 */ always @(posedge clk) if (n2347) n2353 <= 1'b0 ? 1'b0 : n5711;
/* FF  3 16  5 */ always @(posedge clk) if (n197) n307 <= 1'b0 ? 1'b0 : n5712;
/* FF 14  5  0 */ always @(posedge clk) if (n1577) n1571 <= 1'b0 ? 1'b0 : n5713;
/* FF 19 14  5 */ always @(posedge clk) if (n2123) n2516 <= 1'b0 ? 1'b0 : n5714;
/* FF 22 20  4 */ always @(posedge clk) if (n3087) n3092 <= 1'b0 ? 1'b0 : n5715;
/* FF 10 14  7 */ always @(posedge clk) if (n750) n1014 <= 1'b0 ? 1'b0 : n5716;
/* FF  5 18  3 */ always @(posedge clk) if (n657) n534 <= 1'b0 ? 1'b0 : n5717;
/* FF  4 14  7 */ always @(posedge clk) if (n79) n409 <= 1'b0 ? 1'b0 : n5718;
/* FF 19  5  4 */ always @(posedge clk) if (n2230) n2439 <= 1'b0 ? 1'b0 : n5719;
/* FF 10 27  0 */ always @(posedge clk) if (n804) n1093 <= 1'b0 ? 1'b0 : n5720;
/* FF 22 25  7 */ always @(posedge clk) if (n2812) n3131 <= 1'b0 ? 1'b0 : n5721;
/* FF 27 18  0 */ always @(posedge clk) if (n3553) n3657 <= 1'b0 ? 1'b0 : n5722;
/* FF 24 12  7 */ always @(posedge clk) if (n3351) n3360 <= 1'b0 ? 1'b0 : n5723;
/* FF 28 10  6 */ always @(posedge clk) if (n3462) n3747 <= 1'b0 ? 1'b0 : n5724;
/* FF 13 14  6 */ always @(posedge clk) if (n1461) n1468 <= 1'b0 ? 1'b0 : n5725;
/* FF 18  7  3 */ assign \rco[96]  = n5726;
/* FF  9 17  1 */ always @(posedge clk) if (n1030) n884 <= 1'b0 ? 1'b0 : n5727;
/* FF 26 22  1 */ always @(posedge clk) if (n2730) n3570 <= 1'b0 ? 1'b0 : n5728;
/* FF 15  5  3 */ always @(posedge clk) if (n1742) n1728 <= 1'b0 ? 1'b0 : n5729;
/* FF 14 23  7 */ assign n1375 = n5730;
/* FF 20 12  6 */ always @(posedge clk) if (n2682) n2704 <= 1'b0 ? 1'b0 : n5731;
/* FF 14  8  6 */ always @(posedge clk) if (n1741) n1599 <= 1'b0 ? 1'b0 : n5732;
/* FF 17 21  2 */ always @(posedge clk) if (n2347) n2146 <= 1'b0 ? 1'b0 : n5733;
/* FF 19 19  5 */ assign n2553 = n5734;
/* FF 10 13  3 */ always @(posedge clk) if (n629) n1004 <= 1'b0 ? 1'b0 : n5735;
/* FF 24 26  0 */ always @(posedge clk) if (n2613) n3454 <= 1'b0 ? 1'b0 : n5736;
/* FF 23 12  7 */ always @(posedge clk) if (n3031) n3206 <= 1'b0 ? 1'b0 : n5737;
/* FF 28  5  4 */ always @(posedge clk) if (n3488) n3709 <= 1'b0 ? 1'b0 : n5738;
/* FF 16 27  1 */ always @(posedge clk) if (n1) n1311 <= 1'b0 ? 1'b0 : n5739;
/* FF  3 12  3 */ always @(posedge clk) if (n168) n280 <= 1'b0 ? 1'b0 : n5740;
/* FF  7 10  0 */ always @(posedge clk) if (n589) n729 <= 1'b0 ? 1'b0 : n5741;
/* FF 21 17  3 */ assign \rco[65]  = n5742;
/* FF 30 10  5 */ always @(posedge clk) if (n3892) n3463 <= 1'b0 ? 1'b0 : n5743;
/* FF 15 11  4 */ always @(posedge clk) if (n1624) n1767 <= 1'b0 ? 1'b0 : n5744;
/* FF 12  8  4 */ always @(posedge clk) if (n1131) n1280 <= 1'b0 ? 1'b0 : n5745;
/* FF 26 21  5 */ always @(posedge clk) if (n3421) n3240 <= 1'b0 ? 1'b0 : n5746;
/* FF 15  6  7 */ always @(posedge clk) if (n1744) n1740 <= 1'b0 ? 1'b0 : n5747;
/* FF 17  7  7 */ always @(posedge clk) if (n2045) n2053 <= 1'b0 ? 1'b0 : n5748;
/* FF 18 25  3 */ always @(posedge clk) if (n1878) n2380 <= 1'b0 ? 1'b0 : n5749;
/* FF  6 22  1 */ always @(posedge clk) if (n673) n679 <= 1'b0 ? 1'b0 : n5750;
/* FF 20 15  0 */ always @(posedge clk) if (n2715) n2717 <= 1'b0 ? 1'b0 : n5751;
/* FF 23 23  1 */ always @(posedge clk) if (n3104) n3288 <= 1'b0 ? 1'b0 : n5752;
/* FF 11 16  3 */ always @(posedge clk) if (n891) n1162 <= 1'b0 ? 1'b0 : n5753;
/* FF 16  9  0 */ always @(posedge clk) if (n1771) n1923 <= 1'b0 ? 1'b0 : n5754;
/* FF  1 12  1 */ always @(posedge clk) if (n39) n47 <= 1'b0 ? 1'b0 : n5755;
/* FF 13  7  6 */ always @(posedge clk) if (n977) n1429 <= 1'b0 ? 1'b0 : n5756;
/* FF  7  7  6 */ always @(posedge clk) if (n588) n715 <= 1'b0 ? 1'b0 : n5757;
/* FF 13 18  1 */ always @(posedge clk) if (n1205) n1493 <= 1'b0 ? 1'b0 : n5758;
/* FF 27  5  6 */ always @(posedge clk) if (n3594) n3591 <= 1'b0 ? 1'b0 : n5759;
/* FF 18 11  6 */ assign n2230 = n5760;
/* FF 15 20  2 */ always @(posedge clk) if (n1347) n1829 <= 1'b0 ? 1'b0 : n5761;
/* FF 18 20  7 */ assign n2347 = n5762;
/* FF 12 30  0 */ always @(posedge clk) if (n1394) n1407 <= 1'b0 ? 1'b0 : n5763;
/* FF 26  7  1 */ always @(posedge clk) if (n3603) n3482 <= 1'b0 ? 1'b0 : n5764;
/* FF  2 14  2 */ always @(posedge clk) if (n83) n189 <= 1'b0 ? 1'b0 : n5765;
/* FF 16  7  3 */ always @(posedge clk) if (n1743) n1910 <= 1'b0 ? 1'b0 : n5766;
/* FF 19 15  6 */ always @(posedge clk) if (n2715) n2531 <= 1'b0 ? 1'b0 : n5767;
/* FF 23  5  5 */ always @(posedge clk) if (n3158) n3155 <= 1'b0 ? 1'b0 : n5768;
/* FF 22 23  5 */ always @(posedge clk) if (n3104) n2539 <= 1'b0 ? 1'b0 : n5769;
/* FF 24 22  5 */ always @(posedge clk) if (n3422) n2934 <= 1'b0 ? 1'b0 : n5770;
/* FF  5 19  4 */ always @(posedge clk) if (n349) n543 <= 1'b0 ? 1'b0 : n5771;
/* FF  4 13  6 */ assign n76 = n5772;
/* FF 22 24  4 */ always @(posedge clk) if (n3113) n3120 <= 1'b0 ? 1'b0 : n5773;
/* FF 10 26  7 */ assign n1091 = n5774;
/* FF 24 11  6 */ assign \rco[66]  = n3468;
/* FF 28  9  7 */ always @(posedge clk) if (n3621) n3740 <= 1'b0 ? 1'b0 : n5775;
/* FF 27 19  3 */ always @(posedge clk) if (n3553) n3670 <= 1'b0 ? 1'b0 : n5776;
/* FF  9 18  0 */ always @(posedge clk) if (n1030) n892 <= 1'b0 ? 1'b0 : n5777;
/* FF 26  9  0 */ always @(posedge clk) if (n3460) n3498 <= 1'b0 ? 1'b0 : n5778;
/* FF 29 17  1 */ always @(posedge clk) if (n3765) n3857 <= 1'b0 ? 1'b0 : n5779;
/* FF 14 22  0 */ always @(posedge clk) if (n1402) n1687 <= 1'b0 ? 1'b0 : n5780;
/* FF 17  3  4 */ always @(posedge clk) if (n1887) n2029 <= 1'b0 ? 1'b0 : n5781;
/* FF  6 18  6 */ always @(posedge clk) if (n657) n655 <= 1'b0 ? 1'b0 : n5782;
/* FF  5 10  4 */ always @(posedge clk) if (n184) n478 <= 1'b0 ? 1'b0 : n5783;
/* FF 14 11  7 */ always @(posedge clk) if (n1622) n1618 <= 1'b0 ? 1'b0 : n5784;
/* FF 17 22  3 */ always @(posedge clk) if (n1999) n2155 <= 1'b0 ? 1'b0 : n5785;
/* FF 19 29  3 */ always @(posedge clk) if (n2614) n2630 <= 1'b0 ? 1'b0 : n5786;
/* FF 19 16  4 */ always @(posedge clk) if (n2730) n2537 <= 1'b0 ? 1'b0 : n5787;
/* FF 23  6  1 */ always @(posedge clk) if (n3158) n3160 <= 1'b0 ? 1'b0 : n5788;
/* FF 11 28  6 */ always @(posedge clk) if (n1384) n1261 <= 1'b0 ? 1'b0 : n5789;
/* FF 10 12  0 */ always @(posedge clk) if (n996) n997 <= 1'b0 ? 1'b0 : n5790;
/* FF 24 25  1 */ always @(posedge clk) if (n2812) n3447 <= 1'b0 ? 1'b0 : n5791;
/* FF  3 13  4 */ assign \rco[16]  = n407;
/* FF 22 10  0 */ always @(posedge clk) if (n2856) n3022 <= 1'b0 ? 1'b0 : n5792;
/* FF  9 28  3 */ always @(posedge clk) if (n961) n959 <= 1'b0 ? 1'b0 : n5793;
/* FF 21 18  2 */ always @(posedge clk) if (n2757) n2904 <= 1'b0 ? 1'b0 : n5794;
/* FF 15  8  5 */ always @(posedge clk) if (n1741) n1750 <= 1'b0 ? 1'b0 : n5795;
/* FF  3 22  6 */ always @(posedge clk) if (n352) n358 <= 1'b0 ? 1'b0 : n5796;
/* FF 12 15  5 */ always @(posedge clk) if (n1155) n1301 <= 1'b0 ? 1'b0 : n5797;
/* FF 26 20  6 */ assign n1710 = n3686;
/* FF 15  7  4 */ assign n1742 = n5798;
/* FF 18 24  0 */ always @(posedge clk) if (n1878) n2370 <= 1'b0 ? 1'b0 : n5799;
/* FF  6 17  0 */ always @(posedge clk) if (n549) n646 <= 1'b0 ? 1'b0 : n5800;
/* FF 23 20  0 */ always @(posedge clk) if (n3258) n3263 <= 1'b0 ? 1'b0 : n5801;
/* FF  1 13  2 */ always @(posedge clk) if (n83) n61 <= 1'b0 ? 1'b0 : n5802;
/* FF 24  7  5 */ assign n3006 = n5803;
/* FF  9 14  6 */ always @(posedge clk) if (n629) n865 <= 1'b0 ? 1'b0 : n5804;
/* FF 13 19  6 */ assign \rco[99]  = n1675;
/* FF 18 10  1 */ always @(posedge clk) if (n2282) n2274 <= 1'b0 ? 1'b0 : n5805;
/* FF 20 28  0 */ assign n2196 = n5806;
/* FF 18 23  6 */ always @(posedge clk) if (n1999) n2367 <= 1'b0 ? 1'b0 : n5807;
/* FF 12 29  1 */ always @(posedge clk) if (n1532) n1404 <= 1'b0 ? 1'b0 : n5808;
/* FF 14  7  2 */ always @(posedge clk) if (n1743) n1587 <= 1'b0 ? 1'b0 : n5809;
/* FF 16  6  0 */ always @(posedge clk) if (n1744) n1897 <= 1'b0 ? 1'b0 : n5810;
/* FF 19 12  7 */ always @(posedge clk) if (n1936) n2504 <= 1'b0 ? 1'b0 : n5811;
/* FF 23 10  4 */ always @(posedge clk) if (n2697) n3187 <= 1'b0 ? 1'b0 : n5812;
/* FF 22 22  2 */ always @(posedge clk) if (n2961) n3107 <= 1'b0 ? 1'b0 : n5813;
/* FF 24 21  4 */ always @(posedge clk) if (n3411) n3423 <= 1'b0 ? 1'b0 : n5814;
/* FF 19  3  6 */ always @(posedge clk) if (n1887) n2433 <= 1'b0 ? 1'b0 : n5815;
/* FF 22 27  5 */ always @(posedge clk) if (n2970) n3148 <= 1'b0 ? 1'b0 : n5816;
/* FF 24 10  5 */ always @(posedge clk) if (n3352) n3345 <= 1'b0 ? 1'b0 : n5817;
/* FF 28  8  0 */ always @(posedge clk) if (n3605) n3726 <= 1'b0 ? 1'b0 : n5818;
/* FF  3  9  1 */ always @(posedge clk) if (n260) n253 <= 1'b0 ? 1'b0 : n5819;
/* FF 12 19  0 */ always @(posedge clk) if (n1501) n1328 <= 1'b0 ? 1'b0 : n5820;
/* FF 26  8  3 */ always @(posedge clk) if (n3603) n3493 <= 1'b0 ? 1'b0 : n5821;
/* FF 14 17  1 */ always @(posedge clk) if (n1672) n1655 <= 1'b0 ? 1'b0 : n5822;
/* FF 17 12  5 */ always @(posedge clk) if (n2056) n2082 <= 1'b0 ? 1'b0 : n5823;
/* FF 19 26  2 */ assign n2612 = n5824;
/* FF 17 23  4 */ always @(posedge clk) if (n1069) n2163 <= 1'b0 ? 1'b0 : n5825;
/* FF  2 12  7 */ always @(posedge clk) if (n39) n183 <= 1'b0 ? 1'b0 : n5826;
/* FF 23  7  2 */ always @(posedge clk) if (n3006) n3168 <= 1'b0 ? 1'b0 : n5827;
/* FF 11 29  1 */ assign \rco[101]  = n5828;
/* FF 10 15  1 */ always @(posedge clk) if (n750) n1016 <= 1'b0 ? 1'b0 : n5829;
/* FF 16 25  3 */ always @(posedge clk) if (n1557) n2006 <= 1'b0 ? 1'b0 : n5830;
/* FF 21 24  4 */ always @(posedge clk) if (n3113) n2957 <= 1'b0 ? 1'b0 : n5831;
/* FF  3 10  5 */ always @(posedge clk) if (n251) n267 <= 1'b0 ? 1'b0 : n5832;
/* FF 21 19  5 */ always @(posedge clk) if (n2757) n2915 <= 1'b0 ? 1'b0 : n5833;
/* FF 13 23  3 */ always @(posedge clk) if (n1069) n1527 <= 1'b0 ? 1'b0 : n5834;
/* FF 27 14  2 */ always @(posedge clk) if (n3527) n3643 <= 1'b0 ? 1'b0 : n5835;
/* FF 18 14  6 */ assign \rco[34]  = n5836;
/* FF 12 14  6 */ always @(posedge clk) if (n1154) n1294 <= 1'b0 ? 1'b0 : n5837;
/* FF 26 23  7 */ always @(posedge clk) if (n3703) n3582 <= 1'b0 ? 1'b0 : n5838;
/* FF 18 27  1 */ always @(posedge clk) if (n2020) n2394 <= 1'b0 ? 1'b0 : n5839;
/* FF  6 16  3 */ always @(posedge clk) if (n511) n641 <= 1'b0 ? 1'b0 : n5840;
/* FF 20 13  2 */ assign n2306 = n2881;
/* FF  4 11  7 */ always @(posedge clk) if (n184) n392 <= 1'b0 ? 1'b0 : n5841;
/* FF 22 18  7 */ always @(posedge clk) if (n3065) n3086 <= 1'b0 ? 1'b0 : n5842;
/* FF  1 14  3 */ always @(posedge clk) if (n85) n71 <= 1'b0 ? 1'b0 : n5843;
/* FF 22  7  0 */ always @(posedge clk) if (n2841) n2998 <= 1'b0 ? 1'b0 : n5844;
/* FF 10 17  5 */ assign n5845 = n1177;
/* FF  9 15  1 */ always @(posedge clk) if (n645) n868 <= 1'b0 ? 1'b0 : n5846;
/* FF 13  9  4 */ always @(posedge clk) if (n850) n1433 <= 1'b0 ? 1'b0 : n5847;
/* FF 24  6  6 */ always @(posedge clk) if (n3006) n3327 <= 1'b0 ? 1'b0 : n5848;
/* FF 28 12  5 */ always @(posedge clk) if (n3462) n3758 <= 1'b0 ? 1'b0 : n5849;
/* FF 13 20  7 */ always @(posedge clk) if (n1339) n1204 <= 1'b0 ? 1'b0 : n5850;
/* FF 18 13  0 */ always @(posedge clk) if (n2283) n2295 <= 1'b0 ? 1'b0 : n5851;
/* FF 20 19  1 */ always @(posedge clk) if (n2562) n2750 <= 1'b0 ? 1'b0 : n5852;
/* FF 14  6  5 */ always @(posedge clk) if (n1577) n1580 <= 1'b0 ? 1'b0 : n5853;
/* FF 16  5  1 */ always @(posedge clk) if (n1742) n1889 <= 1'b0 ? 1'b0 : n5854;
/* FF 17 19  1 */ always @(posedge clk) if (n1982) n2129 <= 1'b0 ? 1'b0 : n5855;
/* FF 23 11  7 */ always @(posedge clk) if (n3031) n3197 <= 1'b0 ? 1'b0 : n5856;
/* FF 22 17  3 */ always @(posedge clk) if (n3065) n3075 <= 1'b0 ? 1'b0 : n5857;
/* FF 24 20  3 */ always @(posedge clk) if (n3411) n3415 <= 1'b0 ? 1'b0 : n5858;
/* FF 10 28  5 */ always @(posedge clk) if (n821) n1106 <= 1'b0 ? 1'b0 : n5859;
/* FF 24  9  4 */ always @(posedge clk) if (n3352) n3336 <= 1'b0 ? 1'b0 : n5860;
/* FF 13  6  2 */ always @(posedge clk) if (n977) n1417 <= 1'b0 ? 1'b0 : n5861;
/* FF 28 15  1 */ always @(posedge clk) if (n3233) n3391 <= 1'b0 ? 1'b0 : n5862;
/* FF 15 24  3 */ always @(posedge clk) if (n778) n1867 <= 1'b0 ? 1'b0 : n5863;
/* FF 21 23  2 */ always @(posedge clk) if (n2961) n2945 <= 1'b0 ? 1'b0 : n5864;
/* FF 26 11  2 */ assign \rco[69]  = n5865;
/* FF 12 18  3 */ always @(posedge clk) if (n1501) n1323 <= 1'b0 ? 1'b0 : n5866;
/* FF 29 19  7 */ always @(posedge clk) if (n3786) n3867 <= 1'b0 ? 1'b0 : n5867;
/* FF 14 16  2 */ always @(posedge clk) if (n1792) n1648 <= 1'b0 ? 1'b0 : n5868;
/* FF 17 13  6 */ always @(posedge clk) if (n2056) n2092 <= 1'b0 ? 1'b0 : n5869;
/* FF  5 12  2 */ always @(posedge clk) if (n77) n486 <= 1'b0 ? 1'b0 : n5870;
/* FF 17 16  5 */ assign n2112 = n2324;
/* FF  2 15  6 */ always @(posedge clk) if (n197) n201 <= 1'b0 ? 1'b0 : n5871;
/* FF 19 27  1 */ always @(posedge clk) if (n2614) n2617 <= 1'b0 ? 1'b0 : n5872;
/* FF 11 26  0 */ always @(posedge clk) if (n954) n1236 <= 1'b0 ? 1'b0 : n5873;
/* FF 21 25  7 */ always @(posedge clk) if (n2970) n2969 <= 1'b0 ? 1'b0 : n5874;
/* FF  9 11  6 */ always @(posedge clk) if (n988) n848 <= 1'b0 ? 1'b0 : n5875;
/* FF  3 11  6 */ always @(posedge clk) if (n153) n275 <= 1'b0 ? 1'b0 : n5876;
/* FF  7  9  5 */ always @(posedge clk) if (n589) n723 <= 1'b0 ? 1'b0 : n5877;
/* FF 21 20  4 */ always @(posedge clk) if (n3087) n2922 <= 1'b0 ? 1'b0 : n5878;
/* FF 13 24  2 */ assign n1357 = n5879;
/* FF 31 21  4 */ assign \rco[186]  = n5880;
/* FF 27 15  1 */ always @(posedge clk) if (n3233) n3649 <= 1'b0 ? 1'b0 : n5881;
/* FF 15 14  3 */ always @(posedge clk) if (n1791) n1786 <= 1'b0 ? 1'b0 : n5882;
/* FF  3 20  4 */ always @(posedge clk) if (n119) n346 <= 1'b0 ? 1'b0 : n5883;
/* FF 18 17  7 */ always @(posedge clk) if (n1825) n2332 <= 1'b0 ? 1'b0 : n5884;
/* FF 18 26  6 */ always @(posedge clk) if (n2615) n2391 <= 1'b0 ? 1'b0 : n5885;
/* FF  6 19  2 */ assign n657 = n5886;
/* FF 28 19  3 */ always @(posedge clk) if (n3424) n3780 <= 1'b0 ? 1'b0 : n5887;
/* FF 19  9  5 */ always @(posedge clk) if (n2451) n2476 <= 1'b0 ? 1'b0 : n5888;
/* FF  4 10  4 */ always @(posedge clk) if (n251) n383 <= 1'b0 ? 1'b0 : n5889;
/* FF  1 15  4 */ always @(posedge clk) if (n85) n86 <= 1'b0 ? 1'b0 : n5890;
/* FF 22  6  7 */ always @(posedge clk) if (n2841) n2997 <= 1'b0 ? 1'b0 : n5891;
/* FF 10 16  6 */ always @(posedge clk) if (n891) n1028 <= 1'b0 ? 1'b0 : n5892;
/* FF 13 10  5 */ always @(posedge clk) if (n850) n206 <= 1'b0 ? 1'b0 : n5893;
/* FF 13 21  4 */ always @(posedge clk) if (n1356) n1517 <= 1'b0 ? 1'b0 : n5894;
/* FF 18 12  3 */ always @(posedge clk) if (n1936) n2289 <= 1'b0 ? 1'b0 : n5895;
/* FF 21  6  0 */ always @(posedge clk) if (n2247) n2833 <= 1'b0 ? 1'b0 : n5896;
/* FF  6 13  1 */ always @(posedge clk) if (n78) n616 <= 1'b0 ? 1'b0 : n5897;
/* FF 20 18  2 */ always @(posedge clk) if (n2348) n2743 <= 1'b0 ? 1'b0 : n5898;
/* FF 11  6  2 */ always @(posedge clk) if (en_in) n1120 <= 1'b0 ? 1'b0 : n5899;
/* FF 14 12  7 */ always @(posedge clk) if (n1137) n1619 <= 1'b0 ? 1'b0 : n5900;
/* FF 29  2  3 */ assign \rco[50]  = n5901;
/* FF 19 10  1 */ always @(posedge clk) if (n2678) n2480 <= 1'b0 ? 1'b0 : n5902;
/* FF 22 16  0 */ always @(posedge clk) if (n2551) n3070 <= 1'b0 ? 1'b0 : n5903;
/* FF  5 22  7 */ always @(posedge clk) if (n673) n561 <= 1'b0 ? 1'b0 : n5904;
/* FF 28 14  2 */ always @(posedge clk) if (n2085) n3763 <= 1'b0 ? 1'b0 : n5905;
/* FF 15 25  4 */ assign \rco[191]  = n5906;
/* FF  7 13  2 */ assign \rco[156]  = n5907;
/* FF 21  8  3 */ always @(posedge clk) if (n2989) n2843 <= 1'b0 ? 1'b0 : n5908;
/* FF 26 17  4 */ always @(posedge clk) if (n3249) n3550 <= 1'b0 ? 1'b0 : n5909;
/* FF 12 17  2 */ always @(posedge clk) if (n900) n1314 <= 1'b0 ? 1'b0 : n5910;
/* FF 26 10  5 */ always @(posedge clk) if (n3033) n3510 <= 1'b0 ? 1'b0 : n5911;
/* FF 18 30  3 */ always @(posedge clk) if (n1881) n2420 <= 1'b0 ? 1'b0 : n5912;
/* FF 14 19  3 */ assign n777 = n5913;
/* FF 17 14  7 */ always @(posedge clk) if (n1625) n1631 <= 1'b0 ? 1'b0 : n5914;
/* FF 29 20  6 */ always @(posedge clk) if (n3786) n3874 <= 1'b0 ? 1'b0 : n5915;
/* FF  5 13  1 */ always @(posedge clk) if (n402) n493 <= 1'b0 ? 1'b0 : n5916;
/* FF 17 17  6 */ always @(posedge clk) if (n2111) n2120 <= 1'b0 ? 1'b0 : n5917;
/* FF 19 24  0 */ always @(posedge clk) if (n2775) n2594 <= 1'b0 ? 1'b0 : n5918;
/* FF 11 27  3 */ always @(posedge clk) if (n1393) n1250 <= 1'b0 ? 1'b0 : n5919;
/* FF  1 11  1 */ assign \rco[3]  = n175;
/* FF 21 26  6 */ assign n982 = n3142;
/* FF 21 21  7 */ always @(posedge clk) if (n2564) n2933 <= 1'b0 ? 1'b0 : n5920;
/* FF 13 25  1 */ always @(posedge clk) if (n697) n1535 <= 1'b0 ? 1'b0 : n5921;
/* FF 27 12  0 */ always @(posedge clk) if (n3368) n3629 <= 1'b0 ? 1'b0 : n5922;
/* FF 18 16  4 */ always @(posedge clk) if (n2540) n2318 <= 1'b0 ? 1'b0 : n5923;
/* FF  3 21  3 */ assign n5924 = n460;
/* FF 18 29  7 */ always @(posedge clk) if (n1881) n2415 <= 1'b0 ? 1'b0 : n5925;
/* FF 11  9  0 */ assign n1131 = n5926;
/* FF 28 18  0 */ assign n3765 = n5927;
/* FF 19  6  4 */ always @(posedge clk) if (n2241) n2447 <= 1'b0 ? 1'b0 : n5928;
/* FF  4  9  5 */ always @(posedge clk) if (n260) n376 <= 1'b0 ? 1'b0 : n5929;
/* FF  9  9  3 */ always @(posedge clk) if (n983) n830 <= 1'b0 ? 1'b0 : n5930;
/* FF 16 32  6 */ assign \rco[58]  = n5931;
/* FF 13 11  2 */ always @(posedge clk) if (n1137) n1443 <= 1'b0 ? 1'b0 : n5932;
/* FF 13 22  5 */ assign n1521 = n5933;
/* FF 18 15  2 */ always @(posedge clk) if (n1) n2310 <= 1'b0 ? 1'b0 : n5934;
/* FF  6 12  2 */ always @(posedge clk) if (n286) n608 <= 1'b0 ? 1'b0 : n5935;
/* FF 20 17  3 */ always @(posedge clk) if (n2727) n2735 <= 1'b0 ? 1'b0 : n5936;
/* FF 26 14  2 */ always @(posedge clk) if (n3527) n3535 <= 1'b0 ? 1'b0 : n5937;
/* FF 14 15  6 */ always @(posedge clk) if (n1792) n1644 <= 1'b0 ? 1'b0 : n5938;
/* FF  2  9  7 */ always @(posedge clk) if (n153) n164 <= 1'b0 ? 1'b0 : n5939;
/* FF 20  4  7 */ always @(posedge clk) if (n1761) n2220 <= 1'b0 ? 1'b0 : n5940;
/* FF 17 29  3 */ assign \rco[54]  = n5941;
/* FF 16  3  7 */ assign \rco[91]  = n5942;
/* FF 19 11  2 */ always @(posedge clk) if (n2076) n2488 <= 1'b0 ? 1'b0 : n5943;
/* FF 23  9  1 */ always @(posedge clk) if (n2678) n3177 <= 1'b0 ? 1'b0 : n5944;
/* FF 22 19  1 */ assign n5945 = n3260;
/* FF 10  5  2 */ always @(posedge clk) if (en_in) n968 <= 1'b0 ? 1'b0 : n5946;
/* FF 24 18  1 */ always @(posedge clk) if (n3411) n3403 <= 1'b0 ? 1'b0 : n5947;
/* FF  4 20  0 */ assign n439 = n5948;
/* FF 21  9  0 */ always @(posedge clk) if (n2856) n2845 <= 1'b0 ? 1'b0 : n5949;
/* FF  9 27  3 */ always @(posedge clk) if (n804) n949 <= 1'b0 ? 1'b0 : n5950;
/* FF 12 16  5 */ always @(posedge clk) if (n1155) n737 <= 1'b0 ? 1'b0 : n5951;
/* FF 26 13  4 */ always @(posedge clk) if (n3033) n3529 <= 1'b0 ? 1'b0 : n5952;
/* FF 29 21  5 */ always @(posedge clk) if (n3788) n2942 <= 1'b0 ? 1'b0 : n5953;
/* FF 17 15  0 */ always @(posedge clk) if (n2111) n2101 <= 1'b0 ? 1'b0 : n5954;
/* FF 20  7  3 */ always @(posedge clk) if (n2670) n2664 <= 1'b0 ? 1'b0 : n5955;
/* FF  5 14  0 */ always @(posedge clk) if (n402) n504 <= 1'b0 ? 1'b0 : n5956;
/* FF 11 24  2 */ always @(posedge clk) if (n796) n1225 <= 1'b0 ? 1'b0 : n5957;
/* FF 22 13  5 */ always @(posedge clk) if (n2085) n3048 <= 1'b0 ? 1'b0 : n5958;
/* FF 21 27  1 */ always @(posedge clk) if (n2196) n2973 <= 1'b0 ? 1'b0 : n5959;
/* FF 13 15  7 */ always @(posedge clk) if (n739) n1167 <= 1'b0 ? 1'b0 : n5960;
/* FF 27  6  6 */ always @(posedge clk) if (n3488) n3595 <= 1'b0 ? 1'b0 : n5961;
/* FF  7 15  7 */ always @(posedge clk) if (n630) n740 <= 1'b0 ? 1'b0 : n5962;
/* FF 21 22  6 */ always @(posedge clk) if (n2384) n2940 <= 1'b0 ? 1'b0 : n5963;
/* FF 13 26  0 */ always @(posedge clk) if (n1271) n1544 <= 1'b0 ? 1'b0 : n5964;
/* FF 18 19  5 */ always @(posedge clk) if (n1982) n2344 <= 1'b0 ? 1'b0 : n5965;
/* FF  3 18  2 */ always @(posedge clk) if (n215) n320 <= 1'b0 ? 1'b0 : n5966;
/* FF  2 22  0 */ always @(posedge clk) if (n352) n235 <= 1'b0 ? 1'b0 : n5967;
/* FF 18 28  4 */ always @(posedge clk) if (n2020) n2404 <= 1'b0 ? 1'b0 : n5968;
/* FF 11 22  1 */ always @(posedge clk) if (n695) n1207 <= 1'b0 ? 1'b0 : n5969;
/* FF 28 17  1 */ always @(posedge clk) if (n3765) n3767 <= 1'b0 ? 1'b0 : n5970;
/* FF 16 15  2 */ always @(posedge clk) if (n739) n1945 <= 1'b0 ? 1'b0 : n5971;
/* FF  5 16  4 */ always @(posedge clk) if (n511) n522 <= 1'b0 ? 1'b0 : n5972;
/* FF 19  7  7 */ always @(posedge clk) if (n2670) n2459 <= 1'b0 ? 1'b0 : n5973;
/* FF 23 13  6 */ always @(posedge clk) if (n3045) n3214 <= 1'b0 ? 1'b0 : n5974;
/* FF 10 18  0 */ always @(posedge clk) if (n1187) n1033 <= 1'b0 ? 1'b0 : n5975;
/* FF  9 10  2 */ always @(posedge clk) if (n988) n836 <= 1'b0 ? 1'b0 : n5976;
/* FF 13 12  3 */ always @(posedge clk) if (n1137) n1452 <= 1'b0 ? 1'b0 : n5977;
/* FF 15 18  0 */ always @(posedge clk) if (n1355) n1808 <= 1'b0 ? 1'b0 : n5978;
/* FF 20 27  5 */ always @(posedge clk) if (n2195) n2819 <= 1'b0 ? 1'b0 : n5979;
/* FF  6 15  3 */ always @(posedge clk) if (n630) n633 <= 1'b0 ? 1'b0 : n5980;
/* FF 20 16  4 */ assign n1491 = n5981;
/* FF 12 20  2 */ assign n5982 = n1511;
/* FF 14 14  1 */ always @(posedge clk) if (n1791) n1633 <= 1'b0 ? 1'b0 : n5983;
/* FF 17 11  5 */ always @(posedge clk) if (n2076) n2071 <= 1'b0 ? 1'b0 : n5984;
/* FF  1 16  2 */ always @(posedge clk) if (n85) n90 <= 1'b0 ? 1'b0 : n5985;
/* FF 19  8  3 */ always @(posedge clk) if (n2451) n2464 <= 1'b0 ? 1'b0 : n5986;
/* FF 23 14  0 */ assign n3045 = n5987;
/* FF 24 17  0 */ always @(posedge clk) if (n2123) n3394 <= 1'b0 ? 1'b0 : n5988;
/* FF  3 14  4 */ always @(posedge clk) if (n197) n289 <= 1'b0 ? 1'b0 : n5989;
/* FF  7 19  0 */ assign n350 = n5990;
/* FF  9 20  2 */ always @(posedge clk) if (n961) n696 <= 1'b0 ? 1'b0 : n5991;
/* FF 21 10  1 */ assign \rco[51]  = n5992;
/* FF 26 19  6 */ always @(posedge clk) if (n2730) n3561 <= 1'b0 ? 1'b0 : n5993;
/* FF 27  9  4 */ always @(posedge clk) if (n3621) n3614 <= 1'b0 ? 1'b0 : n5994;
/* FF 12 23  4 */ always @(posedge clk) if (n1357) n1362 <= 1'b0 ? 1'b0 : n5995;
/* FF 26 12  7 */ always @(posedge clk) if (n3368) n3524 <= 1'b0 ? 1'b0 : n5996;
/* FF 17  8  1 */ assign n2045 = n5997;
/* FF 20  6  0 */ always @(posedge clk) if (n2247) n2659 <= 1'b0 ? 1'b0 : n5998;
/* FF  4 12  7 */ always @(posedge clk) if (n77) n400 <= 1'b0 ? 1'b0 : n5999;
/* FF 16 16  0 */ always @(posedge clk) if (n2110) n1955 <= 1'b0 ? 1'b0 : n6000;
/* FF 22 12  6 */ always @(posedge clk) if (n3029) n3042 <= 1'b0 ? 1'b0 : n6001;
/* FF 10 22  5 */ assign n246 = n6002;
/* FF 21 28  0 */ always @(posedge clk) if (n2196) n2979 <= 1'b0 ? 1'b0 : n6003;
/* FF 13 16  6 */ always @(posedge clk) if (n922) n1483 <= 1'b0 ? 1'b0 : n6004;
/* FF 27  7  5 */ always @(posedge clk) if (n3459) n3600 <= 1'b0 ? 1'b0 : n6005;
/* FF  9 25  4 */ always @(posedge clk) if (n2) n939 <= 1'b0 ? 1'b0 : n6006;
/* FF 27 10  6 */ assign n3464 = n6007;
/* FF 13 27  7 */ always @(posedge clk) if (n1532) n1556 <= 1'b0 ? 1'b0 : n6008;
/* FF 18 18  2 */ always @(posedge clk) if (n1825) n2336 <= 1'b0 ? 1'b0 : n6009;
/* FF  3 19  1 */ always @(posedge clk) if (n115) n327 <= 1'b0 ? 1'b0 : n6010;
/* FF 20 20  1 */ always @(posedge clk) if (n2562) n2762 <= 1'b0 ? 1'b0 : n6011;
/* FF 23 18  2 */ always @(posedge clk) if (n2573) n3244 <= 1'b0 ? 1'b0 : n6012;
/* FF 14 10  6 */ always @(posedge clk) if (n1622) n1610 <= 1'b0 ? 1'b0 : n6013;
/* FF 11 23  2 */ always @(posedge clk) if (n796) n1216 <= 1'b0 ? 1'b0 : n6014;
/* FF  5 17  7 */ always @(posedge clk) if (n2) n530 <= 1'b0 ? 1'b0 : n6015;
/* FF  4 15  3 */ always @(posedge clk) if (n207) n415 <= 1'b0 ? 1'b0 : n6016;
/* FF  1 10  7 */ always @(posedge clk) if (n37) n34 <= 1'b0 ? 1'b0 : n6017;
/* FF 10 21  1 */ always @(posedge clk) if (n818) n1059 <= 1'b0 ? 1'b0 : n6018;
/* FF 13 13  0 */ assign n1015 = n6019;
/* FF 15 19  3 */ always @(posedge clk) if (n1355) n1820 <= 1'b0 ? 1'b0 : n6020;
/* FF 20 26  6 */ always @(posedge clk) if (n2615) n2810 <= 1'b0 ? 1'b0 : n6021;
/* FF 20 23  5 */ assign n2775 = n6022;
/* FF  6 14  4 */ always @(posedge clk) if (n78) n401 <= 1'b0 ? 1'b0 : n6023;
/* FF 12 27  3 */ always @(posedge clk) if (n1384) n1272 <= 1'b0 ? 1'b0 : n6024;
/* FF 17 20  4 */ always @(posedge clk) if (n1843) n2140 <= 1'b0 ? 1'b0 : n6025;
/* FF  2 11  5 */ always @(posedge clk) if (n168) n173 <= 1'b0 ? 1'b0 : n6026;
/* FF 29  5  6 */ always @(posedge clk) if (n3605) n3824 <= 1'b0 ? 1'b0 : n6027;
/* FF 23 15  3 */ always @(posedge clk) if (n3216) n3225 <= 1'b0 ? 1'b0 : n6028;
/* FF 27 22  0 */ always @(posedge clk) if (n3703) n3695 <= 1'b0 ? 1'b0 : n6029;
/* FF  3 15  7 */ always @(posedge clk) if (n207) n300 <= 1'b0 ? 1'b0 : n6030;
/* FF 21 16  7 */ always @(posedge clk) if (n2551) n2894 <= 1'b0 ? 1'b0 : n6031;
/* FF  7 16  1 */ always @(posedge clk) if (n630) n742 <= 1'b0 ? 1'b0 : n6032;
/* FF  9 21  1 */ always @(posedge clk) if (n818) n915 <= 1'b0 ? 1'b0 : n6033;
/* FF 21 11  6 */ always @(posedge clk) if (n2085) n2863 <= 1'b0 ? 1'b0 : n6034;
/* FF 26 18  1 */ assign n3553 = n6035;
/* FF 12  9  6 */ always @(posedge clk) if (n850) n1284 <= 1'b0 ? 1'b0 : n6036;
/* FF 18 22  7 */ always @(posedge clk) if (n2164) n2360 <= 1'b0 ? 1'b0 : n6037;
/* FF 12 22  7 */ always @(posedge clk) if (n1357) n1354 <= 1'b0 ? 1'b0 : n6038;
/* FF 17  9  2 */ assign \rco[39]  = n2271;
/* FF  6 24  0 */ assign \rco[113]  = n6039;
/* FF 20  5  1 */ always @(posedge clk) if (n2247) n2658 <= 1'b0 ? 1'b0 : n6040;
/* FF 10  9  3 */ always @(posedge clk) if (n983) n979 <= 1'b0 ? 1'b0 : n6041;
/* FF 28 20  3 */ assign \rco[170]  = n6042;
/* FF 22 15  7 */ always @(posedge clk) if (n3216) n3064 <= 1'b0 ? 1'b0 : n6043;
/* FF  7  6  0 */ always @(posedge clk) if (n588) n706 <= 1'b0 ? 1'b0 : n6044;
/* FF  9  7  2 */ always @(posedge clk) if (n588) n825 <= 1'b0 ? 1'b0 : n6045;
/* FF 13 17  5 */ always @(posedge clk) if (n1461) n668 <= 1'b0 ? 1'b0 : n6046;
/* FF  9 26  5 */ always @(posedge clk) if (n954) n943 <= 1'b0 ? 1'b0 : n6047;
/* FF 13 28  6 */ always @(posedge clk) if (n1394) n1566 <= 1'b0 ? 1'b0 : n6048;
/* FF 27 11  5 */ always @(posedge clk) if (n3460) n3626 <= 1'b0 ? 1'b0 : n6049;
/* FF 18 21  3 */ always @(posedge clk) if (n2347) n2352 <= 1'b0 ? 1'b0 : n6050;
/* FF  3 16  0 */ always @(posedge clk) if (n197) n303 <= 1'b0 ? 1'b0 : n6051;
/* FF  6 10  1 */ always @(posedge clk) if (n589) n592 <= 1'b0 ? 1'b0 : n6052;
/* FF 20 11  0 */ assign n6053 = n2865;
/* FF 23 19  1 */ always @(posedge clk) if (n2573) n3251 <= 1'b0 ? 1'b0 : n6054;
/* FF 11 20  3 */ always @(posedge clk) if (n1339) n1192 <= 1'b0 ? 1'b0 : n6055;
/* FF 29  9  3 */ assign \rco[80]  = n6056;
/* FF 17 27  2 */ always @(posedge clk) if (n1) n2190 <= 1'b0 ? 1'b0 : n6057;
/* FF 28 23  7 */ always @(posedge clk) if (n3704) n3813 <= 1'b0 ? 1'b0 : n6058;
/* FF  5 18  6 */ always @(posedge clk) if (n657) n537 <= 1'b0 ? 1'b0 : n6059;
/* FF  4 14  0 */ assign \rco[18]  = n512;
/* FF 19  5  1 */ always @(posedge clk) if (n2230) n2436 <= 1'b0 ? 1'b0 : n6060;
/* FF 22 25  2 */ always @(posedge clk) if (n2812) n3127 <= 1'b0 ? 1'b0 : n6061;
/* FF 10 20  2 */ always @(posedge clk) if (n922) n1050 <= 1'b0 ? 1'b0 : n6062;
/* FF 13 14  1 */ always @(posedge clk) if (n1461) n1463 <= 1'b0 ? 1'b0 : n6063;
/* FF 15 16  2 */ always @(posedge clk) if (n1500) n1795 <= 1'b0 ? 1'b0 : n6064;
/* FF 21 15  3 */ assign n2564 = n6065;
/* FF 20 25  7 */ always @(posedge clk) if (n2612) n2804 <= 1'b0 ? 1'b0 : n6066;
/* FF 26 22  6 */ always @(posedge clk) if (n2730) n3574 <= 1'b0 ? 1'b0 : n6067;
/* FF  6  9  5 */ assign n56 = n728;
/* FF 20 22  6 */ always @(posedge clk) if (n2384) n2782 <= 1'b0 ? 1'b0 : n6068;
/* FF 12 26  0 */ always @(posedge clk) if (n1393) n1385 <= 1'b0 ? 1'b0 : n6069;
/* FF 14  8  3 */ always @(posedge clk) if (n1741) n1596 <= 1'b0 ? 1'b0 : n6070;
/* FF  2 10  2 */ always @(posedge clk) if (n168) n167 <= 1'b0 ? 1'b0 : n6071;
/* FF  1 18  0 */ always @(posedge clk) if (n115) n98 <= 1'b0 ? 1'b0 : n6072;
/* FF 17 21  7 */ always @(posedge clk) if (n2347) n2151 <= 1'b0 ? 1'b0 : n6073;
/* FF 17 24  4 */ always @(posedge clk) if (n2000) n2170 <= 1'b0 ? 1'b0 : n6074;
/* FF 23 12  2 */ always @(posedge clk) if (n3031) n3202 <= 1'b0 ? 1'b0 : n6075;
/* FF 27 23  3 */ assign n3703 = n6076;
/* FF  3 12  6 */ always @(posedge clk) if (n168) n283 <= 1'b0 ? 1'b0 : n6077;
/* FF 21 17  4 */ always @(posedge clk) if (n2519) n2898 <= 1'b0 ? 1'b0 : n6078;
/* FF 18  2  4 */ always @(posedge clk) if (n2207) n2203 <= 1'b0 ? 1'b0 : n6079;
/* FF  7 17  6 */ always @(posedge clk) if (n549) n757 <= 1'b0 ? 1'b0 : n6080;
/* FF  9 22  0 */ always @(posedge clk) if (n819) n923 <= 1'b0 ? 1'b0 : n6081;
/* FF 21 12  7 */ always @(posedge clk) if (n3029) n2873 <= 1'b0 ? 1'b0 : n6082;
/* FF 12  8  1 */ always @(posedge clk) if (n1131) n1279 <= 1'b0 ? 1'b0 : n6083;
/* FF 26 21  0 */ always @(posedge clk) if (n3421) n3562 <= 1'b0 ? 1'b0 : n6084;
/* FF 15  6  2 */ always @(posedge clk) if (n1744) n1735 <= 1'b0 ? 1'b0 : n6085;
/* FF 14 26  0 */ always @(posedge clk) if (n1271) n1711 <= 1'b0 ? 1'b0 : n6086;
/* FF 12 21  6 */ always @(posedge clk) if (n1205) n1345 <= 1'b0 ? 1'b0 : n6087;
/* FF 17 10  3 */ always @(posedge clk) if (n2282) n2062 <= 1'b0 ? 1'b0 : n6088;
/* FF  1 12  4 */ always @(posedge clk) if (n39) n50 <= 1'b0 ? 1'b0 : n6089;
/* FF 22 14  0 */ always @(posedge clk) if (n3045) n3051 <= 1'b0 ? 1'b0 : n6090;
/* FF  7  7  3 */ always @(posedge clk) if (n588) n712 <= 1'b0 ? 1'b0 : n6091;
/* FF 13 18  4 */ always @(posedge clk) if (n1205) n1496 <= 1'b0 ? 1'b0 : n6092;
/* FF 27  5  3 */ always @(posedge clk) if (n3594) n3588 <= 1'b0 ? 1'b0 : n6093;
/* FF 27  8  4 */ always @(posedge clk) if (n3464) n3606 <= 1'b0 ? 1'b0 : n6094;
/* FF 18 20  0 */ assign \rco[158]  = n6095;
/* FF  6 21  0 */ assign n360 = n6096;
/* FF 20 10  3 */ always @(posedge clk) if (n2697) n2686 <= 1'b0 ? 1'b0 : n6097;
/* FF 23 16  0 */ assign n2540 = n6098;
/* FF 11 14  5 */ always @(posedge clk) if (n1154) n1151 <= 1'b0 ? 1'b0 : n6099;
/* FF 16  7  6 */ always @(posedge clk) if (n1743) n1913 <= 1'b0 ? 1'b0 : n6100;
/* FF 11 21  4 */ always @(posedge clk) if (n819) n1200 <= 1'b0 ? 1'b0 : n6101;
/* FF 29 10  2 */ always @(posedge clk) if (n3464) n3834 <= 1'b0 ? 1'b0 : n6102;
/* FF 28 22  4 */ always @(posedge clk) if (n3704) n3803 <= 1'b0 ? 1'b0 : n6103;
/* FF  5 19  1 */ always @(posedge clk) if (n349) n540 <= 1'b0 ? 1'b0 : n6104;
/* FF  4 13  1 */ assign \rco[17]  = n502;
/* FF 22 24  1 */ always @(posedge clk) if (n3113) n3117 <= 1'b0 ? 1'b0 : n6105;
/* FF 10 23  3 */ assign n820 = n6106;
/* FF 30 12  2 */ always @(posedge clk) if (n3892) n3896 <= 1'b0 ? 1'b0 : n6107;
/* FF 15 17  5 */ always @(posedge clk) if (n1500) n758 <= 1'b0 ? 1'b0 : n6108;
/* FF 18  6  1 */ always @(posedge clk) if (n2241) n2232 <= 1'b0 ? 1'b0 : n6109;
/* FF  7 21  3 */ always @(posedge clk) if (n360) n771 <= 1'b0 ? 1'b0 : n6110;
/* FF  6  7  7 */ always @(posedge clk) if (n570) n578 <= 1'b0 ? 1'b0 : n6111;
/* FF 20 24  0 */ always @(posedge clk) if (n2775) n2788 <= 1'b0 ? 1'b0 : n6112;
/* FF  6  8  6 */ always @(posedge clk) if (n570) n585 <= 1'b0 ? 1'b0 : n6113;
/* FF 12 25  1 */ always @(posedge clk) if (n1532) n1377 <= 1'b0 ? 1'b0 : n6114;
/* FF 14 11  2 */ always @(posedge clk) if (n1622) n1614 <= 1'b0 ? 1'b0 : n6115;
/* FF 17 22  6 */ always @(posedge clk) if (n1999) n2158 <= 1'b0 ? 1'b0 : n6116;
/* FF 17 25  7 */ always @(posedge clk) if (n2017) n2183 <= 1'b0 ? 1'b0 : n6117;
/* FF 27 20  2 */ always @(posedge clk) if (n3424) n3677 <= 1'b0 ? 1'b0 : n6118;
/* FF  4 19  5 */ assign n2 = n6119;
/* FF  3 13  1 */ assign n285 = n404;
/* FF 21 18  5 */ always @(posedge clk) if (n2757) n2907 <= 1'b0 ? 1'b0 : n6120;
/* FF 22 10  5 */ always @(posedge clk) if (n2856) n3027 <= 1'b0 ? 1'b0 : n6121;
/* FF 18  5  5 */ always @(posedge clk) if (n2230) n2226 <= 1'b0 ? 1'b0 : n6122;
/* FF  7 22  7 */ always @(posedge clk) if (n695) n565 <= 1'b0 ? 1'b0 : n6123;
/* FF 21 13  4 */ always @(posedge clk) if (n2519) n2878 <= 1'b0 ? 1'b0 : n6124;
/* FF 12 15  0 */ always @(posedge clk) if (n1155) n1296 <= 1'b0 ? 1'b0 : n6125;
/* FF 26 20  3 */ assign n6126 = n3683;
/* FF 18 24  5 */ always @(posedge clk) if (n1878) n2011 <= 1'b0 ? 1'b0 : n6127;
/* FF 14 21  1 */ assign n1671 = n1845;
/* FF 19 30  2 */ always @(posedge clk) if (n2592) n2636 <= 1'b0 ? 1'b0 : n6128;
/* FF 11 17  1 */ always @(posedge clk) if (n900) n1169 <= 1'b0 ? 1'b0 : n6129;
/* FF 10 11  1 */ assign n990 = n1136;
/* FF 16  8  4 */ always @(posedge clk) if (n1625) n1919 <= 1'b0 ? 1'b0 : n6130;
/* FF  1 13  7 */ always @(posedge clk) if (n83) n66 <= 1'b0 ? 1'b0 : n6131;
/* FF 13 19  3 */ assign n1501 = n6132;
/* FF 15 21  2 */ always @(posedge clk) if (n1356) n1838 <= 1'b0 ? 1'b0 : n6133;
/* FF 20 28  5 */ always @(posedge clk) if (n2195) n2826 <= 1'b0 ? 1'b0 : n6134;
/* FF 18 23  1 */ always @(posedge clk) if (n1999) n2363 <= 1'b0 ? 1'b0 : n6135;
/* FF  6 20  3 */ always @(posedge clk) if (n552) n663 <= 1'b0 ? 1'b0 : n6136;
/* FF 20  9  2 */ assign n2679 = n6137;
/* FF 23 17  7 */ always @(posedge clk) if (n2540) n3239 <= 1'b0 ? 1'b0 : n6138;
/* FF 11 15  6 */ always @(posedge clk) if (n733) n1157 <= 1'b0 ? 1'b0 : n6139;
/* FF 26  6  3 */ always @(posedge clk) if (n3459) n3476 <= 1'b0 ? 1'b0 : n6140;
/* FF 14  7  5 */ always @(posedge clk) if (n1743) n587 <= 1'b0 ? 1'b0 : n6141;
/* FF 16  6  5 */ always @(posedge clk) if (n1744) n1902 <= 1'b0 ? 1'b0 : n6142;
/* FF 11 18  5 */ always @(posedge clk) if (n1187) n1184 <= 1'b0 ? 1'b0 : n6143;
/* FF 29 11  5 */ always @(posedge clk) if (n3751) n3844 <= 1'b0 ? 1'b0 : n6144;
/* FF 28 21  5 */ always @(posedge clk) if (n3788) n3796 <= 1'b0 ? 1'b0 : n6145;
/* FF 19  3  3 */ always @(posedge clk) if (n1887) n2430 <= 1'b0 ? 1'b0 : n6146;
/* FF 22 27  0 */ always @(posedge clk) if (n2970) n3143 <= 1'b0 ? 1'b0 : n6147;
/* FF  3  9  6 */ always @(posedge clk) if (n260) n258 <= 1'b0 ? 1'b0 : n6148;
/* FF 15 22  4 */ always @(posedge clk) if (n1835) n1850 <= 1'b0 ? 1'b0 : n6149;
/* FF 18  9  0 */ always @(posedge clk) if (n2055) n2261 <= 1'b0 ? 1'b0 : n6150;
/* FF  7 26  2 */ always @(posedge clk) if (n567) n800 <= 1'b0 ? 1'b0 : n6151;
/* FF  9 19  4 */ always @(posedge clk) if (n454) n905 <= 1'b0 ? 1'b0 : n6152;
/* FF 12 19  7 */ always @(posedge clk) if (n1501) n1334 <= 1'b0 ? 1'b0 : n6153;
/* FF 26  8  4 */ always @(posedge clk) if (n3603) n3494 <= 1'b0 ? 1'b0 : n6154;
/* FF  6 11  7 */ always @(posedge clk) if (n286) n605 <= 1'b0 ? 1'b0 : n6155;
/* FF 12 24  6 */ always @(posedge clk) if (n961) n1373 <= 1'b0 ? 1'b0 : n6156;
/* FF 17 23  1 */ always @(posedge clk) if (n1069) n2161 <= 1'b0 ? 1'b0 : n6157;
/* FF  2 12  0 */ always @(posedge clk) if (n39) n176 <= 1'b0 ? 1'b0 : n6158;
/* FF 19 17  0 */ always @(posedge clk) if (n2727) n2541 <= 1'b0 ? 1'b0 : n6159;
/* FF 17 26  6 */ always @(posedge clk) if (n1557) n2187 <= 1'b0 ? 1'b0 : n6160;
/* FF 22 21  3 */ always @(posedge clk) if (n2564) n3099 <= 1'b0 ? 1'b0 : n6161;
/* FF 24 24  3 */ always @(posedge clk) if (n3112) n3442 <= 1'b0 ? 1'b0 : n6162;
/* FF 27 21  5 */ always @(posedge clk) if (n3421) n3692 <= 1'b0 ? 1'b0 : n6163;
/* FF  4 18  6 */ always @(posedge clk) if (n349) n436 <= 1'b0 ? 1'b0 : n6164;
/* FF  3 10  0 */ always @(posedge clk) if (n251) n262 <= 1'b0 ? 1'b0 : n6165;
/* FF 21 19  2 */ always @(posedge clk) if (n2757) n2912 <= 1'b0 ? 1'b0 : n6166;
/* FF 18  4  6 */ always @(posedge clk) if (n2207) n2219 <= 1'b0 ? 1'b0 : n6167;
/* FF 21 14  5 */ always @(posedge clk) if (n2519) n2885 <= 1'b0 ? 1'b0 : n6168;
/* FF  9 16  6 */ always @(posedge clk) if (n645) n881 <= 1'b0 ? 1'b0 : n6169;
/* FF 12 14  3 */ always @(posedge clk) if (n1154) n1291 <= 1'b0 ? 1'b0 : n6170;
/* FF 26 23  2 */ always @(posedge clk) if (n3703) n3578 <= 1'b0 ? 1'b0 : n6171;
/* FF 18 27  4 */ always @(posedge clk) if (n2020) n2397 <= 1'b0 ? 1'b0 : n6172;
/* FF 14 20  2 */ always @(posedge clk) if (n1347) n1678 <= 1'b0 ? 1'b0 : n6173;
/* FF  5  8  2 */ always @(posedge clk) if (n21) n470 <= 1'b0 ? 1'b0 : n6174;
/* FF 19 31  1 */ always @(posedge clk) if (n2592) n2642 <= 1'b0 ? 1'b0 : n6175;
/* FF 23 21  4 */ always @(posedge clk) if (n3258) n3275 <= 1'b0 ? 1'b0 : n6176;
/* FF 11 30  0 */ always @(posedge clk) if (n1384) n1273 <= 1'b0 ? 1'b0 : n6177;
/* FF 16 23  5 */ always @(posedge clk) if (n2000) n913 <= 1'b0 ? 1'b0 : n6178;
/* FF  1 14  6 */ always @(posedge clk) if (n85) n74 <= 1'b0 ? 1'b0 : n6179;
/* FF 22  8  2 */ always @(posedge clk) if (n2989) n3011 <= 1'b0 ? 1'b0 : n6180;
/* FF 13 20  2 */ always @(posedge clk) if (n1339) n1505 <= 1'b0 ? 1'b0 : n6181;
/* FF 15 10  3 */ always @(posedge clk) if (n1624) n1757 <= 1'b0 ? 1'b0 : n6182;
/* FF 20 19  4 */ always @(posedge clk) if (n2562) n2753 <= 1'b0 ? 1'b0 : n6183;
/* FF  6 23  2 */ always @(posedge clk) if (n360) n689 <= 1'b0 ? 1'b0 : n6184;
/* FF 20  8  5 */ always @(posedge clk) if (n2247) n2673 <= 1'b0 ? 1'b0 : n6185;
/* FF 12 28  3 */ always @(posedge clk) if (n1394) n1397 <= 1'b0 ? 1'b0 : n6186;
/* FF 23 22  6 */ always @(posedge clk) if (n3422) n3285 <= 1'b0 ? 1'b0 : n6187;
/* FF 17 19  6 */ always @(posedge clk) if (n1982) n2134 <= 1'b0 ? 1'b0 : n6188;
/* FF 16  5  4 */ always @(posedge clk) if (n1742) n1892 <= 1'b0 ? 1'b0 : n6189;
/* FF 11 19  6 */ assign n6190 = n1336;
/* FF 29 12  4 */ always @(posedge clk) if (n3751) n3853 <= 1'b0 ? 1'b0 : n6191;
/* FF 16 10  5 */ always @(posedge clk) if (n1771) n1772 <= 1'b0 ? 1'b0 : n6192;
/* FF  5 21  3 */ assign n6193 = n677;
/* FF 27 17  2 */ always @(posedge clk) if (n3249) n3653 <= 1'b0 ? 1'b0 : n6194;
/* FF 15 24  6 */ always @(posedge clk) if (n778) n1869 <= 1'b0 ? 1'b0 : n6195;
/* FF 21 23  7 */ always @(posedge clk) if (n2961) n2950 <= 1'b0 ? 1'b0 : n6196;
/* FF 15 23  7 */ always @(posedge clk) if (n778) n1859 <= 1'b0 ? 1'b0 : n6197;
/* FF 18  8  3 */ always @(posedge clk) if (n2055) n2252 <= 1'b0 ? 1'b0 : n6198;
/* FF 12 18  4 */ always @(posedge clk) if (n1501) n1324 <= 1'b0 ? 1'b0 : n6199;
/* FF 26 11  5 */ always @(posedge clk) if (n3033) n3513 <= 1'b0 ? 1'b0 : n6200;
/* FF 17 16  0 */ assign n2109 = n6201;
/* FF  2 15  1 */ assign \rco[6]  = n302;
/* FF 19 14  1 */ always @(posedge clk) if (n2123) n2512 <= 1'b0 ? 1'b0 : n6202;
/* FF 22 20  0 */ always @(posedge clk) if (n3087) n3088 <= 1'b0 ? 1'b0 : n6203;
/* FF 10 14  3 */ always @(posedge clk) if (n750) n1010 <= 1'b0 ? 1'b0 : n6204;
/* FF 24 23  2 */ always @(posedge clk) if (n3104) n3435 <= 1'b0 ? 1'b0 : n6205;
/* FF 28 10  2 */ always @(posedge clk) if (n3462) n3743 <= 1'b0 ? 1'b0 : n6206;
/* FF 27 18  4 */ always @(posedge clk) if (n3553) n3661 <= 1'b0 ? 1'b0 : n6207;
/* FF  3 11  3 */ always @(posedge clk) if (n153) n273 <= 1'b0 ? 1'b0 : n6208;
/* FF  7  9  2 */ always @(posedge clk) if (n589) n720 <= 1'b0 ? 1'b0 : n6209;
/* FF 21 20  3 */ always @(posedge clk) if (n3087) n2921 <= 1'b0 ? 1'b0 : n6210;
/* FF 18  7  7 */ always @(posedge clk) if (n1761) n2246 <= 1'b0 ? 1'b0 : n6211;
/* FF  7 20  5 */ assign n768 = n6212;
/* FF  9 17  5 */ always @(posedge clk) if (n1030) n888 <= 1'b0 ? 1'b0 : n6213;
/* FF 18 26  3 */ always @(posedge clk) if (n2615) n2388 <= 1'b0 ? 1'b0 : n6214;
/* FF 14 23  3 */ assign \rco[114]  = n6215;
/* FF 20 12  2 */ always @(posedge clk) if (n2682) n2700 <= 1'b0 ? 1'b0 : n6216;
/* FF  5  9  1 */ always @(posedge clk) if (n21) n154 <= 1'b0 ? 1'b0 : n6217;
/* FF 19 28  0 */ always @(posedge clk) if (n2614) n2624 <= 1'b0 ? 1'b0 : n6218;
/* FF  1 15  1 */ assign n83 = n6219;
/* FF 22 11  3 */ assign n3031 = n6220;
/* FF 13 21  1 */ always @(posedge clk) if (n1356) n1514 <= 1'b0 ? 1'b0 : n6221;
/* FF 30 10  1 */ always @(posedge clk) if (n3892) n3886 <= 1'b0 ? 1'b0 : n6222;
/* FF 15 11  0 */ always @(posedge clk) if (n1624) n1763 <= 1'b0 ? 1'b0 : n6223;
/* FF  6 13  4 */ always @(posedge clk) if (n78) n619 <= 1'b0 ? 1'b0 : n6224;
/* FF 20 18  7 */ always @(posedge clk) if (n2348) n2747 <= 1'b0 ? 1'b0 : n6225;
/* FF  6 22  5 */ always @(posedge clk) if (n673) n683 <= 1'b0 ? 1'b0 : n6226;
/* FF 20 15  4 */ always @(posedge clk) if (n2715) n2721 <= 1'b0 ? 1'b0 : n6227;
/* FF 23 23  5 */ always @(posedge clk) if (n3104) n3292 <= 1'b0 ? 1'b0 : n6228;
/* FF 11 13  0 */ always @(posedge clk) if (n733) n1138 <= 1'b0 ? 1'b0 : n6229;
/* FF 11 16  7 */ always @(posedge clk) if (n891) n1166 <= 1'b0 ? 1'b0 : n6230;
/* FF  5 22  2 */ always @(posedge clk) if (n673) n557 <= 1'b0 ? 1'b0 : n6231;
/* FF 13  7  2 */ always @(posedge clk) if (n977) n1425 <= 1'b0 ? 1'b0 : n6232;
/* FF 15 25  1 */ assign \rco[193]  = n6233;
/* FF  7 13  7 */ always @(posedge clk) if (n733) n731 <= 1'b0 ? 1'b0 : n6234;
/* FF 18 11  2 */ assign n6235 = n2495;
/* FF 15 20  6 */ always @(posedge clk) if (n1347) n1833 <= 1'b0 ? 1'b0 : n6236;
/* FF  7 24  0 */ always @(posedge clk) if (n697) n795 <= 1'b0 ? 1'b0 : n6237;
/* FF 12 17  5 */ always @(posedge clk) if (n900) n1317 <= 1'b0 ? 1'b0 : n6238;
/* FF 26 10  2 */ always @(posedge clk) if (n3033) n3507 <= 1'b0 ? 1'b0 : n6239;
/* FF 26  7  5 */ always @(posedge clk) if (n3603) n3455 <= 1'b0 ? 1'b0 : n6240;
/* FF 17 17  3 */ always @(posedge clk) if (n2111) n2117 <= 1'b0 ? 1'b0 : n6241;
/* FF 19 15  2 */ always @(posedge clk) if (n2715) n2527 <= 1'b0 ? 1'b0 : n6242;
/* FF 23  5  1 */ always @(posedge clk) if (n3158) n3151 <= 1'b0 ? 1'b0 : n6243;
/* FF 22 23  1 */ assign n3112 = n6244;
/* FF 24 22  1 */ always @(posedge clk) if (n3422) n3426 <= 1'b0 ? 1'b0 : n6245;
/* FF 28  9  3 */ always @(posedge clk) if (n3621) n3737 <= 1'b0 ? 1'b0 : n6246;
/* FF 27 19  7 */ always @(posedge clk) if (n3553) n3674 <= 1'b0 ? 1'b0 : n6247;
/* FF  4 16  0 */ always @(posedge clk) if (n79) n420 <= 1'b0 ? 1'b0 : n6248;
/* FF 21 21  0 */ always @(posedge clk) if (n2564) n2926 <= 1'b0 ? 1'b0 : n6249;
/* FF  9 18  4 */ always @(posedge clk) if (n1030) n896 <= 1'b0 ? 1'b0 : n6250;
/* FF 18 29  2 */ always @(posedge clk) if (n1881) n2410 <= 1'b0 ? 1'b0 : n6251;
/* FF 14 22  4 */ always @(posedge clk) if (n1402) n1691 <= 1'b0 ? 1'b0 : n6252;
/* FF 17  3  0 */ always @(posedge clk) if (n1887) n2025 <= 1'b0 ? 1'b0 : n6253;
/* FF  6 18  2 */ always @(posedge clk) if (n657) n651 <= 1'b0 ? 1'b0 : n6254;
/* FF  5 10  0 */ assign n184 = n6255;
/* FF 23 27  6 */ always @(posedge clk) if (n2017) n3317 <= 1'b0 ? 1'b0 : n6256;
/* FF 23  6  5 */ always @(posedge clk) if (n3158) n3164 <= 1'b0 ? 1'b0 : n6257;
/* FF 11 28  2 */ always @(posedge clk) if (n1384) n1257 <= 1'b0 ? 1'b0 : n6258;
/* FF 10 12  4 */ always @(posedge clk) if (n996) n1001 <= 1'b0 ? 1'b0 : n6259;
/* FF 24 25  5 */ always @(posedge clk) if (n2812) n3451 <= 1'b0 ? 1'b0 : n6260;
/* FF 16 21  7 */ always @(posedge clk) if (n1835) n1987 <= 1'b0 ? 1'b0 : n6261;
/* FF  1  8  0 */ always @(posedge clk) if (n37) n14 <= 1'b0 ? 1'b0 : n6262;
/* FF 16 26  6 */ always @(posedge clk) if (n1557) n2016 <= 1'b0 ? 1'b0 : n6263;
/* FF 13 22  0 */ assign n695 = n6264;
/* FF 15  8  1 */ always @(posedge clk) if (n1741) n1747 <= 1'b0 ? 1'b0 : n6265;
/* FF  3 22  2 */ always @(posedge clk) if (n352) n355 <= 1'b0 ? 1'b0 : n6266;
/* FF 21  7  4 */ assign n2247 = n6267;
/* FF  2 18  0 */ always @(posedge clk) if (n115) n209 <= 1'b0 ? 1'b0 : n6268;
/* FF  6 12  7 */ always @(posedge clk) if (n286) n613 <= 1'b0 ? 1'b0 : n6269;
/* FF 20 17  6 */ always @(posedge clk) if (n2727) n2738 <= 1'b0 ? 1'b0 : n6270;
/* FF 26 14  7 */ always @(posedge clk) if (n3527) n3540 <= 1'b0 ? 1'b0 : n6271;
/* FF 23 20  4 */ always @(posedge clk) if (n3258) n3267 <= 1'b0 ? 1'b0 : n6272;
/* FF 24  7  1 */ assign n3175 = n3457;
/* FF  9 14  2 */ always @(posedge clk) if (n629) n861 <= 1'b0 ? 1'b0 : n6273;
/* FF  4 20  5 */ always @(posedge clk) if (n215) n443 <= 1'b0 ? 1'b0 : n6274;
/* FF 21  9  5 */ always @(posedge clk) if (n2856) n2689 <= 1'b0 ? 1'b0 : n6275;
/* FF 18 10  5 */ always @(posedge clk) if (n2282) n2278 <= 1'b0 ? 1'b0 : n6276;
/* FF 12 16  2 */ always @(posedge clk) if (n1155) n1306 <= 1'b0 ? 1'b0 : n6277;
/* FF 26 13  3 */ always @(posedge clk) if (n3033) n3528 <= 1'b0 ? 1'b0 : n6278;
/* FF 14 18  1 */ always @(posedge clk) if (n1672) n1662 <= 1'b0 ? 1'b0 : n6279;
/* FF 19 25  4 */ always @(posedge clk) if (n2612) n2608 <= 1'b0 ? 1'b0 : n6280;
/* FF 17 18  2 */ always @(posedge clk) if (n1825) n2127 <= 1'b0 ? 1'b0 : n6281;
/* FF 19 12  3 */ always @(posedge clk) if (n1936) n2500 <= 1'b0 ? 1'b0 : n6282;
/* FF 23 10  0 */ always @(posedge clk) if (n2697) n3183 <= 1'b0 ? 1'b0 : n6283;
/* FF 22 22  6 */ always @(posedge clk) if (n2961) n3110 <= 1'b0 ? 1'b0 : n6284;
/* FF 24 21  0 */ assign n3258 = n6285;
/* FF 28  8  4 */ always @(posedge clk) if (n3605) n3730 <= 1'b0 ? 1'b0 : n6286;
/* FF  7 15  0 */ assign \rco[26]  = n6287;
/* FF  9 24  2 */ always @(posedge clk) if (n820) n934 <= 1'b0 ? 1'b0 : n6288;
/* FF 21 22  1 */ always @(posedge clk) if (n2384) n2936 <= 1'b0 ? 1'b0 : n6289;
/* FF  2 22  5 */ always @(posedge clk) if (n352) n240 <= 1'b0 ? 1'b0 : n6290;
/* FF 18 28  1 */ assign \rco[198]  = n6291;
/* FF 14 17  5 */ always @(posedge clk) if (n1672) n1659 <= 1'b0 ? 1'b0 : n6292;
/* FF 17 12  1 */ always @(posedge clk) if (n2056) n2078 <= 1'b0 ? 1'b0 : n6293;
/* FF 19 26  6 */ assign n2614 = n6294;
/* FF 23 24  7 */ always @(posedge clk) if (n3112) n3303 <= 1'b0 ? 1'b0 : n6295;
/* FF 11 22  4 */ always @(posedge clk) if (n695) n1210 <= 1'b0 ? 1'b0 : n6296;
/* FF 28 17  4 */ always @(posedge clk) if (n3765) n3770 <= 1'b0 ? 1'b0 : n6297;
/* FF 23  7  6 */ always @(posedge clk) if (n3006) n3172 <= 1'b0 ? 1'b0 : n6298;
/* FF 11 29  5 */ always @(posedge clk) if (n1384) n1267 <= 1'b0 ? 1'b0 : n6299;
/* FF 10 15  5 */ always @(posedge clk) if (n750) n1020 <= 1'b0 ? 1'b0 : n6300;
/* FF 16 20  0 */ always @(posedge clk) if (n1843) n1974 <= 1'b0 ? 1'b0 : n6301;
/* FF 21 24  0 */ always @(posedge clk) if (n3113) n2784 <= 1'b0 ? 1'b0 : n6302;
/* FF 15 18  7 */ always @(posedge clk) if (n1355) n1815 <= 1'b0 ? 1'b0 : n6303;
/* FF 18 14  2 */ assign n2304 = n6304;
/* FF  2 21  1 */ always @(posedge clk) if (n126) n228 <= 1'b0 ? 1'b0 : n6305;
/* FF  6 15  6 */ always @(posedge clk) if (n630) n636 <= 1'b0 ? 1'b0 : n6306;
/* FF 20 16  1 */ assign n2726 = n2896;
/* FF 12 20  7 */ assign n1339 = n6307;
/* FF 20 13  6 */ always @(posedge clk) if (n2283) n2710 <= 1'b0 ? 1'b0 : n6308;
/* FF  4 11  3 */ always @(posedge clk) if (n184) n388 <= 1'b0 ? 1'b0 : n6309;
/* FF 22 18  3 */ always @(posedge clk) if (n3065) n3083 <= 1'b0 ? 1'b0 : n6310;
/* FF 10 17  1 */ assign \rco[147]  = n6311;
/* FF  9 15  5 */ always @(posedge clk) if (n645) n872 <= 1'b0 ? 1'b0 : n6312;
/* FF 24  6  2 */ always @(posedge clk) if (n3006) n3323 <= 1'b0 ? 1'b0 : n6313;
/* FF 28 12  1 */ always @(posedge clk) if (n3462) n3754 <= 1'b0 ? 1'b0 : n6314;
/* FF  7 19  5 */ always @(posedge clk) if (n549) n762 <= 1'b0 ? 1'b0 : n6315;
/* FF 21 10  4 */ assign n2697 = n6316;
/* FF 18 13  4 */ always @(posedge clk) if (n2283) n2299 <= 1'b0 ? 1'b0 : n6317;
/* FF  3 24  5 */ assign \rco[124]  = n6318;
/* FF 12 23  3 */ always @(posedge clk) if (n1357) n1361 <= 1'b0 ? 1'b0 : n6319;
/* FF 26 12  0 */ always @(posedge clk) if (n3368) n3517 <= 1'b0 ? 1'b0 : n6320;
/* FF 14 13  0 */ always @(posedge clk) if (n1015) n1626 <= 1'b0 ? 1'b0 : n6321;
/* FF  5 15  4 */ always @(posedge clk) if (n511) n518 <= 1'b0 ? 1'b0 : n6322;
/* FF 23 11  3 */ always @(posedge clk) if (n3031) n3193 <= 1'b0 ? 1'b0 : n6323;
/* FF 11 25  2 */ always @(posedge clk) if (n954) n1233 <= 1'b0 ? 1'b0 : n6324;
/* FF 22 17  7 */ always @(posedge clk) if (n3065) n3079 <= 1'b0 ? 1'b0 : n6325;
/* FF 24 20  7 */ always @(posedge clk) if (n3411) n3419 <= 1'b0 ? 1'b0 : n6326;
/* FF 16 16  5 */ always @(posedge clk) if (n2110) n1960 <= 1'b0 ? 1'b0 : n6327;
/* FF 13  6  6 */ always @(posedge clk) if (n977) n1421 <= 1'b0 ? 1'b0 : n6328;
/* FF  4 22  2 */ assign n456 = n6329;
/* FF 15 13  3 */ always @(posedge clk) if (n1015) n1780 <= 1'b0 ? 1'b0 : n6330;
/* FF 20 20  6 */ always @(posedge clk) if (n2562) n2766 <= 1'b0 ? 1'b0 : n6331;
/* FF 14 16  6 */ always @(posedge clk) if (n1792) n1652 <= 1'b0 ? 1'b0 : n6332;
/* FF 17 13  2 */ always @(posedge clk) if (n2056) n2088 <= 1'b0 ? 1'b0 : n6333;
/* FF  5 12  6 */ always @(posedge clk) if (n77) n490 <= 1'b0 ? 1'b0 : n6334;
/* FF 23 25  0 */ assign n2812 = n6335;
/* FF 11 23  7 */ always @(posedge clk) if (n796) n1220 <= 1'b0 ? 1'b0 : n6336;
/* FF 19 27  5 */ always @(posedge clk) if (n2614) n2621 <= 1'b0 ? 1'b0 : n6337;
/* FF 11 26  4 */ always @(posedge clk) if (n954) n1240 <= 1'b0 ? 1'b0 : n6338;
/* FF 16 19  1 */ assign n1685 = n6339;
/* FF  1 10  2 */ always @(posedge clk) if (n37) n30 <= 1'b0 ? 1'b0 : n6340;
/* FF 21 25  3 */ always @(posedge clk) if (n2970) n2965 <= 1'b0 ? 1'b0 : n6341;
/* FF  9 11  2 */ always @(posedge clk) if (n988) n844 <= 1'b0 ? 1'b0 : n6342;
/* FF 15 19  4 */ always @(posedge clk) if (n1355) n1821 <= 1'b0 ? 1'b0 : n6343;
/* FF 15 14  7 */ always @(posedge clk) if (n1791) n1790 <= 1'b0 ? 1'b0 : n6344;
/* FF  3 20  0 */ always @(posedge clk) if (n119) n342 <= 1'b0 ? 1'b0 : n6345;
/* FF  2 20  2 */ always @(posedge clk) if (n126) n219 <= 1'b0 ? 1'b0 : n6346;
/* FF 20 23  0 */ assign n2384 = n6347;
/* FF  6 14  1 */ always @(posedge clk) if (n78) n624 <= 1'b0 ? 1'b0 : n6348;
/* FF 12 27  6 */ assign n6349 = n1560;
/* FF 18 17  3 */ always @(posedge clk) if (n1825) n2328 <= 1'b0 ? 1'b0 : n6350;
/* FF  6 19  6 */ assign n660 = n6351;
/* FF 11  8  3 */ always @(posedge clk) if (n1131) n1126 <= 1'b0 ? 1'b0 : n6352;
/* FF 29  5  3 */ always @(posedge clk) if (n3605) n3821 <= 1'b0 ? 1'b0 : n6353;
/* FF 19  9  1 */ always @(posedge clk) if (n2451) n2472 <= 1'b0 ? 1'b0 : n6354;
/* FF  4 10  0 */ always @(posedge clk) if (n251) n379 <= 1'b0 ? 1'b0 : n6355;
/* FF 24 16  4 */ always @(posedge clk) if (n3376) n3388 <= 1'b0 ? 1'b0 : n6356;
/* FF 27 22  7 */ always @(posedge clk) if (n3703) n3702 <= 1'b0 ? 1'b0 : n6357;
/* FF 10 16  2 */ always @(posedge clk) if (n891) n1025 <= 1'b0 ? 1'b0 : n6358;
/* FF 13 10  1 */ always @(posedge clk) if (n850) n1435 <= 1'b0 ? 1'b0 : n6359;
/* FF 18  3  6 */ assign \rco[92]  = n6360;
/* FF 15 28  2 */ always @(posedge clk) if (n1402) n1879 <= 1'b0 ? 1'b0 : n6361;
/* FF  7 16  4 */ always @(posedge clk) if (n630) n745 <= 1'b0 ? 1'b0 : n6362;
/* FF 21 11  3 */ always @(posedge clk) if (n2085) n2860 <= 1'b0 ? 1'b0 : n6363;
/* FF 18 12  7 */ always @(posedge clk) if (n1936) n2293 <= 1'b0 ? 1'b0 : n6364;
/* FF 21  6  4 */ always @(posedge clk) if (n2247) n2837 <= 1'b0 ? 1'b0 : n6365;
/* FF 12 22  0 */ always @(posedge clk) if (n1357) n1348 <= 1'b0 ? 1'b0 : n6366;
/* FF 26 15  1 */ always @(posedge clk) if (n3233) n3541 <= 1'b0 ? 1'b0 : n6367;
/* FF 14 12  3 */ assign n6368 = n1775;
/* FF 19 23  6 */ assign \rco[183]  = n6369;
/* FF 19 10  5 */ always @(posedge clk) if (n2678) n1934 <= 1'b0 ? 1'b0 : n6370;
/* FF  4 21  3 */ always @(posedge clk) if (n552) n450 <= 1'b0 ? 1'b0 : n6371;
/* FF  9 26  0 */ always @(posedge clk) if (n954) n942 <= 1'b0 ? 1'b0 : n6372;
/* FF 26 17  0 */ assign n3249 = n6373;
/* FF 12  4  1 */ assign \rco[149]  = n6374;
/* FF  6 10  6 */ always @(posedge clk) if (n589) n597 <= 1'b0 ? 1'b0 : n6375;
/* FF 20 11  7 */ always @(posedge clk) if (n2682) n2695 <= 1'b0 ? 1'b0 : n6376;
/* FF 17 14  3 */ always @(posedge clk) if (n1625) n2097 <= 1'b0 ? 1'b0 : n6377;
/* FF  5 13  5 */ always @(posedge clk) if (n402) n497 <= 1'b0 ? 1'b0 : n6378;
/* FF 19 24  4 */ always @(posedge clk) if (n2775) n2598 <= 1'b0 ? 1'b0 : n6379;
/* FF 11 20  6 */ always @(posedge clk) if (n1339) n1194 <= 1'b0 ? 1'b0 : n6380;
/* FF 29  9  4 */ always @(posedge clk) if (n3464) n3829 <= 1'b0 ? 1'b0 : n6381;
/* FF 28 23  2 */ always @(posedge clk) if (n3704) n3809 <= 1'b0 ? 1'b0 : n6382;
/* FF 11 27  7 */ always @(posedge clk) if (n1393) n1254 <= 1'b0 ? 1'b0 : n6383;
/* FF 21 26  2 */ assign n6384 = n3141;
/* FF 15 16  5 */ always @(posedge clk) if (n1500) n1798 <= 1'b0 ? 1'b0 : n6385;
/* FF 15 15  4 */ assign n1500 = n6386;
/* FF 18 16  0 */ assign \rco[30]  = n6387;
/* FF  6  9  0 */ assign n21 = n6388;
/* FF 20 22  3 */ always @(posedge clk) if (n2384) n2779 <= 1'b0 ? 1'b0 : n6389;
/* FF 12 26  5 */ always @(posedge clk) if (n1393) n1390 <= 1'b0 ? 1'b0 : n6390;
/* FF 17 24  3 */ always @(posedge clk) if (n2000) n2169 <= 1'b0 ? 1'b0 : n6391;
/* FF 19  6  0 */ always @(posedge clk) if (n2241) n2443 <= 1'b0 ? 1'b0 : n6392;
/* FF  4  9  1 */ always @(posedge clk) if (n260) n372 <= 1'b0 ? 1'b0 : n6393;
/* FF 10  6  4 */ always @(posedge clk) if (en_in) n974 <= 1'b0 ? 1'b0 : n6394;
/* FF 24 15  5 */ always @(posedge clk) if (n3233) n3380 <= 1'b0 ? 1'b0 : n6395;
/* FF 10 19  3 */ always @(posedge clk) if (n454) n1044 <= 1'b0 ? 1'b0 : n6396;
/* FF  9  9  7 */ always @(posedge clk) if (n983) n833 <= 1'b0 ? 1'b0 : n6397;
/* FF 13 11  6 */ always @(posedge clk) if (n1137) n1447 <= 1'b0 ? 1'b0 : n6398;
/* FF 18  2  1 */ always @(posedge clk) if (n2207) n2200 <= 1'b0 ? 1'b0 : n6399;
/* FF  7 17  3 */ always @(posedge clk) if (n549) n754 <= 1'b0 ? 1'b0 : n6400;
/* FF 21 12  2 */ always @(posedge clk) if (n3029) n2869 <= 1'b0 ? 1'b0 : n6401;
/* FF 18 15  6 */ always @(posedge clk) if (n1) n2313 <= 1'b0 ? 1'b0 : n6402;
/* FF 14 26  5 */ always @(posedge clk) if (n1271) n1716 <= 1'b0 ? 1'b0 : n6403;
/* FF 14 15  2 */ always @(posedge clk) if (n1792) n1641 <= 1'b0 ? 1'b0 : n6404;
/* FF  2  9  3 */ always @(posedge clk) if (n153) n160 <= 1'b0 ? 1'b0 : n6405;
/* FF 20  4  3 */ always @(posedge clk) if (n1761) n2653 <= 1'b0 ? 1'b0 : n6406;
/* FF 19 20  7 */ always @(posedge clk) if (n2553) n2572 <= 1'b0 ? 1'b0 : n6407;
/* FF 19 11  6 */ always @(posedge clk) if (n2076) n2492 <= 1'b0 ? 1'b0 : n6408;
/* FF 23  9  5 */ always @(posedge clk) if (n2678) n3181 <= 1'b0 ? 1'b0 : n6409;
/* FF 22 19  5 */ assign n6410 = n3262;
/* FF 24 18  5 */ always @(posedge clk) if (n3411) n3406 <= 1'b0 ? 1'b0 : n6411;
/* FF  3 17  4 */ always @(posedge clk) if (n79) n314 <= 1'b0 ? 1'b0 : n6412;
/* FF 14 25  1 */ always @(posedge clk) if (n697) n1702 <= 1'b0 ? 1'b0 : n6413;
/* FF  6 21  7 */ assign n673 = n6414;
/* FF 17  4  5 */ always @(posedge clk) if (n1761) n2035 <= 1'b0 ? 1'b0 : n6415;
/* FF 17 15  4 */ always @(posedge clk) if (n2111) n2105 <= 1'b0 ? 1'b0 : n6416;
/* FF 20 10  4 */ always @(posedge clk) if (n2697) n2687 <= 1'b0 ? 1'b0 : n6417;
/* FF 20  7  7 */ always @(posedge clk) if (n2670) n2668 <= 1'b0 ? 1'b0 : n6418;
/* FF  5 14  4 */ always @(posedge clk) if (n402) n508 <= 1'b0 ? 1'b0 : n6419;
/* FF 11 21  1 */ always @(posedge clk) if (n819) n769 <= 1'b0 ? 1'b0 : n6420;
/* FF 29 10  5 */ always @(posedge clk) if (n3464) n3837 <= 1'b0 ? 1'b0 : n6421;
/* FF 28 22  1 */ always @(posedge clk) if (n3704) n3800 <= 1'b0 ? 1'b0 : n6422;
/* FF 11 24  6 */ always @(posedge clk) if (n796) n1229 <= 1'b0 ? 1'b0 : n6423;
/* FF 16 17  3 */ always @(posedge clk) if (n2110) n1966 <= 1'b0 ? 1'b0 : n6424;
/* FF 21 27  5 */ always @(posedge clk) if (n2196) n2376 <= 1'b0 ? 1'b0 : n6425;
/* FF 27  6  2 */ assign n3594 = n6426;
/* FF 13 15  3 */ always @(posedge clk) if (n739) n1473 <= 1'b0 ? 1'b0 : n6427;
/* FF 30 12  7 */ always @(posedge clk) if (n3892) n3893 <= 1'b0 ? 1'b0 : n6428;
/* FF 15 17  2 */ always @(posedge clk) if (n1500) n1803 <= 1'b0 ? 1'b0 : n6429;
/* FF 18  6  6 */ always @(posedge clk) if (n2241) n2237 <= 1'b0 ? 1'b0 : n6430;
/* FF 18 19  1 */ always @(posedge clk) if (n1982) n2340 <= 1'b0 ? 1'b0 : n6431;
/* FF  3 18  6 */ always @(posedge clk) if (n215) n324 <= 1'b0 ? 1'b0 : n6432;
/* FF  6  8  3 */ always @(posedge clk) if (n570) n583 <= 1'b0 ? 1'b0 : n6433;
/* FF 20 21  2 */ always @(posedge clk) if (n2553) n2770 <= 1'b0 ? 1'b0 : n6434;
/* FF 12 25  4 */ always @(posedge clk) if (n1532) n1380 <= 1'b0 ? 1'b0 : n6435;
/* FF  1 19  4 */ always @(posedge clk) if (n119) n108 <= 1'b0 ? 1'b0 : n6436;
/* FF 17 25  0 */ always @(posedge clk) if (n2017) n2176 <= 1'b0 ? 1'b0 : n6437;
/* FF  5 16  0 */ always @(posedge clk) if (n511) n520 <= 1'b0 ? 1'b0 : n6438;
/* FF 19  7  3 */ always @(posedge clk) if (n2670) n2455 <= 1'b0 ? 1'b0 : n6439;
/* FF 23 13  2 */ always @(posedge clk) if (n3045) n3210 <= 1'b0 ? 1'b0 : n6440;
/* FF 10 25  5 */ always @(posedge clk) if (n567) n803 <= 1'b0 ? 1'b0 : n6441;
/* FF 24 14  6 */ always @(posedge clk) if (n3376) n3374 <= 1'b0 ? 1'b0 : n6442;
/* FF 27 20  5 */ always @(posedge clk) if (n3424) n3680 <= 1'b0 ? 1'b0 : n6443;
/* FF 10 18  4 */ always @(posedge clk) if (n1187) n1037 <= 1'b0 ? 1'b0 : n6444;
/* FF  9 10  6 */ always @(posedge clk) if (n988) n840 <= 1'b0 ? 1'b0 : n6445;
/* FF 18  5  0 */ always @(posedge clk) if (n2230) n2221 <= 1'b0 ? 1'b0 : n6446;
/* FF  7 22  2 */ always @(posedge clk) if (n695) n785 <= 1'b0 ? 1'b0 : n6447;
/* FF 20 27  1 */ always @(posedge clk) if (n2195) n2815 <= 1'b0 ? 1'b0 : n6448;
/* FF 21 13  1 */ always @(posedge clk) if (n2519) n2875 <= 1'b0 ? 1'b0 : n6449;
/* FF 14 21  4 */ assign n1356 = n6450;
/* FF 14 14  5 */ always @(posedge clk) if (n1791) n1130 <= 1'b0 ? 1'b0 : n6451;
/* FF  2  8  0 */ always @(posedge clk) if (n21) n155 <= 1'b0 ? 1'b0 : n6452;
/* FF  1 16  6 */ always @(posedge clk) if (n85) n93 <= 1'b0 ? 1'b0 : n6453;
/* FF  6 26  3 */ always @(posedge clk) if (n567) n699 <= 1'b0 ? 1'b0 : n6454;
/* FF 17 11  1 */ always @(posedge clk) if (n2076) n2067 <= 1'b0 ? 1'b0 : n6455;
/* FF 11 17  6 */ always @(posedge clk) if (n900) n1174 <= 1'b0 ? 1'b0 : n6456;
/* FF 10 11  4 */ always @(posedge clk) if (n996) n992 <= 1'b0 ? 1'b0 : n6457;
/* FF 19  8  7 */ always @(posedge clk) if (n2451) n2468 <= 1'b0 ? 1'b0 : n6458;
/* FF 19 21  0 */ always @(posedge clk) if (n2164) n2576 <= 1'b0 ? 1'b0 : n6459;
/* FF 23 14  4 */ always @(posedge clk) if (n2551) n3218 <= 1'b0 ? 1'b0 : n6460;
/* FF 24 17  4 */ always @(posedge clk) if (n2123) n3398 <= 1'b0 ? 1'b0 : n6461;
/* FF 28  7  1 */ always @(posedge clk) if (n3488) n3720 <= 1'b0 ? 1'b0 : n6462;
/* FF  3 14  0 */ assign \rco[12]  = n410;
/* FF 15 21  7 */ always @(posedge clk) if (n1356) n1686 <= 1'b0 ? 1'b0 : n6463;
/* FF 27  9  0 */ always @(posedge clk) if (n3621) n3610 <= 1'b0 ? 1'b0 : n6464;
/* FF 12 10  3 */ always @(posedge clk) if (n850) n1286 <= 1'b0 ? 1'b0 : n6465;
/* FF 26 19  2 */ always @(posedge clk) if (n2730) n3557 <= 1'b0 ? 1'b0 : n6466;
/* FF 14 24  2 */ assign n697 = n6467;
/* FF 17  5  6 */ assign \rco[179]  = n6468;
/* FF  6 20  4 */ always @(posedge clk) if (n552) n664 <= 1'b0 ? 1'b0 : n6469;
/* FF 20  9  5 */ assign n6470 = n2854;
/* FF 17  8  5 */ assign \rco[93]  = n2260;
/* FF  2  7  6 */ always @(posedge clk) if (n21) n151 <= 1'b0 ? 1'b0 : n6471;
/* FF 23 28  3 */ assign \rco[178]  = n6472;
/* FF 11 18  0 */ always @(posedge clk) if (n1187) n1179 <= 1'b0 ? 1'b0 : n6473;
/* FF 29 11  2 */ always @(posedge clk) if (n3751) n3841 <= 1'b0 ? 1'b0 : n6474;
/* FF 28 21  0 */ always @(posedge clk) if (n3788) n3791 <= 1'b0 ? 1'b0 : n6475;
/* FF  4 12  3 */ always @(posedge clk) if (n77) n396 <= 1'b0 ? 1'b0 : n6476;
/* FF 22 12  2 */ always @(posedge clk) if (n3029) n3038 <= 1'b0 ? 1'b0 : n6477;
/* FF 10 22  1 */ always @(posedge clk) if (n695) n550 <= 1'b0 ? 1'b0 : n6478;
/* FF 21 28  4 */ always @(posedge clk) if (n2196) n2983 <= 1'b0 ? 1'b0 : n6479;
/* FF 13 16  2 */ always @(posedge clk) if (n922) n1479 <= 1'b0 ? 1'b0 : n6480;
/* FF 27  7  1 */ always @(posedge clk) if (n3459) n3174 <= 1'b0 ? 1'b0 : n6481;
/* FF 15 22  3 */ always @(posedge clk) if (n1835) n1849 <= 1'b0 ? 1'b0 : n6482;
/* FF 18  9  7 */ always @(posedge clk) if (n2055) n2268 <= 1'b0 ? 1'b0 : n6483;
/* FF 18 18  6 */ always @(posedge clk) if (n1825) n2337 <= 1'b0 ? 1'b0 : n6484;
/* FF  3 19  5 */ always @(posedge clk) if (n115) n332 <= 1'b0 ? 1'b0 : n6485;
/* FF  6 11  2 */ always @(posedge clk) if (n286) n601 <= 1'b0 ? 1'b0 : n6486;
/* FF 12 24  3 */ always @(posedge clk) if (n961) n1370 <= 1'b0 ? 1'b0 : n6487;
/* FF 14 10  2 */ always @(posedge clk) if (n1622) n1606 <= 1'b0 ? 1'b0 : n6488;
/* FF 19 17  5 */ always @(posedge clk) if (n2727) n2546 <= 1'b0 ? 1'b0 : n6489;
/* FF 17 26  1 */ always @(posedge clk) if (n1557) n2185 <= 1'b0 ? 1'b0 : n6490;
/* FF 22 21  6 */ always @(posedge clk) if (n2564) n3102 <= 1'b0 ? 1'b0 : n6491;
/* FF  5 17  3 */ always @(posedge clk) if (n2) n527 <= 1'b0 ? 1'b0 : n6492;
/* FF  4 15  7 */ always @(posedge clk) if (n207) n419 <= 1'b0 ? 1'b0 : n6493;
/* FF 10 24  6 */ always @(posedge clk) if (n820) n1078 <= 1'b0 ? 1'b0 : n6494;
/* FF 24 13  7 */ always @(posedge clk) if (n3351) n3367 <= 1'b0 ? 1'b0 : n6495;
/* FF 28 11  4 */ always @(posedge clk) if (n3462) n3636 <= 1'b0 ? 1'b0 : n6496;
/* FF 27 21  2 */ always @(posedge clk) if (n3421) n3689 <= 1'b0 ? 1'b0 : n6497;
/* FF 10 21  5 */ always @(posedge clk) if (n818) n365 <= 1'b0 ? 1'b0 : n6498;
/* FF 13 13  4 */ always @(posedge clk) if (n1015) n1459 <= 1'b0 ? 1'b0 : n6499;
/* FF 18  4  3 */ always @(posedge clk) if (n2207) n2216 <= 1'b0 ? 1'b0 : n6500;
/* FF  7 23  1 */ always @(posedge clk) if (n454) n791 <= 1'b0 ? 1'b0 : n6501;
/* FF 20 26  2 */ always @(posedge clk) if (n2615) n2807 <= 1'b0 ? 1'b0 : n6502;
/* FF 21 14  0 */ always @(posedge clk) if (n2519) n2882 <= 1'b0 ? 1'b0 : n6503;
/* FF 14 20  7 */ always @(posedge clk) if (n1347) n1682 <= 1'b0 ? 1'b0 : n6504;
/* FF 17 20  0 */ always @(posedge clk) if (n1843) n2136 <= 1'b0 ? 1'b0 : n6505;
/* FF  2 11  1 */ always @(posedge clk) if (n168) n169 <= 1'b0 ? 1'b0 : n6506;
/* FF 19 18  1 */ always @(posedge clk) if (n2348) n2555 <= 1'b0 ? 1'b0 : n6507;
/* FF 10 10  3 */ always @(posedge clk) if (n983) n986 <= 1'b0 ? 1'b0 : n6508;
/* FF 23 15  7 */ always @(posedge clk) if (n3216) n3229 <= 1'b0 ? 1'b0 : n6509;
/* FF 28  6  2 */ always @(posedge clk) if (n3594) n3713 <= 1'b0 ? 1'b0 : n6510;
/* FF  3 15  3 */ always @(posedge clk) if (n207) n296 <= 1'b0 ? 1'b0 : n6511;
/* FF 21 16  3 */ always @(posedge clk) if (n2551) n2890 <= 1'b0 ? 1'b0 : n6512;
/* FF 15 10  6 */ always @(posedge clk) if (n1624) n1760 <= 1'b0 ? 1'b0 : n6513;
/* FF 26 18  5 */ assign \rco[31]  = n6514;
/* FF 18 22  3 */ assign n6515 = n2591;
/* FF 14 27  3 */ always @(posedge clk) if (n1402) n1720 <= 1'b0 ? 1'b0 : n6516;
/* FF  6 23  5 */ always @(posedge clk) if (n360) n692 <= 1'b0 ? 1'b0 : n6517;
/* FF 20  8  2 */ assign n2671 = n2844;
/* FF 17  9  6 */ assign n2056 = n6518;
/* FF 11 19  3 */ assign n1187 = n6519;
/* FF 29 12  3 */ always @(posedge clk) if (n3751) n3852 <= 1'b0 ? 1'b0 : n6520;
/* FF 22 26  4 */ always @(posedge clk) if (n2613) n3137 <= 1'b0 ? 1'b0 : n6521;
/* FF  9 12  7 */ always @(posedge clk) if (n996) n853 <= 1'b0 ? 1'b0 : n6522;
/* FF 27 17  7 */ always @(posedge clk) if (n3249) n3656 <= 1'b0 ? 1'b0 : n6523;
/* FF 22 15  3 */ always @(posedge clk) if (n3216) n3061 <= 1'b0 ? 1'b0 : n6524;
/* FF  7  6  4 */ always @(posedge clk) if (n588) n709 <= 1'b0 ? 1'b0 : n6525;
/* FF 13 17  1 */ always @(posedge clk) if (n1461) n1485 <= 1'b0 ? 1'b0 : n6526;
/* FF 15 23  0 */ assign \rco[115]  = n6527;
/* FF 18  8  4 */ always @(posedge clk) if (n2055) n2253 <= 1'b0 ? 1'b0 : n6528;
/* FF 18 21  7 */ always @(posedge clk) if (n2347) n2356 <= 1'b0 ? 1'b0 : n6529;
/* FF  3 16  4 */ always @(posedge clk) if (n197) n292 <= 1'b0 ? 1'b0 : n6530;
/* FF 14  5  3 */ always @(posedge clk) if (n1577) n1574 <= 1'b0 ? 1'b0 : n6531;
/* FF 19 14  4 */ always @(posedge clk) if (n2123) n2515 <= 1'b0 ? 1'b0 : n6532;
/* FF 22 20  5 */ always @(posedge clk) if (n3087) n3093 <= 1'b0 ? 1'b0 : n6533;
/* FF  5 18  2 */ always @(posedge clk) if (n657) n533 <= 1'b0 ? 1'b0 : n6534;
/* FF  4 14  4 */ assign n79 = n6535;
/* FF 19  5  5 */ always @(posedge clk) if (n2230) n2440 <= 1'b0 ? 1'b0 : n6536;
/* FF 10 27  7 */ always @(posedge clk) if (n804) n1099 <= 1'b0 ? 1'b0 : n6537;
/* FF 24 12  0 */ always @(posedge clk) if (n3351) n3353 <= 1'b0 ? 1'b0 : n6538;
/* FF 16 24  6 */ always @(posedge clk) if (n1557) n129 <= 1'b0 ? 1'b0 : n6539;
/* FF 22 25  6 */ always @(posedge clk) if (n2812) n3130 <= 1'b0 ? 1'b0 : n6540;
/* FF 10 20  6 */ always @(posedge clk) if (n922) n1053 <= 1'b0 ? 1'b0 : n6541;
/* FF 27 18  3 */ always @(posedge clk) if (n3553) n3660 <= 1'b0 ? 1'b0 : n6542;
/* FF 13 14  5 */ always @(posedge clk) if (n1461) n1467 <= 1'b0 ? 1'b0 : n6543;
/* FF 28 10  7 */ always @(posedge clk) if (n3462) n3748 <= 1'b0 ? 1'b0 : n6544;
/* FF 18  7  2 */ assign n2241 = n6545;
/* FF  7 20  0 */ assign n562 = n6546;
/* FF 20 25  3 */ always @(posedge clk) if (n2612) n2801 <= 1'b0 ? 1'b0 : n6547;
/* FF 26 22  2 */ always @(posedge clk) if (n2730) n3571 <= 1'b0 ? 1'b0 : n6548;
/* FF 15  5  4 */ always @(posedge clk) if (n1742) n1729 <= 1'b0 ? 1'b0 : n6549;
/* FF 14 23  6 */ assign n6550 = n1863;
/* FF 20 12  7 */ always @(posedge clk) if (n2682) n2705 <= 1'b0 ? 1'b0 : n6551;
/* FF 14  8  7 */ always @(posedge clk) if (n1741) n1600 <= 1'b0 ? 1'b0 : n6552;
/* FF 17 21  3 */ always @(posedge clk) if (n2347) n2147 <= 1'b0 ? 1'b0 : n6553;
/* FF  1 18  4 */ always @(posedge clk) if (n115) n101 <= 1'b0 ? 1'b0 : n6554;
/* FF 10 13  2 */ assign n996 = n6555;
/* FF 24 26  1 */ always @(posedge clk) if (n2613) n3453 <= 1'b0 ? 1'b0 : n6556;
/* FF 23 12  6 */ always @(posedge clk) if (n3031) n3205 <= 1'b0 ? 1'b0 : n6557;
/* FF 28  5  3 */ always @(posedge clk) if (n3488) n3708 <= 1'b0 ? 1'b0 : n6558;
/* FF  3 12  2 */ always @(posedge clk) if (n168) n279 <= 1'b0 ? 1'b0 : n6559;
/* FF 21 17  0 */ assign \rco[60]  = n6560;
/* FF 26 24  7 */ always @(posedge clk) if (n2730) n3583 <= 1'b0 ? 1'b0 : n6561;
/* FF 30 10  6 */ always @(posedge clk) if (n3892) n3890 <= 1'b0 ? 1'b0 : n6562;
/* FF 15 11  5 */ always @(posedge clk) if (n1624) n1768 <= 1'b0 ? 1'b0 : n6563;
/* FF 26 21  4 */ always @(posedge clk) if (n3421) n3566 <= 1'b0 ? 1'b0 : n6564;
/* FF 15  6  6 */ always @(posedge clk) if (n1744) n1739 <= 1'b0 ? 1'b0 : n6565;
/* FF 17  7  0 */ always @(posedge clk) if (n2045) n2046 <= 1'b0 ? 1'b0 : n6566;
/* FF 18 25  2 */ always @(posedge clk) if (n1878) n2379 <= 1'b0 ? 1'b0 : n6567;
/* FF  6 22  2 */ always @(posedge clk) if (n673) n680 <= 1'b0 ? 1'b0 : n6568;
/* FF 20 15  3 */ always @(posedge clk) if (n2715) n2720 <= 1'b0 ? 1'b0 : n6569;
/* FF 17 10  7 */ always @(posedge clk) if (n2282) n2066 <= 1'b0 ? 1'b0 : n6570;
/* FF 11 16  2 */ always @(posedge clk) if (n891) n1161 <= 1'b0 ? 1'b0 : n6571;
/* FF  1 12  0 */ always @(posedge clk) if (n39) n46 <= 1'b0 ? 1'b0 : n6572;
/* FF 24  8  5 */ assign n3330 = n6573;
/* FF 13  7  7 */ always @(posedge clk) if (n977) n1430 <= 1'b0 ? 1'b0 : n6574;
/* FF 22 14  4 */ always @(posedge clk) if (n3045) n3055 <= 1'b0 ? 1'b0 : n6575;
/* FF  7  7  7 */ always @(posedge clk) if (n588) n716 <= 1'b0 ? 1'b0 : n6576;
/* FF 13 18  0 */ always @(posedge clk) if (n1205) n1492 <= 1'b0 ? 1'b0 : n6577;
/* FF 27  5  7 */ always @(posedge clk) if (n3594) n3592 <= 1'b0 ? 1'b0 : n6578;
/* FF 30  9  0 */ assign \rco[72]  = n6579;
/* FF 15 20  1 */ always @(posedge clk) if (n1347) n1828 <= 1'b0 ? 1'b0 : n6580;
/* FF 18 11  5 */ assign \rco[41]  = n2496;
/* FF 18 20  4 */ assign n1843 = n6581;
/* FF 26  7  0 */ always @(posedge clk) if (n3603) n3481 <= 1'b0 ? 1'b0 : n6582;
/* FF 11 14  1 */ always @(posedge clk) if (n1154) n1147 <= 1'b0 ? 1'b0 : n6583;
/* FF  2 14  3 */ always @(posedge clk) if (n83) n190 <= 1'b0 ? 1'b0 : n6584;
/* FF 16  7  2 */ always @(posedge clk) if (n1743) n1909 <= 1'b0 ? 1'b0 : n6585;
/* FF 19 15  7 */ always @(posedge clk) if (n2715) n2532 <= 1'b0 ? 1'b0 : n6586;
/* FF 23  5  6 */ always @(posedge clk) if (n3158) n3156 <= 1'b0 ? 1'b0 : n6587;
/* FF 22 23  4 */ assign n3114 = n6588;
/* FF  5 19  5 */ always @(posedge clk) if (n349) n244 <= 1'b0 ? 1'b0 : n6589;
/* FF  4 13  5 */ assign n6590 = n503;
/* FF 19  2  4 */ always @(posedge clk) if (n2207) n2426 <= 1'b0 ? 1'b0 : n6591;
/* FF 10 26  0 */ assign n804 = n6592;
/* FF 24 11  1 */ assign \rco[63]  = n6593;
/* FF 13  4  3 */ assign \rco[165]  = n6594;
/* FF 22 24  5 */ always @(posedge clk) if (n3113) n3121 <= 1'b0 ? 1'b0 : n6595;
/* FF 10 23  7 */ always @(posedge clk) if (n821) n1068 <= 1'b0 ? 1'b0 : n6596;
/* FF 27 19  0 */ always @(posedge clk) if (n3553) n3667 <= 1'b0 ? 1'b0 : n6597;
/* FF 28  9  6 */ always @(posedge clk) if (n3621) n3739 <= 1'b0 ? 1'b0 : n6598;
/* FF  6  7  3 */ always @(posedge clk) if (n570) n574 <= 1'b0 ? 1'b0 : n6599;
/* FF 20 24  4 */ always @(posedge clk) if (n2775) n2792 <= 1'b0 ? 1'b0 : n6600;
/* FF 26  9  3 */ always @(posedge clk) if (n3460) n3501 <= 1'b0 ? 1'b0 : n6601;
/* FF 29 17  6 */ always @(posedge clk) if (n3765) n3859 <= 1'b0 ? 1'b0 : n6602;
/* FF 14 22  1 */ always @(posedge clk) if (n1402) n1688 <= 1'b0 ? 1'b0 : n6603;
/* FF 17  3  5 */ always @(posedge clk) if (n1887) n2030 <= 1'b0 ? 1'b0 : n6604;
/* FF  6 18  7 */ always @(posedge clk) if (n657) n656 <= 1'b0 ? 1'b0 : n6605;
/* FF 14 11  6 */ always @(posedge clk) if (n1622) n1617 <= 1'b0 ? 1'b0 : n6606;
/* FF 17 22  2 */ always @(posedge clk) if (n1999) n2154 <= 1'b0 ? 1'b0 : n6607;
/* FF 19 16  3 */ assign n2536 = n6608;
/* FF 23  6  0 */ always @(posedge clk) if (n3158) n3159 <= 1'b0 ? 1'b0 : n6609;
/* FF 11 28  5 */ always @(posedge clk) if (n1384) n1260 <= 1'b0 ? 1'b0 : n6610;
/* FF 10 12  1 */ always @(posedge clk) if (n996) n998 <= 1'b0 ? 1'b0 : n6611;
/* FF 24 25  0 */ always @(posedge clk) if (n2812) n3446 <= 1'b0 ? 1'b0 : n6612;
/* FF 16 26  3 */ always @(posedge clk) if (n1557) n2010 <= 1'b0 ? 1'b0 : n6613;
/* FF  4 19  1 */ assign \rco[131]  = n6614;
/* FF  3 13  5 */ assign n286 = n6615;
/* FF 21 18  1 */ always @(posedge clk) if (n2757) n2903 <= 1'b0 ? 1'b0 : n6616;
/* FF  9 28  2 */ always @(posedge clk) if (n961) n958 <= 1'b0 ? 1'b0 : n6617;
/* FF 22 10  1 */ always @(posedge clk) if (n2856) n3023 <= 1'b0 ? 1'b0 : n6618;
/* FF 15  8  4 */ always @(posedge clk) if (n1741) n810 <= 1'b0 ? 1'b0 : n6619;
/* FF 26 20  7 */ assign n2602 = n6620;
/* FF 12 15  4 */ always @(posedge clk) if (n1155) n1300 <= 1'b0 ? 1'b0 : n6621;
/* FF 15  7  5 */ assign n1743 = n6622;
/* FF 18 24  1 */ always @(posedge clk) if (n1878) n2371 <= 1'b0 ? 1'b0 : n6623;
/* FF 20 14  0 */ always @(posedge clk) if (n2682) n2712 <= 1'b0 ? 1'b0 : n6624;
/* FF 16  8  0 */ always @(posedge clk) if (n1625) n1915 <= 1'b0 ? 1'b0 : n6625;
/* FF  1 13  3 */ always @(posedge clk) if (n83) n62 <= 1'b0 ? 1'b0 : n6626;
/* FF  5 23  2 */ assign n563 = n6627;
/* FF  9 14  5 */ always @(posedge clk) if (n629) n864 <= 1'b0 ? 1'b0 : n6628;
/* FF 22  9  5 */ always @(posedge clk) if (n2989) n3019 <= 1'b0 ? 1'b0 : n6629;
/* FF 13 19  7 */ assign \rco[110]  = n6630;
/* FF 18 10  2 */ always @(posedge clk) if (n2282) n2275 <= 1'b0 ? 1'b0 : n6631;
/* FF  2 17  1 */ always @(posedge clk) if (n215) n102 <= 1'b0 ? 1'b0 : n6632;
/* FF 20 28  1 */ always @(posedge clk) if (n2195) n2823 <= 1'b0 ? 1'b0 : n6633;
/* FF 18 23  5 */ always @(posedge clk) if (n1999) n2361 <= 1'b0 ? 1'b0 : n6634;
/* FF 14 18  6 */ always @(posedge clk) if (n1672) n1665 <= 1'b0 ? 1'b0 : n6635;
/* FF 12 29  0 */ always @(posedge clk) if (n1532) n1403 <= 1'b0 ? 1'b0 : n6636;
/* FF 11 15  2 */ assign n1154 = n6637;
/* FF 14  7  1 */ always @(posedge clk) if (n1743) n1586 <= 1'b0 ? 1'b0 : n6638;
/* FF 16  6  1 */ always @(posedge clk) if (n1744) n1898 <= 1'b0 ? 1'b0 : n6639;
/* FF 19 12  6 */ always @(posedge clk) if (n1936) n2503 <= 1'b0 ? 1'b0 : n6640;
/* FF 23 10  7 */ always @(posedge clk) if (n2697) n2858 <= 1'b0 ? 1'b0 : n6641;
/* FF 22 22  3 */ always @(posedge clk) if (n2961) n3108 <= 1'b0 ? 1'b0 : n6642;
/* FF 19  3  7 */ always @(posedge clk) if (n1887) n2212 <= 1'b0 ? 1'b0 : n6643;
/* FF 22 27  4 */ always @(posedge clk) if (n2970) n3147 <= 1'b0 ? 1'b0 : n6644;
/* FF 10 29  1 */ always @(posedge clk) if (n821) n1070 <= 1'b0 ? 1'b0 : n6645;
/* FF 24 10  2 */ always @(posedge clk) if (n3352) n3342 <= 1'b0 ? 1'b0 : n6646;
/* FF 13  5  0 */ always @(posedge clk) if (n1577) n1410 <= 1'b0 ? 1'b0 : n6647;
/* FF 28  8  1 */ always @(posedge clk) if (n3605) n3727 <= 1'b0 ? 1'b0 : n6648;
/* FF  3  9  2 */ always @(posedge clk) if (n260) n254 <= 1'b0 ? 1'b0 : n6649;
/* FF  9 19  0 */ always @(posedge clk) if (n454) n901 <= 1'b0 ? 1'b0 : n6650;
/* FF 12 19  3 */ always @(posedge clk) if (n1501) n1331 <= 1'b0 ? 1'b0 : n6651;
/* FF 26  8  0 */ always @(posedge clk) if (n3603) n3490 <= 1'b0 ? 1'b0 : n6652;
/* FF 14 17  0 */ always @(posedge clk) if (n1672) n1654 <= 1'b0 ? 1'b0 : n6653;
/* FF 17 12  4 */ always @(posedge clk) if (n2056) n2081 <= 1'b0 ? 1'b0 : n6654;
/* FF  2 12  4 */ always @(posedge clk) if (n39) n180 <= 1'b0 ? 1'b0 : n6655;
/* FF 23  7  3 */ always @(posedge clk) if (n3006) n3169 <= 1'b0 ? 1'b0 : n6656;
/* FF 11 29  2 */ always @(posedge clk) if (n1384) n1264 <= 1'b0 ? 1'b0 : n6657;
/* FF 10 15  0 */ always @(posedge clk) if (n750) n749 <= 1'b0 ? 1'b0 : n6658;
/* FF 16 25  2 */ always @(posedge clk) if (n1557) n2005 <= 1'b0 ? 1'b0 : n6659;
/* FF 21 24  7 */ always @(posedge clk) if (n3113) n2960 <= 1'b0 ? 1'b0 : n6660;
/* FF  4 18  2 */ always @(posedge clk) if (n349) n432 <= 1'b0 ? 1'b0 : n6661;
/* FF  3 10  4 */ always @(posedge clk) if (n251) n266 <= 1'b0 ? 1'b0 : n6662;
/* FF 21 19  6 */ always @(posedge clk) if (n2757) n2916 <= 1'b0 ? 1'b0 : n6663;
/* FF 13 23  4 */ always @(posedge clk) if (n1069) n1528 <= 1'b0 ? 1'b0 : n6664;
/* FF 27 14  5 */ always @(posedge clk) if (n3527) n3646 <= 1'b0 ? 1'b0 : n6665;
/* FF 15  9  3 */ always @(posedge clk) if (n1624) n1753 <= 1'b0 ? 1'b0 : n6666;
/* FF 18 14  7 */ always @(posedge clk) if (n2045) n2305 <= 1'b0 ? 1'b0 : n6667;
/* FF 12 14  7 */ always @(posedge clk) if (n1154) n1295 <= 1'b0 ? 1'b0 : n6668;
/* FF 26 23  6 */ always @(posedge clk) if (n3703) n3581 <= 1'b0 ? 1'b0 : n6669;
/* FF 18 27  0 */ always @(posedge clk) if (n2020) n2393 <= 1'b0 ? 1'b0 : n6670;
/* FF  6 16  0 */ always @(posedge clk) if (n511) n638 <= 1'b0 ? 1'b0 : n6671;
/* FF 20 13  1 */ assign n2708 = n6672;
/* FF 23 21  0 */ always @(posedge clk) if (n3258) n3271 <= 1'b0 ? 1'b0 : n6673;
/* FF  4 11  6 */ always @(posedge clk) if (n184) n391 <= 1'b0 ? 1'b0 : n6674;
/* FF 16 23  1 */ always @(posedge clk) if (n2000) n1992 <= 1'b0 ? 1'b0 : n6675;
/* FF  1 14  2 */ always @(posedge clk) if (n85) n70 <= 1'b0 ? 1'b0 : n6676;
/* FF 22  7  7 */ always @(posedge clk) if (n2841) n3005 <= 1'b0 ? 1'b0 : n6677;
/* FF 10 17  4 */ always @(posedge clk) if (n629) n1031 <= 1'b0 ? 1'b0 : n6678;
/* FF  9 15  2 */ always @(posedge clk) if (n645) n869 <= 1'b0 ? 1'b0 : n6679;
/* FF 24  6  7 */ always @(posedge clk) if (n3006) n3328 <= 1'b0 ? 1'b0 : n6680;
/* FF 22  8  6 */ always @(posedge clk) if (n2989) n3014 <= 1'b0 ? 1'b0 : n6681;
/* FF 28 12  6 */ always @(posedge clk) if (n3462) n3759 <= 1'b0 ? 1'b0 : n6682;
/* FF 13 20  6 */ always @(posedge clk) if (n1339) n1509 <= 1'b0 ? 1'b0 : n6683;
/* FF 31 17  0 */ always @(posedge clk) if (n3249) n3773 <= 1'b0 ? 1'b0 : n6684;
/* FF 18 13  3 */ always @(posedge clk) if (n2283) n2298 <= 1'b0 ? 1'b0 : n6685;
/* FF 20 19  0 */ always @(posedge clk) if (n2562) n2749 <= 1'b0 ? 1'b0 : n6686;
/* FF 14 13  7 */ always @(posedge clk) if (n1015) n1630 <= 1'b0 ? 1'b0 : n6687;
/* FF 14  6  6 */ always @(posedge clk) if (n1577) n1581 <= 1'b0 ? 1'b0 : n6688;
/* FF 16  5  0 */ always @(posedge clk) if (n1742) n1888 <= 1'b0 ? 1'b0 : n6689;
/* FF 17 19  2 */ always @(posedge clk) if (n1982) n2130 <= 1'b0 ? 1'b0 : n6690;
/* FF 19 13  1 */ always @(posedge clk) if (n2283) n2506 <= 1'b0 ? 1'b0 : n6691;
/* FF 23 11  4 */ always @(posedge clk) if (n3031) n3194 <= 1'b0 ? 1'b0 : n6692;
/* FF 22 17  2 */ always @(posedge clk) if (n3065) n3074 <= 1'b0 ? 1'b0 : n6693;
/* FF 10 28  2 */ always @(posedge clk) if (n821) n1103 <= 1'b0 ? 1'b0 : n6694;
/* FF 24  9  3 */ always @(posedge clk) if (n3352) n3335 <= 1'b0 ? 1'b0 : n6695;
/* FF 13  6  1 */ always @(posedge clk) if (n977) n1416 <= 1'b0 ? 1'b0 : n6696;
/* FF 15 24  2 */ always @(posedge clk) if (n778) n1866 <= 1'b0 ? 1'b0 : n6697;
/* FF 21 23  3 */ always @(posedge clk) if (n2961) n2946 <= 1'b0 ? 1'b0 : n6698;
/* FF 12 18  0 */ always @(posedge clk) if (n1501) n1320 <= 1'b0 ? 1'b0 : n6699;
/* FF 26 11  1 */ assign \rco[68]  = n6700;
/* FF 30 21  2 */ always @(posedge clk) if (n2730) n2549 <= 1'b0 ? 1'b0 : n6701;
/* FF 14 16  3 */ always @(posedge clk) if (n1792) n1649 <= 1'b0 ? 1'b0 : n6702;
/* FF 17 13  7 */ always @(posedge clk) if (n2056) n2093 <= 1'b0 ? 1'b0 : n6703;
/* FF 29 19  0 */ always @(posedge clk) if (n3786) n3861 <= 1'b0 ? 1'b0 : n6704;
/* FF 17 16  4 */ assign n2111 = n6705;
/* FF  2 15  5 */ always @(posedge clk) if (n197) n200 <= 1'b0 ? 1'b0 : n6706;
/* FF 11 26  3 */ always @(posedge clk) if (n954) n1239 <= 1'b0 ? 1'b0 : n6707;
/* FF 21 25  4 */ always @(posedge clk) if (n2970) n2966 <= 1'b0 ? 1'b0 : n6708;
/* FF  9 11  7 */ always @(posedge clk) if (n988) n849 <= 1'b0 ? 1'b0 : n6709;
/* FF  4 17  3 */ always @(posedge clk) if (n2) n427 <= 1'b0 ? 1'b0 : n6710;
/* FF  3 11  7 */ always @(posedge clk) if (n153) n276 <= 1'b0 ? 1'b0 : n6711;
/* FF  7  9  6 */ always @(posedge clk) if (n589) n724 <= 1'b0 ? 1'b0 : n6712;
/* FF 21 20  7 */ always @(posedge clk) if (n3087) n2925 <= 1'b0 ? 1'b0 : n6713;
/* FF 13 24  5 */ assign n961 = n6714;
/* FF 15 14  2 */ always @(posedge clk) if (n1791) n1785 <= 1'b0 ? 1'b0 : n6715;
/* FF 18 17  6 */ always @(posedge clk) if (n1825) n2331 <= 1'b0 ? 1'b0 : n6716;
/* FF 18 26  7 */ always @(posedge clk) if (n2615) n2392 <= 1'b0 ? 1'b0 : n6717;
/* FF  6 19  1 */ assign n6718 = n765;
/* FF 23 26  1 */ always @(posedge clk) if (n2195) n2830 <= 1'b0 ? 1'b0 : n6719;
/* FF 28 19  2 */ always @(posedge clk) if (n3424) n3779 <= 1'b0 ? 1'b0 : n6720;
/* FF 19  9  6 */ always @(posedge clk) if (n2451) n2477 <= 1'b0 ? 1'b0 : n6721;
/* FF  4 10  5 */ always @(posedge clk) if (n251) n384 <= 1'b0 ? 1'b0 : n6722;
/* FF 16 22  2 */ always @(posedge clk) if (n1835) n1988 <= 1'b0 ? 1'b0 : n6723;
/* FF 22  6  0 */ always @(posedge clk) if (n2841) n2990 <= 1'b0 ? 1'b0 : n6724;
/* FF 10 16  7 */ always @(posedge clk) if (n891) n1029 <= 1'b0 ? 1'b0 : n6725;
/* FF 13 10  4 */ always @(posedge clk) if (n850) n1438 <= 1'b0 ? 1'b0 : n6726;
/* FF 22 11  7 */ assign n3029 = n6727;
/* FF 13 21  5 */ always @(posedge clk) if (n1356) n667 <= 1'b0 ? 1'b0 : n6728;
/* FF 18 12  0 */ always @(posedge clk) if (n1936) n2286 <= 1'b0 ? 1'b0 : n6729;
/* FF  2 19  3 */ assign n6730 = n340;
/* FF  6 13  0 */ always @(posedge clk) if (n78) n615 <= 1'b0 ? 1'b0 : n6731;
/* FF 20 18  3 */ always @(posedge clk) if (n2348) n2744 <= 1'b0 ? 1'b0 : n6732;
/* FF 11  6  5 */ always @(posedge clk) if (en_in) \rco[0]  <= 1'b0 ? 1'b0 : n6733;
/* FF 14 12  4 */ assign n1622 = n1776;
/* FF 11 13  4 */ always @(posedge clk) if (n733) n1142 <= 1'b0 ? 1'b0 : n6734;
/* FF 19 10  0 */ always @(posedge clk) if (n2678) n2479 <= 1'b0 ? 1'b0 : n6735;
/* FF 22 16  1 */ always @(posedge clk) if (n2551) n3071 <= 1'b0 ? 1'b0 : n6736;
/* FF  5 22  6 */ always @(posedge clk) if (n673) n560 <= 1'b0 ? 1'b0 : n6737;
/* FF 28 14  3 */ always @(posedge clk) if (n2085) n3764 <= 1'b0 ? 1'b0 : n6738;
/* FF 15 25  5 */ assign \rco[195]  = n6739;
/* FF  7 13  3 */ assign \rco[159]  = n6740;
/* FF 12 17  1 */ always @(posedge clk) if (n900) n1313 <= 1'b0 ? 1'b0 : n6741;
/* FF 18 30  4 */ always @(posedge clk) if (n1881) n2421 <= 1'b0 ? 1'b0 : n6742;
/* FF 14 19  2 */ always @(posedge clk) if (n1672) n1667 <= 1'b0 ? 1'b0 : n6743;
/* FF 17 14  6 */ always @(posedge clk) if (n1625) n2100 <= 1'b0 ? 1'b0 : n6744;
/* FF 29 20  1 */ always @(posedge clk) if (n3786) n3869 <= 1'b0 ? 1'b0 : n6745;
/* FF 17 17  7 */ always @(posedge clk) if (n2111) n2121 <= 1'b0 ? 1'b0 : n6746;
/* FF 11 27  0 */ always @(posedge clk) if (n1393) n1247 <= 1'b0 ? 1'b0 : n6747;
/* FF  1 11  2 */ assign n39 = n6748;
/* FF 21 26  5 */ assign n2971 = n6749;
/* FF  4 16  4 */ always @(posedge clk) if (n79) n424 <= 1'b0 ? 1'b0 : n6750;
/* FF 21 21  4 */ always @(posedge clk) if (n2564) n2930 <= 1'b0 ? 1'b0 : n6751;
/* FF 13 25  6 */ always @(posedge clk) if (n697) n1540 <= 1'b0 ? 1'b0 : n6752;
/* FF 27 12  7 */ always @(posedge clk) if (n3368) n3635 <= 1'b0 ? 1'b0 : n6753;
/* FF 18 16  5 */ always @(posedge clk) if (n2540) n2319 <= 1'b0 ? 1'b0 : n6754;
/* FF 18 29  6 */ always @(posedge clk) if (n1881) n2414 <= 1'b0 ? 1'b0 : n6755;
/* FF 23 27  2 */ always @(posedge clk) if (n2017) n3314 <= 1'b0 ? 1'b0 : n6756;
/* FF 28 18  1 */ always @(posedge clk) if (n3765) n3774 <= 1'b0 ? 1'b0 : n6757;
/* FF 19  6  7 */ always @(posedge clk) if (n2241) n2450 <= 1'b0 ? 1'b0 : n6758;
/* FF  4  9  4 */ always @(posedge clk) if (n260) n375 <= 1'b0 ? 1'b0 : n6759;
/* FF  1  8  4 */ always @(posedge clk) if (n37) n18 <= 1'b0 ? 1'b0 : n6760;
/* FF 10 19  6 */ always @(posedge clk) if (n454) n776 <= 1'b0 ? 1'b0 : n6761;
/* FF  9  9  0 */ always @(posedge clk) if (n983) n827 <= 1'b0 ? 1'b0 : n6762;
/* FF 13 11  3 */ always @(posedge clk) if (n1137) n1444 <= 1'b0 ? 1'b0 : n6763;
/* FF 13 22  4 */ assign n1069 = n6764;
/* FF 18 15  1 */ always @(posedge clk) if (n1) n2309 <= 1'b0 ? 1'b0 : n6765;
/* FF  2 18  4 */ always @(posedge clk) if (n115) n213 <= 1'b0 ? 1'b0 : n6766;
/* FF  6 12  3 */ always @(posedge clk) if (n286) n609 <= 1'b0 ? 1'b0 : n6767;
/* FF 20 17  2 */ always @(posedge clk) if (n2727) n2734 <= 1'b0 ? 1'b0 : n6768;
/* FF 26 14  3 */ always @(posedge clk) if (n3527) n3536 <= 1'b0 ? 1'b0 : n6769;
/* FF 14 15  5 */ always @(posedge clk) if (n1792) n1175 <= 1'b0 ? 1'b0 : n6770;
/* FF  2  9  6 */ always @(posedge clk) if (n153) n163 <= 1'b0 ? 1'b0 : n6771;
/* FF 19 11  3 */ always @(posedge clk) if (n2076) n2489 <= 1'b0 ? 1'b0 : n6772;
/* FF 23  9  2 */ always @(posedge clk) if (n2678) n3178 <= 1'b0 ? 1'b0 : n6773;
/* FF 22 19  0 */ assign n2573 = n6774;
/* FF 21  9  1 */ always @(posedge clk) if (n2856) n2846 <= 1'b0 ? 1'b0 : n6775;
/* FF  9 27  4 */ always @(posedge clk) if (n804) n950 <= 1'b0 ? 1'b0 : n6776;
/* FF 12 16  6 */ always @(posedge clk) if (n1155) n1309 <= 1'b0 ? 1'b0 : n6777;
/* FF 26 13  7 */ always @(posedge clk) if (n3033) n3532 <= 1'b0 ? 1'b0 : n6778;
/* FF 17 15  1 */ always @(posedge clk) if (n2111) n2102 <= 1'b0 ? 1'b0 : n6779;
/* FF 20  7  2 */ always @(posedge clk) if (n2670) n2663 <= 1'b0 ? 1'b0 : n6780;
/* FF 19 25  0 */ always @(posedge clk) if (n2612) n2604 <= 1'b0 ? 1'b0 : n6781;
/* FF 11 24  1 */ always @(posedge clk) if (n796) n1224 <= 1'b0 ? 1'b0 : n6782;
/* FF 22 13  4 */ always @(posedge clk) if (n2085) n3047 <= 1'b0 ? 1'b0 : n6783;
/* FF 21 27  2 */ always @(posedge clk) if (n2196) n2974 <= 1'b0 ? 1'b0 : n6784;
/* FF  4 23  5 */ assign \rco[135]  = n6785;
/* FF  7 15  4 */ assign \rco[23]  = n816;
/* FF  9 24  6 */ always @(posedge clk) if (n820) n938 <= 1'b0 ? 1'b0 : n6786;
/* FF 13 26  7 */ always @(posedge clk) if (n1271) n1550 <= 1'b0 ? 1'b0 : n6787;
/* FF 21 22  5 */ always @(posedge clk) if (n2384) n2589 <= 1'b0 ? 1'b0 : n6788;
/* FF 27 13  0 */ always @(posedge clk) if (n3460) n3637 <= 1'b0 ? 1'b0 : n6789;
/* FF 15 12  0 */ always @(posedge clk) if (n1625) n1762 <= 1'b0 ? 1'b0 : n6790;
/* FF 18 19  4 */ always @(posedge clk) if (n1982) n2343 <= 1'b0 ? 1'b0 : n6791;
/* FF  2 22  1 */ always @(posedge clk) if (n352) n236 <= 1'b0 ? 1'b0 : n6792;
/* FF 18 28  5 */ always @(posedge clk) if (n2020) n2405 <= 1'b0 ? 1'b0 : n6793;
/* FF 23 24  3 */ always @(posedge clk) if (n3112) n3299 <= 1'b0 ? 1'b0 : n6794;
/* FF 11 22  0 */ always @(posedge clk) if (n695) n1206 <= 1'b0 ? 1'b0 : n6795;
/* FF 28 17  0 */ always @(posedge clk) if (n3765) n3766 <= 1'b0 ? 1'b0 : n6796;
/* FF 16 15  5 */ always @(posedge clk) if (n739) n812 <= 1'b0 ? 1'b0 : n6797;
/* FF 19  7  4 */ always @(posedge clk) if (n2670) n2456 <= 1'b0 ? 1'b0 : n6798;
/* FF 23 13  7 */ always @(posedge clk) if (n3045) n3215 <= 1'b0 ? 1'b0 : n6799;
/* FF 16 20  4 */ always @(posedge clk) if (n1843) n1978 <= 1'b0 ? 1'b0 : n6800;
/* FF 10 18  1 */ always @(posedge clk) if (n1187) n1034 <= 1'b0 ? 1'b0 : n6801;
/* FF  9 10  1 */ always @(posedge clk) if (n988) n835 <= 1'b0 ? 1'b0 : n6802;
/* FF 13 12  2 */ always @(posedge clk) if (n1137) n1451 <= 1'b0 ? 1'b0 : n6803;
/* FF 15 18  3 */ always @(posedge clk) if (n1355) n1811 <= 1'b0 ? 1'b0 : n6804;
/* FF 20 27  4 */ always @(posedge clk) if (n2195) n2818 <= 1'b0 ? 1'b0 : n6805;
/* FF  2 21  5 */ always @(posedge clk) if (n126) n232 <= 1'b0 ? 1'b0 : n6806;
/* FF  6 15  2 */ always @(posedge clk) if (n630) n632 <= 1'b0 ? 1'b0 : n6807;
/* FF 12 20  3 */ assign \rco[118]  = n1512;
/* FF 14 14  2 */ always @(posedge clk) if (n1791) n1634 <= 1'b0 ? 1'b0 : n6808;
/* FF 17 11  6 */ always @(posedge clk) if (n2076) n2072 <= 1'b0 ? 1'b0 : n6809;
/* FF 17 30  1 */ always @(posedge clk) if (n2020) n2198 <= 1'b0 ? 1'b0 : n6810;
/* FF 19  8  2 */ always @(posedge clk) if (n2451) n2463 <= 1'b0 ? 1'b0 : n6811;
/* FF 23 14  3 */ always @(posedge clk) if (n2551) n3217 <= 1'b0 ? 1'b0 : n6812;
/* FF  3 14  7 */ assign \rco[8]  = n6813;
/* FF  7 19  1 */ always @(posedge clk) if (n549) n336 <= 1'b0 ? 1'b0 : n6814;
/* FF  9 20  5 */ always @(posedge clk) if (n961) n909 <= 1'b0 ? 1'b0 : n6815;
/* FF 21 10  0 */ assign \rco[52]  = n6816;
/* FF 12 10  4 */ always @(posedge clk) if (n850) n1287 <= 1'b0 ? 1'b0 : n6817;
/* FF 26 19  5 */ always @(posedge clk) if (n2730) n3560 <= 1'b0 ? 1'b0 : n6818;
/* FF 27  9  5 */ always @(posedge clk) if (n3621) n3615 <= 1'b0 ? 1'b0 : n6819;
/* FF 12 23  7 */ always @(posedge clk) if (n1357) n1365 <= 1'b0 ? 1'b0 : n6820;
/* FF 26 12  4 */ always @(posedge clk) if (n3368) n3521 <= 1'b0 ? 1'b0 : n6821;
/* FF 29 22  3 */ always @(posedge clk) if (n3788) n3882 <= 1'b0 ? 1'b0 : n6822;
/* FF 17  8  0 */ always @(posedge clk) if (n1741) n1603 <= 1'b0 ? 1'b0 : n6823;
/* FF 20  6  1 */ always @(posedge clk) if (n2247) n2660 <= 1'b0 ? 1'b0 : n6824;
/* FF  5 15  0 */ assign n511 = n6825;
/* FF 19 22  1 */ always @(posedge clk) if (n2164) n2585 <= 1'b0 ? 1'b0 : n6826;
/* FF 16 16  1 */ always @(posedge clk) if (n2110) n1956 <= 1'b0 ? 1'b0 : n6827;
/* FF 22 12  7 */ always @(posedge clk) if (n3029) n3043 <= 1'b0 ? 1'b0 : n6828;
/* FF 21 28  3 */ always @(posedge clk) if (n2196) n2982 <= 1'b0 ? 1'b0 : n6829;
/* FF  4 22  6 */ assign n455 = n6830;
/* FF  9 25  5 */ always @(posedge clk) if (n2) n940 <= 1'b0 ? 1'b0 : n6831;
/* FF 13 27  0 */ assign n1271 = n6832;
/* FF 20 20  2 */ always @(posedge clk) if (n2562) n2763 <= 1'b0 ? 1'b0 : n6833;
/* FF 23 18  5 */ always @(posedge clk) if (n2573) n1409 <= 1'b0 ? 1'b0 : n6834;
/* FF 14 10  7 */ always @(posedge clk) if (n1622) n1611 <= 1'b0 ? 1'b0 : n6835;
/* FF 23 25  4 */ always @(posedge clk) if (n2613) n3306 <= 1'b0 ? 1'b0 : n6836;
/* FF 11 23  3 */ always @(posedge clk) if (n796) n1217 <= 1'b0 ? 1'b0 : n6837;
/* FF  5 17  4 */ always @(posedge clk) if (n2) n528 <= 1'b0 ? 1'b0 : n6838;
/* FF  4 15  2 */ always @(posedge clk) if (n207) n414 <= 1'b0 ? 1'b0 : n6839;
/* FF 19  4  5 */ assign \rco[146]  = n6840;
/* FF 16 19  5 */ always @(posedge clk) if (n1402) n1972 <= 1'b0 ? 1'b0 : n6841;
/* FF 10 21  0 */ always @(posedge clk) if (n818) n1058 <= 1'b0 ? 1'b0 : n6842;
/* FF 13 13  1 */ always @(posedge clk) if (n1015) n1456 <= 1'b0 ? 1'b0 : n6843;
/* FF 15 19  0 */ always @(posedge clk) if (n1355) n1817 <= 1'b0 ? 1'b0 : n6844;
/* FF 20 26  7 */ always @(posedge clk) if (n2615) n2811 <= 1'b0 ? 1'b0 : n6845;
/* FF  2 20  6 */ always @(posedge clk) if (n126) n222 <= 1'b0 ? 1'b0 : n6846;
/* FF  6 14  5 */ always @(posedge clk) if (n78) n627 <= 1'b0 ? 1'b0 : n6847;
/* FF 20 23  4 */ assign n2003 = n2953;
/* FF 12 27  2 */ assign n1393 = n6848;
/* FF 17 20  7 */ always @(posedge clk) if (n1843) n2143 <= 1'b0 ? 1'b0 : n6849;
/* FF  2 11  4 */ always @(posedge clk) if (n168) n172 <= 1'b0 ? 1'b0 : n6850;
/* FF 11  8  7 */ always @(posedge clk) if (n1131) n1129 <= 1'b0 ? 1'b0 : n6851;
/* FF 29  5  7 */ always @(posedge clk) if (n3605) n3618 <= 1'b0 ? 1'b0 : n6852;
/* FF 23 15  0 */ always @(posedge clk) if (n3216) n3222 <= 1'b0 ? 1'b0 : n6853;
/* FF 24 16  0 */ always @(posedge clk) if (n3376) n3384 <= 1'b0 ? 1'b0 : n6854;
/* FF 27 22  3 */ always @(posedge clk) if (n3703) n3698 <= 1'b0 ? 1'b0 : n6855;
/* FF  3 15  4 */ always @(posedge clk) if (n207) n297 <= 1'b0 ? 1'b0 : n6856;
/* FF 21 16  6 */ always @(posedge clk) if (n2551) n2893 <= 1'b0 ? 1'b0 : n6857;
/* FF 18  3  2 */ assign \rco[89]  = n6858;
/* FF  7 16  0 */ always @(posedge clk) if (n630) n741 <= 1'b0 ? 1'b0 : n6859;
/* FF  9 21  6 */ always @(posedge clk) if (n818) n920 <= 1'b0 ? 1'b0 : n6860;
/* FF 21 11  7 */ always @(posedge clk) if (n2085) n2864 <= 1'b0 ? 1'b0 : n6861;
/* FF 26 18  2 */ assign n6862 = n3665;
/* FF 12 22  4 */ always @(posedge clk) if (n1357) n1352 <= 1'b0 ? 1'b0 : n6863;
/* FF 26 15  5 */ always @(posedge clk) if (n3233) n3545 <= 1'b0 ? 1'b0 : n6864;
/* FF 17  9  3 */ assign n1761 = n6865;
/* FF 20  5  0 */ always @(posedge clk) if (n2247) n2657 <= 1'b0 ? 1'b0 : n6866;
/* FF 19 23  2 */ assign n6867 = n2786;
/* FF 28 20  4 */ assign n3788 = n6868;
/* FF  4 24  0 */ assign \rco[125]  = n6869;
/* FF 22 15  6 */ always @(posedge clk) if (n3216) n3063 <= 1'b0 ? 1'b0 : n6870;
/* FF  7  6  3 */ always @(posedge clk) if (n588) n708 <= 1'b0 ? 1'b0 : n6871;
/* FF  9  7  3 */ always @(posedge clk) if (n588) n826 <= 1'b0 ? 1'b0 : n6872;
/* FF  4 21  7 */ always @(posedge clk) if (n552) n453 <= 1'b0 ? 1'b0 : n6873;
/* FF 13 28  1 */ always @(posedge clk) if (n1394) n1562 <= 1'b0 ? 1'b0 : n6874;
/* FF 27 11  2 */ always @(posedge clk) if (n3460) n3623 <= 1'b0 ? 1'b0 : n6875;
/* FF 18 21  2 */ always @(posedge clk) if (n2347) n2351 <= 1'b0 ? 1'b0 : n6876;
/* FF  6 10  2 */ always @(posedge clk) if (n589) n593 <= 1'b0 ? 1'b0 : n6877;
/* FF 20 11  3 */ always @(posedge clk) if (n2682) n2691 <= 1'b0 ? 1'b0 : n6878;
/* FF 23 19  6 */ always @(posedge clk) if (n2573) n3256 <= 1'b0 ? 1'b0 : n6879;
/* FF 11 20  2 */ always @(posedge clk) if (n1339) n1191 <= 1'b0 ? 1'b0 : n6880;
/* FF 29  9  0 */ assign \rco[75]  = n6881;
/* FF 17 27  3 */ always @(posedge clk) if (n1) n2191 <= 1'b0 ? 1'b0 : n6882;
/* FF 28 23  6 */ always @(posedge clk) if (n3704) n3812 <= 1'b0 ? 1'b0 : n6883;
/* FF  5 18  5 */ always @(posedge clk) if (n657) n536 <= 1'b0 ? 1'b0 : n6884;
/* FF  4 14  1 */ assign n207 = n6885;
/* FF 19  5  2 */ always @(posedge clk) if (n2230) n2437 <= 1'b0 ? 1'b0 : n6886;
/* FF 10 20  3 */ always @(posedge clk) if (n922) n1051 <= 1'b0 ? 1'b0 : n6887;
/* FF 13 14  0 */ always @(posedge clk) if (n1461) n1462 <= 1'b0 ? 1'b0 : n6888;
/* FF 15 16  1 */ always @(posedge clk) if (n1500) n1794 <= 1'b0 ? 1'b0 : n6889;
/* FF 21 15  4 */ assign n6890 = n3068;
/* FF 20 25  6 */ always @(posedge clk) if (n2612) n2803 <= 1'b0 ? 1'b0 : n6891;
/* FF 26 22  7 */ always @(posedge clk) if (n2730) n3575 <= 1'b0 ? 1'b0 : n6892;
/* FF  6  9  4 */ always @(posedge clk) if (n570) n590 <= 1'b0 ? 1'b0 : n6893;
/* FF 20 22  7 */ always @(posedge clk) if (n2384) n2783 <= 1'b0 ? 1'b0 : n6894;
/* FF 12 26  1 */ always @(posedge clk) if (n1393) n1386 <= 1'b0 ? 1'b0 : n6895;
/* FF 14  8  0 */ always @(posedge clk) if (n1741) n1593 <= 1'b0 ? 1'b0 : n6896;
/* FF 17 21  4 */ always @(posedge clk) if (n2347) n2148 <= 1'b0 ? 1'b0 : n6897;
/* FF 17 24  7 */ always @(posedge clk) if (n2000) n2165 <= 1'b0 ? 1'b0 : n6898;
/* FF 23 12  1 */ always @(posedge clk) if (n3031) n3201 <= 1'b0 ? 1'b0 : n6899;
/* FF 24 15  1 */ always @(posedge clk) if (n3233) n2122 <= 1'b0 ? 1'b0 : n6900;
/* FF  3 12  5 */ always @(posedge clk) if (n168) n282 <= 1'b0 ? 1'b0 : n6901;
/* FF 21 17  5 */ always @(posedge clk) if (n2519) n2899 <= 1'b0 ? 1'b0 : n6902;
/* FF 18  2  5 */ always @(posedge clk) if (n2207) n2204 <= 1'b0 ? 1'b0 : n6903;
/* FF 21 12  6 */ always @(posedge clk) if (n3029) n2872 <= 1'b0 ? 1'b0 : n6904;
/* FF 26 21  3 */ always @(posedge clk) if (n3421) n3565 <= 1'b0 ? 1'b0 : n6905;
/* FF 14 26  1 */ always @(posedge clk) if (n1271) n1712 <= 1'b0 ? 1'b0 : n6906;
/* FF 12 21  5 */ always @(posedge clk) if (n1205) n1344 <= 1'b0 ? 1'b0 : n6907;
/* FF 17 10  2 */ always @(posedge clk) if (n2282) n2061 <= 1'b0 ? 1'b0 : n6908;
/* FF 19 20  3 */ always @(posedge clk) if (n2553) n2568 <= 1'b0 ? 1'b0 : n6909;
/* FF  9 32  1 */ assign \rco[108]  = n1115;
/* FF  1 12  7 */ always @(posedge clk) if (n39) n53 <= 1'b0 ? 1'b0 : n6910;
/* FF 22 14  1 */ always @(posedge clk) if (n3045) n3052 <= 1'b0 ? 1'b0 : n6911;
/* FF  7  7  0 */ assign n570 = n6912;
/* FF 27  8  3 */ always @(posedge clk) if (n3464) n3348 <= 1'b0 ? 1'b0 : n6913;
/* FF 18 20  1 */ assign \rco[157]  = n6914;
/* FF  3 17  0 */ always @(posedge clk) if (n79) n310 <= 1'b0 ? 1'b0 : n6915;
/* FF 14 25  5 */ always @(posedge clk) if (n697) n1706 <= 1'b0 ? 1'b0 : n6916;
/* FF  6 21  3 */ assign n671 = n6917;
/* FF 17  4  1 */ always @(posedge clk) if (n1761) n2032 <= 1'b0 ? 1'b0 : n6918;
/* FF 23 16  7 */ assign n807 = n6919;
/* FF 11 14  4 */ always @(posedge clk) if (n1154) n1150 <= 1'b0 ? 1'b0 : n6920;
/* FF 20 10  0 */ always @(posedge clk) if (n2697) n2683 <= 1'b0 ? 1'b0 : n6921;
/* FF 14  4  5 */ assign \rco[86]  = n6922;
/* FF 11 21  5 */ always @(posedge clk) if (n819) n1201 <= 1'b0 ? 1'b0 : n6923;
/* FF 29 10  1 */ always @(posedge clk) if (n3464) n3833 <= 1'b0 ? 1'b0 : n6924;
/* FF 28 22  5 */ always @(posedge clk) if (n3704) n3804 <= 1'b0 ? 1'b0 : n6925;
/* FF 16 12  0 */ assign \rco[43]  = n6926;
/* FF  5 19  2 */ always @(posedge clk) if (n349) n541 <= 1'b0 ? 1'b0 : n6927;
/* FF  4 13  0 */ assign \rco[14]  = n501;
/* FF 16 17  7 */ always @(posedge clk) if (n2110) n1970 <= 1'b0 ? 1'b0 : n6928;
/* FF 10 23  2 */ assign n6929 = n1222;
/* FF 30 12  3 */ always @(posedge clk) if (n3892) n3897 <= 1'b0 ? 1'b0 : n6930;
/* FF 15 17  6 */ always @(posedge clk) if (n1500) n1806 <= 1'b0 ? 1'b0 : n6931;
/* FF 18  6  2 */ always @(posedge clk) if (n2241) n2233 <= 1'b0 ? 1'b0 : n6932;
/* FF  7 21  4 */ always @(posedge clk) if (n360) n772 <= 1'b0 ? 1'b0 : n6933;
/* FF  6  7  6 */ always @(posedge clk) if (n570) n577 <= 1'b0 ? 1'b0 : n6934;
/* FF 20 24  1 */ always @(posedge clk) if (n2775) n2789 <= 1'b0 ? 1'b0 : n6935;
/* FF 26  9  6 */ always @(posedge clk) if (n3460) n3461 <= 1'b0 ? 1'b0 : n6936;
/* FF  6  8  7 */ always @(posedge clk) if (n570) n586 <= 1'b0 ? 1'b0 : n6937;
/* FF 20 21  6 */ always @(posedge clk) if (n2553) n2774 <= 1'b0 ? 1'b0 : n6938;
/* FF 12 25  0 */ always @(posedge clk) if (n1532) n1376 <= 1'b0 ? 1'b0 : n6939;
/* FF 14 11  1 */ always @(posedge clk) if (n1622) n1613 <= 1'b0 ? 1'b0 : n6940;
/* FF 17 22  5 */ always @(posedge clk) if (n1999) n2157 <= 1'b0 ? 1'b0 : n6941;
/* FF  1 19  0 */ always @(posedge clk) if (n119) n104 <= 1'b0 ? 1'b0 : n6942;
/* FF 17 25  4 */ always @(posedge clk) if (n2017) n2180 <= 1'b0 ? 1'b0 : n6943;
/* FF 10 25  1 */ always @(posedge clk) if (n567) n1081 <= 1'b0 ? 1'b0 : n6944;
/* FF 24 14  2 */ always @(posedge clk) if (n3376) n3371 <= 1'b0 ? 1'b0 : n6945;
/* FF 27 20  1 */ always @(posedge clk) if (n3424) n3676 <= 1'b0 ? 1'b0 : n6946;
/* FF  4 19  4 */ assign \rco[123]  = n547;
/* FF  3 13  2 */ assign n277 = n405;
/* FF 21 18  4 */ always @(posedge clk) if (n2757) n2906 <= 1'b0 ? 1'b0 : n6947;
/* FF 22 10  6 */ always @(posedge clk) if (n2856) n3028 <= 1'b0 ? 1'b0 : n6948;
/* FF 18  5  4 */ always @(posedge clk) if (n2230) n2225 <= 1'b0 ? 1'b0 : n6949;
/* FF  7 22  6 */ always @(posedge clk) if (n695) n789 <= 1'b0 ? 1'b0 : n6950;
/* FF 21 13  5 */ always @(posedge clk) if (n2519) n2879 <= 1'b0 ? 1'b0 : n6951;
/* FF 26 20  0 */ assign \rco[169]  = n6952;
/* FF 12 15  3 */ always @(posedge clk) if (n1155) n1299 <= 1'b0 ? 1'b0 : n6953;
/* FF 14 21  0 */ assign n1196 = n1844;
/* FF 19 30  5 */ always @(posedge clk) if (n2592) n2627 <= 1'b0 ? 1'b0 : n6954;
/* FF 19 21  4 */ always @(posedge clk) if (n2164) n2580 <= 1'b0 ? 1'b0 : n6955;
/* FF 11 17  2 */ always @(posedge clk) if (n900) n1170 <= 1'b0 ? 1'b0 : n6956;
/* FF 10 11  0 */ always @(posedge clk) if (n996) n989 <= 1'b0 ? 1'b0 : n6957;
/* FF 16  8  5 */ always @(posedge clk) if (n1625) n1920 <= 1'b0 ? 1'b0 : n6958;
/* FF  1 13  4 */ always @(posedge clk) if (n83) n63 <= 1'b0 ? 1'b0 : n6959;
/* FF 28  7  5 */ always @(posedge clk) if (n3488) n2676 <= 1'b0 ? 1'b0 : n6960;
/* FF 16 29  2 */ assign \rco[117]  = n6961;
/* FF 22  9  0 */ assign n2989 = n6962;
/* FF 15 21  3 */ always @(posedge clk) if (n1356) n1839 <= 1'b0 ? 1'b0 : n6963;
/* FF 20 28  6 */ always @(posedge clk) if (n2195) n2827 <= 1'b0 ? 1'b0 : n6964;
/* FF 18 23  0 */ always @(posedge clk) if (n1999) n2362 <= 1'b0 ? 1'b0 : n6965;
/* FF 20  9  1 */ assign n1933 = n2852;
/* FF 23 17  0 */ assign n3065 = n6966;
/* FF 11 15  7 */ always @(posedge clk) if (n733) n1158 <= 1'b0 ? 1'b0 : n6967;
/* FF 26  6  4 */ always @(posedge clk) if (n3459) n3477 <= 1'b0 ? 1'b0 : n6968;
/* FF 14  7  4 */ always @(posedge clk) if (n1743) n1589 <= 1'b0 ? 1'b0 : n6969;
/* FF 11 18  4 */ always @(posedge clk) if (n1187) n1183 <= 1'b0 ? 1'b0 : n6970;
/* FF 29 11  6 */ always @(posedge clk) if (n3751) n3845 <= 1'b0 ? 1'b0 : n6971;
/* FF 28 21  4 */ always @(posedge clk) if (n3788) n3795 <= 1'b0 ? 1'b0 : n6972;
/* FF  5 20  3 */ always @(posedge clk) if (n552) n548 <= 1'b0 ? 1'b0 : n6973;
/* FF 19  3  0 */ always @(posedge clk) if (n1887) n2427 <= 1'b0 ? 1'b0 : n6974;
/* FF  3  9  7 */ always @(posedge clk) if (n260) n259 <= 1'b0 ? 1'b0 : n6975;
/* FF 15 22  7 */ always @(posedge clk) if (n1835) n1852 <= 1'b0 ? 1'b0 : n6976;
/* FF 18  9  3 */ always @(posedge clk) if (n2055) n2264 <= 1'b0 ? 1'b0 : n6977;
/* FF  9 19  5 */ always @(posedge clk) if (n454) n906 <= 1'b0 ? 1'b0 : n6978;
/* FF 12 19  6 */ always @(posedge clk) if (n1501) n1333 <= 1'b0 ? 1'b0 : n6979;
/* FF 26  8  5 */ always @(posedge clk) if (n3603) n3495 <= 1'b0 ? 1'b0 : n6980;
/* FF  6 11  6 */ always @(posedge clk) if (n286) n604 <= 1'b0 ? 1'b0 : n6981;
/* FF 12 24  7 */ always @(posedge clk) if (n961) n945 <= 1'b0 ? 1'b0 : n6982;
/* FF 17 23  2 */ always @(posedge clk) if (n1069) n1695 <= 1'b0 ? 1'b0 : n6983;
/* FF  2 12  1 */ always @(posedge clk) if (n39) n177 <= 1'b0 ? 1'b0 : n6984;
/* FF 19 17  1 */ always @(posedge clk) if (n2727) n2542 <= 1'b0 ? 1'b0 : n6985;
/* FF 22 21  2 */ always @(posedge clk) if (n2564) n3098 <= 1'b0 ? 1'b0 : n6986;
/* FF 24 24  4 */ always @(posedge clk) if (n3112) n3443 <= 1'b0 ? 1'b0 : n6987;
/* FF 10 24  2 */ always @(posedge clk) if (n820) n1074 <= 1'b0 ? 1'b0 : n6988;
/* FF 24 13  3 */ always @(posedge clk) if (n3351) n3364 <= 1'b0 ? 1'b0 : n6989;
/* FF 27 21  6 */ always @(posedge clk) if (n3421) n3693 <= 1'b0 ? 1'b0 : n6990;
/* FF  4 18  7 */ always @(posedge clk) if (n349) n437 <= 1'b0 ? 1'b0 : n6991;
/* FF  3 10  3 */ always @(posedge clk) if (n251) n265 <= 1'b0 ? 1'b0 : n6992;
/* FF  7  8  4 */ always @(posedge clk) if (n588) n717 <= 1'b0 ? 1'b0 : n6993;
/* FF 21 19  3 */ always @(posedge clk) if (n2757) n2913 <= 1'b0 ? 1'b0 : n6994;
/* FF  9 16  1 */ always @(posedge clk) if (n645) n876 <= 1'b0 ? 1'b0 : n6995;
/* FF 12 14  0 */ always @(posedge clk) if (n1154) n1288 <= 1'b0 ? 1'b0 : n6996;
/* FF 26 23  1 */ always @(posedge clk) if (n3703) n3577 <= 1'b0 ? 1'b0 : n6997;
/* FF 14 20  3 */ always @(posedge clk) if (n1347) n1679 <= 1'b0 ? 1'b0 : n6998;
/* FF 19 31  6 */ always @(posedge clk) if (n2592) n2647 <= 1'b0 ? 1'b0 : n6999;
/* FF 23 21  5 */ always @(posedge clk) if (n3258) n3276 <= 1'b0 ? 1'b0 : n7000;
/* FF 19 18  5 */ always @(posedge clk) if (n2348) n2559 <= 1'b0 ? 1'b0 : n7001;
/* FF 16 23  4 */ always @(posedge clk) if (n2000) n1995 <= 1'b0 ? 1'b0 : n7002;
/* FF  1 14  5 */ always @(posedge clk) if (n85) n73 <= 1'b0 ? 1'b0 : n7003;
/* FF 28  6  6 */ always @(posedge clk) if (n3594) n3716 <= 1'b0 ? 1'b0 : n7004;
/* FF 15 10  2 */ always @(posedge clk) if (n1624) n1756 <= 1'b0 ? 1'b0 : n7005;
/* FF 20 19  7 */ always @(posedge clk) if (n2562) n2756 <= 1'b0 ? 1'b0 : n7006;
/* FF 17  6  3 */ always @(posedge clk) if (n2045) n2041 <= 1'b0 ? 1'b0 : n7007;
/* FF  6 23  1 */ always @(posedge clk) if (n360) n688 <= 1'b0 ? 1'b0 : n7008;
/* FF 20  8  6 */ always @(posedge clk) if (n2247) n2674 <= 1'b0 ? 1'b0 : n7009;
/* FF 12 28  4 */ always @(posedge clk) if (n1394) n1398 <= 1'b0 ? 1'b0 : n7010;
/* FF 23 22  1 */ always @(posedge clk) if (n3422) n3280 <= 1'b0 ? 1'b0 : n7011;
/* FF 14  6  3 */ assign n1577 = n7012;
/* FF 17 19  7 */ always @(posedge clk) if (n1982) n2135 <= 1'b0 ? 1'b0 : n7013;
/* FF 11 19  7 */ assign n912 = n7014;
/* FF 29 12  7 */ always @(posedge clk) if (n3751) n3855 <= 1'b0 ? 1'b0 : n7015;
/* FF 16 10  2 */ always @(posedge clk) if (n1771) n1928 <= 1'b0 ? 1'b0 : n7016;
/* FF  5 21  0 */ assign n7017 = n675;
/* FF 22 26  0 */ always @(posedge clk) if (n2613) n3133 <= 1'b0 ? 1'b0 : n7018;
/* FF  9 12  3 */ always @(posedge clk) if (n996) n852 <= 1'b0 ? 1'b0 : n7019;
/* FF 27 17  3 */ always @(posedge clk) if (n3249) n3651 <= 1'b0 ? 1'b0 : n7020;
/* FF 15 24  5 */ always @(posedge clk) if (n778) n1868 <= 1'b0 ? 1'b0 : n7021;
/* FF 15 23  4 */ always @(posedge clk) if (n778) n1856 <= 1'b0 ? 1'b0 : n7022;
/* FF 18  8  0 */ always @(posedge clk) if (n2055) n2249 <= 1'b0 ? 1'b0 : n7023;
/* FF 12 18  5 */ always @(posedge clk) if (n1501) n1325 <= 1'b0 ? 1'b0 : n7024;
/* FF 26 11  4 */ always @(posedge clk) if (n3033) n3512 <= 1'b0 ? 1'b0 : n7025;
/* FF 17 16  3 */ assign \rco[28]  = n2323;
/* FF  2 15  0 */ always @(posedge clk) if (n197) n196 <= 1'b0 ? 1'b0 : n7026;
/* FF 19 14  0 */ assign n2511 = n7027;
/* FF 22 20  1 */ always @(posedge clk) if (n3087) n3089 <= 1'b0 ? 1'b0 : n7028;
/* FF 10 14  4 */ always @(posedge clk) if (n750) n1011 <= 1'b0 ? 1'b0 : n7029;
/* FF 24 23  5 */ always @(posedge clk) if (n3104) n3438 <= 1'b0 ? 1'b0 : n7030;
/* FF 10 27  3 */ always @(posedge clk) if (n804) n1096 <= 1'b0 ? 1'b0 : n7031;
/* FF 24 12  4 */ always @(posedge clk) if (n3351) n3357 <= 1'b0 ? 1'b0 : n7032;
/* FF 16 24  2 */ assign n338 = n2174;
/* FF 27 18  7 */ always @(posedge clk) if (n3553) n2521 <= 1'b0 ? 1'b0 : n7033;
/* FF 28 10  3 */ always @(posedge clk) if (n3462) n3744 <= 1'b0 ? 1'b0 : n7034;
/* FF  3 11  0 */ always @(posedge clk) if (n153) n270 <= 1'b0 ? 1'b0 : n7035;
/* FF  7  9  3 */ always @(posedge clk) if (n589) n721 <= 1'b0 ? 1'b0 : n7036;
/* FF 21 20  2 */ always @(posedge clk) if (n3087) n2920 <= 1'b0 ? 1'b0 : n7037;
/* FF 18  7  6 */ always @(posedge clk) if (n1761) n2245 <= 1'b0 ? 1'b0 : n7038;
/* FF  9 17  2 */ always @(posedge clk) if (n1030) n885 <= 1'b0 ? 1'b0 : n7039;
/* FF 15  5  0 */ always @(posedge clk) if (n1742) n1725 <= 1'b0 ? 1'b0 : n7040;
/* FF 14 23  2 */ assign n335 = n1861;
/* FF 20 12  3 */ always @(posedge clk) if (n2682) n2701 <= 1'b0 ? 1'b0 : n7041;
/* FF 19 19  6 */ assign \rco[162]  = n2760;
/* FF  1 15  2 */ assign \rco[4]  = n203;
/* FF 16 27  4 */ always @(posedge clk) if (n1) n2018 <= 1'b0 ? 1'b0 : n7042;
/* FF 22 11  2 */ assign n2085 = n3198;
/* FF 30 10  2 */ always @(posedge clk) if (n3892) n3887 <= 1'b0 ? 1'b0 : n7043;
/* FF 15 11  1 */ always @(posedge clk) if (n1624) n1764 <= 1'b0 ? 1'b0 : n7044;
/* FF  6 13  7 */ always @(posedge clk) if (n78) n622 <= 1'b0 ? 1'b0 : n7045;
/* FF 20 18  4 */ always @(posedge clk) if (n2348) n2745 <= 1'b0 ? 1'b0 : n7046;
/* FF 17  7  4 */ always @(posedge clk) if (n2045) n2050 <= 1'b0 ? 1'b0 : n7047;
/* FF  6 22  6 */ always @(posedge clk) if (n673) n684 <= 1'b0 ? 1'b0 : n7048;
/* FF 20 15  7 */ always @(posedge clk) if (n2715) n2724 <= 1'b0 ? 1'b0 : n7049;
/* FF 23 23  2 */ always @(posedge clk) if (n3104) n3289 <= 1'b0 ? 1'b0 : n7050;
/* FF 11 13  1 */ always @(posedge clk) if (n733) n1139 <= 1'b0 ? 1'b0 : n7051;
/* FF 11 16  6 */ always @(posedge clk) if (n891) n1165 <= 1'b0 ? 1'b0 : n7052;
/* FF  5 22  1 */ always @(posedge clk) if (n673) n556 <= 1'b0 ? 1'b0 : n7053;
/* FF  9 13  0 */ always @(posedge clk) if (n629) n855 <= 1'b0 ? 1'b0 : n7054;
/* FF 13  7  3 */ always @(posedge clk) if (n977) n1426 <= 1'b0 ? 1'b0 : n7055;
/* FF 15 25  2 */ assign \rco[184]  = n7056;
/* FF 18 11  1 */ assign n1624 = n7057;
/* FF 15 20  5 */ always @(posedge clk) if (n1347) n1832 <= 1'b0 ? 1'b0 : n7058;
/* FF 12 17  4 */ always @(posedge clk) if (n900) n1316 <= 1'b0 ? 1'b0 : n7059;
/* FF 26 10  3 */ always @(posedge clk) if (n3033) n3508 <= 1'b0 ? 1'b0 : n7060;
/* FF 26  7  4 */ always @(posedge clk) if (n3603) n3485 <= 1'b0 ? 1'b0 : n7061;
/* FF 17 17  0 */ always @(posedge clk) if (n2111) n2114 <= 1'b0 ? 1'b0 : n7062;
/* FF  5 24  0 */ always @(posedge clk) if (n360) n566 <= 1'b0 ? 1'b0 : n7063;
/* FF 19 15  3 */ always @(posedge clk) if (n2715) n2528 <= 1'b0 ? 1'b0 : n7064;
/* FF 22 23  0 */ assign n2229 = n3295;
/* FF 23  5  2 */ always @(posedge clk) if (n3158) n3152 <= 1'b0 ? 1'b0 : n7065;
/* FF 24 22  6 */ always @(posedge clk) if (n3422) n3430 <= 1'b0 ? 1'b0 : n7066;
/* FF 10 26  4 */ assign n821 = n7067;
/* FF 24 11  5 */ assign n7068 = n3467;
/* FF 27 19  4 */ always @(posedge clk) if (n3553) n3671 <= 1'b0 ? 1'b0 : n7069;
/* FF 28  9  2 */ always @(posedge clk) if (n3621) n3736 <= 1'b0 ? 1'b0 : n7070;
/* FF  4 16  1 */ always @(posedge clk) if (n79) n421 <= 1'b0 ? 1'b0 : n7071;
/* FF 21 21  1 */ always @(posedge clk) if (n2564) n2927 <= 1'b0 ? 1'b0 : n7072;
/* FF  9 18  3 */ always @(posedge clk) if (n1030) n895 <= 1'b0 ? 1'b0 : n7073;
/* FF 14 22  5 */ always @(posedge clk) if (n1402) n1692 <= 1'b0 ? 1'b0 : n7074;
/* FF 17  3  1 */ always @(posedge clk) if (n1887) n2026 <= 1'b0 ? 1'b0 : n7075;
/* FF  6 18  3 */ always @(posedge clk) if (n657) n652 <= 1'b0 ? 1'b0 : n7076;
/* FF 19 29  0 */ assign n1881 = n7077;
/* FF 19 16  7 */ assign n1951 = n7078;
/* FF 23  6  4 */ always @(posedge clk) if (n3158) n3163 <= 1'b0 ? 1'b0 : n7079;
/* FF 11 28  1 */ always @(posedge clk) if (n1384) n1256 <= 1'b0 ? 1'b0 : n7080;
/* FF 10 12  5 */ always @(posedge clk) if (n996) n1002 <= 1'b0 ? 1'b0 : n7081;
/* FF 24 25  4 */ always @(posedge clk) if (n2812) n3450 <= 1'b0 ? 1'b0 : n7082;
/* FF  1  8  3 */ always @(posedge clk) if (n37) n17 <= 1'b0 ? 1'b0 : n7083;
/* FF 27  1  0 */ assign \rco[79]  = n7084;
/* FF 15  8  0 */ always @(posedge clk) if (n1741) n1746 <= 1'b0 ? 1'b0 : n7085;
/* FF  3 22  5 */ always @(posedge clk) if (n352) n247 <= 1'b0 ? 1'b0 : n7086;
/* FF  2 18  1 */ always @(posedge clk) if (n115) n210 <= 1'b0 ? 1'b0 : n7087;
/* FF  6 12  4 */ always @(posedge clk) if (n286) n610 <= 1'b0 ? 1'b0 : n7088;
/* FF 20 17  5 */ always @(posedge clk) if (n2727) n2737 <= 1'b0 ? 1'b0 : n7089;
/* FF 23 20  3 */ always @(posedge clk) if (n3258) n3266 <= 1'b0 ? 1'b0 : n7090;
/* FF 24  7  0 */ assign \rco[82]  = n7091;
/* FF  9 14  1 */ always @(posedge clk) if (n629) n860 <= 1'b0 ? 1'b0 : n7092;
/* FF  4 20  6 */ always @(posedge clk) if (n215) n444 <= 1'b0 ? 1'b0 : n7093;
/* FF 18 10  6 */ always @(posedge clk) if (n2282) n2279 <= 1'b0 ? 1'b0 : n7094;
/* FF 26 13  2 */ assign n3527 = n7095;
/* FF 12 16  3 */ always @(posedge clk) if (n1155) n1307 <= 1'b0 ? 1'b0 : n7096;
/* FF 14 18  2 */ always @(posedge clk) if (n1672) n1663 <= 1'b0 ? 1'b0 : n7097;
/* FF 19 25  5 */ always @(posedge clk) if (n2612) n2609 <= 1'b0 ? 1'b0 : n7098;
/* FF 17 18  1 */ always @(posedge clk) if (n1825) n2126 <= 1'b0 ? 1'b0 : n7099;
/* FF 19 12  2 */ always @(posedge clk) if (n1936) n2499 <= 1'b0 ? 1'b0 : n7100;
/* FF 23 10  3 */ always @(posedge clk) if (n2697) n3186 <= 1'b0 ? 1'b0 : n7101;
/* FF 22 22  7 */ always @(posedge clk) if (n2961) n3111 <= 1'b0 ? 1'b0 : n7102;
/* FF 24 10  6 */ always @(posedge clk) if (n3352) n3346 <= 1'b0 ? 1'b0 : n7103;
/* FF 28  8  5 */ always @(posedge clk) if (n3605) n2681 <= 1'b0 ? 1'b0 : n7104;
/* FF  7 15  1 */ assign n739 = n7105;
/* FF 21 22  0 */ always @(posedge clk) if (n2384) n2935 <= 1'b0 ? 1'b0 : n7106;
/* FF 14 28  7 */ always @(posedge clk) if (n1402) n1722 <= 1'b0 ? 1'b0 : n7107;
/* FF  2 22  6 */ always @(posedge clk) if (n352) n241 <= 1'b0 ? 1'b0 : n7108;
/* FF 14 17  4 */ always @(posedge clk) if (n1672) n1658 <= 1'b0 ? 1'b0 : n7109;
/* FF 17 12  0 */ always @(posedge clk) if (n2056) n2077 <= 1'b0 ? 1'b0 : n7110;
/* FF 19 26  1 */ assign n2020 = n7111;
/* FF  5 11  0 */ always @(posedge clk) if (n184) n481 <= 1'b0 ? 1'b0 : n7112;
/* FF 23 24  6 */ always @(posedge clk) if (n3112) n3302 <= 1'b0 ? 1'b0 : n7113;
/* FF 23  7  7 */ always @(posedge clk) if (n3006) n3173 <= 1'b0 ? 1'b0 : n7114;
/* FF 11 29  6 */ always @(posedge clk) if (n1384) n1268 <= 1'b0 ? 1'b0 : n7115;
/* FF 10 15  4 */ always @(posedge clk) if (n750) n1019 <= 1'b0 ? 1'b0 : n7116;
/* FF 16 20  1 */ always @(posedge clk) if (n1843) n1975 <= 1'b0 ? 1'b0 : n7117;
/* FF 21 24  3 */ always @(posedge clk) if (n3113) n2956 <= 1'b0 ? 1'b0 : n7118;
/* FF 15 18  6 */ always @(posedge clk) if (n1355) n1814 <= 1'b0 ? 1'b0 : n7119;
/* FF 13 23  0 */ always @(posedge clk) if (n1069) n1524 <= 1'b0 ? 1'b0 : n7120;
/* FF 27 14  1 */ always @(posedge clk) if (n3527) n3642 <= 1'b0 ? 1'b0 : n7121;
/* FF 18 14  3 */ assign n7122 = n2524;
/* FF 32  7  2 */ assign \rco[49]  = n7123;
/* FF  2 21  0 */ always @(posedge clk) if (n126) n227 <= 1'b0 ? 1'b0 : n7124;
/* FF 20 16  2 */ assign n2727 = n7125;
/* FF  6 15  5 */ always @(posedge clk) if (n630) n635 <= 1'b0 ? 1'b0 : n7126;
/* FF  6 16  4 */ always @(posedge clk) if (n511) n642 <= 1'b0 ? 1'b0 : n7127;
/* FF 20 13  5 */ always @(posedge clk) if (n2283) n2709 <= 1'b0 ? 1'b0 : n7128;
/* FF  4 11  2 */ always @(posedge clk) if (n184) n387 <= 1'b0 ? 1'b0 : n7129;
/* FF 22 18  4 */ always @(posedge clk) if (n3065) n3084 <= 1'b0 ? 1'b0 : n7130;
/* FF 22  7  3 */ always @(posedge clk) if (n2841) n3001 <= 1'b0 ? 1'b0 : n7131;
/* FF 10 17  0 */ assign \rco[148]  = n7132;
/* FF  9 15  6 */ always @(posedge clk) if (n645) n873 <= 1'b0 ? 1'b0 : n7133;
/* FF 13  9  1 */ always @(posedge clk) if (n850) n1431 <= 1'b0 ? 1'b0 : n7134;
/* FF 24  6  3 */ always @(posedge clk) if (n3006) n3324 <= 1'b0 ? 1'b0 : n7135;
/* FF 28 12  2 */ always @(posedge clk) if (n3462) n3755 <= 1'b0 ? 1'b0 : n7136;
/* FF 30 11  6 */ assign n3892 = n7137;
/* FF 18 13  7 */ always @(posedge clk) if (n2283) n2302 <= 1'b0 ? 1'b0 : n7138;
/* FF 12 23  2 */ always @(posedge clk) if (n1357) n1360 <= 1'b0 ? 1'b0 : n7139;
/* FF 26 12  1 */ always @(posedge clk) if (n3368) n3518 <= 1'b0 ? 1'b0 : n7140;
/* FF 14 13  3 */ always @(posedge clk) if (n1015) n1627 <= 1'b0 ? 1'b0 : n7141;
/* FF  5 15  5 */ always @(posedge clk) if (n511) n519 <= 1'b0 ? 1'b0 : n7142;
/* FF 19 22  4 */ always @(posedge clk) if (n2164) n2588 <= 1'b0 ? 1'b0 : n7143;
/* FF 19 13  5 */ always @(posedge clk) if (n2283) n2509 <= 1'b0 ? 1'b0 : n7144;
/* FF 23 11  0 */ always @(posedge clk) if (n3031) n3190 <= 1'b0 ? 1'b0 : n7145;
/* FF 11 25  3 */ always @(posedge clk) if (n954) n1234 <= 1'b0 ? 1'b0 : n7146;
/* FF 22 17  6 */ always @(posedge clk) if (n3065) n3078 <= 1'b0 ? 1'b0 : n7147;
/* FF 24 20  0 */ always @(posedge clk) if (n3411) n3414 <= 1'b0 ? 1'b0 : n7148;
/* FF 16 16  6 */ always @(posedge clk) if (n2110) n1961 <= 1'b0 ? 1'b0 : n7149;
/* FF 10 28  6 */ always @(posedge clk) if (n821) n1107 <= 1'b0 ? 1'b0 : n7150;
/* FF 24  9  7 */ always @(posedge clk) if (n3352) n3339 <= 1'b0 ? 1'b0 : n7151;
/* FF 13  6  5 */ always @(posedge clk) if (n977) n1420 <= 1'b0 ? 1'b0 : n7152;
/* FF  4 22  3 */ assign \rco[136]  = n7153;
/* FF 15 13  4 */ always @(posedge clk) if (n1015) n1781 <= 1'b0 ? 1'b0 : n7154;
/* FF 20 20  7 */ always @(posedge clk) if (n2562) n2767 <= 1'b0 ? 1'b0 : n7155;
/* FF 29 19  4 */ always @(posedge clk) if (n3786) n3865 <= 1'b0 ? 1'b0 : n7156;
/* FF 14 16  7 */ always @(posedge clk) if (n1792) n1653 <= 1'b0 ? 1'b0 : n7157;
/* FF 17 13  3 */ always @(posedge clk) if (n2056) n2089 <= 1'b0 ? 1'b0 : n7158;
/* FF  5 12  1 */ always @(posedge clk) if (n77) n485 <= 1'b0 ? 1'b0 : n7159;
/* FF 19 27  2 */ always @(posedge clk) if (n2614) n2618 <= 1'b0 ? 1'b0 : n7160;
/* FF 11 23  4 */ always @(posedge clk) if (n796) n1218 <= 1'b0 ? 1'b0 : n7161;
/* FF 23 25  1 */ always @(posedge clk) if (n2613) n2797 <= 1'b0 ? 1'b0 : n7162;
/* FF 11 26  7 */ always @(posedge clk) if (n954) n1242 <= 1'b0 ? 1'b0 : n7163;
/* FF 16 19  0 */ assign \rco[138]  = n7164;
/* FF  1 10  1 */ always @(posedge clk) if (n37) n29 <= 1'b0 ? 1'b0 : n7165;
/* FF 21 25  0 */ always @(posedge clk) if (n2970) n2962 <= 1'b0 ? 1'b0 : n7166;
/* FF  9 11  3 */ always @(posedge clk) if (n988) n845 <= 1'b0 ? 1'b0 : n7167;
/* FF 15 19  5 */ always @(posedge clk) if (n1355) n1822 <= 1'b0 ? 1'b0 : n7168;
/* FF 13 24  1 */ assign n7169 = n1700;
/* FF 15 14  6 */ always @(posedge clk) if (n1791) n1789 <= 1'b0 ? 1'b0 : n7170;
/* FF  3 20  7 */ always @(posedge clk) if (n119) n348 <= 1'b0 ? 1'b0 : n7171;
/* FF  2 20  3 */ always @(posedge clk) if (n126) n220 <= 1'b0 ? 1'b0 : n7172;
/* FF  6 14  2 */ always @(posedge clk) if (n78) n625 <= 1'b0 ? 1'b0 : n7173;
/* FF 18 17  2 */ always @(posedge clk) if (n1825) n2327 <= 1'b0 ? 1'b0 : n7174;
/* FF 20 23  3 */ assign n2785 = n2952;
/* FF  6 19  5 */ assign n659 = n7175;
/* FF 11  8  2 */ always @(posedge clk) if (n1131) n1125 <= 1'b0 ? 1'b0 : n7176;
/* FF 29  5  0 */ always @(posedge clk) if (n3605) n3818 <= 1'b0 ? 1'b0 : n7177;
/* FF 19  9  2 */ always @(posedge clk) if (n2451) n2473 <= 1'b0 ? 1'b0 : n7178;
/* FF  4 10  1 */ always @(posedge clk) if (n251) n380 <= 1'b0 ? 1'b0 : n7179;
/* FF 24 16  5 */ always @(posedge clk) if (n3376) n3389 <= 1'b0 ? 1'b0 : n7180;
/* FF 27 22  6 */ always @(posedge clk) if (n3703) n3701 <= 1'b0 ? 1'b0 : n7181;
/* FF 22  6  4 */ always @(posedge clk) if (n2841) n2994 <= 1'b0 ? 1'b0 : n7182;
/* FF 10 16  3 */ always @(posedge clk) if (n891) n1026 <= 1'b0 ? 1'b0 : n7183;
/* FF 13 10  0 */ always @(posedge clk) if (n850) n1434 <= 1'b0 ? 1'b0 : n7184;
/* FF 18  3  5 */ assign n2207 = n7185;
/* FF 31 22  5 */ assign \rco[185]  = n7186;
/* FF 18 12  4 */ always @(posedge clk) if (n1936) n2290 <= 1'b0 ? 1'b0 : n7187;
/* FF 21  6  3 */ always @(posedge clk) if (n2247) n2836 <= 1'b0 ? 1'b0 : n7188;
/* FF 26 15  0 */ assign n3233 = n7189;
/* FF 11  6  1 */ always @(posedge clk) if (en_in) n1119 <= 1'b0 ? 1'b0 : n7190;
/* FF 12 22  1 */ always @(posedge clk) if (n1357) n1349 <= 1'b0 ? 1'b0 : n7191;
/* FF 14 12  0 */ assign n7192 = n1773;
/* FF 19 23  7 */ assign n2017 = n7193;
/* FF 19 10  4 */ always @(posedge clk) if (n2678) n2483 <= 1'b0 ? 1'b0 : n7194;
/* FF  4 21  2 */ always @(posedge clk) if (n552) n449 <= 1'b0 ? 1'b0 : n7195;
/* FF 26 17  3 */ always @(posedge clk) if (n3249) n3549 <= 1'b0 ? 1'b0 : n7196;
/* FF  6 10  7 */ always @(posedge clk) if (n589) n598 <= 1'b0 ? 1'b0 : n7197;
/* FF 18 30  0 */ always @(posedge clk) if (n1881) n2417 <= 1'b0 ? 1'b0 : n7198;
/* FF 14 19  6 */ always @(posedge clk) if (n1672) n1670 <= 1'b0 ? 1'b0 : n7199;
/* FF 17 14  2 */ always @(posedge clk) if (n1625) n2096 <= 1'b0 ? 1'b0 : n7200;
/* FF 20 11  6 */ always @(posedge clk) if (n2682) n2694 <= 1'b0 ? 1'b0 : n7201;
/* FF  5 13  2 */ always @(posedge clk) if (n402) n494 <= 1'b0 ? 1'b0 : n7202;
/* FF 19 24  3 */ always @(posedge clk) if (n2775) n2597 <= 1'b0 ? 1'b0 : n7203;
/* FF 11 20  5 */ always @(posedge clk) if (n1339) n137 <= 1'b0 ? 1'b0 : n7204;
/* FF 29  9  5 */ always @(posedge clk) if (n3464) n3830 <= 1'b0 ? 1'b0 : n7205;
/* FF 29 20  5 */ always @(posedge clk) if (n3786) n3873 <= 1'b0 ? 1'b0 : n7206;
/* FF 11 27  4 */ always @(posedge clk) if (n1393) n1251 <= 1'b0 ? 1'b0 : n7207;
/* FF 21 26  1 */ assign \rco[174]  = n7208;
/* FF 15 16  4 */ always @(posedge clk) if (n1500) n1797 <= 1'b0 ? 1'b0 : n7209;
/* FF 13 25  2 */ always @(posedge clk) if (n697) n1536 <= 1'b0 ? 1'b0 : n7210;
/* FF 27 12  3 */ always @(posedge clk) if (n3368) n3632 <= 1'b0 ? 1'b0 : n7211;
/* FF 15 15  5 */ assign n7212 = n1953;
/* FF  3 21  0 */ assign n7213 = n458;
/* FF 18 16  1 */ always @(posedge clk) if (n2540) n2315 <= 1'b0 ? 1'b0 : n7214;
/* FF  6  9  3 */ assign n589 = n7215;
/* FF 20 22  0 */ always @(posedge clk) if (n2384) n2776 <= 1'b0 ? 1'b0 : n7216;
/* FF 17 24  2 */ always @(posedge clk) if (n2000) n2168 <= 1'b0 ? 1'b0 : n7217;
/* FF 19  6  3 */ always @(posedge clk) if (n2241) n2446 <= 1'b0 ? 1'b0 : n7218;
/* FF  4  9  0 */ always @(posedge clk) if (n260) n371 <= 1'b0 ? 1'b0 : n7219;
/* FF 10  6  5 */ always @(posedge clk) if (en_in) n975 <= 1'b0 ? 1'b0 : n7220;
/* FF 24 15  4 */ always @(posedge clk) if (n3233) n3379 <= 1'b0 ? 1'b0 : n7221;
/* FF 27 23  5 */ assign n3704 = n7222;
/* FF 10 19  2 */ assign n117 = n7223;
/* FF  9  9  4 */ always @(posedge clk) if (n983) n831 <= 1'b0 ? 1'b0 : n7224;
/* FF 13 11  7 */ always @(posedge clk) if (n1137) n1448 <= 1'b0 ? 1'b0 : n7225;
/* FF 18  2  2 */ always @(posedge clk) if (n2207) n2201 <= 1'b0 ? 1'b0 : n7226;
/* FF 18 15  5 */ always @(posedge clk) if (n1) n2312 <= 1'b0 ? 1'b0 : n7227;
/* FF 14 26  6 */ always @(posedge clk) if (n1271) n1717 <= 1'b0 ? 1'b0 : n7228;
/* FF 12 21  0 */ assign \rco[120]  = n7229;
/* FF 14 15  1 */ always @(posedge clk) if (n1792) n1640 <= 1'b0 ? 1'b0 : n7230;
/* FF  2  9  2 */ always @(posedge clk) if (n153) n159 <= 1'b0 ? 1'b0 : n7231;
/* FF 20  4  4 */ always @(posedge clk) if (n1761) n2654 <= 1'b0 ? 1'b0 : n7232;
/* FF 19 20  6 */ always @(posedge clk) if (n2553) n2571 <= 1'b0 ? 1'b0 : n7233;
/* FF 19 11  7 */ always @(posedge clk) if (n2076) n2075 <= 1'b0 ? 1'b0 : n7234;
/* FF 23  9  6 */ always @(posedge clk) if (n2678) n3182 <= 1'b0 ? 1'b0 : n7235;
/* FF 22 19  4 */ always @(posedge clk) if (n2757) n2758 <= 1'b0 ? 1'b0 : n7236;
/* FF 10  5  1 */ always @(posedge clk) if (en_in) n967 <= 1'b0 ? 1'b0 : n7237;
/* FF 24 18  2 */ always @(posedge clk) if (n3411) n3404 <= 1'b0 ? 1'b0 : n7238;
/* FF  9 27  0 */ always @(posedge clk) if (n804) n946 <= 1'b0 ? 1'b0 : n7239;
/* FF 26 16  0 */ always @(posedge clk) if (n3249) n2333 <= 1'b0 ? 1'b0 : n7240;
/* FF  3 17  5 */ always @(posedge clk) if (n79) n103 <= 1'b0 ? 1'b0 : n7241;
/* FF 14 25  0 */ always @(posedge clk) if (n697) n1701 <= 1'b0 ? 1'b0 : n7242;
/* FF  6 21  6 */ assign n7243 = n782;
/* FF 17  4  4 */ always @(posedge clk) if (n1761) n2034 <= 1'b0 ? 1'b0 : n7244;
/* FF 17 15  5 */ always @(posedge clk) if (n2111) n2106 <= 1'b0 ? 1'b0 : n7245;
/* FF 20 10  5 */ always @(posedge clk) if (n2697) n2494 <= 1'b0 ? 1'b0 : n7246;
/* FF 20  7  6 */ always @(posedge clk) if (n2670) n2667 <= 1'b0 ? 1'b0 : n7247;
/* FF  5 14  3 */ always @(posedge clk) if (n402) n507 <= 1'b0 ? 1'b0 : n7248;
/* FF 29 21  6 */ always @(posedge clk) if (n3788) n3880 <= 1'b0 ? 1'b0 : n7249;
/* FF 11 21  2 */ always @(posedge clk) if (n819) n1198 <= 1'b0 ? 1'b0 : n7250;
/* FF 29 10  4 */ always @(posedge clk) if (n3464) n3836 <= 1'b0 ? 1'b0 : n7251;
/* FF 11 24  5 */ always @(posedge clk) if (n796) n1228 <= 1'b0 ? 1'b0 : n7252;
/* FF 16 17  2 */ always @(posedge clk) if (n2110) n1965 <= 1'b0 ? 1'b0 : n7253;
/* FF 22 13  0 */ assign \rco[53]  = n7254;
/* FF 21 27  6 */ always @(posedge clk) if (n2196) n2977 <= 1'b0 ? 1'b0 : n7255;
/* FF  9  5  1 */ assign \rco[151]  = n7256;
/* FF 13 15  4 */ always @(posedge clk) if (n739) n1474 <= 1'b0 ? 1'b0 : n7257;
/* FF 27  6  5 */ assign \rco[78]  = n7258;
/* FF 30 12  4 */ always @(posedge clk) if (n3892) n3898 <= 1'b0 ? 1'b0 : n7259;
/* FF 15 17  3 */ always @(posedge clk) if (n1500) n1804 <= 1'b0 ? 1'b0 : n7260;
/* FF 13 26  3 */ always @(posedge clk) if (n1271) n1547 <= 1'b0 ? 1'b0 : n7261;
/* FF 18  6  7 */ always @(posedge clk) if (n2241) n2238 <= 1'b0 ? 1'b0 : n7262;
/* FF 27 13  4 */ always @(posedge clk) if (n3460) n3628 <= 1'b0 ? 1'b0 : n7263;
/* FF 18 19  0 */ always @(posedge clk) if (n1982) n2339 <= 1'b0 ? 1'b0 : n7264;
/* FF  3 18  1 */ always @(posedge clk) if (n215) n319 <= 1'b0 ? 1'b0 : n7265;
/* FF  6  8  0 */ always @(posedge clk) if (n570) n580 <= 1'b0 ? 1'b0 : n7266;
/* FF 20 21  1 */ always @(posedge clk) if (n2553) n2769 <= 1'b0 ? 1'b0 : n7267;
/* FF  1 19  5 */ always @(posedge clk) if (n119) n109 <= 1'b0 ? 1'b0 : n7268;
/* FF 17 25  1 */ always @(posedge clk) if (n2017) n2177 <= 1'b0 ? 1'b0 : n7269;
/* FF 16 15  1 */ always @(posedge clk) if (n739) n1944 <= 1'b0 ? 1'b0 : n7270;
/* FF 19  7  0 */ always @(posedge clk) if (n2670) n2452 <= 1'b0 ? 1'b0 : n7271;
/* FF 23 13  3 */ always @(posedge clk) if (n3045) n3211 <= 1'b0 ? 1'b0 : n7272;
/* FF 10 25  4 */ always @(posedge clk) if (n567) n1084 <= 1'b0 ? 1'b0 : n7273;
/* FF 24 14  7 */ always @(posedge clk) if (n3376) n3375 <= 1'b0 ? 1'b0 : n7274;
/* FF 27 20  4 */ always @(posedge clk) if (n3424) n3679 <= 1'b0 ? 1'b0 : n7275;
/* FF 10 18  5 */ always @(posedge clk) if (n1187) n1038 <= 1'b0 ? 1'b0 : n7276;
/* FF  9 10  5 */ always @(posedge clk) if (n988) n839 <= 1'b0 ? 1'b0 : n7277;
/* FF 13 12  6 */ always @(posedge clk) if (n1137) n1455 <= 1'b0 ? 1'b0 : n7278;
/* FF 18  5  3 */ always @(posedge clk) if (n2230) n2224 <= 1'b0 ? 1'b0 : n7279;
/* FF 20 27  0 */ always @(posedge clk) if (n2195) n2814 <= 1'b0 ? 1'b0 : n7280;
/* FF 14 21  7 */ assign n1683 = n7281;
/* FF 14 14  6 */ always @(posedge clk) if (n1791) n1637 <= 1'b0 ? 1'b0 : n7282;
/* FF  2  8  1 */ always @(posedge clk) if (n21) n156 <= 1'b0 ? 1'b0 : n7283;
/* FF  1 16  1 */ always @(posedge clk) if (n85) n89 <= 1'b0 ? 1'b0 : n7284;
/* FF  6 26  4 */ always @(posedge clk) if (n567) n700 <= 1'b0 ? 1'b0 : n7285;
/* FF 17 11  2 */ always @(posedge clk) if (n2076) n2068 <= 1'b0 ? 1'b0 : n7286;
/* FF 19 21  1 */ always @(posedge clk) if (n2164) n2577 <= 1'b0 ? 1'b0 : n7287;
/* FF 19  8  6 */ always @(posedge clk) if (n2451) n2467 <= 1'b0 ? 1'b0 : n7288;
/* FF 23 14  7 */ always @(posedge clk) if (n2551) n3221 <= 1'b0 ? 1'b0 : n7289;
/* FF 24 17  3 */ always @(posedge clk) if (n2123) n3397 <= 1'b0 ? 1'b0 : n7290;
/* FF 28  7  0 */ always @(posedge clk) if (n3488) n3719 <= 1'b0 ? 1'b0 : n7291;
/* FF  3 14  3 */ assign n260 = n7292;
/* FF  9 20  1 */ assign n454 = n7293;
/* FF 27  9  1 */ always @(posedge clk) if (n3621) n3611 <= 1'b0 ? 1'b0 : n7294;
/* FF 12 10  0 */ assign n850 = n7295;
/* FF 26 19  1 */ always @(posedge clk) if (n2730) n3556 <= 1'b0 ? 1'b0 : n7296;
/* FF 14 24  3 */ assign n1697 = n7297;
/* FF 17  5  7 */ assign \rco[182]  = n7298;
/* FF  6 20  5 */ always @(posedge clk) if (n552) n665 <= 1'b0 ? 1'b0 : n7299;
/* FF 20  9  4 */ assign n1460 = n7300;
/* FF 17  8  4 */ assign n2054 = n2259;
/* FF 11 18  3 */ always @(posedge clk) if (n1187) n1182 <= 1'b0 ? 1'b0 : n7301;
/* FF 29 11  3 */ always @(posedge clk) if (n3751) n3842 <= 1'b0 ? 1'b0 : n7302;
/* FF  4 12  4 */ always @(posedge clk) if (n77) n397 <= 1'b0 ? 1'b0 : n7303;
/* FF 22 12  3 */ always @(posedge clk) if (n3029) n3039 <= 1'b0 ? 1'b0 : n7304;
/* FF 10 22  2 */ assign n780 = n7305;
/* FF 21 28  7 */ always @(posedge clk) if (n2196) n2986 <= 1'b0 ? 1'b0 : n7306;
/* FF 13 16  5 */ always @(posedge clk) if (n922) n1482 <= 1'b0 ? 1'b0 : n7307;
/* FF 27  7  6 */ always @(posedge clk) if (n3459) n3601 <= 1'b0 ? 1'b0 : n7308;
/* FF 15 22  2 */ always @(posedge clk) if (n1835) n1848 <= 1'b0 ? 1'b0 : n7309;
/* FF 27 10  5 */ assign \rco[59]  = n3750;
/* FF 13 27  4 */ always @(posedge clk) if (n1532) n1553 <= 1'b0 ? 1'b0 : n7310;
/* FF 18  9  6 */ always @(posedge clk) if (n2055) n2267 <= 1'b0 ? 1'b0 : n7311;
/* FF 18 18  7 */ always @(posedge clk) if (n1825) n2338 <= 1'b0 ? 1'b0 : n7312;
/* FF  3 19  2 */ assign n329 = n7313;
/* FF  6 11  1 */ always @(posedge clk) if (n286) n600 <= 1'b0 ? 1'b0 : n7314;
/* FF 23 18  1 */ always @(posedge clk) if (n2573) n3243 <= 1'b0 ? 1'b0 : n7315;
/* FF 14 10  3 */ always @(posedge clk) if (n1622) n1607 <= 1'b0 ? 1'b0 : n7316;
/* FF 19 17  6 */ always @(posedge clk) if (n2727) n2547 <= 1'b0 ? 1'b0 : n7317;
/* FF  5 17  0 */ always @(posedge clk) if (n2) n524 <= 1'b0 ? 1'b0 : n7318;
/* FF  4 15  6 */ always @(posedge clk) if (n207) n418 <= 1'b0 ? 1'b0 : n7319;
/* FF 10 24  7 */ always @(posedge clk) if (n820) n1079 <= 1'b0 ? 1'b0 : n7320;
/* FF 24 13  6 */ always @(posedge clk) if (n3351) n3366 <= 1'b0 ? 1'b0 : n7321;
/* FF 28 11  7 */ assign n3752 = n7322;
/* FF 27 21  3 */ always @(posedge clk) if (n3421) n3690 <= 1'b0 ? 1'b0 : n7323;
/* FF 10 21  4 */ always @(posedge clk) if (n818) n1062 <= 1'b0 ? 1'b0 : n7324;
/* FF 18  4  0 */ always @(posedge clk) if (n2207) n2213 <= 1'b0 ? 1'b0 : n7325;
/* FF 20 26  3 */ always @(posedge clk) if (n2615) n2808 <= 1'b0 ? 1'b0 : n7326;
/* FF 14 20  4 */ always @(posedge clk) if (n1347) n1680 <= 1'b0 ? 1'b0 : n7327;
/* FF 17 20  3 */ always @(posedge clk) if (n1843) n2139 <= 1'b0 ? 1'b0 : n7328;
/* FF  2 11  0 */ assign n168 = n7329;
/* FF 19 18  0 */ always @(posedge clk) if (n2348) n2554 <= 1'b0 ? 1'b0 : n7330;
/* FF 23 15  4 */ always @(posedge clk) if (n3216) n3226 <= 1'b0 ? 1'b0 : n7331;
/* FF 28  6  3 */ always @(posedge clk) if (n3594) n3714 <= 1'b0 ? 1'b0 : n7332;
/* FF  3 15  0 */ always @(posedge clk) if (n207) n293 <= 1'b0 ? 1'b0 : n7333;
/* FF 21 16  2 */ always @(posedge clk) if (n2551) n2889 <= 1'b0 ? 1'b0 : n7334;
/* FF  9 21  2 */ always @(posedge clk) if (n818) n916 <= 1'b0 ? 1'b0 : n7335;
/* FF 26 18  6 */ assign \rco[35]  = n7336;
/* FF 18 22  4 */ assign n1999 = n7337;
/* FF 20  8  3 */ assign n2670 = n7338;
/* FF  6 23  4 */ always @(posedge clk) if (n360) n691 <= 1'b0 ? 1'b0 : n7339;
/* FF 17  9  7 */ assign \rco[97]  = n7340;
/* FF 11 19  0 */ assign \rco[126]  = n7341;
/* FF 29 12  2 */ always @(posedge clk) if (n3751) n3851 <= 1'b0 ? 1'b0 : n7342;
/* FF 28 20  0 */ assign \rco[171]  = n7343;
/* FF 22 26  5 */ always @(posedge clk) if (n2613) n3138 <= 1'b0 ? 1'b0 : n7344;
/* FF 22 15  2 */ always @(posedge clk) if (n3216) n3060 <= 1'b0 ? 1'b0 : n7345;
/* FF 13 17  6 */ always @(posedge clk) if (n1461) n1489 <= 1'b0 ? 1'b0 : n7346;
/* FF 15 23  1 */ always @(posedge clk) if (n778) n1853 <= 1'b0 ? 1'b0 : n7347;
/* FF 13 28  5 */ always @(posedge clk) if (n1394) n1558 <= 1'b0 ? 1'b0 : n7348;
/* FF 18  8  5 */ always @(posedge clk) if (n2055) n2254 <= 1'b0 ? 1'b0 : n7349;
/* FF 27 11  6 */ always @(posedge clk) if (n3460) n3627 <= 1'b0 ? 1'b0 : n7350;
/* FF 18 21  6 */ always @(posedge clk) if (n2347) n2355 <= 1'b0 ? 1'b0 : n7351;
/* FF  3 16  3 */ always @(posedge clk) if (n197) n306 <= 1'b0 ? 1'b0 : n7352;
/* FF 23 19  2 */ always @(posedge clk) if (n2573) n3252 <= 1'b0 ? 1'b0 : n7353;
/* FF 14  5  2 */ always @(posedge clk) if (n1577) n1573 <= 1'b0 ? 1'b0 : n7354;
/* FF 19 14  7 */ always @(posedge clk) if (n2123) n2518 <= 1'b0 ? 1'b0 : n7355;
/* FF  5 18  1 */ always @(posedge clk) if (n657) n532 <= 1'b0 ? 1'b0 : n7356;
/* FF  4 14  5 */ assign n195 = n7357;
/* FF 19  5  6 */ always @(posedge clk) if (n2230) n2441 <= 1'b0 ? 1'b0 : n7358;
/* FF 10 27  6 */ always @(posedge clk) if (n804) n1098 <= 1'b0 ? 1'b0 : n7359;
/* FF 22 25  1 */ always @(posedge clk) if (n2812) n3126 <= 1'b0 ? 1'b0 : n7360;
/* FF 16 24  7 */ always @(posedge clk) if (n1557) n2001 <= 1'b0 ? 1'b0 : n7361;
/* FF 24 12  1 */ always @(posedge clk) if (n3351) n3354 <= 1'b0 ? 1'b0 : n7362;
/* FF 10 20  7 */ always @(posedge clk) if (n922) n1054 <= 1'b0 ? 1'b0 : n7363;
/* FF 27 18  2 */ always @(posedge clk) if (n3553) n3659 <= 1'b0 ? 1'b0 : n7364;
/* FF 13 14  4 */ always @(posedge clk) if (n1461) n1466 <= 1'b0 ? 1'b0 : n7365;
/* FF 28 10  4 */ always @(posedge clk) if (n3462) n3745 <= 1'b0 ? 1'b0 : n7366;
/* FF 18  7  1 */ assign n2057 = n2460;
/* FF 20 25  2 */ always @(posedge clk) if (n2612) n2800 <= 1'b0 ? 1'b0 : n7367;
/* FF 26 22  3 */ always @(posedge clk) if (n2730) n3572 <= 1'b0 ? 1'b0 : n7368;
/* FF 15  5  5 */ always @(posedge clk) if (n1742) n1583 <= 1'b0 ? 1'b0 : n7369;
/* FF 14 23  5 */ assign n7370 = n1862;
/* FF 14  8  4 */ always @(posedge clk) if (n1741) n1597 <= 1'b0 ? 1'b0 : n7371;
/* FF 17 21  0 */ always @(posedge clk) if (n2347) n2144 <= 1'b0 ? 1'b0 : n7372;
/* FF 19 19  3 */ assign n2562 = n7373;
/* FF 23 12  5 */ always @(posedge clk) if (n3031) n2706 <= 1'b0 ? 1'b0 : n7374;
/* FF 28  5  2 */ always @(posedge clk) if (n3488) n3707 <= 1'b0 ? 1'b0 : n7375;
/* FF  3 12  1 */ always @(posedge clk) if (n168) n278 <= 1'b0 ? 1'b0 : n7376;
/* FF 21 17  1 */ assign \rco[61]  = n7377;
/* FF 30 10  7 */ always @(posedge clk) if (n3892) n3891 <= 1'b0 ? 1'b0 : n7378;
/* FF 12  8  6 */ always @(posedge clk) if (n1131) n1281 <= 1'b0 ? 1'b0 : n7379;
/* FF 26 21  7 */ always @(posedge clk) if (n3421) n3568 <= 1'b0 ? 1'b0 : n7380;
/* FF 15  6  1 */ always @(posedge clk) if (n1744) n1734 <= 1'b0 ? 1'b0 : n7381;
/* FF 17  7  1 */ always @(posedge clk) if (n2045) n2047 <= 1'b0 ? 1'b0 : n7382;
/* FF 18 25  5 */ always @(posedge clk) if (n1878) n2382 <= 1'b0 ? 1'b0 : n7383;
/* FF  6 22  3 */ always @(posedge clk) if (n673) n681 <= 1'b0 ? 1'b0 : n7384;
/* FF 20 15  2 */ always @(posedge clk) if (n2715) n2719 <= 1'b0 ? 1'b0 : n7385;
/* FF 17 10  6 */ always @(posedge clk) if (n2282) n2065 <= 1'b0 ? 1'b0 : n7386;
/* FF 11 16  1 */ always @(posedge clk) if (n891) n1160 <= 1'b0 ? 1'b0 : n7387;
/* FF  1 12  3 */ always @(posedge clk) if (n39) n49 <= 1'b0 ? 1'b0 : n7388;
/* FF  9 13  5 */ always @(posedge clk) if (n629) n858 <= 1'b0 ? 1'b0 : n7389;
/* FF 22 14  5 */ always @(posedge clk) if (n3045) n2729 <= 1'b0 ? 1'b0 : n7390;
/* FF  7  7  4 */ always @(posedge clk) if (n588) n713 <= 1'b0 ? 1'b0 : n7391;
/* FF 13 18  7 */ always @(posedge clk) if (n1205) n1499 <= 1'b0 ? 1'b0 : n7392;
/* FF 27  5  0 */ always @(posedge clk) if (n3594) n3585 <= 1'b0 ? 1'b0 : n7393;
/* FF 18 11  4 */ assign n1936 = n7394;
/* FF 15 20  0 */ always @(posedge clk) if (n1347) n1827 <= 1'b0 ? 1'b0 : n7395;
/* FF 27  8  7 */ always @(posedge clk) if (n3464) n3609 <= 1'b0 ? 1'b0 : n7396;
/* FF 18 20  5 */ assign n736 = n7397;
/* FF 23 16  3 */ assign n2123 = n7398;
/* FF 11 14  0 */ always @(posedge clk) if (n1154) n1146 <= 1'b0 ? 1'b0 : n7399;
/* FF  2 14  4 */ always @(posedge clk) if (n83) n191 <= 1'b0 ? 1'b0 : n7400;
/* FF 16  7  5 */ always @(posedge clk) if (n1743) n1912 <= 1'b0 ? 1'b0 : n7401;
/* FF 19 15  4 */ always @(posedge clk) if (n2715) n2529 <= 1'b0 ? 1'b0 : n7402;
/* FF 23  5  7 */ always @(posedge clk) if (n3158) n3157 <= 1'b0 ? 1'b0 : n7403;
/* FF 16 12  4 */ always @(posedge clk) if (n1771) n1939 <= 1'b0 ? 1'b0 : n7404;
/* FF  5 19  6 */ always @(posedge clk) if (n349) n544 <= 1'b0 ? 1'b0 : n7405;
/* FF  4 13  4 */ assign n78 = n7406;
/* FF 22 24  2 */ always @(posedge clk) if (n3113) n3118 <= 1'b0 ? 1'b0 : n7407;
/* FF 10 26  1 */ assign n567 = n7408;
/* FF 24 11  0 */ assign \rco[64]  = n7409;
/* FF 28  9  5 */ always @(posedge clk) if (n3621) n3516 <= 1'b0 ? 1'b0 : n7410;
/* FF 27 19  1 */ always @(posedge clk) if (n3553) n3668 <= 1'b0 ? 1'b0 : n7411;
/* FF 10 23  6 */ always @(posedge clk) if (n821) n1067 <= 1'b0 ? 1'b0 : n7412;
/* FF  7 21  0 */ assign n118 = n7413;
/* FF  6  7  2 */ always @(posedge clk) if (n570) n573 <= 1'b0 ? 1'b0 : n7414;
/* FF 20 24  5 */ always @(posedge clk) if (n2775) n2793 <= 1'b0 ? 1'b0 : n7415;
/* FF 26  9  2 */ always @(posedge clk) if (n3460) n3500 <= 1'b0 ? 1'b0 : n7416;
/* FF 14 22  2 */ always @(posedge clk) if (n1402) n1689 <= 1'b0 ? 1'b0 : n7417;
/* FF 17  3  6 */ always @(posedge clk) if (n1887) n2031 <= 1'b0 ? 1'b0 : n7418;
/* FF 14 11  5 */ always @(posedge clk) if (n1622) n614 <= 1'b0 ? 1'b0 : n7419;
/* FF  2 13  6 */ always @(posedge clk) if (n83) n186 <= 1'b0 ? 1'b0 : n7420;
/* FF 17 22  1 */ always @(posedge clk) if (n1999) n2153 <= 1'b0 ? 1'b0 : n7421;
/* FF 19 16  2 */ assign n2535 = n7422;
/* FF 23  6  3 */ always @(posedge clk) if (n3158) n3162 <= 1'b0 ? 1'b0 : n7423;
/* FF 11 28  4 */ always @(posedge clk) if (n1384) n1259 <= 1'b0 ? 1'b0 : n7424;
/* FF 16 26  0 */ always @(posedge clk) if (n1557) n2012 <= 1'b0 ? 1'b0 : n7425;
/* FF  4 19  0 */ assign n7426 = n546;
/* FF  3 13  6 */ assign \rco[19]  = n7427;
/* FF 21 18  0 */ always @(posedge clk) if (n2757) n2902 <= 1'b0 ? 1'b0 : n7428;
/* FF 22 10  2 */ always @(posedge clk) if (n2856) n3024 <= 1'b0 ? 1'b0 : n7429;
/* FF  9 23  4 */ always @(posedge clk) if (n819) n929 <= 1'b0 ? 1'b0 : n7430;
/* FF 12 15  7 */ always @(posedge clk) if (n1155) n1303 <= 1'b0 ? 1'b0 : n7431;
/* FF 26 20  4 */ assign n3432 = n3684;
/* FF 18 24  6 */ always @(posedge clk) if (n1878) n2375 <= 1'b0 ? 1'b0 : n7432;
/* FF 20 14  1 */ always @(posedge clk) if (n2682) n2713 <= 1'b0 ? 1'b0 : n7433;
/* FF 19 30  1 */ always @(posedge clk) if (n2592) n2635 <= 1'b0 ? 1'b0 : n7434;
/* FF 16  8  1 */ always @(posedge clk) if (n1625) n1916 <= 1'b0 ? 1'b0 : n7435;
/* FF  1 13  0 */ assign n59 = n7436;
/* FF 24  7  7 */ assign n1601 = n7437;
/* FF  9 14  4 */ always @(posedge clk) if (n629) n863 <= 1'b0 ? 1'b0 : n7438;
/* FF 22  9  4 */ always @(posedge clk) if (n2989) n3018 <= 1'b0 ? 1'b0 : n7439;
/* FF 13 19  0 */ assign \rco[143]  = n7440;
/* FF 18 10  3 */ always @(posedge clk) if (n2282) n2276 <= 1'b0 ? 1'b0 : n7441;
/* FF  2 17  0 */ always @(posedge clk) if (n215) n208 <= 1'b0 ? 1'b0 : n7442;
/* FF 20 28  2 */ assign \rco[192]  = n7443;
/* FF 18 23  4 */ always @(posedge clk) if (n1999) n2366 <= 1'b0 ? 1'b0 : n7444;
/* FF 26  6  0 */ always @(posedge clk) if (n3459) n3473 <= 1'b0 ? 1'b0 : n7445;
/* FF 11 15  3 */ assign n1155 = n7446;
/* FF 23 17  4 */ always @(posedge clk) if (n2540) n3236 <= 1'b0 ? 1'b0 : n7447;
/* FF 14  7  0 */ always @(posedge clk) if (n1743) n1585 <= 1'b0 ? 1'b0 : n7448;
/* FF 16  6  6 */ always @(posedge clk) if (n1744) n1903 <= 1'b0 ? 1'b0 : n7449;
/* FF 19 12  5 */ always @(posedge clk) if (n1936) n2502 <= 1'b0 ? 1'b0 : n7450;
/* FF 23 10  6 */ always @(posedge clk) if (n2697) n3189 <= 1'b0 ? 1'b0 : n7451;
/* FF 19  3  4 */ always @(posedge clk) if (n1887) n2431 <= 1'b0 ? 1'b0 : n7452;
/* FF 22 27  3 */ always @(posedge clk) if (n2970) n3146 <= 1'b0 ? 1'b0 : n7453;
/* FF 10 29  0 */ always @(posedge clk) if (n821) n1109 <= 1'b0 ? 1'b0 : n7454;
/* FF 24 10  3 */ always @(posedge clk) if (n3352) n3343 <= 1'b0 ? 1'b0 : n7455;
/* FF 13  5  1 */ always @(posedge clk) if (n1577) n1411 <= 1'b0 ? 1'b0 : n7456;
/* FF 28  8  2 */ always @(posedge clk) if (n3605) n3728 <= 1'b0 ? 1'b0 : n7457;
/* FF  3  9  3 */ always @(posedge clk) if (n260) n255 <= 1'b0 ? 1'b0 : n7458;
/* FF  7 26  1 */ always @(posedge clk) if (n567) n799 <= 1'b0 ? 1'b0 : n7459;
/* FF  9 19  1 */ always @(posedge clk) if (n454) n902 <= 1'b0 ? 1'b0 : n7460;
/* FF 12 19  2 */ always @(posedge clk) if (n1501) n1330 <= 1'b0 ? 1'b0 : n7461;
/* FF 26  8  1 */ always @(posedge clk) if (n3603) n3491 <= 1'b0 ? 1'b0 : n7462;
/* FF 14 17  3 */ always @(posedge clk) if (n1672) n1657 <= 1'b0 ? 1'b0 : n7463;
/* FF 17 12  7 */ always @(posedge clk) if (n2056) n2084 <= 1'b0 ? 1'b0 : n7464;
/* FF  2 12  5 */ always @(posedge clk) if (n39) n181 <= 1'b0 ? 1'b0 : n7465;
/* FF 23  7  0 */ always @(posedge clk) if (n3006) n3166 <= 1'b0 ? 1'b0 : n7466;
/* FF 11 29  3 */ always @(posedge clk) if (n1384) n1265 <= 1'b0 ? 1'b0 : n7467;
/* FF 24 24  0 */ always @(posedge clk) if (n3112) n3439 <= 1'b0 ? 1'b0 : n7468;
/* FF 16 25  1 */ always @(posedge clk) if (n1557) n2004 <= 1'b0 ? 1'b0 : n7469;
/* FF 21 24  6 */ always @(posedge clk) if (n3113) n2959 <= 1'b0 ? 1'b0 : n7470;
/* FF  4 18  3 */ always @(posedge clk) if (n349) n433 <= 1'b0 ? 1'b0 : n7471;
/* FF  3 10  7 */ always @(posedge clk) if (n251) n269 <= 1'b0 ? 1'b0 : n7472;
/* FF 21 19  7 */ always @(posedge clk) if (n2757) n2917 <= 1'b0 ? 1'b0 : n7473;
/* FF 13 23  5 */ always @(posedge clk) if (n1069) n1529 <= 1'b0 ? 1'b0 : n7474;
/* FF 27 14  4 */ always @(posedge clk) if (n3527) n3645 <= 1'b0 ? 1'b0 : n7475;
/* FF  9 16  5 */ always @(posedge clk) if (n645) n880 <= 1'b0 ? 1'b0 : n7476;
/* FF 12 14  4 */ always @(posedge clk) if (n1154) n1292 <= 1'b0 ? 1'b0 : n7477;
/* FF 26 23  5 */ always @(posedge clk) if (n3703) n2951 <= 1'b0 ? 1'b0 : n7478;
/* FF 18 27  7 */ always @(posedge clk) if (n2020) n2399 <= 1'b0 ? 1'b0 : n7479;
/* FF  6 16  1 */ always @(posedge clk) if (n511) n639 <= 1'b0 ? 1'b0 : n7480;
/* FF  5  8  1 */ always @(posedge clk) if (n21) n469 <= 1'b0 ? 1'b0 : n7481;
/* FF 20 13  0 */ assign n2707 = n7482;
/* FF 19 31  2 */ always @(posedge clk) if (n2592) n2643 <= 1'b0 ? 1'b0 : n7483;
/* FF 23 21  1 */ always @(posedge clk) if (n3258) n3272 <= 1'b0 ? 1'b0 : n7484;
/* FF 16 23  0 */ always @(posedge clk) if (n2000) n1991 <= 1'b0 ? 1'b0 : n7485;
/* FF  1 14  1 */ always @(posedge clk) if (n85) n69 <= 1'b0 ? 1'b0 : n7486;
/* FF 22  7  6 */ always @(posedge clk) if (n2841) n3004 <= 1'b0 ? 1'b0 : n7487;
/* FF 10 17  7 */ assign n817 = n7488;
/* FF  9 15  3 */ always @(posedge clk) if (n645) n870 <= 1'b0 ? 1'b0 : n7489;
/* FF 24  6  4 */ always @(posedge clk) if (n3006) n3325 <= 1'b0 ? 1'b0 : n7490;
/* FF 22  8  7 */ always @(posedge clk) if (n2989) n3015 <= 1'b0 ? 1'b0 : n7491;
/* FF 13 20  1 */ always @(posedge clk) if (n1339) n1504 <= 1'b0 ? 1'b0 : n7492;
/* FF 18 13  2 */ always @(posedge clk) if (n2283) n2297 <= 1'b0 ? 1'b0 : n7493;
/* FF 20 19  3 */ always @(posedge clk) if (n2562) n2752 <= 1'b0 ? 1'b0 : n7494;
/* FF 14 13  6 */ always @(posedge clk) if (n1015) n1629 <= 1'b0 ? 1'b0 : n7495;
/* FF 12 28  0 */ assign \rco[103]  = n7496;
/* FF 23 22  5 */ always @(posedge clk) if (n3422) n3284 <= 1'b0 ? 1'b0 : n7497;
/* FF 14  6  7 */ always @(posedge clk) if (n1577) n1582 <= 1'b0 ? 1'b0 : n7498;
/* FF 16  5  7 */ always @(posedge clk) if (n1742) n1895 <= 1'b0 ? 1'b0 : n7499;
/* FF 17 19  3 */ always @(posedge clk) if (n1982) n2131 <= 1'b0 ? 1'b0 : n7500;
/* FF 19 13  2 */ always @(posedge clk) if (n2283) n2507 <= 1'b0 ? 1'b0 : n7501;
/* FF 23 11  5 */ always @(posedge clk) if (n3031) n3195 <= 1'b0 ? 1'b0 : n7502;
/* FF 16 10  6 */ always @(posedge clk) if (n1771) n1931 <= 1'b0 ? 1'b0 : n7503;
/* FF  5 21  4 */ assign n553 = n7504;
/* FF 10 28  3 */ always @(posedge clk) if (n821) n1104 <= 1'b0 ? 1'b0 : n7505;
/* FF 24  9  2 */ always @(posedge clk) if (n3352) n3334 <= 1'b0 ? 1'b0 : n7506;
/* FF 13  6  0 */ always @(posedge clk) if (n977) n1415 <= 1'b0 ? 1'b0 : n7507;
/* FF 15 24  1 */ always @(posedge clk) if (n778) n1865 <= 1'b0 ? 1'b0 : n7508;
/* FF 21 23  4 */ always @(posedge clk) if (n2961) n2947 <= 1'b0 ? 1'b0 : n7509;
/* FF 26 11  0 */ assign \rco[67]  = n7510;
/* FF 12 18  1 */ always @(posedge clk) if (n1501) n1321 <= 1'b0 ? 1'b0 : n7511;
/* FF 29 19  1 */ always @(posedge clk) if (n3786) n3862 <= 1'b0 ? 1'b0 : n7512;
/* FF 14 16  0 */ always @(posedge clk) if (n1792) n1646 <= 1'b0 ? 1'b0 : n7513;
/* FF 17 13  4 */ always @(posedge clk) if (n2056) n2090 <= 1'b0 ? 1'b0 : n7514;
/* FF 17 16  7 */ assign \rco[29]  = n7515;
/* FF  2 15  4 */ always @(posedge clk) if (n197) n199 <= 1'b0 ? 1'b0 : n7516;
/* FF 11 26  2 */ always @(posedge clk) if (n954) n1238 <= 1'b0 ? 1'b0 : n7517;
/* FF 10 14  0 */ always @(posedge clk) if (n750) n1007 <= 1'b0 ? 1'b0 : n7518;
/* FF 24 23  1 */ always @(posedge clk) if (n3104) n3434 <= 1'b0 ? 1'b0 : n7519;
/* FF 21 25  5 */ always @(posedge clk) if (n2970) n2967 <= 1'b0 ? 1'b0 : n7520;
/* FF  4 17  2 */ always @(posedge clk) if (n2) n426 <= 1'b0 ? 1'b0 : n7521;
/* FF  3 11  4 */ always @(posedge clk) if (n153) n274 <= 1'b0 ? 1'b0 : n7522;
/* FF  7  9  7 */ always @(posedge clk) if (n589) n725 <= 1'b0 ? 1'b0 : n7523;
/* FF 21 20  6 */ always @(posedge clk) if (n3087) n2924 <= 1'b0 ? 1'b0 : n7524;
/* FF  9 17  6 */ always @(posedge clk) if (n1030) n889 <= 1'b0 ? 1'b0 : n7525;
/* FF 18 26  0 */ always @(posedge clk) if (n2615) n2385 <= 1'b0 ? 1'b0 : n7526;
/* FF  6 19  0 */ always @(posedge clk) if (n657) n123 <= 1'b0 ? 1'b0 : n7527;
/* FF 23 26  0 */ always @(posedge clk) if (n2195) n3311 <= 1'b0 ? 1'b0 : n7528;
/* FF 28 19  5 */ always @(posedge clk) if (n3424) n3782 <= 1'b0 ? 1'b0 : n7529;
/* FF 19  9  7 */ always @(posedge clk) if (n2451) n2478 <= 1'b0 ? 1'b0 : n7530;
/* FF 16 22  3 */ always @(posedge clk) if (n1835) n1989 <= 1'b0 ? 1'b0 : n7531;
/* FF 22  6  1 */ always @(posedge clk) if (n2841) n2991 <= 1'b0 ? 1'b0 : n7532;
/* FF 10 16  4 */ always @(posedge clk) if (n891) n1027 <= 1'b0 ? 1'b0 : n7533;
/* FF 22 11  6 */ assign n7534 = n3199;
/* FF 13 21  2 */ always @(posedge clk) if (n1356) n1515 <= 1'b0 ? 1'b0 : n7535;
/* FF 18 12  1 */ always @(posedge clk) if (n1936) n2287 <= 1'b0 ? 1'b0 : n7536;
/* FF  2 19  2 */ assign n216 = n7537;
/* FF  6 13  3 */ always @(posedge clk) if (n78) n618 <= 1'b0 ? 1'b0 : n7538;
/* FF 20 18  0 */ always @(posedge clk) if (n2348) n2741 <= 1'b0 ? 1'b0 : n7539;
/* FF 11  6  4 */ always @(posedge clk) if (en_in) n1122 <= 1'b0 ? 1'b0 : n7540;
/* FF 14 12  5 */ assign n1137 = n7541;
/* FF 23 23  6 */ always @(posedge clk) if (n3104) n3293 <= 1'b0 ? 1'b0 : n7542;
/* FF 11 13  5 */ always @(posedge clk) if (n733) n1143 <= 1'b0 ? 1'b0 : n7543;
/* FF 19 10  3 */ always @(posedge clk) if (n2678) n2482 <= 1'b0 ? 1'b0 : n7544;
/* FF 16  9  7 */ always @(posedge clk) if (n1771) n1925 <= 1'b0 ? 1'b0 : n7545;
/* FF  5 22  5 */ always @(posedge clk) if (n673) n226 <= 1'b0 ? 1'b0 : n7546;
/* FF 28 14  0 */ always @(posedge clk) if (n2085) n3761 <= 1'b0 ? 1'b0 : n7547;
/* FF 15 25  6 */ always @(posedge clk) if (n1878) n1875 <= 1'b0 ? 1'b0 : n7548;
/* FF  3  7  1 */ always @(posedge clk) if (n21) n250 <= 1'b0 ? 1'b0 : n7549;
/* FF  7 13  4 */ assign \rco[160]  = n7550;
/* FF 21  8  5 */ always @(posedge clk) if (n2989) n2840 <= 1'b0 ? 1'b0 : n7551;
/* FF 26 17  6 */ always @(posedge clk) if (n3249) n3552 <= 1'b0 ? 1'b0 : n7552;
/* FF 12 17  0 */ always @(posedge clk) if (n900) n1312 <= 1'b0 ? 1'b0 : n7553;
/* FF 18 30  5 */ always @(posedge clk) if (n1881) n1872 <= 1'b0 ? 1'b0 : n7554;
/* FF 14 19  1 */ assign n1592 = n7555;
/* FF 17 14  5 */ always @(posedge clk) if (n1625) n2099 <= 1'b0 ? 1'b0 : n7556;
/* FF 29 20  0 */ always @(posedge clk) if (n3786) n3868 <= 1'b0 ? 1'b0 : n7557;
/* FF 17 17  4 */ always @(posedge clk) if (n2111) n2118 <= 1'b0 ? 1'b0 : n7558;
/* FF 11 27  1 */ always @(posedge clk) if (n1393) n1248 <= 1'b0 ? 1'b0 : n7559;
/* FF 24 22  2 */ always @(posedge clk) if (n3422) n3427 <= 1'b0 ? 1'b0 : n7560;
/* FF  1 11  3 */ always @(posedge clk) if (n37) n40 <= 1'b0 ? 1'b0 : n7561;
/* FF 31 10  2 */ assign \rco[71]  = n7562;
/* FF 21 26  4 */ always @(posedge clk) if (n2017) n2044 <= 1'b0 ? 1'b0 : n7563;
/* FF  4 16  5 */ always @(posedge clk) if (n79) n425 <= 1'b0 ? 1'b0 : n7564;
/* FF 21 21  5 */ always @(posedge clk) if (n2564) n2931 <= 1'b0 ? 1'b0 : n7565;
/* FF 13 25  7 */ always @(posedge clk) if (n697) n698 <= 1'b0 ? 1'b0 : n7566;
/* FF 27 12  6 */ always @(posedge clk) if (n3368) n3634 <= 1'b0 ? 1'b0 : n7567;
/* FF  9 18  7 */ always @(posedge clk) if (n1030) n899 <= 1'b0 ? 1'b0 : n7568;
/* FF 18 29  1 */ always @(posedge clk) if (n1881) n2409 <= 1'b0 ? 1'b0 : n7569;
/* FF  5 10  3 */ always @(posedge clk) if (n184) n477 <= 1'b0 ? 1'b0 : n7570;
/* FF 19 29  4 */ always @(posedge clk) if (n2614) n2631 <= 1'b0 ? 1'b0 : n7571;
/* FF 11  9  2 */ always @(posedge clk) if (n1131) n1132 <= 1'b0 ? 1'b0 : n7572;
/* FF 23 27  3 */ always @(posedge clk) if (n2017) n3315 <= 1'b0 ? 1'b0 : n7573;
/* FF 19  6  6 */ always @(posedge clk) if (n2241) n2449 <= 1'b0 ? 1'b0 : n7574;
/* FF 10 19  5 */ always @(posedge clk) if (n454) n1046 <= 1'b0 ? 1'b0 : n7575;
/* FF  9  9  1 */ always @(posedge clk) if (n983) n828 <= 1'b0 ? 1'b0 : n7576;
/* FF 13 22  3 */ assign \rco[112]  = n7577;
/* FF 18 15  0 */ assign n2308 = n7578;
/* FF  3 22  1 */ always @(posedge clk) if (n352) n354 <= 1'b0 ? 1'b0 : n7579;
/* FF 21  7  1 */ assign \rco[44]  = n3007;
/* FF  2 18  5 */ always @(posedge clk) if (n115) n214 <= 1'b0 ? 1'b0 : n7580;
/* FF  6 12  0 */ always @(posedge clk) if (n286) n606 <= 1'b0 ? 1'b0 : n7581;
/* FF 20 17  1 */ always @(posedge clk) if (n2727) n2733 <= 1'b0 ? 1'b0 : n7582;
/* FF 26 14  4 */ always @(posedge clk) if (n3527) n3537 <= 1'b0 ? 1'b0 : n7583;
/* FF 14 15  4 */ always @(posedge clk) if (n1792) n1643 <= 1'b0 ? 1'b0 : n7584;
/* FF 23 20  7 */ always @(posedge clk) if (n3258) n3270 <= 1'b0 ? 1'b0 : n7585;
/* FF 16  3  1 */ assign \rco[90]  = n7586;
/* FF 19 11  0 */ always @(posedge clk) if (n2076) n2486 <= 1'b0 ? 1'b0 : n7587;
/* FF 23  9  3 */ always @(posedge clk) if (n2678) n3179 <= 1'b0 ? 1'b0 : n7588;
/* FF  4 20  2 */ assign n440 = n7589;
/* FF 21  9  6 */ always @(posedge clk) if (n2856) n2850 <= 1'b0 ? 1'b0 : n7590;
/* FF  9 27  5 */ always @(posedge clk) if (n804) n951 <= 1'b0 ? 1'b0 : n7591;
/* FF  7 25  4 */ always @(posedge clk) if (n567) n797 <= 1'b0 ? 1'b0 : n7592;
/* FF 21  4  5 */ assign \rco[46]  = n7593;
/* FF 12 16  7 */ always @(posedge clk) if (n1155) n1310 <= 1'b0 ? 1'b0 : n7594;
/* FF 26 13  6 */ always @(posedge clk) if (n3033) n3531 <= 1'b0 ? 1'b0 : n7595;
/* FF 29 21  3 */ always @(posedge clk) if (n3788) n3878 <= 1'b0 ? 1'b0 : n7596;
/* FF 17 15  2 */ always @(posedge clk) if (n2111) n2103 <= 1'b0 ? 1'b0 : n7597;
/* FF 19 25  1 */ always @(posedge clk) if (n2612) n2605 <= 1'b0 ? 1'b0 : n7598;
/* FF 11 24  0 */ always @(posedge clk) if (n796) n1223 <= 1'b0 ? 1'b0 : n7599;
/* FF 24 21  3 */ assign n3411 = n7600;
/* FF 22 13  7 */ always @(posedge clk) if (n2085) n3044 <= 1'b0 ? 1'b0 : n7601;
/* FF 21 27  3 */ always @(posedge clk) if (n2196) n2975 <= 1'b0 ? 1'b0 : n7602;
/* FF  7 15  5 */ assign \rco[25]  = n7603;
/* FF  9 24  1 */ always @(posedge clk) if (n820) n933 <= 1'b0 ? 1'b0 : n7604;
/* FF 13 26  6 */ always @(posedge clk) if (n1271) n1549 <= 1'b0 ? 1'b0 : n7605;
/* FF 21 22  4 */ always @(posedge clk) if (n2384) n2939 <= 1'b0 ? 1'b0 : n7606;
/* FF 14 28  3 */ always @(posedge clk) if (n1402) n1721 <= 1'b0 ? 1'b0 : n7607;
/* FF  2 22  2 */ always @(posedge clk) if (n352) n237 <= 1'b0 ? 1'b0 : n7608;
/* FF 18 28  2 */ always @(posedge clk) if (n2020) n2402 <= 1'b0 ? 1'b0 : n7609;
/* FF 19 26  5 */ assign n2195 = n7610;
/* FF 23 24  2 */ always @(posedge clk) if (n3112) n3298 <= 1'b0 ? 1'b0 : n7611;
/* FF 11 22  3 */ always @(posedge clk) if (n695) n1209 <= 1'b0 ? 1'b0 : n7612;
/* FF 28 17  7 */ always @(posedge clk) if (n3765) n3772 <= 1'b0 ? 1'b0 : n7613;
/* FF 16 15  4 */ always @(posedge clk) if (n739) n1947 <= 1'b0 ? 1'b0 : n7614;
/* FF 19  7  5 */ always @(posedge clk) if (n2670) n2457 <= 1'b0 ? 1'b0 : n7615;
/* FF 16 20  5 */ always @(posedge clk) if (n1843) n1979 <= 1'b0 ? 1'b0 : n7616;
/* FF 10 18  2 */ always @(posedge clk) if (n1187) n1035 <= 1'b0 ? 1'b0 : n7617;
/* FF  9 10  0 */ always @(posedge clk) if (n988) n834 <= 1'b0 ? 1'b0 : n7618;
/* FF 15 18  2 */ always @(posedge clk) if (n1355) n1810 <= 1'b0 ? 1'b0 : n7619;
/* FF 20 27  7 */ always @(posedge clk) if (n2195) n2821 <= 1'b0 ? 1'b0 : n7620;
/* FF  2 21  4 */ always @(posedge clk) if (n126) n231 <= 1'b0 ? 1'b0 : n7621;
/* FF 20 16  6 */ assign n2715 = n7622;
/* FF  6 15  1 */ always @(posedge clk) if (n630) n631 <= 1'b0 ? 1'b0 : n7623;
/* FF 12 20  4 */ assign n922 = n7624;
/* FF 14 14  3 */ always @(posedge clk) if (n1791) n1635 <= 1'b0 ? 1'b0 : n7625;
/* FF 17 11  7 */ always @(posedge clk) if (n2076) n2073 <= 1'b0 ? 1'b0 : n7626;
/* FF 17 30  0 */ always @(posedge clk) if (n2020) n2197 <= 1'b0 ? 1'b0 : n7627;
/* FF 19  8  1 */ always @(posedge clk) if (n2451) n2462 <= 1'b0 ? 1'b0 : n7628;
/* FF 23 14  2 */ assign n3216 = n7629;
/* FF 22 18  0 */ always @(posedge clk) if (n3065) n3080 <= 1'b0 ? 1'b0 : n7630;
/* FF  3 14  6 */ assign \rco[7]  = n411;
/* FF  7 19  6 */ always @(posedge clk) if (n549) n763 <= 1'b0 ? 1'b0 : n7631;
/* FF  9 20  4 */ assign n818 = n7632;
/* FF 21 10  7 */ assign \rco[74]  = n7633;
/* FF 26 19  4 */ always @(posedge clk) if (n2730) n3559 <= 1'b0 ? 1'b0 : n7634;
/* FF 27  9  6 */ always @(posedge clk) if (n3621) n3616 <= 1'b0 ? 1'b0 : n7635;
/* FF 12 23  6 */ always @(posedge clk) if (n1357) n1364 <= 1'b0 ? 1'b0 : n7636;
/* FF 26 12  5 */ always @(posedge clk) if (n3368) n3522 <= 1'b0 ? 1'b0 : n7637;
/* FF 17  8  3 */ assign n1584 = n2258;
/* FF  5 15  1 */ always @(posedge clk) if (n511) n515 <= 1'b0 ? 1'b0 : n7638;

endmodule

